VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 112.465 219.150 113.275 219.290 ;
        RECT 112.275 218.980 113.275 219.150 ;
        RECT 112.465 217.920 113.275 218.980 ;
        RECT 112.465 217.770 113.275 217.910 ;
        RECT 112.275 217.600 113.275 217.770 ;
        RECT 112.465 212.400 113.275 217.600 ;
        RECT 112.465 212.250 113.275 212.390 ;
        RECT 112.275 212.080 113.275 212.250 ;
        RECT 112.465 208.720 113.275 212.080 ;
        RECT 112.305 208.455 112.415 208.575 ;
        RECT 112.465 208.110 113.145 208.250 ;
        RECT 112.275 207.940 113.145 208.110 ;
        RECT 112.465 207.765 113.145 207.940 ;
        RECT 112.465 206.420 113.375 207.765 ;
        RECT 112.550 205.970 113.335 206.400 ;
        RECT 112.305 205.695 112.415 205.815 ;
        RECT 112.465 204.145 113.375 205.490 ;
        RECT 112.465 203.970 113.145 204.145 ;
        RECT 112.275 203.800 113.145 203.970 ;
        RECT 112.465 203.660 113.145 203.800 ;
        RECT 112.465 203.510 113.145 203.650 ;
        RECT 112.275 203.340 113.145 203.510 ;
        RECT 112.465 200.135 113.145 203.340 ;
        RECT 112.465 199.225 113.365 200.135 ;
        RECT 112.465 197.690 113.145 199.225 ;
        RECT 112.465 196.340 113.375 197.690 ;
        RECT 112.465 194.945 113.375 196.290 ;
        RECT 112.465 194.770 113.145 194.945 ;
        RECT 112.275 194.600 113.145 194.770 ;
        RECT 112.465 194.460 113.145 194.600 ;
        RECT 112.310 194.140 112.420 194.300 ;
        RECT 112.550 193.090 113.335 193.520 ;
        RECT 112.310 192.760 112.420 192.920 ;
        RECT 112.465 192.010 113.145 192.150 ;
        RECT 112.275 191.840 113.145 192.010 ;
        RECT 112.465 191.665 113.145 191.840 ;
        RECT 112.465 190.320 113.375 191.665 ;
        RECT 112.465 189.260 113.245 190.310 ;
        RECT 112.275 189.090 113.245 189.260 ;
        RECT 112.465 188.940 113.245 189.090 ;
        RECT 112.310 188.620 112.420 188.780 ;
        RECT 112.465 187.870 113.145 188.010 ;
        RECT 112.275 187.700 113.145 187.870 ;
        RECT 112.465 186.190 113.145 187.700 ;
        RECT 112.465 185.260 113.375 186.190 ;
        RECT 112.305 184.995 112.415 185.115 ;
        RECT 112.465 183.730 113.275 184.790 ;
        RECT 112.275 183.560 113.275 183.730 ;
        RECT 112.465 183.420 113.275 183.560 ;
      LAYER nwell ;
        RECT 113.665 183.225 116.495 219.485 ;
      LAYER pwell ;
        RECT 116.885 219.150 117.695 219.290 ;
        RECT 117.905 219.150 118.715 219.290 ;
        RECT 116.885 218.980 118.715 219.150 ;
        RECT 116.885 217.920 117.695 218.980 ;
        RECT 117.905 217.920 118.715 218.980 ;
        RECT 116.785 216.565 117.695 217.910 ;
        RECT 117.015 216.390 117.695 216.565 ;
        RECT 117.905 216.520 118.815 217.870 ;
        RECT 117.015 216.220 117.885 216.390 ;
        RECT 117.015 216.080 117.695 216.220 ;
        RECT 117.740 215.760 117.850 215.920 ;
        RECT 116.785 214.735 117.695 215.150 ;
        RECT 117.905 214.985 118.585 216.520 ;
        RECT 116.785 214.565 117.885 214.735 ;
        RECT 116.785 214.220 117.695 214.565 ;
        RECT 117.015 211.250 117.695 214.220 ;
        RECT 117.905 214.075 118.805 214.985 ;
        RECT 116.885 210.870 117.695 211.010 ;
        RECT 117.905 210.870 118.585 214.075 ;
        RECT 116.885 210.700 118.585 210.870 ;
        RECT 116.885 207.340 117.695 210.700 ;
        RECT 117.905 210.560 118.585 210.700 ;
        RECT 117.905 210.410 118.715 210.550 ;
        RECT 117.715 210.240 118.715 210.410 ;
        RECT 116.885 207.190 117.695 207.330 ;
        RECT 116.885 207.020 117.885 207.190 ;
        RECT 116.885 205.960 117.695 207.020 ;
        RECT 117.905 206.880 118.715 210.240 ;
        RECT 117.745 206.615 117.855 206.735 ;
        RECT 117.990 205.970 118.775 206.400 ;
        RECT 116.785 204.560 117.695 205.910 ;
        RECT 117.905 205.810 118.585 205.950 ;
        RECT 117.715 205.640 118.585 205.810 ;
        RECT 117.015 203.025 117.695 204.560 ;
        RECT 116.795 202.115 117.695 203.025 ;
        RECT 117.015 198.910 117.695 202.115 ;
        RECT 117.015 198.740 117.885 198.910 ;
        RECT 117.015 198.600 117.695 198.740 ;
        RECT 116.785 198.175 117.695 198.590 ;
        RECT 116.785 198.005 117.885 198.175 ;
        RECT 116.785 197.660 117.695 198.005 ;
        RECT 117.015 194.690 117.695 197.660 ;
        RECT 117.905 196.845 118.585 205.640 ;
        RECT 117.905 196.610 118.715 196.750 ;
        RECT 117.715 196.440 118.715 196.610 ;
        RECT 117.905 195.380 118.715 196.440 ;
        RECT 117.905 195.230 118.685 195.370 ;
        RECT 117.715 195.060 118.685 195.230 ;
        RECT 117.740 194.140 117.850 194.300 ;
        RECT 117.905 194.000 118.685 195.060 ;
        RECT 117.905 193.850 118.685 193.990 ;
        RECT 117.715 193.680 118.685 193.850 ;
        RECT 116.825 193.090 117.610 193.520 ;
        RECT 116.785 192.055 117.695 192.975 ;
        RECT 117.905 192.620 118.685 193.680 ;
        RECT 117.905 192.470 118.685 192.610 ;
        RECT 117.715 192.300 118.685 192.470 ;
        RECT 117.015 189.710 117.695 192.055 ;
        RECT 117.905 191.240 118.685 192.300 ;
        RECT 117.905 191.090 118.685 191.230 ;
        RECT 117.715 190.920 118.685 191.090 ;
        RECT 117.905 189.860 118.685 190.920 ;
        RECT 117.015 189.540 117.885 189.710 ;
        RECT 117.015 189.510 117.695 189.540 ;
        RECT 117.740 189.080 117.850 189.240 ;
        RECT 117.905 188.795 118.815 189.830 ;
        RECT 117.715 188.625 118.815 188.795 ;
        RECT 117.905 188.480 118.815 188.625 ;
        RECT 116.785 186.030 117.695 188.470 ;
        RECT 117.905 188.330 118.815 188.390 ;
        RECT 117.715 188.160 118.815 188.330 ;
        RECT 116.785 185.860 117.885 186.030 ;
        RECT 116.785 185.720 117.695 185.860 ;
        RECT 117.740 185.400 117.850 185.560 ;
        RECT 117.905 184.940 118.815 188.160 ;
        RECT 116.885 183.730 117.695 184.790 ;
        RECT 117.905 183.730 118.715 184.790 ;
        RECT 116.885 183.560 118.715 183.730 ;
        RECT 116.885 183.420 117.695 183.560 ;
        RECT 117.905 183.420 118.715 183.560 ;
      LAYER nwell ;
        RECT 119.105 183.225 121.935 219.485 ;
      LAYER pwell ;
        RECT 122.325 219.150 123.135 219.290 ;
        RECT 123.345 219.150 124.155 219.290 ;
        RECT 122.325 218.980 124.155 219.150 ;
        RECT 122.325 217.920 123.135 218.980 ;
        RECT 123.345 217.920 124.155 218.980 ;
        RECT 122.225 216.565 123.135 217.910 ;
        RECT 123.345 217.770 124.025 217.910 ;
        RECT 123.155 217.600 124.025 217.770 ;
        RECT 122.455 216.390 123.135 216.565 ;
        RECT 122.455 216.220 123.325 216.390 ;
        RECT 122.455 216.080 123.135 216.220 ;
        RECT 123.180 215.760 123.290 215.920 ;
        RECT 122.455 215.010 123.135 215.040 ;
        RECT 122.455 214.840 123.325 215.010 ;
        RECT 122.455 212.495 123.135 214.840 ;
        RECT 122.225 211.575 123.135 212.495 ;
        RECT 123.345 214.395 124.025 217.600 ;
        RECT 123.345 213.485 124.245 214.395 ;
        RECT 123.345 211.950 124.025 213.485 ;
        RECT 123.180 211.160 123.290 211.320 ;
        RECT 123.345 210.600 124.255 211.950 ;
        RECT 122.455 210.410 123.135 210.440 ;
        RECT 123.345 210.410 124.155 210.550 ;
        RECT 122.455 210.240 124.155 210.410 ;
        RECT 122.455 207.895 123.135 210.240 ;
        RECT 122.225 206.975 123.135 207.895 ;
        RECT 123.345 206.880 124.155 210.240 ;
        RECT 122.455 203.670 123.135 206.640 ;
        RECT 123.185 206.615 123.295 206.735 ;
        RECT 123.430 205.970 124.215 206.400 ;
        RECT 123.345 205.810 124.025 205.950 ;
        RECT 123.155 205.640 124.025 205.810 ;
        RECT 122.225 203.325 123.135 203.670 ;
        RECT 122.225 203.155 123.325 203.325 ;
        RECT 122.225 202.740 123.135 203.155 ;
        RECT 122.325 202.590 123.135 202.730 ;
        RECT 122.325 202.420 123.325 202.590 ;
        RECT 123.345 202.435 124.025 205.640 ;
        RECT 122.325 200.900 123.135 202.420 ;
        RECT 123.345 201.525 124.245 202.435 ;
        RECT 122.455 200.750 123.135 200.890 ;
        RECT 122.455 200.580 123.325 200.750 ;
        RECT 122.455 197.375 123.135 200.580 ;
        RECT 123.345 199.990 124.025 201.525 ;
        RECT 123.345 198.640 124.255 199.990 ;
        RECT 123.345 198.445 124.025 198.590 ;
        RECT 123.155 198.275 124.025 198.445 ;
        RECT 122.235 196.465 123.135 197.375 ;
        RECT 122.455 194.930 123.135 196.465 ;
        RECT 123.345 196.745 124.025 198.275 ;
        RECT 123.345 195.380 124.255 196.745 ;
        RECT 123.345 195.230 124.155 195.370 ;
        RECT 123.155 195.060 124.155 195.230 ;
        RECT 122.225 193.580 123.135 194.930 ;
        RECT 122.265 193.090 123.050 193.520 ;
        RECT 122.225 192.655 123.135 193.070 ;
        RECT 122.225 192.485 123.325 192.655 ;
        RECT 123.345 192.620 124.155 195.060 ;
        RECT 122.225 192.140 123.135 192.485 ;
        RECT 123.185 192.355 123.295 192.475 ;
        RECT 122.455 189.170 123.135 192.140 ;
        RECT 123.345 192.010 124.025 192.040 ;
        RECT 123.155 191.840 124.025 192.010 ;
        RECT 123.345 189.495 124.025 191.840 ;
        RECT 122.355 188.790 123.135 188.930 ;
        RECT 122.355 188.620 123.325 188.790 ;
        RECT 122.355 187.560 123.135 188.620 ;
        RECT 123.345 188.575 124.255 189.495 ;
        RECT 123.345 188.330 124.255 188.390 ;
        RECT 123.155 188.160 124.255 188.330 ;
        RECT 122.225 186.605 123.135 187.550 ;
        RECT 122.425 185.115 123.105 186.605 ;
        RECT 123.345 185.390 124.255 188.160 ;
        RECT 122.425 184.945 123.325 185.115 ;
        RECT 122.425 184.800 123.105 184.945 ;
        RECT 122.325 183.730 123.135 184.790 ;
        RECT 123.345 183.730 124.155 184.790 ;
        RECT 122.325 183.560 124.155 183.730 ;
        RECT 122.325 183.420 123.135 183.560 ;
        RECT 123.345 183.420 124.155 183.560 ;
      LAYER nwell ;
        RECT 124.545 183.225 127.375 219.485 ;
      LAYER pwell ;
        RECT 127.765 219.150 128.575 219.290 ;
        RECT 128.785 219.150 129.595 219.290 ;
        RECT 127.765 218.980 129.595 219.150 ;
        RECT 127.765 217.920 128.575 218.980 ;
        RECT 128.785 217.920 129.595 218.980 ;
        RECT 127.665 216.565 128.575 217.910 ;
        RECT 128.785 217.770 129.595 217.910 ;
        RECT 128.595 217.600 129.595 217.770 ;
        RECT 127.895 216.390 128.575 216.565 ;
        RECT 128.785 216.540 129.595 217.600 ;
        RECT 128.785 216.390 129.465 216.420 ;
        RECT 127.895 216.220 129.465 216.390 ;
        RECT 127.895 216.080 128.575 216.220 ;
        RECT 128.625 215.815 128.735 215.935 ;
        RECT 127.665 215.195 128.575 215.610 ;
        RECT 127.665 215.025 128.765 215.195 ;
        RECT 127.665 214.680 128.575 215.025 ;
        RECT 127.895 211.710 128.575 214.680 ;
        RECT 128.785 213.875 129.465 216.220 ;
        RECT 128.785 212.955 129.695 213.875 ;
        RECT 128.785 211.835 129.695 212.755 ;
        RECT 127.895 211.330 128.575 211.470 ;
        RECT 127.895 211.160 128.765 211.330 ;
        RECT 127.895 207.955 128.575 211.160 ;
        RECT 128.785 209.490 129.465 211.835 ;
        RECT 128.595 209.320 129.465 209.490 ;
        RECT 128.785 209.290 129.465 209.320 ;
        RECT 128.785 209.030 129.595 209.170 ;
        RECT 128.595 208.860 129.595 209.030 ;
        RECT 127.675 207.045 128.575 207.955 ;
        RECT 127.895 205.510 128.575 207.045 ;
        RECT 128.785 206.420 129.595 208.860 ;
        RECT 128.870 205.970 129.655 206.400 ;
        RECT 127.665 204.160 128.575 205.510 ;
        RECT 128.785 204.895 129.695 205.930 ;
        RECT 128.595 204.725 129.695 204.895 ;
        RECT 128.785 204.580 129.695 204.725 ;
        RECT 127.665 203.695 128.575 204.110 ;
        RECT 127.665 203.525 128.765 203.695 ;
        RECT 127.665 203.180 128.575 203.525 ;
        RECT 127.895 200.210 128.575 203.180 ;
        RECT 128.785 200.750 129.695 204.500 ;
        RECT 128.595 200.580 129.695 200.750 ;
        RECT 128.785 200.440 129.695 200.580 ;
        RECT 127.665 198.955 128.575 199.875 ;
        RECT 127.895 196.610 128.575 198.955 ;
        RECT 128.785 199.415 129.695 200.335 ;
        RECT 128.785 197.070 129.465 199.415 ;
        RECT 128.595 196.900 129.465 197.070 ;
        RECT 128.785 196.870 129.465 196.900 ;
        RECT 128.785 196.610 129.595 196.750 ;
        RECT 127.895 196.440 129.595 196.610 ;
        RECT 127.895 196.410 128.575 196.440 ;
        RECT 127.765 196.150 128.575 196.290 ;
        RECT 127.765 195.980 128.765 196.150 ;
        RECT 127.765 193.540 128.575 195.980 ;
        RECT 128.785 195.380 129.595 196.440 ;
        RECT 128.785 194.420 129.695 195.370 ;
        RECT 127.705 193.090 128.490 193.520 ;
        RECT 127.665 190.175 128.575 192.780 ;
        RECT 128.815 192.015 129.495 194.420 ;
        RECT 128.595 191.845 129.495 192.015 ;
        RECT 128.815 191.700 129.495 191.845 ;
        RECT 128.785 191.545 129.695 191.690 ;
        RECT 128.595 191.375 129.695 191.545 ;
        RECT 128.785 190.340 129.695 191.375 ;
        RECT 127.665 190.160 128.765 190.175 ;
        RECT 128.785 190.160 129.565 190.310 ;
        RECT 127.665 190.005 129.565 190.160 ;
        RECT 127.665 189.860 128.575 190.005 ;
        RECT 128.595 189.990 129.565 190.005 ;
        RECT 128.620 189.540 128.730 189.700 ;
        RECT 128.785 188.940 129.565 189.990 ;
        RECT 127.665 185.570 128.575 188.790 ;
        RECT 128.785 185.570 129.695 188.790 ;
        RECT 127.665 185.400 129.695 185.570 ;
        RECT 127.665 185.340 128.575 185.400 ;
        RECT 128.785 185.340 129.695 185.400 ;
        RECT 128.625 184.995 128.735 185.115 ;
        RECT 127.765 183.730 128.575 184.790 ;
        RECT 128.785 183.730 129.595 184.790 ;
        RECT 127.765 183.560 129.595 183.730 ;
        RECT 127.765 183.420 128.575 183.560 ;
        RECT 128.785 183.420 129.595 183.560 ;
      LAYER nwell ;
        RECT 129.985 183.225 132.815 219.485 ;
      LAYER pwell ;
        RECT 133.205 219.150 134.015 219.290 ;
        RECT 134.225 219.150 135.035 219.290 ;
        RECT 133.205 218.980 135.035 219.150 ;
        RECT 133.205 217.920 134.015 218.980 ;
        RECT 134.225 217.920 135.035 218.980 ;
        RECT 133.105 216.520 134.015 217.870 ;
        RECT 134.225 217.495 135.135 217.910 ;
        RECT 134.035 217.325 135.135 217.495 ;
        RECT 133.335 214.985 134.015 216.520 ;
        RECT 133.115 214.075 134.015 214.985 ;
        RECT 133.335 210.870 134.015 214.075 ;
        RECT 134.225 216.980 135.135 217.325 ;
        RECT 134.225 214.010 134.905 216.980 ;
        RECT 134.225 213.630 134.905 213.770 ;
        RECT 134.035 213.460 134.905 213.630 ;
        RECT 133.335 210.700 134.205 210.870 ;
        RECT 133.335 210.560 134.015 210.700 ;
        RECT 133.205 210.410 134.015 210.550 ;
        RECT 133.205 210.240 134.205 210.410 ;
        RECT 134.225 210.255 134.905 213.460 ;
        RECT 133.205 207.800 134.015 210.240 ;
        RECT 134.225 209.345 135.125 210.255 ;
        RECT 134.225 207.810 134.905 209.345 ;
        RECT 134.065 207.535 134.175 207.655 ;
        RECT 133.335 207.190 134.015 207.330 ;
        RECT 133.335 207.020 134.205 207.190 ;
        RECT 133.335 198.225 134.015 207.020 ;
        RECT 134.225 206.460 135.135 207.810 ;
        RECT 134.310 205.970 135.095 206.400 ;
        RECT 134.225 205.810 134.905 205.950 ;
        RECT 134.035 205.640 134.905 205.810 ;
        RECT 134.225 202.435 134.905 205.640 ;
        RECT 134.225 201.525 135.125 202.435 ;
        RECT 134.225 199.990 134.905 201.525 ;
        RECT 134.225 198.640 135.135 199.990 ;
        RECT 134.065 198.335 134.175 198.455 ;
        RECT 133.105 197.115 134.015 198.035 ;
        RECT 133.335 194.770 134.015 197.115 ;
        RECT 134.225 196.765 135.135 198.130 ;
        RECT 134.225 195.235 134.905 196.765 ;
        RECT 134.035 195.065 134.905 195.235 ;
        RECT 134.225 194.920 134.905 195.065 ;
        RECT 133.335 194.600 134.205 194.770 ;
        RECT 133.335 194.570 134.015 194.600 ;
        RECT 134.060 194.140 134.170 194.300 ;
        RECT 134.225 193.850 135.135 193.910 ;
        RECT 134.035 193.680 135.135 193.850 ;
        RECT 133.145 193.090 133.930 193.520 ;
        RECT 133.305 192.935 133.985 193.060 ;
        RECT 133.305 192.765 134.205 192.935 ;
        RECT 133.305 191.735 133.985 192.765 ;
        RECT 133.105 190.780 134.015 191.735 ;
        RECT 134.225 190.910 135.135 193.680 ;
        RECT 133.205 190.630 134.015 190.770 ;
        RECT 133.205 190.625 134.205 190.630 ;
        RECT 134.225 190.625 135.135 190.770 ;
        RECT 133.205 190.460 135.135 190.625 ;
        RECT 133.205 188.020 134.015 190.460 ;
        RECT 134.035 190.455 135.135 190.460 ;
        RECT 134.225 189.420 135.135 190.455 ;
        RECT 134.065 189.135 134.175 189.255 ;
        RECT 134.225 188.790 135.135 188.850 ;
        RECT 134.035 188.620 135.135 188.790 ;
        RECT 134.065 187.755 134.175 187.875 ;
        RECT 133.105 186.495 134.015 187.530 ;
        RECT 133.105 186.325 134.205 186.495 ;
        RECT 133.105 186.180 134.015 186.325 ;
        RECT 133.235 185.110 134.015 186.170 ;
        RECT 134.225 185.400 135.135 188.620 ;
        RECT 134.065 185.110 134.175 185.115 ;
        RECT 133.235 184.940 134.205 185.110 ;
        RECT 133.235 184.800 134.015 184.940 ;
        RECT 133.205 183.730 134.015 184.790 ;
        RECT 134.225 183.730 135.035 184.790 ;
        RECT 133.205 183.560 135.035 183.730 ;
        RECT 133.205 183.420 134.015 183.560 ;
        RECT 134.225 183.420 135.035 183.560 ;
      LAYER nwell ;
        RECT 135.425 183.225 138.255 219.485 ;
      LAYER pwell ;
        RECT 138.645 219.150 139.455 219.290 ;
        RECT 139.665 219.150 140.475 219.290 ;
        RECT 138.645 218.980 140.475 219.150 ;
        RECT 138.645 217.920 139.455 218.980 ;
        RECT 139.665 217.920 140.475 218.980 ;
        RECT 138.545 216.565 139.455 217.910 ;
        RECT 139.665 217.770 140.345 217.910 ;
        RECT 139.475 217.600 140.345 217.770 ;
        RECT 138.775 216.390 139.455 216.565 ;
        RECT 138.775 216.220 139.645 216.390 ;
        RECT 138.775 216.080 139.455 216.220 ;
        RECT 138.545 215.655 139.455 216.070 ;
        RECT 138.545 215.485 139.645 215.655 ;
        RECT 138.545 215.140 139.455 215.485 ;
        RECT 138.775 212.170 139.455 215.140 ;
        RECT 139.665 214.395 140.345 217.600 ;
        RECT 139.665 213.485 140.565 214.395 ;
        RECT 139.665 211.950 140.345 213.485 ;
        RECT 138.645 211.790 139.455 211.930 ;
        RECT 138.645 211.620 139.645 211.790 ;
        RECT 138.645 210.560 139.455 211.620 ;
        RECT 139.665 210.600 140.575 211.950 ;
        RECT 138.775 201.670 139.455 210.465 ;
        RECT 139.665 209.535 140.575 210.455 ;
        RECT 139.665 207.190 140.345 209.535 ;
        RECT 139.475 207.020 140.345 207.190 ;
        RECT 139.665 206.990 140.345 207.020 ;
        RECT 139.505 206.615 139.615 206.735 ;
        RECT 139.750 205.970 140.535 206.400 ;
        RECT 139.665 205.535 140.575 205.950 ;
        RECT 139.475 205.365 140.575 205.535 ;
        RECT 139.665 205.020 140.575 205.365 ;
        RECT 139.665 202.050 140.345 205.020 ;
        RECT 139.505 201.670 139.615 201.675 ;
        RECT 138.775 201.500 139.645 201.670 ;
        RECT 138.775 201.360 139.455 201.500 ;
        RECT 138.545 200.335 139.455 201.255 ;
        RECT 139.475 201.205 139.645 201.210 ;
        RECT 139.475 201.040 140.345 201.205 ;
        RECT 138.775 197.990 139.455 200.335 ;
        RECT 139.665 200.300 140.345 201.040 ;
        RECT 139.665 199.370 140.575 200.300 ;
        RECT 139.665 197.990 140.575 199.040 ;
        RECT 138.775 197.820 140.575 197.990 ;
        RECT 138.775 197.790 139.455 197.820 ;
        RECT 139.665 197.690 140.575 197.820 ;
        RECT 138.645 197.530 139.455 197.670 ;
        RECT 139.665 197.530 140.345 197.670 ;
        RECT 138.645 197.360 140.345 197.530 ;
        RECT 138.645 196.300 139.455 197.360 ;
        RECT 138.745 196.145 139.425 196.290 ;
        RECT 138.745 195.975 139.645 196.145 ;
        RECT 138.745 194.485 139.425 195.975 ;
        RECT 138.545 193.540 139.455 194.485 ;
        RECT 139.665 194.155 140.345 197.360 ;
        RECT 138.585 193.090 139.370 193.520 ;
        RECT 139.665 193.245 140.565 194.155 ;
        RECT 138.545 192.930 139.455 192.990 ;
        RECT 138.545 192.760 139.645 192.930 ;
        RECT 138.545 189.540 139.455 192.760 ;
        RECT 139.665 191.710 140.345 193.245 ;
        RECT 139.665 190.360 140.575 191.710 ;
        RECT 139.505 190.055 139.615 190.175 ;
        RECT 139.475 189.705 139.645 189.710 ;
        RECT 139.475 189.540 140.345 189.705 ;
        RECT 138.545 189.250 139.455 189.310 ;
        RECT 138.545 189.080 139.645 189.250 ;
        RECT 138.545 185.860 139.455 189.080 ;
        RECT 139.665 188.800 140.345 189.540 ;
        RECT 139.665 187.870 140.575 188.800 ;
        RECT 139.665 187.410 140.445 187.550 ;
        RECT 139.475 187.240 140.445 187.410 ;
        RECT 139.665 186.180 140.445 187.240 ;
        RECT 139.500 185.400 139.610 185.560 ;
        RECT 139.665 185.120 140.445 186.170 ;
        RECT 139.475 184.950 140.445 185.120 ;
        RECT 139.665 184.800 140.445 184.950 ;
        RECT 138.645 183.730 139.455 184.790 ;
        RECT 139.665 183.730 140.475 184.790 ;
        RECT 138.645 183.560 140.475 183.730 ;
        RECT 138.645 183.420 139.455 183.560 ;
        RECT 139.665 183.420 140.475 183.560 ;
      LAYER nwell ;
        RECT 140.865 183.225 143.695 219.485 ;
      LAYER pwell ;
        RECT 144.085 219.150 144.895 219.290 ;
        RECT 145.105 219.150 145.915 219.290 ;
        RECT 144.085 218.980 145.915 219.150 ;
        RECT 144.085 217.920 144.895 218.980 ;
        RECT 145.105 217.920 145.915 218.980 ;
        RECT 144.085 217.770 144.895 217.910 ;
        RECT 145.105 217.770 145.915 217.910 ;
        RECT 144.085 217.600 145.915 217.770 ;
        RECT 144.085 214.240 144.895 217.600 ;
        RECT 144.945 213.975 145.055 214.095 ;
        RECT 143.985 212.380 144.895 213.730 ;
        RECT 145.105 212.400 145.915 217.600 ;
        RECT 144.215 210.845 144.895 212.380 ;
        RECT 144.950 212.080 145.060 212.240 ;
        RECT 145.105 211.330 145.785 211.470 ;
        RECT 144.915 211.160 145.785 211.330 ;
        RECT 143.995 209.935 144.895 210.845 ;
        RECT 144.215 206.730 144.895 209.935 ;
        RECT 145.105 210.985 145.785 211.160 ;
        RECT 145.105 209.640 146.015 210.985 ;
        RECT 145.105 206.730 146.015 209.500 ;
        RECT 144.215 206.560 146.015 206.730 ;
        RECT 144.215 206.420 144.895 206.560 ;
        RECT 145.105 206.500 146.015 206.560 ;
        RECT 144.215 206.270 144.895 206.410 ;
        RECT 144.215 206.100 145.085 206.270 ;
        RECT 144.215 202.895 144.895 206.100 ;
        RECT 145.190 205.970 145.975 206.400 ;
        RECT 144.950 205.640 145.060 205.800 ;
        RECT 145.105 204.890 145.785 204.920 ;
        RECT 144.915 204.720 145.785 204.890 ;
        RECT 143.995 201.985 144.895 202.895 ;
        RECT 144.215 200.450 144.895 201.985 ;
        RECT 145.105 202.375 145.785 204.720 ;
        RECT 145.105 201.455 146.015 202.375 ;
        RECT 144.950 201.040 145.060 201.200 ;
        RECT 143.985 199.100 144.895 200.450 ;
        RECT 145.105 199.085 146.015 200.430 ;
        RECT 145.105 198.910 145.785 199.085 ;
        RECT 144.915 198.740 145.785 198.910 ;
        RECT 143.985 197.810 144.895 198.740 ;
        RECT 145.105 198.600 145.785 198.740 ;
        RECT 145.105 198.450 145.785 198.480 ;
        RECT 144.915 198.280 145.785 198.450 ;
        RECT 144.215 197.070 144.895 197.810 ;
        RECT 144.215 196.905 145.085 197.070 ;
        RECT 144.915 196.900 145.085 196.905 ;
        RECT 144.215 196.610 144.895 196.750 ;
        RECT 144.215 196.440 145.085 196.610 ;
        RECT 144.215 196.265 144.895 196.440 ;
        RECT 143.985 194.920 144.895 196.265 ;
        RECT 145.105 195.935 145.785 198.280 ;
        RECT 145.105 195.015 146.015 195.935 ;
        RECT 143.985 194.770 144.895 194.900 ;
        RECT 143.985 194.760 145.085 194.770 ;
        RECT 145.105 194.760 145.885 194.910 ;
        RECT 143.985 194.600 145.885 194.760 ;
        RECT 143.985 193.550 144.895 194.600 ;
        RECT 144.915 194.590 145.885 194.600 ;
        RECT 145.105 193.540 145.885 194.590 ;
        RECT 144.025 193.090 144.810 193.520 ;
        RECT 145.190 193.090 145.975 193.520 ;
        RECT 143.985 192.930 144.895 192.990 ;
        RECT 143.985 192.760 145.085 192.930 ;
        RECT 143.985 189.990 144.895 192.760 ;
        RECT 145.105 190.805 146.015 192.150 ;
        RECT 145.105 190.630 145.785 190.805 ;
        RECT 144.915 190.460 145.785 190.630 ;
        RECT 145.105 190.320 145.785 190.460 ;
        RECT 145.105 190.170 145.915 190.310 ;
        RECT 144.915 190.000 145.915 190.170 ;
        RECT 144.215 189.710 144.895 189.740 ;
        RECT 144.215 189.540 145.085 189.710 ;
        RECT 144.215 187.195 144.895 189.540 ;
        RECT 145.105 188.940 145.915 190.000 ;
        RECT 145.105 187.870 145.885 188.930 ;
        RECT 144.915 187.700 145.885 187.870 ;
        RECT 145.105 187.560 145.885 187.700 ;
        RECT 143.985 186.275 144.895 187.195 ;
        RECT 145.105 186.490 145.885 187.550 ;
        RECT 144.915 186.320 145.885 186.490 ;
        RECT 145.105 186.180 145.885 186.320 ;
        RECT 144.115 185.120 144.895 186.170 ;
        RECT 145.105 185.120 145.885 186.170 ;
        RECT 144.115 184.950 145.885 185.120 ;
        RECT 144.115 184.800 144.895 184.950 ;
        RECT 145.105 184.800 145.885 184.950 ;
        RECT 144.085 183.730 144.895 184.790 ;
        RECT 145.105 183.730 145.915 184.790 ;
        RECT 144.085 183.560 145.915 183.730 ;
        RECT 144.085 183.420 144.895 183.560 ;
        RECT 145.105 183.420 145.915 183.560 ;
      LAYER nwell ;
        RECT 146.305 183.225 147.910 219.485 ;
      LAYER pwell ;
        RECT 100.450 167.190 106.550 176.980 ;
        RECT 100.450 167.160 106.560 167.190 ;
        RECT 100.650 166.760 101.810 167.160 ;
        RECT 103.770 165.080 106.560 167.160 ;
      LAYER nwell ;
        RECT 101.660 162.970 106.500 165.080 ;
        RECT 107.780 164.740 117.970 176.990 ;
      LAYER pwell ;
        RECT 120.330 167.140 126.430 176.930 ;
        RECT 120.330 167.110 126.440 167.140 ;
        RECT 120.530 166.710 121.690 167.110 ;
        RECT 123.650 165.030 126.440 167.110 ;
      LAYER nwell ;
        RECT 121.540 162.920 126.380 165.030 ;
        RECT 127.660 164.690 137.850 176.940 ;
      LAYER pwell ;
        RECT 140.360 167.190 146.460 176.980 ;
        RECT 140.360 167.160 146.470 167.190 ;
        RECT 140.560 166.760 141.720 167.160 ;
        RECT 143.680 165.080 146.470 167.160 ;
      LAYER nwell ;
        RECT 141.570 162.970 146.410 165.080 ;
        RECT 147.690 164.740 157.880 176.990 ;
      LAYER pwell ;
        RECT 100.450 152.190 106.550 161.980 ;
        RECT 100.450 152.160 106.560 152.190 ;
        RECT 100.650 151.760 101.810 152.160 ;
        RECT 103.770 150.080 106.560 152.160 ;
      LAYER nwell ;
        RECT 101.660 147.970 106.500 150.080 ;
        RECT 107.780 149.740 117.970 161.990 ;
      LAYER pwell ;
        RECT 120.330 152.190 126.430 161.980 ;
        RECT 120.330 152.160 126.440 152.190 ;
        RECT 120.530 151.760 121.690 152.160 ;
        RECT 123.650 150.080 126.440 152.160 ;
      LAYER nwell ;
        RECT 121.540 147.970 126.380 150.080 ;
        RECT 127.660 149.740 137.850 161.990 ;
      LAYER pwell ;
        RECT 140.410 152.140 146.510 161.930 ;
        RECT 140.410 152.110 146.520 152.140 ;
        RECT 140.610 151.710 141.770 152.110 ;
        RECT 143.730 150.030 146.520 152.110 ;
      LAYER nwell ;
        RECT 141.620 147.920 146.460 150.030 ;
        RECT 147.740 149.690 157.930 161.940 ;
      LAYER pwell ;
        RECT 100.450 137.140 106.550 146.930 ;
        RECT 100.450 137.110 106.560 137.140 ;
        RECT 100.650 136.710 101.810 137.110 ;
        RECT 103.770 135.030 106.560 137.110 ;
      LAYER nwell ;
        RECT 101.660 132.920 106.500 135.030 ;
        RECT 107.780 134.690 117.970 146.940 ;
      LAYER pwell ;
        RECT 120.330 137.140 126.430 146.930 ;
        RECT 120.330 137.110 126.440 137.140 ;
        RECT 120.530 136.710 121.690 137.110 ;
        RECT 123.650 135.030 126.440 137.110 ;
      LAYER nwell ;
        RECT 121.540 132.920 126.380 135.030 ;
        RECT 127.660 134.690 137.850 146.940 ;
      LAYER pwell ;
        RECT 140.360 137.140 146.460 146.930 ;
        RECT 140.360 137.110 146.470 137.140 ;
        RECT 140.560 136.710 141.720 137.110 ;
        RECT 143.680 135.030 146.470 137.110 ;
      LAYER nwell ;
        RECT 141.570 132.920 146.410 135.030 ;
        RECT 147.690 134.690 157.880 146.940 ;
      LAYER pwell ;
        RECT 100.450 122.140 106.550 131.930 ;
        RECT 100.450 122.110 106.560 122.140 ;
        RECT 100.650 121.710 101.810 122.110 ;
        RECT 103.770 120.030 106.560 122.110 ;
      LAYER nwell ;
        RECT 101.660 117.920 106.500 120.030 ;
        RECT 107.780 119.690 117.970 131.940 ;
      LAYER pwell ;
        RECT 120.330 122.200 126.430 131.990 ;
        RECT 120.330 122.170 126.440 122.200 ;
        RECT 120.530 121.770 121.690 122.170 ;
        RECT 123.650 120.090 126.440 122.170 ;
      LAYER nwell ;
        RECT 121.540 117.980 126.380 120.090 ;
        RECT 127.660 119.750 137.850 132.000 ;
      LAYER pwell ;
        RECT 140.360 122.200 146.460 131.990 ;
        RECT 140.360 122.170 146.470 122.200 ;
        RECT 140.560 121.770 141.720 122.170 ;
        RECT 143.680 120.090 146.470 122.170 ;
      LAYER nwell ;
        RECT 141.570 117.980 146.410 120.090 ;
        RECT 147.690 119.750 157.880 132.000 ;
      LAYER pwell ;
        RECT 100.400 107.200 106.500 116.990 ;
        RECT 100.400 107.170 106.510 107.200 ;
        RECT 100.600 106.770 101.760 107.170 ;
        RECT 103.720 105.090 106.510 107.170 ;
      LAYER nwell ;
        RECT 101.610 102.980 106.450 105.090 ;
        RECT 107.730 104.750 117.920 117.000 ;
      LAYER pwell ;
        RECT 120.330 107.200 126.430 116.990 ;
        RECT 120.330 107.170 126.440 107.200 ;
        RECT 120.530 106.770 121.690 107.170 ;
        RECT 123.650 105.090 126.440 107.170 ;
      LAYER nwell ;
        RECT 121.540 102.980 126.380 105.090 ;
        RECT 127.660 104.750 137.850 117.000 ;
      LAYER pwell ;
        RECT 140.360 107.200 146.460 116.990 ;
        RECT 140.360 107.170 146.470 107.200 ;
        RECT 140.560 106.770 141.720 107.170 ;
        RECT 143.680 105.090 146.470 107.170 ;
      LAYER nwell ;
        RECT 141.570 102.980 146.410 105.090 ;
        RECT 147.690 104.750 157.880 117.000 ;
      LAYER li1 ;
        RECT 112.275 219.210 112.445 219.295 ;
        RECT 114.995 219.210 115.165 219.295 ;
        RECT 117.715 219.210 117.885 219.295 ;
        RECT 120.435 219.210 120.605 219.295 ;
        RECT 123.155 219.210 123.325 219.295 ;
        RECT 125.875 219.210 126.045 219.295 ;
        RECT 128.595 219.210 128.765 219.295 ;
        RECT 131.315 219.210 131.485 219.295 ;
        RECT 134.035 219.210 134.205 219.295 ;
        RECT 136.755 219.210 136.925 219.295 ;
        RECT 139.475 219.210 139.645 219.295 ;
        RECT 142.195 219.210 142.365 219.295 ;
        RECT 144.915 219.210 145.085 219.295 ;
        RECT 147.635 219.210 147.805 219.295 ;
        RECT 112.275 218.690 113.735 219.210 ;
        RECT 112.275 218.000 113.195 218.690 ;
        RECT 113.905 218.520 116.255 219.210 ;
        RECT 116.425 218.690 119.175 219.210 ;
        RECT 113.365 218.000 116.795 218.520 ;
        RECT 116.965 218.000 118.635 218.690 ;
        RECT 119.345 218.520 121.695 219.210 ;
        RECT 121.865 218.690 124.615 219.210 ;
        RECT 118.805 218.000 122.235 218.520 ;
        RECT 122.405 218.000 124.075 218.690 ;
        RECT 124.785 218.520 127.135 219.210 ;
        RECT 127.305 218.690 130.055 219.210 ;
        RECT 124.245 218.000 127.675 218.520 ;
        RECT 127.845 218.000 129.515 218.690 ;
        RECT 130.225 218.520 132.575 219.210 ;
        RECT 132.745 218.690 135.495 219.210 ;
        RECT 129.685 218.000 133.115 218.520 ;
        RECT 133.285 218.000 134.955 218.690 ;
        RECT 135.665 218.520 138.015 219.210 ;
        RECT 138.185 218.690 140.935 219.210 ;
        RECT 135.125 218.000 138.555 218.520 ;
        RECT 138.725 218.000 140.395 218.690 ;
        RECT 141.105 218.520 143.455 219.210 ;
        RECT 143.625 218.690 146.375 219.210 ;
        RECT 140.565 218.000 143.995 218.520 ;
        RECT 144.165 218.000 145.835 218.690 ;
        RECT 146.545 218.520 147.805 219.210 ;
        RECT 146.005 218.000 147.805 218.520 ;
        RECT 112.275 217.830 112.445 218.000 ;
        RECT 114.995 217.830 115.165 218.000 ;
        RECT 112.275 216.245 112.990 217.830 ;
        RECT 114.560 217.825 115.165 217.830 ;
        RECT 117.715 217.825 117.885 218.000 ;
        RECT 114.560 217.565 116.315 217.825 ;
        RECT 116.875 217.565 117.885 217.825 ;
        RECT 118.540 217.780 119.375 217.830 ;
        RECT 114.560 216.965 115.165 217.565 ;
        RECT 115.335 217.220 117.545 217.390 ;
        RECT 115.335 217.135 116.240 217.220 ;
        RECT 116.970 217.135 117.545 217.220 ;
        RECT 117.715 217.280 117.885 217.565 ;
        RECT 118.105 217.770 119.375 217.780 ;
        RECT 120.435 217.825 120.605 218.000 ;
        RECT 123.155 217.825 123.325 218.000 ;
        RECT 125.875 217.825 126.045 218.000 ;
        RECT 128.595 217.830 128.765 218.000 ;
        RECT 131.315 217.830 131.485 218.000 ;
        RECT 128.595 217.825 130.055 217.830 ;
        RECT 118.105 217.660 120.220 217.770 ;
        RECT 118.105 217.605 118.665 217.660 ;
        RECT 119.245 217.615 120.220 217.660 ;
        RECT 118.105 217.450 118.625 217.605 ;
        RECT 117.715 217.110 118.495 217.280 ;
        RECT 116.475 216.965 116.805 217.050 ;
        RECT 117.715 216.965 117.885 217.110 ;
        RECT 114.560 216.635 115.925 216.965 ;
        RECT 116.095 216.795 117.165 216.965 ;
        RECT 112.275 215.905 113.820 216.245 ;
        RECT 112.275 212.485 112.990 215.905 ;
        RECT 114.560 214.560 115.165 216.635 ;
        RECT 116.095 216.420 116.265 216.795 ;
        RECT 115.335 216.250 116.265 216.420 ;
        RECT 116.445 216.160 116.815 216.515 ;
        RECT 116.995 216.420 117.165 216.795 ;
        RECT 117.335 216.635 117.885 216.965 ;
        RECT 118.795 216.940 119.125 217.490 ;
        RECT 119.295 217.440 120.220 217.615 ;
        RECT 120.435 217.565 121.755 217.825 ;
        RECT 122.315 217.565 123.325 217.825 ;
        RECT 123.585 217.570 124.045 217.740 ;
        RECT 120.435 217.270 120.605 217.565 ;
        RECT 123.155 217.400 123.325 217.565 ;
        RECT 119.425 217.100 120.605 217.270 ;
        RECT 120.775 217.220 122.985 217.390 ;
        RECT 120.775 217.135 121.680 217.220 ;
        RECT 122.410 217.135 122.985 217.220 ;
        RECT 116.995 216.250 117.545 216.420 ;
        RECT 117.715 216.350 117.885 216.635 ;
        RECT 118.100 216.930 119.125 216.940 ;
        RECT 120.435 216.965 120.605 217.100 ;
        RECT 123.155 217.070 123.705 217.400 ;
        RECT 123.875 217.305 124.045 217.570 ;
        RECT 124.215 217.475 124.865 217.825 ;
        RECT 125.035 217.570 125.705 217.740 ;
        RECT 125.035 217.305 125.205 217.570 ;
        RECT 125.875 217.565 127.195 217.825 ;
        RECT 127.755 217.565 130.055 217.825 ;
        RECT 125.875 217.400 126.045 217.565 ;
        RECT 123.875 217.075 125.205 217.305 ;
        RECT 125.375 217.070 126.045 217.400 ;
        RECT 126.215 217.220 128.425 217.390 ;
        RECT 126.215 217.135 127.120 217.220 ;
        RECT 127.850 217.135 128.425 217.220 ;
        RECT 128.595 217.310 130.055 217.565 ;
        RECT 121.915 216.965 122.245 217.050 ;
        RECT 123.155 216.965 123.325 217.070 ;
        RECT 118.100 216.740 120.265 216.930 ;
        RECT 118.100 216.610 118.625 216.740 ;
        RECT 119.330 216.590 120.265 216.740 ;
        RECT 120.435 216.635 121.365 216.965 ;
        RECT 121.535 216.795 122.605 216.965 ;
        RECT 117.715 216.140 118.415 216.350 ;
        RECT 115.335 214.895 117.545 215.065 ;
        RECT 115.335 214.730 116.305 214.895 ;
        RECT 116.975 214.810 117.545 214.895 ;
        RECT 116.475 214.640 116.805 214.725 ;
        RECT 117.715 214.640 117.885 216.140 ;
        RECT 118.795 215.865 119.125 216.570 ;
        RECT 119.330 216.035 119.705 216.590 ;
        RECT 120.435 216.360 120.605 216.635 ;
        RECT 121.535 216.420 121.705 216.795 ;
        RECT 119.935 216.045 120.605 216.360 ;
        RECT 120.775 216.250 121.705 216.420 ;
        RECT 121.885 216.160 122.255 216.515 ;
        RECT 122.435 216.420 122.605 216.795 ;
        RECT 122.775 216.635 123.325 216.965 ;
        RECT 125.875 216.965 126.045 217.070 ;
        RECT 127.355 216.965 127.685 217.050 ;
        RECT 128.595 216.965 129.515 217.310 ;
        RECT 130.225 217.270 131.485 217.830 ;
        RECT 132.545 217.780 133.380 217.830 ;
        RECT 132.545 217.770 133.815 217.780 ;
        RECT 131.700 217.660 133.815 217.770 ;
        RECT 131.700 217.615 132.675 217.660 ;
        RECT 131.700 217.440 132.625 217.615 ;
        RECT 133.255 217.605 133.815 217.660 ;
        RECT 130.225 217.140 132.495 217.270 ;
        RECT 123.585 216.715 125.705 216.900 ;
        RECT 123.155 216.460 123.325 216.635 ;
        RECT 125.875 216.635 126.805 216.965 ;
        RECT 126.975 216.795 128.045 216.965 ;
        RECT 122.435 216.250 122.985 216.420 ;
        RECT 123.155 216.210 123.785 216.460 ;
        RECT 123.955 216.265 124.905 216.545 ;
        RECT 125.875 216.475 126.045 216.635 ;
        RECT 125.415 216.210 126.045 216.475 ;
        RECT 126.975 216.420 127.145 216.795 ;
        RECT 126.215 216.250 127.145 216.420 ;
        RECT 118.165 215.695 120.135 215.865 ;
        RECT 118.165 215.080 118.335 215.695 ;
        RECT 118.505 215.205 119.795 215.525 ;
        RECT 118.505 215.060 118.835 215.205 ;
        RECT 114.560 214.425 116.305 214.560 ;
        RECT 116.475 214.470 117.145 214.640 ;
        RECT 113.310 214.390 116.305 214.425 ;
        RECT 113.310 214.075 115.165 214.390 ;
        RECT 116.475 214.220 116.805 214.245 ;
        RECT 114.560 212.485 115.165 214.075 ;
        RECT 112.275 212.310 112.445 212.485 ;
        RECT 114.995 212.310 115.165 212.485 ;
        RECT 112.275 210.660 113.735 212.310 ;
        RECT 113.905 212.020 115.165 212.310 ;
        RECT 115.335 214.050 116.805 214.220 ;
        RECT 115.335 212.360 115.505 214.050 ;
        RECT 116.975 213.885 117.145 214.470 ;
        RECT 117.315 214.325 117.885 214.640 ;
        RECT 118.165 214.675 118.335 214.910 ;
        RECT 119.045 214.845 119.765 215.035 ;
        RECT 119.965 214.980 120.135 215.695 ;
        RECT 119.935 214.675 120.265 214.755 ;
        RECT 118.165 214.505 120.265 214.675 ;
        RECT 117.315 214.310 118.385 214.325 ;
        RECT 117.715 213.955 118.385 214.310 ;
        RECT 118.565 214.045 118.865 214.505 ;
        RECT 120.435 214.500 120.605 216.045 ;
        RECT 120.775 214.670 121.455 214.955 ;
        RECT 120.435 214.335 121.065 214.500 ;
        RECT 119.045 214.165 119.375 214.335 ;
        RECT 119.635 214.230 121.065 214.335 ;
        RECT 119.635 214.165 120.605 214.230 ;
        RECT 116.975 213.880 117.545 213.885 ;
        RECT 115.675 213.710 117.545 213.880 ;
        RECT 115.675 212.755 115.845 213.710 ;
        RECT 116.015 213.370 116.985 213.540 ;
        RECT 116.015 212.720 116.185 213.370 ;
        RECT 117.180 213.355 117.545 213.710 ;
        RECT 117.205 213.165 117.375 213.170 ;
        RECT 116.385 212.890 117.545 213.165 ;
        RECT 116.015 212.530 117.545 212.720 ;
        RECT 115.335 212.190 116.360 212.360 ;
        RECT 117.715 212.350 117.885 213.955 ;
        RECT 118.565 213.845 118.895 214.045 ;
        RECT 119.115 213.995 119.375 214.165 ;
        RECT 119.115 213.825 120.160 213.995 ;
        RECT 119.115 213.635 119.285 213.825 ;
        RECT 118.165 213.465 119.285 213.635 ;
        RECT 118.165 212.960 118.335 213.465 ;
        RECT 119.455 213.295 119.820 213.655 ;
        RECT 118.535 213.125 119.820 213.295 ;
        RECT 118.535 212.770 118.755 213.125 ;
        RECT 118.165 212.600 118.335 212.765 ;
        RECT 118.925 212.715 119.520 212.955 ;
        RECT 119.990 212.890 120.160 213.825 ;
        RECT 118.165 212.545 118.605 212.600 ;
        RECT 119.710 212.545 120.265 212.680 ;
        RECT 118.165 212.430 120.265 212.545 ;
        RECT 120.435 212.440 120.605 214.165 ;
        RECT 121.235 214.210 121.455 214.670 ;
        RECT 121.625 214.380 122.185 215.070 ;
        RECT 122.355 214.670 122.985 214.955 ;
        RECT 122.355 214.210 122.525 214.670 ;
        RECT 123.155 214.515 123.325 216.210 ;
        RECT 123.915 216.040 125.280 216.095 ;
        RECT 123.605 215.925 125.705 216.040 ;
        RECT 123.605 215.870 124.045 215.925 ;
        RECT 123.605 215.705 123.775 215.870 ;
        RECT 125.150 215.790 125.705 215.925 ;
        RECT 123.605 215.005 123.775 215.510 ;
        RECT 123.975 215.345 124.195 215.700 ;
        RECT 124.365 215.515 124.960 215.755 ;
        RECT 123.975 215.175 125.260 215.345 ;
        RECT 123.605 214.835 124.725 215.005 ;
        RECT 124.555 214.645 124.725 214.835 ;
        RECT 124.895 214.815 125.260 215.175 ;
        RECT 125.430 214.645 125.600 215.580 ;
        RECT 123.155 214.500 123.825 214.515 ;
        RECT 122.695 214.230 123.825 214.500 ;
        RECT 121.235 214.000 122.525 214.210 ;
        RECT 123.155 214.145 123.825 214.230 ;
        RECT 124.005 214.425 124.335 214.625 ;
        RECT 124.555 214.475 125.600 214.645 ;
        RECT 125.875 215.020 126.045 216.210 ;
        RECT 127.325 216.160 127.695 216.515 ;
        RECT 127.875 216.420 128.045 216.795 ;
        RECT 128.215 216.635 129.515 216.965 ;
        RECT 128.595 216.620 129.515 216.635 ;
        RECT 129.685 217.100 132.495 217.140 ;
        RECT 129.685 216.620 131.485 217.100 ;
        RECT 132.795 216.940 133.125 217.490 ;
        RECT 133.295 217.450 133.815 217.605 ;
        RECT 134.035 217.400 134.205 218.000 ;
        RECT 136.755 217.825 136.925 218.000 ;
        RECT 139.475 217.825 139.645 218.000 ;
        RECT 142.195 217.830 142.365 218.000 ;
        RECT 144.915 217.830 145.085 218.000 ;
        RECT 147.635 217.830 147.805 218.000 ;
        RECT 134.375 217.655 136.585 217.825 ;
        RECT 134.375 217.570 134.945 217.655 ;
        RECT 135.615 217.490 136.585 217.655 ;
        RECT 136.755 217.565 138.075 217.825 ;
        RECT 138.635 217.565 139.645 217.825 ;
        RECT 139.905 217.570 140.365 217.740 ;
        RECT 135.115 217.400 135.445 217.485 ;
        RECT 134.035 217.280 134.605 217.400 ;
        RECT 133.425 217.110 134.605 217.280 ;
        RECT 134.035 217.070 134.605 217.110 ;
        RECT 134.775 217.230 135.445 217.400 ;
        RECT 136.755 217.320 136.925 217.565 ;
        RECT 139.475 217.400 139.645 217.565 ;
        RECT 132.795 216.930 133.820 216.940 ;
        RECT 127.875 216.250 128.425 216.420 ;
        RECT 128.595 215.880 128.765 216.620 ;
        RECT 128.935 216.050 129.565 216.335 ;
        RECT 128.595 215.610 129.225 215.880 ;
        RECT 126.215 215.355 128.425 215.525 ;
        RECT 126.215 215.190 127.185 215.355 ;
        RECT 127.855 215.270 128.425 215.355 ;
        RECT 127.355 215.100 127.685 215.185 ;
        RECT 128.595 215.100 128.765 215.610 ;
        RECT 129.395 215.590 129.565 216.050 ;
        RECT 129.735 215.760 130.295 216.450 ;
        RECT 131.315 216.360 131.485 216.620 ;
        RECT 131.655 216.740 133.820 216.930 ;
        RECT 131.655 216.590 132.590 216.740 ;
        RECT 133.295 216.610 133.820 216.740 ;
        RECT 130.465 216.050 131.145 216.335 ;
        RECT 130.465 215.590 130.685 216.050 ;
        RECT 131.315 216.045 131.985 216.360 ;
        RECT 131.315 215.880 131.485 216.045 ;
        RECT 132.215 216.035 132.590 216.590 ;
        RECT 130.855 215.610 131.485 215.880 ;
        RECT 132.795 215.865 133.125 216.570 ;
        RECT 134.035 216.350 134.205 217.070 ;
        RECT 134.775 216.645 134.945 217.230 ;
        RECT 135.615 217.150 136.925 217.320 ;
        RECT 135.115 216.980 135.445 217.005 ;
        RECT 135.115 216.810 136.585 216.980 ;
        RECT 133.505 216.140 134.205 216.350 ;
        RECT 129.395 215.380 130.685 215.590 ;
        RECT 125.875 214.850 127.185 215.020 ;
        RECT 127.355 214.930 128.025 215.100 ;
        RECT 120.775 213.430 122.985 213.830 ;
        RECT 120.775 212.960 121.455 213.240 ;
        RECT 121.235 212.565 121.455 212.960 ;
        RECT 121.625 212.735 122.185 213.430 ;
        RECT 122.355 212.960 122.985 213.240 ;
        RECT 122.355 212.565 122.525 212.960 ;
        RECT 118.475 212.375 119.840 212.430 ;
        RECT 113.905 211.850 115.925 212.020 ;
        RECT 113.905 210.930 115.165 211.850 ;
        RECT 115.515 211.440 115.925 211.615 ;
        RECT 116.170 211.610 116.360 212.190 ;
        RECT 116.735 211.620 116.905 212.330 ;
        RECT 117.180 212.260 117.885 212.350 ;
        RECT 120.435 212.260 121.065 212.440 ;
        RECT 117.180 212.010 118.345 212.260 ;
        RECT 117.180 211.840 117.885 212.010 ;
        RECT 118.515 211.925 119.465 212.205 ;
        RECT 119.975 212.115 121.065 212.260 ;
        RECT 121.235 212.115 122.525 212.565 ;
        RECT 123.155 212.440 123.325 214.145 ;
        RECT 124.005 213.965 124.305 214.425 ;
        RECT 124.555 214.305 124.815 214.475 ;
        RECT 125.875 214.305 126.045 214.850 ;
        RECT 127.355 214.680 127.685 214.705 ;
        RECT 124.485 214.135 124.815 214.305 ;
        RECT 125.075 214.135 126.045 214.305 ;
        RECT 123.605 213.795 125.705 213.965 ;
        RECT 123.605 213.560 123.775 213.795 ;
        RECT 125.375 213.715 125.705 213.795 ;
        RECT 124.485 213.435 125.205 213.625 ;
        RECT 123.605 212.775 123.775 213.390 ;
        RECT 123.945 213.265 124.275 213.410 ;
        RECT 123.945 212.945 125.235 213.265 ;
        RECT 125.405 212.775 125.575 213.490 ;
        RECT 123.605 212.605 125.575 212.775 ;
        RECT 122.695 212.330 123.325 212.440 ;
        RECT 122.695 212.120 123.855 212.330 ;
        RECT 122.695 212.115 123.325 212.120 ;
        RECT 119.975 211.995 120.605 212.115 ;
        RECT 121.915 212.010 122.245 212.115 ;
        RECT 116.735 211.440 117.510 211.620 ;
        RECT 115.515 211.375 117.510 211.440 ;
        RECT 117.715 211.400 117.885 211.840 ;
        RECT 118.145 211.570 120.265 211.755 ;
        RECT 120.435 211.400 120.605 211.995 ;
        RECT 120.775 211.840 121.745 211.945 ;
        RECT 122.415 211.840 122.985 211.945 ;
        RECT 120.775 211.560 122.985 211.840 ;
        RECT 115.515 211.100 116.905 211.375 ;
        RECT 117.715 211.070 118.265 211.400 ;
        RECT 118.435 211.165 119.765 211.395 ;
        RECT 117.715 210.930 117.885 211.070 ;
        RECT 112.275 208.800 113.215 210.660 ;
        RECT 113.905 210.490 116.255 210.930 ;
        RECT 113.385 209.110 116.255 210.490 ;
        RECT 116.425 210.470 117.885 210.930 ;
        RECT 118.435 210.900 118.605 211.165 ;
        RECT 118.145 210.730 118.605 210.900 ;
        RECT 118.775 210.645 119.425 210.995 ;
        RECT 119.595 210.900 119.765 211.165 ;
        RECT 119.935 211.070 120.605 211.400 ;
        RECT 119.595 210.730 120.265 210.900 ;
        RECT 120.435 210.470 120.605 211.070 ;
        RECT 123.155 211.360 123.325 212.115 ;
        RECT 124.235 211.900 124.565 212.605 ;
        RECT 125.875 212.480 126.045 214.135 ;
        RECT 126.215 214.510 127.685 214.680 ;
        RECT 126.215 212.820 126.385 214.510 ;
        RECT 127.855 214.345 128.025 214.930 ;
        RECT 128.195 214.770 128.765 215.100 ;
        RECT 128.935 214.810 131.145 215.210 ;
        RECT 127.855 214.340 128.425 214.345 ;
        RECT 126.555 214.170 128.425 214.340 ;
        RECT 126.555 213.215 126.725 214.170 ;
        RECT 126.895 213.830 127.865 214.000 ;
        RECT 126.895 213.180 127.065 213.830 ;
        RECT 128.060 213.815 128.425 214.170 ;
        RECT 128.595 213.820 128.765 214.770 ;
        RECT 128.935 214.340 129.565 214.620 ;
        RECT 129.395 213.945 129.565 214.340 ;
        RECT 129.735 214.115 130.295 214.810 ;
        RECT 130.465 214.340 131.145 214.620 ;
        RECT 130.465 213.945 130.685 214.340 ;
        RECT 128.085 213.625 128.255 213.630 ;
        RECT 127.265 213.350 128.425 213.625 ;
        RECT 128.595 213.495 129.225 213.820 ;
        RECT 129.395 213.495 130.685 213.945 ;
        RECT 131.315 214.335 131.485 215.610 ;
        RECT 131.785 215.695 133.755 215.865 ;
        RECT 131.785 214.980 131.955 215.695 ;
        RECT 132.125 215.205 133.415 215.525 ;
        RECT 133.085 215.060 133.415 215.205 ;
        RECT 133.585 215.080 133.755 215.695 ;
        RECT 134.035 215.110 134.205 216.140 ;
        RECT 134.375 216.640 134.945 216.645 ;
        RECT 134.375 216.470 136.245 216.640 ;
        RECT 134.375 216.115 134.740 216.470 ;
        RECT 134.935 216.130 135.905 216.300 ;
        RECT 134.545 215.925 134.715 215.930 ;
        RECT 134.375 215.650 135.535 215.925 ;
        RECT 135.735 215.480 135.905 216.130 ;
        RECT 136.075 215.515 136.245 216.470 ;
        RECT 134.375 215.290 135.905 215.480 ;
        RECT 136.415 215.120 136.585 216.810 ;
        RECT 132.155 214.845 132.875 215.035 ;
        RECT 131.655 214.675 131.985 214.755 ;
        RECT 133.585 214.675 133.755 214.910 ;
        RECT 131.655 214.505 133.755 214.675 ;
        RECT 134.035 214.600 134.740 215.110 ;
        RECT 131.315 214.165 132.285 214.335 ;
        RECT 132.545 214.165 132.875 214.335 ;
        RECT 131.315 213.820 131.485 214.165 ;
        RECT 132.545 213.995 132.805 214.165 ;
        RECT 133.055 214.045 133.355 214.505 ;
        RECT 134.035 214.325 134.205 214.600 ;
        RECT 135.015 214.380 135.185 215.090 ;
        RECT 130.855 213.495 131.485 213.820 ;
        RECT 126.895 212.990 128.425 213.180 ;
        RECT 126.215 212.650 127.240 212.820 ;
        RECT 128.595 212.810 128.765 213.495 ;
        RECT 129.675 213.390 130.005 213.495 ;
        RECT 128.935 213.220 129.505 213.325 ;
        RECT 130.175 213.220 131.145 213.325 ;
        RECT 128.935 212.940 131.145 213.220 ;
        RECT 124.770 211.880 125.145 212.435 ;
        RECT 125.875 212.425 126.805 212.480 ;
        RECT 125.375 212.310 126.805 212.425 ;
        RECT 125.375 212.110 126.045 212.310 ;
        RECT 123.540 211.730 124.065 211.860 ;
        RECT 124.770 211.730 125.705 211.880 ;
        RECT 123.540 211.540 125.705 211.730 ;
        RECT 123.540 211.530 124.565 211.540 ;
        RECT 123.155 211.190 123.935 211.360 ;
        RECT 123.155 210.470 123.325 211.190 ;
        RECT 123.545 210.865 124.065 211.020 ;
        RECT 124.235 210.980 124.565 211.530 ;
        RECT 125.875 211.370 126.045 212.110 ;
        RECT 126.395 211.900 126.805 212.075 ;
        RECT 127.050 212.070 127.240 212.650 ;
        RECT 127.615 212.080 127.785 212.790 ;
        RECT 128.060 212.300 128.765 212.810 ;
        RECT 128.935 212.490 131.145 212.770 ;
        RECT 128.935 212.385 129.505 212.490 ;
        RECT 130.175 212.385 131.145 212.490 ;
        RECT 128.595 212.215 128.765 212.300 ;
        RECT 129.675 212.215 130.005 212.320 ;
        RECT 131.315 212.260 131.485 213.495 ;
        RECT 131.760 213.825 132.805 213.995 ;
        RECT 133.025 213.845 133.355 214.045 ;
        RECT 133.535 213.955 134.205 214.325 ;
        RECT 134.410 214.200 135.185 214.380 ;
        RECT 135.560 214.950 136.585 215.120 ;
        RECT 136.755 216.965 136.925 217.150 ;
        RECT 137.095 217.220 139.305 217.390 ;
        RECT 137.095 217.135 138.000 217.220 ;
        RECT 138.730 217.135 139.305 217.220 ;
        RECT 139.475 217.070 140.025 217.400 ;
        RECT 140.195 217.305 140.365 217.570 ;
        RECT 140.535 217.475 141.185 217.825 ;
        RECT 141.355 217.570 142.025 217.740 ;
        RECT 141.355 217.305 141.525 217.570 ;
        RECT 142.195 217.400 143.455 217.830 ;
        RECT 140.195 217.075 141.525 217.305 ;
        RECT 141.695 217.070 143.455 217.400 ;
        RECT 138.235 216.965 138.565 217.050 ;
        RECT 139.475 216.965 139.645 217.070 ;
        RECT 136.755 216.635 137.685 216.965 ;
        RECT 137.855 216.795 138.925 216.965 ;
        RECT 136.755 215.480 136.925 216.635 ;
        RECT 137.855 216.420 138.025 216.795 ;
        RECT 137.095 216.250 138.025 216.420 ;
        RECT 138.205 216.160 138.575 216.515 ;
        RECT 138.755 216.420 138.925 216.795 ;
        RECT 139.095 216.635 139.645 216.965 ;
        RECT 139.905 216.715 142.025 216.900 ;
        RECT 139.475 216.460 139.645 216.635 ;
        RECT 138.755 216.250 139.305 216.420 ;
        RECT 139.475 216.210 140.105 216.460 ;
        RECT 140.275 216.265 141.225 216.545 ;
        RECT 142.195 216.475 143.455 217.070 ;
        RECT 141.735 216.210 143.455 216.475 ;
        RECT 137.095 215.815 139.305 215.985 ;
        RECT 137.095 215.650 138.065 215.815 ;
        RECT 138.735 215.730 139.305 215.815 ;
        RECT 138.235 215.560 138.565 215.645 ;
        RECT 139.475 215.560 139.645 216.210 ;
        RECT 140.235 216.040 141.600 216.095 ;
        RECT 139.925 215.925 142.025 216.040 ;
        RECT 139.925 215.870 140.365 215.925 ;
        RECT 139.925 215.705 140.095 215.870 ;
        RECT 141.470 215.790 142.025 215.925 ;
        RECT 142.195 216.010 143.455 216.210 ;
        RECT 143.625 216.245 145.630 217.830 ;
        RECT 143.625 216.180 146.460 216.245 ;
        RECT 136.755 215.310 138.065 215.480 ;
        RECT 138.235 215.390 138.905 215.560 ;
        RECT 135.560 214.370 135.750 214.950 ;
        RECT 136.755 214.780 136.925 215.310 ;
        RECT 138.235 215.140 138.565 215.165 ;
        RECT 135.995 214.610 136.925 214.780 ;
        RECT 135.995 214.200 136.405 214.375 ;
        RECT 134.410 214.135 136.405 214.200 ;
        RECT 131.760 212.890 131.930 213.825 ;
        RECT 132.100 213.295 132.465 213.655 ;
        RECT 132.635 213.635 132.805 213.825 ;
        RECT 132.635 213.465 133.755 213.635 ;
        RECT 132.100 213.125 133.385 213.295 ;
        RECT 132.400 212.715 132.995 212.955 ;
        RECT 133.165 212.770 133.385 213.125 ;
        RECT 133.585 212.960 133.755 213.465 ;
        RECT 134.035 213.260 134.205 213.955 ;
        RECT 135.015 213.860 136.405 214.135 ;
        RECT 134.465 213.430 134.925 213.600 ;
        RECT 134.035 212.930 134.585 213.260 ;
        RECT 134.755 213.165 134.925 213.430 ;
        RECT 135.095 213.335 135.745 213.685 ;
        RECT 135.915 213.430 136.585 213.600 ;
        RECT 135.915 213.165 136.085 213.430 ;
        RECT 136.755 213.260 136.925 214.610 ;
        RECT 134.755 212.935 136.085 213.165 ;
        RECT 136.255 212.940 136.925 213.260 ;
        RECT 137.095 214.970 138.565 215.140 ;
        RECT 137.095 213.280 137.265 214.970 ;
        RECT 138.735 214.805 138.905 215.390 ;
        RECT 139.075 215.230 139.645 215.560 ;
        RECT 138.735 214.800 139.305 214.805 ;
        RECT 137.435 214.630 139.305 214.800 ;
        RECT 137.435 213.675 137.605 214.630 ;
        RECT 137.775 214.290 138.745 214.460 ;
        RECT 137.775 213.640 137.945 214.290 ;
        RECT 138.940 214.275 139.305 214.630 ;
        RECT 139.475 214.515 139.645 215.230 ;
        RECT 139.925 215.005 140.095 215.510 ;
        RECT 140.295 215.345 140.515 215.700 ;
        RECT 140.685 215.515 141.280 215.755 ;
        RECT 140.295 215.175 141.580 215.345 ;
        RECT 139.925 214.835 141.045 215.005 ;
        RECT 140.875 214.645 141.045 214.835 ;
        RECT 141.215 214.815 141.580 215.175 ;
        RECT 141.750 214.645 141.920 215.580 ;
        RECT 139.475 214.145 140.145 214.515 ;
        RECT 140.325 214.425 140.655 214.625 ;
        RECT 140.875 214.475 141.920 214.645 ;
        RECT 138.965 214.085 139.135 214.090 ;
        RECT 138.145 213.810 139.305 214.085 ;
        RECT 137.775 213.450 139.305 213.640 ;
        RECT 137.095 213.110 138.120 213.280 ;
        RECT 139.475 213.270 139.645 214.145 ;
        RECT 140.325 213.965 140.625 214.425 ;
        RECT 140.875 214.305 141.135 214.475 ;
        RECT 142.195 214.320 143.975 216.010 ;
        RECT 144.145 215.905 146.460 216.180 ;
        RECT 144.145 214.320 145.630 215.905 ;
        RECT 147.200 214.425 147.805 217.830 ;
        RECT 142.195 214.305 142.365 214.320 ;
        RECT 140.805 214.135 141.135 214.305 ;
        RECT 141.395 214.135 142.365 214.305 ;
        RECT 139.925 213.795 142.025 213.965 ;
        RECT 139.925 213.560 140.095 213.795 ;
        RECT 141.695 213.715 142.025 213.795 ;
        RECT 140.805 213.435 141.525 213.625 ;
        RECT 136.255 212.930 137.685 212.940 ;
        RECT 131.655 212.545 132.210 212.680 ;
        RECT 133.585 212.600 133.755 212.765 ;
        RECT 133.315 212.545 133.755 212.600 ;
        RECT 131.655 212.430 133.755 212.545 ;
        RECT 132.080 212.375 133.445 212.430 ;
        RECT 134.035 212.320 134.205 212.930 ;
        RECT 136.755 212.770 137.685 212.930 ;
        RECT 134.465 212.575 136.585 212.760 ;
        RECT 134.035 212.260 134.665 212.320 ;
        RECT 131.315 212.215 131.945 212.260 ;
        RECT 127.615 211.900 128.390 212.080 ;
        RECT 126.395 211.835 128.390 211.900 ;
        RECT 128.595 211.890 129.225 212.215 ;
        RECT 126.395 211.560 127.785 211.835 ;
        RECT 124.865 211.200 126.045 211.370 ;
        RECT 123.545 210.810 124.105 210.865 ;
        RECT 124.735 210.855 125.660 211.030 ;
        RECT 124.685 210.810 125.660 210.855 ;
        RECT 123.545 210.700 125.660 210.810 ;
        RECT 125.875 210.960 126.045 211.200 ;
        RECT 126.215 211.130 126.885 211.300 ;
        RECT 123.545 210.690 124.815 210.700 ;
        RECT 123.980 210.640 124.815 210.690 ;
        RECT 125.875 210.630 126.545 210.960 ;
        RECT 126.715 210.865 126.885 211.130 ;
        RECT 127.055 211.035 127.705 211.385 ;
        RECT 127.875 211.130 128.335 211.300 ;
        RECT 127.875 210.865 128.045 211.130 ;
        RECT 128.595 210.960 128.765 211.890 ;
        RECT 129.395 211.765 130.685 212.215 ;
        RECT 130.855 211.995 131.945 212.215 ;
        RECT 130.855 211.890 131.485 211.995 ;
        RECT 132.455 211.925 133.405 212.205 ;
        RECT 133.575 212.070 134.665 212.260 ;
        RECT 134.835 212.125 135.785 212.405 ;
        RECT 136.755 212.335 136.925 212.770 ;
        RECT 136.295 212.070 136.925 212.335 ;
        RECT 133.575 212.010 134.205 212.070 ;
        RECT 129.395 211.370 129.565 211.765 ;
        RECT 128.935 211.090 129.565 211.370 ;
        RECT 126.715 210.635 128.045 210.865 ;
        RECT 128.215 210.630 128.765 210.960 ;
        RECT 129.735 210.900 130.295 211.595 ;
        RECT 130.465 211.370 130.685 211.765 ;
        RECT 131.315 211.400 131.485 211.890 ;
        RECT 131.655 211.570 133.775 211.755 ;
        RECT 134.035 211.400 134.205 212.010 ;
        RECT 134.795 211.900 136.160 211.955 ;
        RECT 134.485 211.785 136.585 211.900 ;
        RECT 134.485 211.730 134.925 211.785 ;
        RECT 134.485 211.565 134.655 211.730 ;
        RECT 136.030 211.650 136.585 211.785 ;
        RECT 136.755 211.850 136.925 212.070 ;
        RECT 137.275 212.360 137.685 212.535 ;
        RECT 137.930 212.530 138.120 213.110 ;
        RECT 138.495 212.540 138.665 213.250 ;
        RECT 138.940 212.760 139.645 213.270 ;
        RECT 138.495 212.360 139.270 212.540 ;
        RECT 137.275 212.295 139.270 212.360 ;
        RECT 139.475 212.330 139.645 212.760 ;
        RECT 139.925 212.775 140.095 213.390 ;
        RECT 140.265 213.265 140.595 213.410 ;
        RECT 140.265 212.945 141.555 213.265 ;
        RECT 141.725 212.775 141.895 213.490 ;
        RECT 139.925 212.605 141.895 212.775 ;
        RECT 142.195 213.130 142.365 214.135 ;
        RECT 143.425 213.640 144.260 213.690 ;
        RECT 143.425 213.630 144.695 213.640 ;
        RECT 142.580 213.520 144.695 213.630 ;
        RECT 142.580 213.475 143.555 213.520 ;
        RECT 142.580 213.300 143.505 213.475 ;
        RECT 144.135 213.465 144.695 213.520 ;
        RECT 142.195 212.960 143.375 213.130 ;
        RECT 137.275 212.020 138.665 212.295 ;
        RECT 139.475 212.120 140.175 212.330 ;
        RECT 139.475 211.850 139.645 212.120 ;
        RECT 140.555 211.900 140.885 212.605 ;
        RECT 141.090 211.880 141.465 212.435 ;
        RECT 142.195 212.425 142.365 212.960 ;
        RECT 143.675 212.800 144.005 213.350 ;
        RECT 144.175 213.310 144.695 213.465 ;
        RECT 144.915 213.140 145.630 214.320 ;
        RECT 145.950 214.075 147.805 214.425 ;
        RECT 144.305 212.970 145.630 213.140 ;
        RECT 143.675 212.790 144.700 212.800 ;
        RECT 142.535 212.600 144.700 212.790 ;
        RECT 142.535 212.450 143.470 212.600 ;
        RECT 144.175 212.470 144.700 212.600 ;
        RECT 144.915 212.485 145.630 212.970 ;
        RECT 147.200 212.485 147.805 214.075 ;
        RECT 141.695 212.220 142.365 212.425 ;
        RECT 141.695 212.110 142.865 212.220 ;
        RECT 142.195 211.905 142.865 212.110 ;
        RECT 130.465 211.090 131.145 211.370 ;
        RECT 131.315 211.070 131.985 211.400 ;
        RECT 132.155 211.165 133.485 211.395 ;
        RECT 125.875 210.470 126.045 210.630 ;
        RECT 116.425 209.280 119.175 210.470 ;
        RECT 113.385 208.800 116.775 209.110 ;
        RECT 112.275 207.695 112.445 208.800 ;
        RECT 112.615 207.910 113.165 208.080 ;
        RECT 112.275 207.365 112.825 207.695 ;
        RECT 112.995 207.535 113.165 207.910 ;
        RECT 113.345 207.815 113.715 208.170 ;
        RECT 113.895 207.910 114.825 208.080 ;
        RECT 113.895 207.535 114.065 207.910 ;
        RECT 114.995 207.695 116.775 208.800 ;
        RECT 112.995 207.365 114.065 207.535 ;
        RECT 114.235 207.420 116.775 207.695 ;
        RECT 116.945 208.820 119.175 209.280 ;
        RECT 119.345 209.900 120.605 210.470 ;
        RECT 120.775 210.070 121.455 210.355 ;
        RECT 119.345 209.630 121.065 209.900 ;
        RECT 116.945 207.420 118.655 208.820 ;
        RECT 119.345 208.650 120.605 209.630 ;
        RECT 121.235 209.610 121.455 210.070 ;
        RECT 121.625 209.780 122.185 210.470 ;
        RECT 122.355 210.070 122.985 210.355 ;
        RECT 122.355 209.610 122.525 210.070 ;
        RECT 123.155 209.900 124.615 210.470 ;
        RECT 122.695 209.630 124.615 209.900 ;
        RECT 121.235 209.400 122.525 209.610 ;
        RECT 120.775 208.830 122.985 209.230 ;
        RECT 114.235 207.365 115.165 207.420 ;
        RECT 112.275 206.765 112.445 207.365 ;
        RECT 113.355 207.280 113.685 207.365 ;
        RECT 114.995 207.250 115.165 207.365 ;
        RECT 117.715 207.250 118.655 207.420 ;
        RECT 112.615 207.110 113.190 207.195 ;
        RECT 113.920 207.110 114.825 207.195 ;
        RECT 112.615 206.940 114.825 207.110 ;
        RECT 114.995 206.765 116.255 207.250 ;
        RECT 112.275 206.505 113.285 206.765 ;
        RECT 113.845 206.560 116.255 206.765 ;
        RECT 116.425 206.960 118.655 207.250 ;
        RECT 118.825 207.840 120.605 208.650 ;
        RECT 120.775 208.360 121.455 208.640 ;
        RECT 121.235 207.965 121.455 208.360 ;
        RECT 121.625 208.135 122.185 208.830 ;
        RECT 123.155 208.820 124.615 209.630 ;
        RECT 124.785 210.035 126.045 210.470 ;
        RECT 126.215 210.275 128.335 210.460 ;
        RECT 124.785 209.770 126.505 210.035 ;
        RECT 127.015 209.825 127.965 210.105 ;
        RECT 128.595 210.100 128.765 210.630 ;
        RECT 128.935 210.500 131.145 210.900 ;
        RECT 131.315 210.470 131.485 211.070 ;
        RECT 132.155 210.900 132.325 211.165 ;
        RECT 131.655 210.730 132.325 210.900 ;
        RECT 132.495 210.645 133.145 210.995 ;
        RECT 133.315 210.900 133.485 211.165 ;
        RECT 133.655 211.070 134.205 211.400 ;
        RECT 133.315 210.730 133.775 210.900 ;
        RECT 134.035 210.470 134.205 211.070 ;
        RECT 134.485 210.865 134.655 211.370 ;
        RECT 134.855 211.205 135.075 211.560 ;
        RECT 135.245 211.375 135.840 211.615 ;
        RECT 134.855 211.035 136.140 211.205 ;
        RECT 134.485 210.695 135.605 210.865 ;
        RECT 135.435 210.505 135.605 210.695 ;
        RECT 135.775 210.675 136.140 211.035 ;
        RECT 136.310 210.505 136.480 211.440 ;
        RECT 129.395 210.120 130.685 210.330 ;
        RECT 128.595 210.020 129.225 210.100 ;
        RECT 128.135 209.830 129.225 210.020 ;
        RECT 128.135 209.770 128.765 209.830 ;
        RECT 122.355 208.360 122.985 208.640 ;
        RECT 122.355 207.965 122.525 208.360 ;
        RECT 118.825 207.515 121.065 207.840 ;
        RECT 121.235 207.515 122.525 207.965 ;
        RECT 123.155 207.840 124.095 208.820 ;
        RECT 124.785 208.650 126.045 209.770 ;
        RECT 126.640 209.600 128.005 209.655 ;
        RECT 126.215 209.485 128.315 209.600 ;
        RECT 126.215 209.350 126.770 209.485 ;
        RECT 127.875 209.430 128.315 209.485 ;
        RECT 122.695 207.515 124.095 207.840 ;
        RECT 118.825 206.960 120.605 207.515 ;
        RECT 121.915 207.410 122.245 207.515 ;
        RECT 120.775 207.240 121.745 207.345 ;
        RECT 122.415 207.240 122.985 207.345 ;
        RECT 120.775 206.960 122.985 207.240 ;
        RECT 123.155 206.960 124.095 207.515 ;
        RECT 124.265 207.865 126.045 208.650 ;
        RECT 126.320 208.205 126.490 209.140 ;
        RECT 126.960 209.075 127.555 209.315 ;
        RECT 128.145 209.265 128.315 209.430 ;
        RECT 127.725 208.905 127.945 209.260 ;
        RECT 128.595 209.090 128.765 209.770 ;
        RECT 129.395 209.660 129.565 210.120 ;
        RECT 128.935 209.375 129.565 209.660 ;
        RECT 129.735 209.260 130.295 209.950 ;
        RECT 130.465 209.660 130.685 210.120 ;
        RECT 131.315 210.100 132.575 210.470 ;
        RECT 130.855 209.830 132.575 210.100 ;
        RECT 130.465 209.375 131.145 209.660 ;
        RECT 131.315 209.090 132.575 209.830 ;
        RECT 132.745 210.375 134.205 210.470 ;
        RECT 132.745 210.005 134.705 210.375 ;
        RECT 134.885 210.285 135.215 210.485 ;
        RECT 135.435 210.335 136.480 210.505 ;
        RECT 136.755 211.160 138.015 211.850 ;
        RECT 138.185 211.360 139.645 211.850 ;
        RECT 139.860 211.730 140.385 211.860 ;
        RECT 141.090 211.730 142.025 211.880 ;
        RECT 139.860 211.540 142.025 211.730 ;
        RECT 139.860 211.530 140.885 211.540 ;
        RECT 138.185 211.330 140.255 211.360 ;
        RECT 138.725 211.190 140.255 211.330 ;
        RECT 136.755 210.640 138.555 211.160 ;
        RECT 138.725 210.640 139.645 211.190 ;
        RECT 139.865 210.865 140.385 211.020 ;
        RECT 140.555 210.980 140.885 211.530 ;
        RECT 142.195 211.370 142.365 211.905 ;
        RECT 143.095 211.895 143.470 212.450 ;
        RECT 143.675 211.725 144.005 212.430 ;
        RECT 144.915 212.210 145.085 212.485 ;
        RECT 144.385 212.000 145.085 212.210 ;
        RECT 141.185 211.200 142.365 211.370 ;
        RECT 139.865 210.810 140.425 210.865 ;
        RECT 141.055 210.855 141.980 211.030 ;
        RECT 141.005 210.810 141.980 210.855 ;
        RECT 139.865 210.700 141.980 210.810 ;
        RECT 139.865 210.690 141.135 210.700 ;
        RECT 140.300 210.640 141.135 210.690 ;
        RECT 136.755 210.380 136.925 210.640 ;
        RECT 139.475 210.380 139.645 210.640 ;
        RECT 132.745 209.260 134.205 210.005 ;
        RECT 134.885 209.825 135.185 210.285 ;
        RECT 135.435 210.165 135.695 210.335 ;
        RECT 136.755 210.165 137.670 210.380 ;
        RECT 135.365 209.995 135.695 210.165 ;
        RECT 135.955 210.110 137.670 210.165 ;
        RECT 135.955 209.995 136.925 210.110 ;
        RECT 134.485 209.655 136.585 209.825 ;
        RECT 134.485 209.420 134.655 209.655 ;
        RECT 136.255 209.575 136.585 209.655 ;
        RECT 135.365 209.295 136.085 209.485 ;
        RECT 136.755 209.480 136.925 209.995 ;
        RECT 137.840 209.940 138.825 210.380 ;
        RECT 138.995 210.080 139.645 210.380 ;
        RECT 139.815 210.190 142.025 210.470 ;
        RECT 139.815 210.085 140.385 210.190 ;
        RECT 141.055 210.085 142.025 210.190 ;
        RECT 142.195 210.195 142.365 211.200 ;
        RECT 142.665 211.555 144.635 211.725 ;
        RECT 142.665 210.840 142.835 211.555 ;
        RECT 143.005 211.065 144.295 211.385 ;
        RECT 143.965 210.920 144.295 211.065 ;
        RECT 144.465 210.940 144.635 211.555 ;
        RECT 144.915 210.915 145.085 212.000 ;
        RECT 145.255 211.130 145.805 211.300 ;
        RECT 143.035 210.705 143.755 210.895 ;
        RECT 142.535 210.535 142.865 210.615 ;
        RECT 144.465 210.535 144.635 210.770 ;
        RECT 142.535 210.365 144.635 210.535 ;
        RECT 144.915 210.585 145.465 210.915 ;
        RECT 145.635 210.755 145.805 211.130 ;
        RECT 145.985 211.035 146.355 211.390 ;
        RECT 146.535 211.130 147.465 211.300 ;
        RECT 146.535 210.755 146.705 211.130 ;
        RECT 147.635 210.915 147.805 212.485 ;
        RECT 145.635 210.585 146.705 210.755 ;
        RECT 146.875 210.585 147.805 210.915 ;
        RECT 137.100 209.910 138.825 209.940 ;
        RECT 139.475 209.915 139.645 210.080 ;
        RECT 142.195 210.025 143.165 210.195 ;
        RECT 143.425 210.025 143.755 210.195 ;
        RECT 140.555 209.915 140.885 210.020 ;
        RECT 142.195 209.915 142.365 210.025 ;
        RECT 137.100 209.650 139.280 209.910 ;
        RECT 126.660 208.735 127.945 208.905 ;
        RECT 126.660 208.375 127.025 208.735 ;
        RECT 128.145 208.565 128.315 209.070 ;
        RECT 127.195 208.395 128.315 208.565 ;
        RECT 127.195 208.205 127.365 208.395 ;
        RECT 126.320 208.035 127.365 208.205 ;
        RECT 127.105 207.865 127.365 208.035 ;
        RECT 127.585 207.985 127.915 208.185 ;
        RECT 128.595 208.075 130.055 209.090 ;
        RECT 124.265 207.695 126.845 207.865 ;
        RECT 127.105 207.695 127.435 207.865 ;
        RECT 124.265 206.960 126.045 207.695 ;
        RECT 127.615 207.525 127.915 207.985 ;
        RECT 128.095 207.880 130.055 208.075 ;
        RECT 130.225 207.880 133.095 209.090 ;
        RECT 133.265 208.190 134.205 209.260 ;
        RECT 134.485 208.635 134.655 209.250 ;
        RECT 134.825 209.125 135.155 209.270 ;
        RECT 134.825 208.805 136.115 209.125 ;
        RECT 136.285 208.635 136.455 209.350 ;
        RECT 134.485 208.465 136.455 208.635 ;
        RECT 136.755 209.225 137.655 209.480 ;
        RECT 136.755 208.610 136.930 209.225 ;
        RECT 137.840 209.215 138.825 209.650 ;
        RECT 139.475 209.590 140.105 209.915 ;
        RECT 139.475 209.480 139.645 209.590 ;
        RECT 138.995 209.220 139.645 209.480 ;
        RECT 137.840 209.040 138.065 209.215 ;
        RECT 137.100 208.780 138.065 209.040 ;
        RECT 133.265 207.980 134.735 208.190 ;
        RECT 133.265 207.880 134.205 207.980 ;
        RECT 128.095 207.705 129.535 207.880 ;
        RECT 130.225 207.710 131.485 207.880 ;
        RECT 126.215 207.355 128.315 207.525 ;
        RECT 126.215 207.275 126.545 207.355 ;
        RECT 116.425 206.730 117.885 206.960 ;
        RECT 113.845 206.505 116.795 206.560 ;
        RECT 112.275 206.330 112.445 206.505 ;
        RECT 114.995 206.330 116.795 206.505 ;
        RECT 112.275 206.040 113.170 206.330 ;
        RECT 113.830 206.040 116.795 206.330 ;
        RECT 116.965 206.330 117.885 206.730 ;
        RECT 120.435 206.330 120.605 206.960 ;
        RECT 116.965 206.040 118.610 206.330 ;
        RECT 119.270 206.040 120.605 206.330 ;
        RECT 120.955 206.515 122.345 206.790 ;
        RECT 120.955 206.450 122.950 206.515 ;
        RECT 120.955 206.275 121.365 206.450 ;
        RECT 112.275 205.405 112.445 206.040 ;
        RECT 114.995 205.405 115.165 206.040 ;
        RECT 117.715 205.870 117.885 206.040 ;
        RECT 120.435 205.870 121.365 206.040 ;
        RECT 116.225 205.820 117.060 205.870 ;
        RECT 116.225 205.810 117.495 205.820 ;
        RECT 115.380 205.700 117.495 205.810 ;
        RECT 115.380 205.655 116.355 205.700 ;
        RECT 115.380 205.480 116.305 205.655 ;
        RECT 116.935 205.645 117.495 205.700 ;
        RECT 112.275 205.145 113.285 205.405 ;
        RECT 113.845 205.310 115.165 205.405 ;
        RECT 113.845 205.145 116.175 205.310 ;
        RECT 112.275 204.545 112.445 205.145 ;
        RECT 114.995 205.140 116.175 205.145 ;
        RECT 112.615 204.800 114.825 204.970 ;
        RECT 112.615 204.715 113.190 204.800 ;
        RECT 113.920 204.715 114.825 204.800 ;
        RECT 113.355 204.545 113.685 204.630 ;
        RECT 114.995 204.545 115.165 205.140 ;
        RECT 116.475 204.980 116.805 205.530 ;
        RECT 116.975 205.490 117.495 205.645 ;
        RECT 117.715 205.565 118.395 205.870 ;
        RECT 117.715 205.320 117.885 205.565 ;
        RECT 118.565 205.555 119.125 205.870 ;
        RECT 120.435 205.860 120.605 205.870 ;
        RECT 119.625 205.565 120.605 205.860 ;
        RECT 121.610 205.700 121.800 206.280 ;
        RECT 117.105 205.150 117.885 205.320 ;
        RECT 116.475 204.970 117.500 204.980 ;
        RECT 115.335 204.780 117.500 204.970 ;
        RECT 115.335 204.630 116.270 204.780 ;
        RECT 116.975 204.650 117.500 204.780 ;
        RECT 117.715 204.965 117.885 205.150 ;
        RECT 118.065 205.140 120.265 205.385 ;
        RECT 118.065 205.135 119.125 205.140 ;
        RECT 117.715 204.705 118.410 204.965 ;
        RECT 112.275 204.215 112.825 204.545 ;
        RECT 112.995 204.375 114.065 204.545 ;
        RECT 112.275 203.140 112.445 204.215 ;
        RECT 112.995 204.000 113.165 204.375 ;
        RECT 112.615 203.830 113.165 204.000 ;
        RECT 113.345 203.740 113.715 204.095 ;
        RECT 113.895 204.000 114.065 204.375 ;
        RECT 114.235 204.400 115.165 204.545 ;
        RECT 114.235 204.215 115.665 204.400 ;
        RECT 114.995 204.085 115.665 204.215 ;
        RECT 113.895 203.830 114.825 204.000 ;
        RECT 112.705 203.310 113.165 203.480 ;
        RECT 112.275 202.810 112.825 203.140 ;
        RECT 112.995 203.045 113.165 203.310 ;
        RECT 113.335 203.215 113.985 203.565 ;
        RECT 114.155 203.310 114.825 203.480 ;
        RECT 114.155 203.045 114.325 203.310 ;
        RECT 114.995 203.140 115.165 204.085 ;
        RECT 115.895 204.075 116.270 204.630 ;
        RECT 116.475 203.905 116.805 204.610 ;
        RECT 117.715 204.390 117.885 204.705 ;
        RECT 118.875 204.525 119.125 205.135 ;
        RECT 120.435 204.965 120.605 205.565 ;
        RECT 119.625 204.705 120.605 204.965 ;
        RECT 117.185 204.180 117.885 204.390 ;
        RECT 118.065 204.275 120.260 204.525 ;
        RECT 117.715 204.105 117.885 204.180 ;
        RECT 112.995 202.815 114.325 203.045 ;
        RECT 114.495 202.810 115.165 203.140 ;
        RECT 115.465 203.735 117.435 203.905 ;
        RECT 115.465 203.020 115.635 203.735 ;
        RECT 115.805 203.245 117.095 203.565 ;
        RECT 116.765 203.100 117.095 203.245 ;
        RECT 117.265 203.120 117.435 203.735 ;
        RECT 117.715 203.845 118.445 204.105 ;
        RECT 117.715 203.245 117.885 203.845 ;
        RECT 118.080 203.415 118.705 203.675 ;
        RECT 115.835 202.885 116.555 203.075 ;
        RECT 117.715 202.985 118.365 203.245 ;
        RECT 112.275 202.200 112.445 202.810 ;
        RECT 112.705 202.455 114.825 202.640 ;
        RECT 114.995 202.375 115.165 202.810 ;
        RECT 115.335 202.715 115.665 202.795 ;
        RECT 117.265 202.715 117.435 202.950 ;
        RECT 115.335 202.545 117.435 202.715 ;
        RECT 112.275 201.950 112.905 202.200 ;
        RECT 113.075 202.005 114.025 202.285 ;
        RECT 114.995 202.215 115.965 202.375 ;
        RECT 114.535 202.205 115.965 202.215 ;
        RECT 116.225 202.205 116.555 202.375 ;
        RECT 114.535 201.950 115.165 202.205 ;
        RECT 116.225 202.035 116.485 202.205 ;
        RECT 116.735 202.085 117.035 202.545 ;
        RECT 117.715 202.385 117.885 202.985 ;
        RECT 118.535 202.815 118.705 203.415 ;
        RECT 118.080 202.555 118.705 202.815 ;
        RECT 117.715 202.365 118.365 202.385 ;
        RECT 112.275 200.255 112.445 201.950 ;
        RECT 113.035 201.780 114.400 201.835 ;
        RECT 112.725 201.665 114.825 201.780 ;
        RECT 112.725 201.610 113.165 201.665 ;
        RECT 112.725 201.445 112.895 201.610 ;
        RECT 114.270 201.530 114.825 201.665 ;
        RECT 112.725 200.745 112.895 201.250 ;
        RECT 113.095 201.085 113.315 201.440 ;
        RECT 113.485 201.255 114.080 201.495 ;
        RECT 113.095 200.915 114.380 201.085 ;
        RECT 112.725 200.575 113.845 200.745 ;
        RECT 113.675 200.385 113.845 200.575 ;
        RECT 114.015 200.555 114.380 200.915 ;
        RECT 114.550 200.385 114.720 201.320 ;
        RECT 112.275 199.885 112.945 200.255 ;
        RECT 113.125 200.165 113.455 200.365 ;
        RECT 113.675 200.215 114.720 200.385 ;
        RECT 114.995 200.300 115.165 201.950 ;
        RECT 115.440 201.865 116.485 202.035 ;
        RECT 116.705 201.885 117.035 202.085 ;
        RECT 117.215 202.125 118.365 202.365 ;
        RECT 117.215 201.995 117.885 202.125 ;
        RECT 115.440 200.930 115.610 201.865 ;
        RECT 115.780 201.335 116.145 201.695 ;
        RECT 116.315 201.675 116.485 201.865 ;
        RECT 116.315 201.505 117.435 201.675 ;
        RECT 115.780 201.165 117.065 201.335 ;
        RECT 116.080 200.755 116.675 200.995 ;
        RECT 116.845 200.810 117.065 201.165 ;
        RECT 117.265 201.000 117.435 201.505 ;
        RECT 117.715 201.525 117.885 201.995 ;
        RECT 118.535 201.955 118.705 202.555 ;
        RECT 118.080 201.695 118.705 201.955 ;
        RECT 117.715 201.280 118.365 201.525 ;
        RECT 115.335 200.585 115.890 200.720 ;
        RECT 117.265 200.640 117.435 200.805 ;
        RECT 116.995 200.585 117.435 200.640 ;
        RECT 115.335 200.470 117.435 200.585 ;
        RECT 117.715 200.665 117.885 201.280 ;
        RECT 118.535 201.110 118.705 201.695 ;
        RECT 118.080 200.835 118.705 201.110 ;
        RECT 115.760 200.415 117.125 200.470 ;
        RECT 117.715 200.420 118.365 200.665 ;
        RECT 117.715 200.300 117.885 200.420 ;
        RECT 112.275 198.070 112.445 199.885 ;
        RECT 113.125 199.705 113.425 200.165 ;
        RECT 113.675 200.045 113.935 200.215 ;
        RECT 114.995 200.045 115.625 200.300 ;
        RECT 113.605 199.875 113.935 200.045 ;
        RECT 114.195 200.035 115.625 200.045 ;
        RECT 114.195 199.875 115.165 200.035 ;
        RECT 116.135 199.965 117.085 200.245 ;
        RECT 117.255 200.050 117.885 200.300 ;
        RECT 118.535 200.250 118.705 200.835 ;
        RECT 112.725 199.535 114.825 199.705 ;
        RECT 112.725 199.300 112.895 199.535 ;
        RECT 114.495 199.455 114.825 199.535 ;
        RECT 114.995 199.440 115.165 199.875 ;
        RECT 117.715 199.810 117.885 200.050 ;
        RECT 118.080 199.990 118.705 200.250 ;
        RECT 115.335 199.610 117.455 199.795 ;
        RECT 117.715 199.560 118.365 199.810 ;
        RECT 117.715 199.440 117.885 199.560 ;
        RECT 113.605 199.175 114.325 199.365 ;
        RECT 112.725 198.515 112.895 199.130 ;
        RECT 113.065 199.005 113.395 199.150 ;
        RECT 113.065 198.685 114.355 199.005 ;
        RECT 114.525 198.515 114.695 199.230 ;
        RECT 112.725 198.345 114.695 198.515 ;
        RECT 114.995 199.110 115.665 199.440 ;
        RECT 115.835 199.205 117.165 199.435 ;
        RECT 112.275 197.860 112.975 198.070 ;
        RECT 112.275 197.100 112.445 197.860 ;
        RECT 113.355 197.640 113.685 198.345 ;
        RECT 113.890 197.620 114.265 198.175 ;
        RECT 114.995 198.165 115.165 199.110 ;
        RECT 115.835 198.940 116.005 199.205 ;
        RECT 115.335 198.770 116.005 198.940 ;
        RECT 116.175 198.685 116.825 199.035 ;
        RECT 116.995 198.940 117.165 199.205 ;
        RECT 117.335 199.110 117.885 199.440 ;
        RECT 118.535 199.390 118.705 199.990 ;
        RECT 118.080 199.130 118.705 199.390 ;
        RECT 117.715 198.950 117.885 199.110 ;
        RECT 116.995 198.770 117.455 198.940 ;
        RECT 117.715 198.700 118.365 198.950 ;
        RECT 115.335 198.335 117.545 198.505 ;
        RECT 115.335 198.170 116.305 198.335 ;
        RECT 116.975 198.250 117.545 198.335 ;
        RECT 114.495 198.000 115.165 198.165 ;
        RECT 116.475 198.080 116.805 198.165 ;
        RECT 117.715 198.090 117.885 198.700 ;
        RECT 118.535 198.530 118.705 199.130 ;
        RECT 118.080 198.270 118.705 198.530 ;
        RECT 118.535 198.095 118.705 198.270 ;
        RECT 118.875 198.265 119.125 204.275 ;
        RECT 120.435 204.105 120.605 204.705 ;
        RECT 119.635 203.845 120.605 204.105 ;
        RECT 119.295 203.415 120.260 203.675 ;
        RECT 120.430 203.500 120.605 203.845 ;
        RECT 120.775 205.530 121.800 205.700 ;
        RECT 122.175 206.270 122.950 206.450 ;
        RECT 123.155 206.330 123.325 206.960 ;
        RECT 125.875 206.330 126.045 206.960 ;
        RECT 122.175 205.560 122.345 206.270 ;
        RECT 123.155 206.050 124.050 206.330 ;
        RECT 122.620 206.040 124.050 206.050 ;
        RECT 124.710 206.040 126.045 206.330 ;
        RECT 126.345 206.335 126.515 207.050 ;
        RECT 126.715 206.995 127.435 207.185 ;
        RECT 128.145 207.120 128.315 207.355 ;
        RECT 127.645 206.825 127.975 206.970 ;
        RECT 126.685 206.505 127.975 206.825 ;
        RECT 128.145 206.335 128.315 206.950 ;
        RECT 126.345 206.165 128.315 206.335 ;
        RECT 128.595 206.500 129.535 207.705 ;
        RECT 129.705 207.240 131.485 207.710 ;
        RECT 134.035 207.250 134.205 207.880 ;
        RECT 135.115 207.760 135.445 208.465 ;
        RECT 136.755 208.365 137.655 208.610 ;
        RECT 135.650 207.740 136.025 208.295 ;
        RECT 136.755 208.285 136.930 208.365 ;
        RECT 136.255 207.970 136.930 208.285 ;
        RECT 137.825 208.180 138.065 208.780 ;
        RECT 136.755 207.750 136.930 207.970 ;
        RECT 137.100 207.920 138.065 208.180 ;
        RECT 134.420 207.590 134.945 207.720 ;
        RECT 135.650 207.590 136.585 207.740 ;
        RECT 134.420 207.400 136.585 207.590 ;
        RECT 136.755 207.505 137.655 207.750 ;
        RECT 134.420 207.390 135.445 207.400 ;
        RECT 129.705 206.945 132.295 207.240 ;
        RECT 129.705 206.500 131.485 206.945 ;
        RECT 132.795 206.935 133.355 207.250 ;
        RECT 133.525 207.220 134.205 207.250 ;
        RECT 133.525 207.050 134.815 207.220 ;
        RECT 133.525 206.945 134.205 207.050 ;
        RECT 131.655 206.520 133.855 206.765 ;
        RECT 128.595 206.330 128.765 206.500 ;
        RECT 131.315 206.345 131.485 206.500 ;
        RECT 132.795 206.515 133.855 206.520 ;
        RECT 131.315 206.330 132.295 206.345 ;
        RECT 122.620 205.540 123.325 206.040 ;
        RECT 125.875 205.985 126.045 206.040 ;
        RECT 123.585 205.610 124.045 205.780 ;
        RECT 120.775 203.840 120.945 205.530 ;
        RECT 123.155 205.440 123.325 205.540 ;
        RECT 121.455 205.170 122.985 205.360 ;
        RECT 121.115 204.180 121.285 205.135 ;
        RECT 121.455 204.520 121.625 205.170 ;
        RECT 123.155 205.110 123.705 205.440 ;
        RECT 123.875 205.345 124.045 205.610 ;
        RECT 124.215 205.515 124.865 205.865 ;
        RECT 125.035 205.610 125.705 205.780 ;
        RECT 125.875 205.670 126.545 205.985 ;
        RECT 125.035 205.345 125.205 205.610 ;
        RECT 125.875 205.440 126.045 205.670 ;
        RECT 126.775 205.440 127.150 205.995 ;
        RECT 127.355 205.460 127.685 206.165 ;
        RECT 128.595 206.040 129.490 206.330 ;
        RECT 130.150 206.085 132.295 206.330 ;
        RECT 130.150 206.040 131.485 206.085 ;
        RECT 128.595 205.890 128.765 206.040 ;
        RECT 128.065 205.860 128.765 205.890 ;
        RECT 128.065 205.680 129.575 205.860 ;
        RECT 128.595 205.590 129.575 205.680 ;
        RECT 123.875 205.115 125.205 205.345 ;
        RECT 125.375 205.110 126.045 205.440 ;
        RECT 121.825 204.725 122.985 205.000 ;
        RECT 121.965 204.720 122.135 204.725 ;
        RECT 121.455 204.350 122.425 204.520 ;
        RECT 122.620 204.180 122.985 204.535 ;
        RECT 121.115 204.010 122.985 204.180 ;
        RECT 122.415 204.005 122.985 204.010 ;
        RECT 123.155 204.500 123.325 205.110 ;
        RECT 123.585 204.755 125.705 204.940 ;
        RECT 125.875 204.930 126.045 205.110 ;
        RECT 126.215 205.290 127.150 205.440 ;
        RECT 127.855 205.290 128.380 205.420 ;
        RECT 126.215 205.100 128.380 205.290 ;
        RECT 127.355 205.090 128.380 205.100 ;
        RECT 125.875 204.760 127.055 204.930 ;
        RECT 123.155 204.250 123.785 204.500 ;
        RECT 123.955 204.305 124.905 204.585 ;
        RECT 125.875 204.515 126.045 204.760 ;
        RECT 125.415 204.250 126.045 204.515 ;
        RECT 126.260 204.415 127.185 204.590 ;
        RECT 127.355 204.540 127.685 205.090 ;
        RECT 128.595 204.920 128.765 205.590 ;
        RECT 129.755 205.520 130.005 205.870 ;
        RECT 131.315 205.860 131.485 206.040 ;
        RECT 132.795 205.905 133.045 206.515 ;
        RECT 134.035 206.345 134.205 206.945 ;
        RECT 134.425 206.725 134.945 206.880 ;
        RECT 135.115 206.840 135.445 207.390 ;
        RECT 136.755 207.230 136.930 207.505 ;
        RECT 137.825 207.320 138.065 207.920 ;
        RECT 135.745 207.060 136.930 207.230 ;
        RECT 137.100 207.060 138.065 207.320 ;
        RECT 136.755 206.890 136.930 207.060 ;
        RECT 134.425 206.670 134.985 206.725 ;
        RECT 135.615 206.715 136.540 206.890 ;
        RECT 135.565 206.670 136.540 206.715 ;
        RECT 134.425 206.560 136.540 206.670 ;
        RECT 136.755 206.645 137.655 206.890 ;
        RECT 134.425 206.550 135.695 206.560 ;
        RECT 134.860 206.500 135.695 206.550 ;
        RECT 133.510 206.330 134.205 206.345 ;
        RECT 136.755 206.330 136.930 206.645 ;
        RECT 137.825 206.475 138.065 207.060 ;
        RECT 133.510 206.085 134.930 206.330 ;
        RECT 134.035 206.040 134.930 206.085 ;
        RECT 135.590 206.045 136.930 206.330 ;
        RECT 137.100 206.215 138.065 206.475 ;
        RECT 135.590 206.040 137.655 206.045 ;
        RECT 130.175 205.530 131.485 205.860 ;
        RECT 131.660 205.655 133.855 205.905 ;
        RECT 131.315 205.485 131.485 205.530 ;
        RECT 128.935 205.350 129.575 205.420 ;
        RECT 128.935 205.180 130.345 205.350 ;
        RECT 128.935 205.090 129.575 205.180 ;
        RECT 127.985 204.750 129.575 204.920 ;
        RECT 128.595 204.680 129.575 204.750 ;
        RECT 127.855 204.425 128.375 204.580 ;
        RECT 126.260 204.370 127.235 204.415 ;
        RECT 127.815 204.370 128.375 204.425 ;
        RECT 126.260 204.260 128.375 204.370 ;
        RECT 120.775 203.670 122.245 203.840 ;
        RECT 121.915 203.645 122.245 203.670 ;
        RECT 119.295 202.815 119.535 203.415 ;
        RECT 120.430 203.330 121.745 203.500 ;
        RECT 122.415 203.420 122.585 204.005 ;
        RECT 123.155 203.580 123.325 204.250 ;
        RECT 123.915 204.080 125.280 204.135 ;
        RECT 123.605 203.965 125.705 204.080 ;
        RECT 123.605 203.910 124.045 203.965 ;
        RECT 123.605 203.745 123.775 203.910 ;
        RECT 125.150 203.830 125.705 203.965 ;
        RECT 120.430 203.245 120.605 203.330 ;
        RECT 119.705 202.985 120.605 203.245 ;
        RECT 121.915 203.250 122.585 203.420 ;
        RECT 122.755 203.250 123.325 203.580 ;
        RECT 121.915 203.165 122.245 203.250 ;
        RECT 119.295 202.555 120.260 202.815 ;
        RECT 120.430 202.650 120.605 202.985 ;
        RECT 120.775 202.995 121.745 203.160 ;
        RECT 122.415 202.995 122.985 203.080 ;
        RECT 120.775 202.825 122.985 202.995 ;
        RECT 123.155 202.650 123.325 203.250 ;
        RECT 123.605 203.045 123.775 203.550 ;
        RECT 123.975 203.385 124.195 203.740 ;
        RECT 124.365 203.555 124.960 203.795 ;
        RECT 123.975 203.215 125.260 203.385 ;
        RECT 123.605 202.875 124.725 203.045 ;
        RECT 124.555 202.685 124.725 202.875 ;
        RECT 124.895 202.855 125.260 203.215 ;
        RECT 125.430 202.685 125.600 203.620 ;
        RECT 119.295 201.955 119.535 202.555 ;
        RECT 120.430 202.385 121.695 202.650 ;
        RECT 119.705 202.125 121.695 202.385 ;
        RECT 119.295 201.695 120.260 201.955 ;
        RECT 120.430 201.730 121.695 202.125 ;
        RECT 121.865 202.555 123.325 202.650 ;
        RECT 121.865 202.185 123.825 202.555 ;
        RECT 124.005 202.465 124.335 202.665 ;
        RECT 124.555 202.515 125.600 202.685 ;
        RECT 125.875 203.520 126.045 204.250 ;
        RECT 127.105 204.250 128.375 204.260 ;
        RECT 127.105 204.200 127.940 204.250 ;
        RECT 126.215 203.855 128.425 204.025 ;
        RECT 126.215 203.690 127.185 203.855 ;
        RECT 127.855 203.770 128.425 203.855 ;
        RECT 128.595 203.890 128.765 204.680 ;
        RECT 129.755 204.660 130.005 205.010 ;
        RECT 130.175 205.000 130.345 205.180 ;
        RECT 131.315 205.225 132.285 205.485 ;
        RECT 130.175 204.670 131.130 205.000 ;
        RECT 131.315 204.625 131.490 205.225 ;
        RECT 131.660 204.795 132.625 205.055 ;
        RECT 128.935 204.060 129.585 204.390 ;
        RECT 127.355 203.600 127.685 203.685 ;
        RECT 128.595 203.600 129.225 203.890 ;
        RECT 125.875 203.350 127.185 203.520 ;
        RECT 127.355 203.430 128.025 203.600 ;
        RECT 121.865 201.900 123.325 202.185 ;
        RECT 124.005 202.005 124.305 202.465 ;
        RECT 124.555 202.345 124.815 202.515 ;
        RECT 125.875 202.345 126.045 203.350 ;
        RECT 127.355 203.180 127.685 203.205 ;
        RECT 124.485 202.175 124.815 202.345 ;
        RECT 125.075 202.175 126.045 202.345 ;
        RECT 119.295 201.095 119.535 201.695 ;
        RECT 120.430 201.525 122.215 201.730 ;
        RECT 119.705 201.265 122.215 201.525 ;
        RECT 119.295 200.835 120.260 201.095 ;
        RECT 120.430 200.980 122.215 201.265 ;
        RECT 122.385 200.980 123.325 201.900 ;
        RECT 123.605 201.835 125.705 202.005 ;
        RECT 123.605 201.600 123.775 201.835 ;
        RECT 125.375 201.755 125.705 201.835 ;
        RECT 124.485 201.475 125.205 201.665 ;
        RECT 119.295 200.250 119.535 200.835 ;
        RECT 120.430 200.665 120.605 200.980 ;
        RECT 119.705 200.420 120.605 200.665 ;
        RECT 120.775 200.550 121.445 200.720 ;
        RECT 120.430 200.380 120.605 200.420 ;
        RECT 119.295 199.990 120.260 200.250 ;
        RECT 120.430 200.050 121.105 200.380 ;
        RECT 121.275 200.285 121.445 200.550 ;
        RECT 121.615 200.455 122.265 200.805 ;
        RECT 122.435 200.550 122.895 200.720 ;
        RECT 122.435 200.285 122.605 200.550 ;
        RECT 123.155 200.380 123.325 200.980 ;
        RECT 123.605 200.815 123.775 201.430 ;
        RECT 123.945 201.305 124.275 201.450 ;
        RECT 123.945 200.985 125.235 201.305 ;
        RECT 125.405 200.815 125.575 201.530 ;
        RECT 123.605 200.645 125.575 200.815 ;
        RECT 125.875 200.980 126.045 202.175 ;
        RECT 126.215 203.010 127.685 203.180 ;
        RECT 126.215 201.320 126.385 203.010 ;
        RECT 127.855 202.845 128.025 203.430 ;
        RECT 128.195 203.560 129.225 203.600 ;
        RECT 128.195 203.270 128.765 203.560 ;
        RECT 129.415 203.345 129.585 204.060 ;
        RECT 129.755 203.920 130.005 204.430 ;
        RECT 131.315 204.370 132.215 204.625 ;
        RECT 130.195 204.365 132.215 204.370 ;
        RECT 130.195 204.040 131.490 204.365 ;
        RECT 132.385 204.195 132.625 204.795 ;
        RECT 131.315 203.765 131.490 204.040 ;
        RECT 131.660 203.935 132.625 204.195 ;
        RECT 127.855 202.840 128.425 202.845 ;
        RECT 126.555 202.670 128.425 202.840 ;
        RECT 126.555 201.715 126.725 202.670 ;
        RECT 126.895 202.330 127.865 202.500 ;
        RECT 126.895 201.680 127.065 202.330 ;
        RECT 128.060 202.315 128.425 202.670 ;
        RECT 128.595 202.815 128.765 203.270 ;
        RECT 128.935 203.015 129.585 203.345 ;
        RECT 129.755 203.340 131.070 203.710 ;
        RECT 131.315 203.505 132.215 203.765 ;
        RECT 128.595 202.485 129.225 202.815 ;
        RECT 127.405 202.125 127.575 202.130 ;
        RECT 127.265 201.850 128.425 202.125 ;
        RECT 126.895 201.490 128.425 201.680 ;
        RECT 128.595 201.320 128.765 202.485 ;
        RECT 129.415 202.260 129.585 203.015 ;
        RECT 129.755 202.840 131.070 203.170 ;
        RECT 131.315 202.905 131.490 203.505 ;
        RECT 132.385 203.335 132.625 203.935 ;
        RECT 131.660 203.075 132.625 203.335 ;
        RECT 131.315 202.645 132.215 202.905 ;
        RECT 129.755 202.300 131.070 202.630 ;
        RECT 129.095 202.090 129.585 202.260 ;
        RECT 128.950 201.590 129.585 201.920 ;
        RECT 129.755 201.710 129.965 202.130 ;
        RECT 131.315 202.045 131.490 202.645 ;
        RECT 132.385 202.475 132.625 203.075 ;
        RECT 131.660 202.215 132.625 202.475 ;
        RECT 130.135 201.780 131.145 202.030 ;
        RECT 131.315 201.800 132.215 202.045 ;
        RECT 129.395 201.540 129.585 201.590 ;
        RECT 130.135 201.540 130.425 201.780 ;
        RECT 131.315 201.610 131.490 201.800 ;
        RECT 132.385 201.630 132.625 202.215 ;
        RECT 126.215 201.150 127.240 201.320 ;
        RECT 128.595 201.310 129.225 201.320 ;
        RECT 125.875 200.810 126.805 200.980 ;
        RECT 121.275 200.055 122.605 200.285 ;
        RECT 122.775 200.370 123.325 200.380 ;
        RECT 122.775 200.160 123.855 200.370 ;
        RECT 122.775 200.050 123.325 200.160 ;
        RECT 119.295 199.390 119.535 199.990 ;
        RECT 120.430 199.805 120.605 200.050 ;
        RECT 119.705 199.560 120.605 199.805 ;
        RECT 120.775 199.695 122.895 199.880 ;
        RECT 120.430 199.455 120.605 199.560 ;
        RECT 119.295 199.130 120.260 199.390 ;
        RECT 120.430 199.190 121.065 199.455 ;
        RECT 121.575 199.245 122.525 199.525 ;
        RECT 123.155 199.440 123.325 200.050 ;
        RECT 124.235 199.940 124.565 200.645 ;
        RECT 124.770 199.920 125.145 200.475 ;
        RECT 125.875 200.465 126.045 200.810 ;
        RECT 125.375 200.150 126.045 200.465 ;
        RECT 123.540 199.770 124.065 199.900 ;
        RECT 124.770 199.770 125.705 199.920 ;
        RECT 123.540 199.580 125.705 199.770 ;
        RECT 123.540 199.570 124.565 199.580 ;
        RECT 122.695 199.400 123.325 199.440 ;
        RECT 122.695 199.230 123.935 199.400 ;
        RECT 122.695 199.190 123.325 199.230 ;
        RECT 119.295 198.530 119.535 199.130 ;
        RECT 120.430 198.945 120.605 199.190 ;
        RECT 121.200 199.020 122.565 199.075 ;
        RECT 119.705 198.700 120.605 198.945 ;
        RECT 120.775 198.905 122.875 199.020 ;
        RECT 120.775 198.770 121.330 198.905 ;
        RECT 122.435 198.850 122.875 198.905 ;
        RECT 119.295 198.270 120.260 198.530 ;
        RECT 119.295 198.095 119.520 198.270 ;
        RECT 117.715 198.080 118.365 198.090 ;
        RECT 114.495 197.850 116.305 198.000 ;
        RECT 116.475 197.910 117.145 198.080 ;
        RECT 114.995 197.830 116.305 197.850 ;
        RECT 112.660 197.470 113.185 197.600 ;
        RECT 113.890 197.470 114.825 197.620 ;
        RECT 112.660 197.280 114.825 197.470 ;
        RECT 112.660 197.270 113.685 197.280 ;
        RECT 112.275 196.930 113.055 197.100 ;
        RECT 112.275 196.205 112.445 196.930 ;
        RECT 112.665 196.605 113.185 196.760 ;
        RECT 113.355 196.720 113.685 197.270 ;
        RECT 114.995 197.110 115.165 197.830 ;
        RECT 116.475 197.660 116.805 197.685 ;
        RECT 113.985 196.940 115.165 197.110 ;
        RECT 112.665 196.550 113.225 196.605 ;
        RECT 113.855 196.595 114.780 196.770 ;
        RECT 113.805 196.550 114.780 196.595 ;
        RECT 112.665 196.440 114.780 196.550 ;
        RECT 112.665 196.430 113.935 196.440 ;
        RECT 113.100 196.380 113.935 196.430 ;
        RECT 114.995 196.205 115.165 196.940 ;
        RECT 112.275 195.945 113.285 196.205 ;
        RECT 113.845 195.945 115.165 196.205 ;
        RECT 112.275 195.345 112.445 195.945 ;
        RECT 112.615 195.600 114.825 195.770 ;
        RECT 112.615 195.515 113.190 195.600 ;
        RECT 113.920 195.515 114.825 195.600 ;
        RECT 114.995 195.460 115.165 195.945 ;
        RECT 115.335 197.490 116.805 197.660 ;
        RECT 115.335 195.800 115.505 197.490 ;
        RECT 116.975 197.325 117.145 197.910 ;
        RECT 117.315 197.830 118.365 198.080 ;
        RECT 117.315 197.750 117.885 197.830 ;
        RECT 116.975 197.320 117.545 197.325 ;
        RECT 115.675 197.150 117.545 197.320 ;
        RECT 115.675 196.195 115.845 197.150 ;
        RECT 116.015 196.810 116.985 196.980 ;
        RECT 116.015 196.160 116.185 196.810 ;
        RECT 117.180 196.795 117.545 197.150 ;
        RECT 117.715 197.230 117.885 197.750 ;
        RECT 118.535 197.660 119.520 198.095 ;
        RECT 120.430 198.085 120.605 198.700 ;
        RECT 119.705 197.830 120.605 198.085 ;
        RECT 118.080 197.400 120.260 197.660 ;
        RECT 118.535 197.370 120.260 197.400 ;
        RECT 117.715 196.930 118.365 197.230 ;
        RECT 118.535 196.930 119.520 197.370 ;
        RECT 120.435 197.285 120.605 197.830 ;
        RECT 120.880 197.625 121.050 198.560 ;
        RECT 121.520 198.495 122.115 198.735 ;
        RECT 122.705 198.685 122.875 198.850 ;
        RECT 122.285 198.325 122.505 198.680 ;
        RECT 123.155 198.500 123.325 199.190 ;
        RECT 123.545 198.905 124.065 199.060 ;
        RECT 124.235 199.020 124.565 199.570 ;
        RECT 125.875 199.410 126.045 200.150 ;
        RECT 126.395 200.400 126.805 200.575 ;
        RECT 127.050 200.570 127.240 201.150 ;
        RECT 127.615 200.580 127.785 201.290 ;
        RECT 128.060 201.150 129.225 201.310 ;
        RECT 129.395 201.280 130.425 201.540 ;
        RECT 130.595 201.280 131.490 201.610 ;
        RECT 131.660 201.370 132.625 201.630 ;
        RECT 129.395 201.170 129.965 201.280 ;
        RECT 128.060 200.800 128.765 201.150 ;
        RECT 129.755 200.960 129.965 201.170 ;
        RECT 131.315 201.185 131.490 201.280 ;
        RECT 127.615 200.400 128.390 200.580 ;
        RECT 126.395 200.335 128.390 200.400 ;
        RECT 126.395 200.060 127.785 200.335 ;
        RECT 126.215 199.610 128.425 199.890 ;
        RECT 126.215 199.505 127.185 199.610 ;
        RECT 127.855 199.505 128.425 199.610 ;
        RECT 128.595 199.795 128.765 200.800 ;
        RECT 128.935 200.790 129.565 200.860 ;
        RECT 130.135 200.790 131.145 201.045 ;
        RECT 128.935 200.520 131.145 200.790 ;
        RECT 131.315 200.940 132.215 201.185 ;
        RECT 128.935 200.070 131.145 200.350 ;
        RECT 128.935 199.965 129.505 200.070 ;
        RECT 130.175 199.965 131.145 200.070 ;
        RECT 131.315 200.325 131.490 200.940 ;
        RECT 132.385 200.770 132.625 201.370 ;
        RECT 131.660 200.510 132.625 200.770 ;
        RECT 131.315 200.080 132.215 200.325 ;
        RECT 129.675 199.795 130.005 199.900 ;
        RECT 131.315 199.795 131.490 200.080 ;
        RECT 132.385 199.910 132.625 200.510 ;
        RECT 128.595 199.470 129.225 199.795 ;
        RECT 124.865 199.335 126.045 199.410 ;
        RECT 127.355 199.335 127.685 199.440 ;
        RECT 128.595 199.335 128.765 199.470 ;
        RECT 124.865 199.240 126.505 199.335 ;
        RECT 123.545 198.850 124.105 198.905 ;
        RECT 124.735 198.895 125.660 199.070 ;
        RECT 124.685 198.850 125.660 198.895 ;
        RECT 123.545 198.740 125.660 198.850 ;
        RECT 125.875 199.010 126.505 199.240 ;
        RECT 123.545 198.730 124.815 198.740 ;
        RECT 123.980 198.680 124.815 198.730 ;
        RECT 121.220 198.155 122.505 198.325 ;
        RECT 121.220 197.795 121.585 198.155 ;
        RECT 122.705 197.985 122.875 198.490 ;
        RECT 121.755 197.815 122.875 197.985 ;
        RECT 123.155 198.170 123.830 198.500 ;
        RECT 124.685 198.445 124.855 198.450 ;
        RECT 121.755 197.625 121.925 197.815 ;
        RECT 120.880 197.455 121.925 197.625 ;
        RECT 121.665 197.285 121.925 197.455 ;
        RECT 122.145 197.405 122.475 197.605 ;
        RECT 123.155 197.495 123.325 198.170 ;
        RECT 124.005 198.145 124.855 198.445 ;
        RECT 125.025 198.250 125.685 198.420 ;
        RECT 123.520 197.975 123.895 198.000 ;
        RECT 125.025 197.975 125.255 198.250 ;
        RECT 125.875 198.080 126.045 199.010 ;
        RECT 126.675 198.885 127.965 199.335 ;
        RECT 128.135 199.010 128.765 199.335 ;
        RECT 126.675 198.490 126.895 198.885 ;
        RECT 126.215 198.210 126.895 198.490 ;
        RECT 123.520 197.760 125.255 197.975 ;
        RECT 120.435 197.200 121.405 197.285 ;
        RECT 119.690 197.115 121.405 197.200 ;
        RECT 121.665 197.115 121.995 197.285 ;
        RECT 119.690 196.930 120.605 197.115 ;
        RECT 122.175 196.945 122.475 197.405 ;
        RECT 122.655 197.125 123.325 197.495 ;
        RECT 124.045 197.740 125.255 197.760 ;
        RECT 125.425 197.750 126.045 198.080 ;
        RECT 127.065 198.020 127.625 198.715 ;
        RECT 127.795 198.490 127.965 198.885 ;
        RECT 127.795 198.210 128.425 198.490 ;
        RECT 123.510 197.310 123.850 197.480 ;
        RECT 124.045 197.420 124.375 197.740 ;
        RECT 117.715 196.670 117.885 196.930 ;
        RECT 120.435 196.670 120.605 196.930 ;
        RECT 120.775 196.775 122.875 196.945 ;
        RECT 120.775 196.695 121.105 196.775 ;
        RECT 116.525 196.605 116.695 196.610 ;
        RECT 116.385 196.330 117.545 196.605 ;
        RECT 116.015 195.970 117.545 196.160 ;
        RECT 117.715 196.150 119.175 196.670 ;
        RECT 115.335 195.630 116.360 195.800 ;
        RECT 117.715 195.790 118.635 196.150 ;
        RECT 119.345 195.980 120.605 196.670 ;
        RECT 113.355 195.345 113.685 195.430 ;
        RECT 114.995 195.345 115.925 195.460 ;
        RECT 112.275 195.015 112.825 195.345 ;
        RECT 112.995 195.175 114.065 195.345 ;
        RECT 112.275 193.450 112.445 195.015 ;
        RECT 112.995 194.800 113.165 195.175 ;
        RECT 112.615 194.630 113.165 194.800 ;
        RECT 113.345 194.540 113.715 194.895 ;
        RECT 113.895 194.800 114.065 195.175 ;
        RECT 114.235 195.290 115.925 195.345 ;
        RECT 114.235 195.015 115.165 195.290 ;
        RECT 113.895 194.630 114.825 194.800 ;
        RECT 114.995 193.450 115.165 195.015 ;
        RECT 115.515 194.880 115.925 195.055 ;
        RECT 116.170 195.050 116.360 195.630 ;
        RECT 116.735 195.060 116.905 195.770 ;
        RECT 117.180 195.460 118.635 195.790 ;
        RECT 118.805 195.460 120.605 195.980 ;
        RECT 120.905 195.755 121.075 196.470 ;
        RECT 121.275 196.415 121.995 196.605 ;
        RECT 122.705 196.540 122.875 196.775 ;
        RECT 123.155 196.720 123.325 197.125 ;
        RECT 123.655 197.250 123.850 197.310 ;
        RECT 124.545 197.265 125.660 197.550 ;
        RECT 124.545 197.250 124.715 197.265 ;
        RECT 123.655 197.080 124.715 197.250 ;
        RECT 125.875 197.220 126.045 197.750 ;
        RECT 126.215 197.620 128.425 198.020 ;
        RECT 128.595 197.680 128.765 199.010 ;
        RECT 129.395 199.345 130.685 199.795 ;
        RECT 130.855 199.470 131.490 199.795 ;
        RECT 131.660 199.650 132.625 199.910 ;
        RECT 129.395 198.950 129.565 199.345 ;
        RECT 128.935 198.670 129.565 198.950 ;
        RECT 129.735 198.480 130.295 199.175 ;
        RECT 130.465 198.950 130.685 199.345 ;
        RECT 131.315 199.465 131.490 199.470 ;
        RECT 132.400 199.475 132.625 199.650 ;
        RECT 132.795 199.645 133.045 205.655 ;
        RECT 134.035 205.485 134.205 206.040 ;
        RECT 134.465 205.610 134.925 205.780 ;
        RECT 133.475 205.440 134.205 205.485 ;
        RECT 133.475 205.225 134.585 205.440 ;
        RECT 134.035 205.110 134.585 205.225 ;
        RECT 134.755 205.345 134.925 205.610 ;
        RECT 135.095 205.515 135.745 205.865 ;
        RECT 136.755 205.785 137.655 206.040 ;
        RECT 135.915 205.610 136.585 205.780 ;
        RECT 135.915 205.345 136.085 205.610 ;
        RECT 136.755 205.440 136.930 205.785 ;
        RECT 137.825 205.615 138.065 206.215 ;
        RECT 134.755 205.115 136.085 205.345 ;
        RECT 136.255 205.185 136.930 205.440 ;
        RECT 137.100 205.355 138.065 205.615 ;
        RECT 136.255 205.110 137.655 205.185 ;
        RECT 133.215 204.795 133.840 205.055 ;
        RECT 133.215 204.195 133.385 204.795 ;
        RECT 134.035 204.625 134.205 205.110 ;
        RECT 134.465 204.755 136.585 204.940 ;
        RECT 136.755 204.925 137.655 205.110 ;
        RECT 133.555 204.500 134.205 204.625 ;
        RECT 133.555 204.365 134.665 204.500 ;
        RECT 134.035 204.250 134.665 204.365 ;
        RECT 134.835 204.305 135.785 204.585 ;
        RECT 136.755 204.515 136.930 204.925 ;
        RECT 137.825 204.755 138.065 205.355 ;
        RECT 136.295 204.325 136.930 204.515 ;
        RECT 137.100 204.495 138.065 204.755 ;
        RECT 136.295 204.250 137.655 204.325 ;
        RECT 133.215 203.935 133.840 204.195 ;
        RECT 133.215 203.335 133.385 203.935 ;
        RECT 134.035 203.765 134.205 204.250 ;
        RECT 134.795 204.080 136.160 204.135 ;
        RECT 133.555 203.505 134.205 203.765 ;
        RECT 134.485 203.965 136.585 204.080 ;
        RECT 134.485 203.910 134.925 203.965 ;
        RECT 134.485 203.745 134.655 203.910 ;
        RECT 136.030 203.830 136.585 203.965 ;
        RECT 136.755 204.065 137.655 204.250 ;
        RECT 133.215 203.075 133.840 203.335 ;
        RECT 133.215 202.490 133.385 203.075 ;
        RECT 134.035 202.905 134.205 203.505 ;
        RECT 133.555 202.660 134.205 202.905 ;
        RECT 134.485 203.045 134.655 203.550 ;
        RECT 134.855 203.385 135.075 203.740 ;
        RECT 135.245 203.555 135.840 203.795 ;
        RECT 134.855 203.215 136.140 203.385 ;
        RECT 134.485 202.875 135.605 203.045 ;
        RECT 135.435 202.685 135.605 202.875 ;
        RECT 135.775 202.855 136.140 203.215 ;
        RECT 136.310 202.685 136.480 203.620 ;
        RECT 134.035 202.555 134.205 202.660 ;
        RECT 133.215 202.215 133.840 202.490 ;
        RECT 133.215 201.630 133.385 202.215 ;
        RECT 134.035 202.185 134.705 202.555 ;
        RECT 134.885 202.465 135.215 202.665 ;
        RECT 135.435 202.515 136.480 202.685 ;
        RECT 136.755 203.465 136.930 204.065 ;
        RECT 137.825 203.895 138.065 204.495 ;
        RECT 137.100 203.635 138.065 203.895 ;
        RECT 136.755 203.205 137.725 203.465 ;
        RECT 136.755 202.605 136.925 203.205 ;
        RECT 138.235 203.035 138.485 209.045 ;
        RECT 138.655 209.040 138.825 209.215 ;
        RECT 138.655 208.780 139.280 209.040 ;
        RECT 138.655 208.180 138.825 208.780 ;
        RECT 139.475 208.610 139.645 209.220 ;
        RECT 140.275 209.465 141.565 209.915 ;
        RECT 141.735 209.590 142.365 209.915 ;
        RECT 143.425 209.855 143.685 210.025 ;
        RECT 143.935 209.905 144.235 210.365 ;
        RECT 144.915 210.185 145.085 210.585 ;
        RECT 145.995 210.500 146.325 210.585 ;
        RECT 140.275 209.070 140.445 209.465 ;
        RECT 139.815 208.790 140.445 209.070 ;
        RECT 138.995 208.360 139.645 208.610 ;
        RECT 140.615 208.600 141.175 209.295 ;
        RECT 141.345 209.070 141.565 209.465 ;
        RECT 141.345 208.790 142.025 209.070 ;
        RECT 138.655 207.920 139.280 208.180 ;
        RECT 138.655 207.320 138.825 207.920 ;
        RECT 139.475 207.800 139.645 208.360 ;
        RECT 139.815 208.200 142.025 208.600 ;
        RECT 142.195 208.120 142.365 209.590 ;
        RECT 142.640 209.685 143.685 209.855 ;
        RECT 143.905 209.705 144.235 209.905 ;
        RECT 144.415 209.985 145.085 210.185 ;
        RECT 145.255 210.330 145.830 210.415 ;
        RECT 146.560 210.330 147.465 210.415 ;
        RECT 145.255 210.160 147.465 210.330 ;
        RECT 147.635 209.985 147.805 210.585 ;
        RECT 144.415 209.815 145.925 209.985 ;
        RECT 144.915 209.725 145.925 209.815 ;
        RECT 146.485 209.725 147.805 209.985 ;
        RECT 142.640 208.750 142.810 209.685 ;
        RECT 142.980 209.155 143.345 209.515 ;
        RECT 143.515 209.495 143.685 209.685 ;
        RECT 143.515 209.325 144.635 209.495 ;
        RECT 142.980 208.985 144.265 209.155 ;
        RECT 143.280 208.575 143.875 208.815 ;
        RECT 144.045 208.630 144.265 208.985 ;
        RECT 144.465 208.820 144.635 209.325 ;
        RECT 142.535 208.405 143.090 208.540 ;
        RECT 144.465 208.460 144.635 208.625 ;
        RECT 144.195 208.405 144.635 208.460 ;
        RECT 142.535 208.290 144.635 208.405 ;
        RECT 144.915 208.490 145.085 209.725 ;
        RECT 145.255 209.380 146.665 209.550 ;
        RECT 147.635 209.540 147.805 209.725 ;
        RECT 145.255 209.060 145.825 209.380 ;
        RECT 145.255 208.660 145.825 208.890 ;
        RECT 145.995 208.805 146.325 209.210 ;
        RECT 146.495 209.030 146.665 209.380 ;
        RECT 146.835 209.210 147.805 209.540 ;
        RECT 146.495 208.780 147.465 209.030 ;
        RECT 142.960 208.235 144.325 208.290 ;
        RECT 144.915 208.120 145.485 208.490 ;
        RECT 140.275 207.820 141.565 208.030 ;
        RECT 139.475 207.750 140.105 207.800 ;
        RECT 138.995 207.530 140.105 207.750 ;
        RECT 138.995 207.500 139.645 207.530 ;
        RECT 138.655 207.060 139.280 207.320 ;
        RECT 138.655 206.475 138.825 207.060 ;
        RECT 139.475 206.890 139.645 207.500 ;
        RECT 140.275 207.360 140.445 207.820 ;
        RECT 139.815 207.075 140.445 207.360 ;
        RECT 140.615 206.960 141.175 207.650 ;
        RECT 141.345 207.360 141.565 207.820 ;
        RECT 142.195 207.855 142.825 208.120 ;
        RECT 144.455 208.070 145.485 208.120 ;
        RECT 142.195 207.800 142.365 207.855 ;
        RECT 141.735 207.530 142.365 207.800 ;
        RECT 143.335 207.785 144.285 208.065 ;
        RECT 144.455 207.870 145.085 208.070 ;
        RECT 145.655 207.900 145.825 208.660 ;
        RECT 145.995 208.340 147.125 208.590 ;
        RECT 141.345 207.075 142.025 207.360 ;
        RECT 142.195 207.260 142.365 207.530 ;
        RECT 142.535 207.430 144.655 207.615 ;
        RECT 144.915 207.560 145.085 207.870 ;
        RECT 145.255 207.730 145.825 207.900 ;
        RECT 145.995 207.940 147.125 208.140 ;
        RECT 145.995 207.895 146.325 207.940 ;
        RECT 147.295 207.770 147.465 208.780 ;
        RECT 144.915 207.260 145.825 207.560 ;
        RECT 145.995 207.320 146.275 207.710 ;
        RECT 146.445 207.600 147.465 207.770 ;
        RECT 138.995 206.645 139.645 206.890 ;
        RECT 138.655 206.200 139.280 206.475 ;
        RECT 139.475 206.330 139.645 206.645 ;
        RECT 142.195 206.930 142.865 207.260 ;
        RECT 143.035 207.025 144.365 207.255 ;
        RECT 142.195 206.330 142.365 206.930 ;
        RECT 143.035 206.760 143.205 207.025 ;
        RECT 142.535 206.590 143.205 206.760 ;
        RECT 143.375 206.505 144.025 206.855 ;
        RECT 144.195 206.760 144.365 207.025 ;
        RECT 144.535 207.110 145.825 207.260 ;
        RECT 146.445 207.150 146.615 207.600 ;
        RECT 147.635 207.430 147.805 209.210 ;
        RECT 144.535 206.930 145.085 207.110 ;
        RECT 145.995 206.980 146.615 207.150 ;
        RECT 146.785 207.115 147.805 207.430 ;
        RECT 144.195 206.590 144.655 206.760 ;
        RECT 138.655 205.615 138.825 206.200 ;
        RECT 139.475 206.040 140.370 206.330 ;
        RECT 141.030 206.040 142.365 206.330 ;
        RECT 144.915 206.330 145.085 206.930 ;
        RECT 145.265 206.810 145.825 206.940 ;
        RECT 146.835 206.810 147.465 206.940 ;
        RECT 145.265 206.500 147.465 206.810 ;
        RECT 147.635 206.330 147.805 207.115 ;
        RECT 142.535 206.070 143.205 206.240 ;
        RECT 139.475 206.030 139.645 206.040 ;
        RECT 138.995 205.785 139.645 206.030 ;
        RECT 142.195 205.900 142.365 206.040 ;
        RECT 138.655 205.355 139.280 205.615 ;
        RECT 139.475 205.440 139.645 205.785 ;
        RECT 139.815 205.695 142.025 205.865 ;
        RECT 139.815 205.610 140.385 205.695 ;
        RECT 141.055 205.530 142.025 205.695 ;
        RECT 142.195 205.570 142.865 205.900 ;
        RECT 143.035 205.805 143.205 206.070 ;
        RECT 143.375 205.975 144.025 206.325 ;
        RECT 144.195 206.070 144.655 206.240 ;
        RECT 144.195 205.805 144.365 206.070 ;
        RECT 144.915 206.040 145.810 206.330 ;
        RECT 146.470 206.040 147.805 206.330 ;
        RECT 144.915 205.900 145.085 206.040 ;
        RECT 143.035 205.575 144.365 205.805 ;
        RECT 144.535 205.570 145.085 205.900 ;
        RECT 140.555 205.440 140.885 205.525 ;
        RECT 138.655 204.755 138.825 205.355 ;
        RECT 139.475 205.185 140.045 205.440 ;
        RECT 138.995 205.110 140.045 205.185 ;
        RECT 140.215 205.270 140.885 205.440 ;
        RECT 142.195 205.360 142.365 205.570 ;
        RECT 138.995 204.925 139.645 205.110 ;
        RECT 138.655 204.495 139.280 204.755 ;
        RECT 138.655 203.895 138.825 204.495 ;
        RECT 139.475 204.325 139.645 204.925 ;
        RECT 140.215 204.685 140.385 205.270 ;
        RECT 141.055 205.190 142.365 205.360 ;
        RECT 142.535 205.215 144.655 205.400 ;
        RECT 140.555 205.020 140.885 205.045 ;
        RECT 140.555 204.850 142.025 205.020 ;
        RECT 138.995 204.065 139.645 204.325 ;
        RECT 139.815 204.680 140.385 204.685 ;
        RECT 139.815 204.510 141.685 204.680 ;
        RECT 139.815 204.155 140.180 204.510 ;
        RECT 140.375 204.170 141.345 204.340 ;
        RECT 138.655 203.635 139.280 203.895 ;
        RECT 139.475 203.465 139.645 204.065 ;
        RECT 140.665 203.965 140.835 203.970 ;
        RECT 139.815 203.690 140.975 203.965 ;
        RECT 141.175 203.520 141.345 204.170 ;
        RECT 141.515 203.555 141.685 204.510 ;
        RECT 138.915 203.205 139.645 203.465 ;
        RECT 139.815 203.330 141.345 203.520 ;
        RECT 139.475 203.150 139.645 203.205 ;
        RECT 141.855 203.160 142.025 204.850 ;
        RECT 137.100 202.785 139.295 203.035 ;
        RECT 134.035 202.045 134.205 202.185 ;
        RECT 133.555 201.800 134.205 202.045 ;
        RECT 134.885 202.005 135.185 202.465 ;
        RECT 135.435 202.345 135.695 202.515 ;
        RECT 136.755 202.345 137.735 202.605 ;
        RECT 135.365 202.175 135.695 202.345 ;
        RECT 135.955 202.175 136.925 202.345 ;
        RECT 133.215 201.370 133.840 201.630 ;
        RECT 133.215 200.770 133.385 201.370 ;
        RECT 134.035 201.190 134.205 201.800 ;
        RECT 134.485 201.835 136.585 202.005 ;
        RECT 134.485 201.600 134.655 201.835 ;
        RECT 136.255 201.755 136.585 201.835 ;
        RECT 136.755 201.745 136.925 202.175 ;
        RECT 138.235 202.175 138.485 202.785 ;
        RECT 139.475 202.640 140.180 203.150 ;
        RECT 139.475 202.605 139.645 202.640 ;
        RECT 138.950 202.345 139.645 202.605 ;
        RECT 140.455 202.420 140.625 203.130 ;
        RECT 138.235 202.170 139.295 202.175 ;
        RECT 137.095 201.925 139.295 202.170 ;
        RECT 135.365 201.475 136.085 201.665 ;
        RECT 133.555 200.940 134.205 201.190 ;
        RECT 133.215 200.510 133.840 200.770 ;
        RECT 133.215 199.910 133.385 200.510 ;
        RECT 134.035 200.370 134.205 200.940 ;
        RECT 134.485 200.815 134.655 201.430 ;
        RECT 134.825 201.305 135.155 201.450 ;
        RECT 134.825 200.985 136.115 201.305 ;
        RECT 136.285 200.815 136.455 201.530 ;
        RECT 134.485 200.645 136.455 200.815 ;
        RECT 136.755 201.450 137.735 201.745 ;
        RECT 136.755 200.715 136.925 201.450 ;
        RECT 138.235 201.440 138.795 201.755 ;
        RECT 139.475 201.745 139.645 202.345 ;
        RECT 139.850 202.240 140.625 202.420 ;
        RECT 141.000 202.990 142.025 203.160 ;
        RECT 142.195 204.975 142.365 205.190 ;
        RECT 142.195 204.710 142.825 204.975 ;
        RECT 143.335 204.765 144.285 205.045 ;
        RECT 144.915 204.960 145.085 205.570 ;
        RECT 144.455 204.710 145.085 204.960 ;
        RECT 141.000 202.410 141.190 202.990 ;
        RECT 142.195 202.820 142.365 204.710 ;
        RECT 142.960 204.540 144.325 204.595 ;
        RECT 142.535 204.425 144.635 204.540 ;
        RECT 142.535 204.290 143.090 204.425 ;
        RECT 144.195 204.370 144.635 204.425 ;
        RECT 142.640 203.145 142.810 204.080 ;
        RECT 143.280 204.015 143.875 204.255 ;
        RECT 144.465 204.205 144.635 204.370 ;
        RECT 144.915 204.380 145.085 204.710 ;
        RECT 145.255 204.550 145.885 204.835 ;
        RECT 144.045 203.845 144.265 204.200 ;
        RECT 144.915 204.110 145.545 204.380 ;
        RECT 142.980 203.675 144.265 203.845 ;
        RECT 142.980 203.315 143.345 203.675 ;
        RECT 144.465 203.505 144.635 204.010 ;
        RECT 143.515 203.335 144.635 203.505 ;
        RECT 143.515 203.145 143.685 203.335 ;
        RECT 142.640 202.975 143.685 203.145 ;
        RECT 141.435 202.805 142.365 202.820 ;
        RECT 143.425 202.805 143.685 202.975 ;
        RECT 143.905 202.925 144.235 203.125 ;
        RECT 144.915 203.015 145.085 204.110 ;
        RECT 145.715 204.090 145.885 204.550 ;
        RECT 146.055 204.260 146.615 204.950 ;
        RECT 146.785 204.550 147.465 204.835 ;
        RECT 146.785 204.090 147.005 204.550 ;
        RECT 147.635 204.380 147.805 206.040 ;
        RECT 147.175 204.110 147.805 204.380 ;
        RECT 145.715 203.880 147.005 204.090 ;
        RECT 145.255 203.310 147.465 203.710 ;
        RECT 141.435 202.650 143.165 202.805 ;
        RECT 142.195 202.635 143.165 202.650 ;
        RECT 143.425 202.635 143.755 202.805 ;
        RECT 141.435 202.240 141.845 202.415 ;
        RECT 139.850 202.175 141.845 202.240 ;
        RECT 140.455 201.900 141.845 202.175 ;
        RECT 138.965 201.440 139.645 201.745 ;
        RECT 137.095 200.990 139.305 201.270 ;
        RECT 137.095 200.885 138.065 200.990 ;
        RECT 138.735 200.885 139.305 200.990 ;
        RECT 139.475 201.105 139.645 201.440 ;
        RECT 139.475 200.865 140.155 201.105 ;
        RECT 138.235 200.715 138.565 200.820 ;
        RECT 139.475 200.715 139.645 200.865 ;
        RECT 140.325 200.855 140.885 201.210 ;
        RECT 134.035 200.330 134.735 200.370 ;
        RECT 133.555 200.160 134.735 200.330 ;
        RECT 133.555 200.080 134.205 200.160 ;
        RECT 133.215 199.650 133.840 199.910 ;
        RECT 133.215 199.475 133.385 199.650 ;
        RECT 131.315 199.210 132.215 199.465 ;
        RECT 130.465 198.670 131.145 198.950 ;
        RECT 131.315 198.580 131.485 199.210 ;
        RECT 132.400 199.040 133.385 199.475 ;
        RECT 134.035 199.470 134.205 200.080 ;
        RECT 135.115 199.940 135.445 200.645 ;
        RECT 135.650 199.920 136.025 200.475 ;
        RECT 136.755 200.465 137.385 200.715 ;
        RECT 136.255 200.390 137.385 200.465 ;
        RECT 136.255 200.150 136.925 200.390 ;
        RECT 134.420 199.770 134.945 199.900 ;
        RECT 135.650 199.770 136.585 199.920 ;
        RECT 134.420 199.580 136.585 199.770 ;
        RECT 134.420 199.570 135.445 199.580 ;
        RECT 133.555 199.400 134.205 199.470 ;
        RECT 133.555 199.230 134.815 199.400 ;
        RECT 133.555 199.210 134.205 199.230 ;
        RECT 131.660 198.780 133.840 199.040 ;
        RECT 131.660 198.750 133.385 198.780 ;
        RECT 128.935 198.080 131.145 198.480 ;
        RECT 131.315 198.310 132.230 198.580 ;
        RECT 132.400 198.310 133.385 198.750 ;
        RECT 134.035 198.610 134.205 199.210 ;
        RECT 134.425 198.905 134.945 199.060 ;
        RECT 135.115 199.020 135.445 199.570 ;
        RECT 136.755 199.410 136.925 200.150 ;
        RECT 137.555 200.265 138.845 200.715 ;
        RECT 139.015 200.390 139.645 200.715 ;
        RECT 141.055 200.695 141.400 201.085 ;
        RECT 142.195 200.925 142.365 202.635 ;
        RECT 143.935 202.465 144.235 202.925 ;
        RECT 144.415 202.645 145.085 203.015 ;
        RECT 145.255 202.840 145.885 203.120 ;
        RECT 142.535 202.295 144.635 202.465 ;
        RECT 142.535 202.215 142.865 202.295 ;
        RECT 142.665 201.275 142.835 201.990 ;
        RECT 143.035 201.935 143.755 202.125 ;
        RECT 144.465 202.060 144.635 202.295 ;
        RECT 144.915 202.320 145.085 202.645 ;
        RECT 145.715 202.445 145.885 202.840 ;
        RECT 146.055 202.615 146.615 203.310 ;
        RECT 146.785 202.840 147.465 203.120 ;
        RECT 146.785 202.445 147.005 202.840 ;
        RECT 144.915 201.995 145.545 202.320 ;
        RECT 145.715 201.995 147.005 202.445 ;
        RECT 147.635 202.320 147.805 204.110 ;
        RECT 147.175 201.995 147.805 202.320 ;
        RECT 143.965 201.765 144.295 201.910 ;
        RECT 143.005 201.445 144.295 201.765 ;
        RECT 144.465 201.275 144.635 201.890 ;
        RECT 142.665 201.105 144.635 201.275 ;
        RECT 141.055 200.685 141.225 200.695 ;
        RECT 139.825 200.515 141.225 200.685 ;
        RECT 139.825 200.405 140.155 200.515 ;
        RECT 137.555 199.870 137.775 200.265 ;
        RECT 137.095 199.590 137.775 199.870 ;
        RECT 135.745 199.240 136.925 199.410 ;
        RECT 137.945 199.400 138.505 200.095 ;
        RECT 138.675 199.870 138.845 200.265 ;
        RECT 139.475 200.175 139.645 200.390 ;
        RECT 139.475 199.960 140.155 200.175 ;
        RECT 140.325 200.080 140.885 200.345 ;
        RECT 138.675 199.590 139.305 199.870 ;
        RECT 134.425 198.850 134.985 198.905 ;
        RECT 135.615 198.895 136.540 199.070 ;
        RECT 135.565 198.850 136.540 198.895 ;
        RECT 134.425 198.740 136.540 198.850 ;
        RECT 134.425 198.730 135.695 198.740 ;
        RECT 134.860 198.680 135.695 198.730 ;
        RECT 133.555 198.310 134.205 198.610 ;
        RECT 129.395 197.700 130.685 197.910 ;
        RECT 126.675 197.240 127.965 197.450 ;
        RECT 122.205 196.245 122.535 196.390 ;
        RECT 121.245 195.925 122.535 196.245 ;
        RECT 122.705 195.755 122.875 196.370 ;
        RECT 120.905 195.585 122.875 195.755 ;
        RECT 123.155 196.320 123.820 196.720 ;
        RECT 124.185 196.690 124.715 197.080 ;
        RECT 123.155 195.730 123.325 196.320 ;
        RECT 124.185 196.260 124.565 196.690 ;
        RECT 124.885 196.395 125.195 197.090 ;
        RECT 125.875 197.085 126.505 197.220 ;
        RECT 125.405 196.950 126.505 197.085 ;
        RECT 125.405 196.400 126.045 196.950 ;
        RECT 126.675 196.780 126.895 197.240 ;
        RECT 126.215 196.495 126.895 196.780 ;
        RECT 123.495 196.090 124.015 196.150 ;
        RECT 124.820 196.090 125.605 196.220 ;
        RECT 123.495 195.915 125.605 196.090 ;
        RECT 125.875 196.210 126.045 196.400 ;
        RECT 127.065 196.380 127.625 197.070 ;
        RECT 127.795 196.780 127.965 197.240 ;
        RECT 128.595 197.410 129.225 197.680 ;
        RECT 128.595 197.220 128.765 197.410 ;
        RECT 129.395 197.240 129.565 197.700 ;
        RECT 128.135 196.950 128.765 197.220 ;
        RECT 128.935 196.955 129.565 197.240 ;
        RECT 127.795 196.495 128.425 196.780 ;
        RECT 128.595 196.670 128.765 196.950 ;
        RECT 129.735 196.840 130.295 197.530 ;
        RECT 130.465 197.240 130.685 197.700 ;
        RECT 131.315 197.680 131.485 198.310 ;
        RECT 134.035 198.050 134.205 198.310 ;
        RECT 136.755 198.600 136.925 199.240 ;
        RECT 137.095 199.000 139.305 199.400 ;
        RECT 139.475 198.910 139.645 199.960 ;
        RECT 141.055 199.830 141.225 200.515 ;
        RECT 142.195 200.610 142.865 200.925 ;
        RECT 142.195 200.210 142.365 200.610 ;
        RECT 143.095 200.380 143.470 200.935 ;
        RECT 143.675 200.400 144.005 201.105 ;
        RECT 144.915 200.830 145.085 201.995 ;
        RECT 145.995 201.890 146.325 201.995 ;
        RECT 145.255 201.720 145.825 201.825 ;
        RECT 146.495 201.720 147.465 201.825 ;
        RECT 145.255 201.440 147.465 201.720 ;
        RECT 144.385 200.620 145.085 200.830 ;
        RECT 141.395 199.880 142.365 200.210 ;
        RECT 142.535 200.230 143.470 200.380 ;
        RECT 144.175 200.230 144.700 200.360 ;
        RECT 142.535 200.040 144.700 200.230 ;
        RECT 139.815 199.490 140.385 199.790 ;
        RECT 140.555 199.660 141.225 199.830 ;
        RECT 142.195 199.870 142.365 199.880 ;
        RECT 143.675 200.030 144.700 200.040 ;
        RECT 144.915 200.345 145.085 200.620 ;
        RECT 147.635 200.345 147.805 201.995 ;
        RECT 144.915 200.085 145.925 200.345 ;
        RECT 146.485 200.085 147.805 200.345 ;
        RECT 141.405 199.490 142.025 199.710 ;
        RECT 139.815 199.175 142.025 199.490 ;
        RECT 142.195 199.700 143.375 199.870 ;
        RECT 142.195 198.910 142.365 199.700 ;
        RECT 142.580 199.355 143.505 199.530 ;
        RECT 143.675 199.480 144.005 200.030 ;
        RECT 144.915 199.860 145.085 200.085 ;
        RECT 144.305 199.690 145.085 199.860 ;
        RECT 144.175 199.365 144.695 199.520 ;
        RECT 142.580 199.310 143.555 199.355 ;
        RECT 144.135 199.310 144.695 199.365 ;
        RECT 142.580 199.200 144.695 199.310 ;
        RECT 143.425 199.190 144.695 199.200 ;
        RECT 144.915 199.485 145.085 199.690 ;
        RECT 145.255 199.740 147.465 199.910 ;
        RECT 145.255 199.655 145.830 199.740 ;
        RECT 146.560 199.655 147.465 199.740 ;
        RECT 145.995 199.485 146.325 199.570 ;
        RECT 147.635 199.485 147.805 200.085 ;
        RECT 143.425 199.140 144.260 199.190 ;
        RECT 144.915 199.155 145.465 199.485 ;
        RECT 145.635 199.315 146.705 199.485 ;
        RECT 137.555 198.620 138.845 198.830 ;
        RECT 136.755 198.330 137.385 198.600 ;
        RECT 136.755 198.050 136.925 198.330 ;
        RECT 137.555 198.160 137.775 198.620 ;
        RECT 130.855 197.495 131.485 197.680 ;
        RECT 131.655 197.770 133.865 198.050 ;
        RECT 131.655 197.665 132.625 197.770 ;
        RECT 133.295 197.665 133.865 197.770 ;
        RECT 134.035 197.780 134.840 198.050 ;
        RECT 135.800 197.780 136.925 198.050 ;
        RECT 137.095 197.875 137.775 198.160 ;
        RECT 132.795 197.495 133.125 197.600 ;
        RECT 134.035 197.495 134.205 197.780 ;
        RECT 130.855 197.410 131.945 197.495 ;
        RECT 130.465 196.955 131.145 197.240 ;
        RECT 131.315 197.170 131.945 197.410 ;
        RECT 131.315 196.670 131.485 197.170 ;
        RECT 128.595 196.210 130.055 196.670 ;
        RECT 125.875 195.730 127.135 196.210 ;
        RECT 117.180 195.280 117.885 195.460 ;
        RECT 116.735 194.880 117.510 195.060 ;
        RECT 115.515 194.815 117.510 194.880 ;
        RECT 117.715 194.850 117.885 195.280 ;
        RECT 120.435 195.405 120.605 195.460 ;
        RECT 118.055 195.030 118.605 195.200 ;
        RECT 115.515 194.540 116.905 194.815 ;
        RECT 117.715 194.520 118.265 194.850 ;
        RECT 118.435 194.705 118.605 195.030 ;
        RECT 118.785 194.940 119.155 195.270 ;
        RECT 119.335 195.030 120.265 195.200 ;
        RECT 120.435 195.090 121.105 195.405 ;
        RECT 119.335 194.705 119.505 195.030 ;
        RECT 120.435 194.850 120.605 195.090 ;
        RECT 121.335 194.860 121.710 195.415 ;
        RECT 121.915 194.880 122.245 195.585 ;
        RECT 123.155 195.460 123.960 195.730 ;
        RECT 124.920 195.460 127.135 195.730 ;
        RECT 123.155 195.310 123.325 195.460 ;
        RECT 122.625 195.290 123.325 195.310 ;
        RECT 125.875 195.290 127.135 195.460 ;
        RECT 122.625 195.100 124.615 195.290 ;
        RECT 118.435 194.535 119.505 194.705 ;
        RECT 117.715 193.470 117.885 194.520 ;
        RECT 118.860 194.420 119.190 194.535 ;
        RECT 119.675 194.520 120.605 194.850 ;
        RECT 120.775 194.710 121.710 194.860 ;
        RECT 122.415 194.710 122.940 194.840 ;
        RECT 120.775 194.520 122.940 194.710 ;
        RECT 120.435 194.350 120.605 194.520 ;
        RECT 121.915 194.510 122.940 194.520 ;
        RECT 118.055 194.250 118.560 194.340 ;
        RECT 119.360 194.250 120.265 194.350 ;
        RECT 118.055 194.080 120.265 194.250 ;
        RECT 120.435 194.180 121.615 194.350 ;
        RECT 118.055 193.650 118.605 193.820 ;
        RECT 117.715 193.450 118.265 193.470 ;
        RECT 112.275 193.160 113.170 193.450 ;
        RECT 113.830 193.160 116.330 193.450 ;
        RECT 116.990 193.160 118.265 193.450 ;
        RECT 112.275 191.595 112.445 193.160 ;
        RECT 114.995 192.435 115.165 193.160 ;
        RECT 117.715 193.140 118.265 193.160 ;
        RECT 118.435 193.325 118.605 193.650 ;
        RECT 118.785 193.560 119.155 193.890 ;
        RECT 119.335 193.650 120.265 193.820 ;
        RECT 119.335 193.325 119.505 193.650 ;
        RECT 120.435 193.470 120.605 194.180 ;
        RECT 120.820 193.835 121.745 194.010 ;
        RECT 121.915 193.960 122.245 194.510 ;
        RECT 123.155 194.340 124.615 195.100 ;
        RECT 122.545 194.170 124.615 194.340 ;
        RECT 123.155 194.080 124.615 194.170 ;
        RECT 124.785 194.830 127.135 195.290 ;
        RECT 127.305 196.150 130.055 196.210 ;
        RECT 127.305 195.460 129.515 196.150 ;
        RECT 130.225 195.980 131.485 196.670 ;
        RECT 132.115 197.045 133.405 197.495 ;
        RECT 133.575 197.190 134.205 197.495 ;
        RECT 134.375 197.420 136.485 197.595 ;
        RECT 134.375 197.360 134.895 197.420 ;
        RECT 135.700 197.290 136.485 197.420 ;
        RECT 136.755 197.590 136.925 197.780 ;
        RECT 137.945 197.760 138.505 198.450 ;
        RECT 138.675 198.160 138.845 198.620 ;
        RECT 139.475 198.700 140.465 198.910 ;
        RECT 141.055 198.700 142.365 198.910 ;
        RECT 139.475 198.600 139.645 198.700 ;
        RECT 139.015 198.330 139.645 198.600 ;
        RECT 138.675 197.875 139.305 198.160 ;
        RECT 139.475 198.030 139.645 198.330 ;
        RECT 139.815 198.280 142.025 198.530 ;
        RECT 139.815 198.200 140.445 198.280 ;
        RECT 141.045 198.200 142.025 198.280 ;
        RECT 142.195 198.230 142.365 198.700 ;
        RECT 142.535 198.620 144.745 198.935 ;
        RECT 142.535 198.400 143.155 198.620 ;
        RECT 143.335 198.280 144.005 198.450 ;
        RECT 144.175 198.320 144.745 198.620 ;
        RECT 139.475 197.800 140.465 198.030 ;
        RECT 139.475 197.590 139.645 197.800 ;
        RECT 140.635 197.780 140.885 198.110 ;
        RECT 142.195 198.030 143.165 198.230 ;
        RECT 141.055 197.900 143.165 198.030 ;
        RECT 141.055 197.800 142.365 197.900 ;
        RECT 133.575 197.170 134.700 197.190 ;
        RECT 132.115 196.650 132.335 197.045 ;
        RECT 131.655 196.370 132.335 196.650 ;
        RECT 132.505 196.180 133.065 196.875 ;
        RECT 133.235 196.650 133.405 197.045 ;
        RECT 134.035 196.790 134.700 197.170 ;
        RECT 135.065 196.820 135.445 197.250 ;
        RECT 133.235 196.370 133.865 196.650 ;
        RECT 129.685 195.460 131.485 195.980 ;
        RECT 131.655 195.780 133.865 196.180 ;
        RECT 127.305 195.000 128.765 195.460 ;
        RECT 131.315 195.380 131.485 195.460 ;
        RECT 132.115 195.400 133.405 195.610 ;
        RECT 129.095 195.120 131.145 195.290 ;
        RECT 129.095 195.015 129.440 195.120 ;
        RECT 130.175 195.015 131.145 195.120 ;
        RECT 131.315 195.110 131.945 195.380 ;
        RECT 122.415 193.845 122.935 194.000 ;
        RECT 120.820 193.790 121.795 193.835 ;
        RECT 122.375 193.790 122.935 193.845 ;
        RECT 120.820 193.680 122.935 193.790 ;
        RECT 121.665 193.670 122.935 193.680 ;
        RECT 121.665 193.620 122.500 193.670 ;
        RECT 118.435 193.155 119.505 193.325 ;
        RECT 119.675 193.450 120.605 193.470 ;
        RECT 123.155 193.450 124.095 194.080 ;
        RECT 124.785 193.910 127.655 194.830 ;
        RECT 119.675 193.160 121.770 193.450 ;
        RECT 122.430 193.160 124.095 193.450 ;
        RECT 115.335 192.710 117.545 192.990 ;
        RECT 115.335 192.605 116.305 192.710 ;
        RECT 116.975 192.605 117.545 192.710 ;
        RECT 116.475 192.435 116.805 192.540 ;
        RECT 117.715 192.435 117.885 193.140 ;
        RECT 118.860 193.040 119.190 193.155 ;
        RECT 119.675 193.140 120.605 193.160 ;
        RECT 118.055 192.870 118.560 192.960 ;
        RECT 119.360 192.870 120.265 192.970 ;
        RECT 118.055 192.700 120.265 192.870 ;
        RECT 114.995 192.110 115.625 192.435 ;
        RECT 112.615 191.810 113.165 191.980 ;
        RECT 112.275 191.265 112.825 191.595 ;
        RECT 112.995 191.435 113.165 191.810 ;
        RECT 113.345 191.715 113.715 192.070 ;
        RECT 113.895 191.810 114.825 191.980 ;
        RECT 113.895 191.435 114.065 191.810 ;
        RECT 114.995 191.595 115.165 192.110 ;
        RECT 112.995 191.265 114.065 191.435 ;
        RECT 114.235 191.265 115.165 191.595 ;
        RECT 115.795 191.985 117.085 192.435 ;
        RECT 117.255 192.110 117.885 192.435 ;
        RECT 118.055 192.270 118.605 192.440 ;
        RECT 115.795 191.590 116.015 191.985 ;
        RECT 115.335 191.310 116.015 191.590 ;
        RECT 112.275 190.665 112.445 191.265 ;
        RECT 113.355 191.180 113.685 191.265 ;
        RECT 112.615 191.010 113.190 191.095 ;
        RECT 113.920 191.010 114.825 191.095 ;
        RECT 112.615 190.840 114.825 191.010 ;
        RECT 114.995 190.665 115.165 191.265 ;
        RECT 116.185 191.120 116.745 191.815 ;
        RECT 116.915 191.590 117.085 191.985 ;
        RECT 117.715 192.090 117.885 192.110 ;
        RECT 117.715 191.760 118.265 192.090 ;
        RECT 118.435 191.945 118.605 192.270 ;
        RECT 118.785 192.180 119.155 192.510 ;
        RECT 120.435 192.480 120.605 193.140 ;
        RECT 120.775 192.815 122.985 192.985 ;
        RECT 120.775 192.650 121.745 192.815 ;
        RECT 122.415 192.730 122.985 192.815 ;
        RECT 123.155 192.700 124.095 193.160 ;
        RECT 124.265 193.620 127.655 193.910 ;
        RECT 127.825 194.825 128.765 195.000 ;
        RECT 129.675 194.845 130.005 194.950 ;
        RECT 127.825 194.445 129.165 194.825 ;
        RECT 129.335 194.675 130.345 194.845 ;
        RECT 131.315 194.805 131.485 195.110 ;
        RECT 132.115 194.940 132.335 195.400 ;
        RECT 127.825 193.935 128.765 194.445 ;
        RECT 129.335 194.275 129.505 194.675 ;
        RECT 128.985 194.105 129.505 194.275 ;
        RECT 129.675 194.125 130.005 194.505 ;
        RECT 130.175 194.355 130.345 194.675 ;
        RECT 130.515 194.525 131.485 194.805 ;
        RECT 131.655 194.655 132.335 194.940 ;
        RECT 132.505 194.540 133.065 195.230 ;
        RECT 133.235 194.940 133.405 195.400 ;
        RECT 134.035 195.380 134.205 196.790 ;
        RECT 135.065 196.430 135.595 196.820 ;
        RECT 134.535 196.260 135.595 196.430 ;
        RECT 135.765 196.420 136.075 197.115 ;
        RECT 136.755 197.110 138.015 197.590 ;
        RECT 136.285 196.900 138.015 197.110 ;
        RECT 138.185 197.160 139.645 197.590 ;
        RECT 139.905 197.330 140.365 197.500 ;
        RECT 138.185 197.070 140.025 197.160 ;
        RECT 136.285 196.425 138.555 196.900 ;
        RECT 134.535 196.200 134.730 196.260 ;
        RECT 134.390 196.030 134.730 196.200 ;
        RECT 135.425 196.245 135.595 196.260 ;
        RECT 136.755 196.380 138.555 196.425 ;
        RECT 138.725 196.830 140.025 197.070 ;
        RECT 140.195 197.065 140.365 197.330 ;
        RECT 140.535 197.235 141.185 197.585 ;
        RECT 141.355 197.330 142.025 197.500 ;
        RECT 141.355 197.065 141.525 197.330 ;
        RECT 142.195 197.160 142.365 197.800 ;
        RECT 143.335 197.595 143.505 198.280 ;
        RECT 144.915 198.150 145.085 199.155 ;
        RECT 145.635 198.940 145.805 199.315 ;
        RECT 145.255 198.770 145.805 198.940 ;
        RECT 145.985 198.680 146.355 199.035 ;
        RECT 146.535 198.940 146.705 199.315 ;
        RECT 146.875 199.155 147.805 199.485 ;
        RECT 146.535 198.770 147.465 198.940 ;
        RECT 143.675 197.765 144.235 198.030 ;
        RECT 144.405 197.940 145.085 198.150 ;
        RECT 145.255 198.110 145.885 198.395 ;
        RECT 144.405 197.935 145.545 197.940 ;
        RECT 144.405 197.595 144.735 197.705 ;
        RECT 143.335 197.425 144.735 197.595 ;
        RECT 144.915 197.670 145.545 197.935 ;
        RECT 143.335 197.415 143.505 197.425 ;
        RECT 140.195 196.835 141.525 197.065 ;
        RECT 141.695 196.830 142.365 197.160 ;
        RECT 143.160 197.025 143.505 197.415 ;
        RECT 143.675 196.900 144.235 197.255 ;
        RECT 144.915 197.245 145.085 197.670 ;
        RECT 145.715 197.650 145.885 198.110 ;
        RECT 146.055 197.820 146.615 198.510 ;
        RECT 146.785 198.110 147.465 198.395 ;
        RECT 146.785 197.650 147.005 198.110 ;
        RECT 147.635 197.940 147.805 199.155 ;
        RECT 147.175 197.670 147.805 197.940 ;
        RECT 145.715 197.440 147.005 197.650 ;
        RECT 144.405 197.005 145.085 197.245 ;
        RECT 138.725 196.380 139.645 196.830 ;
        RECT 139.905 196.475 142.025 196.660 ;
        RECT 134.925 195.770 135.255 196.090 ;
        RECT 135.425 195.960 136.540 196.245 ;
        RECT 134.925 195.750 136.135 195.770 ;
        RECT 136.755 195.760 136.925 196.380 ;
        RECT 139.475 196.220 139.645 196.380 ;
        RECT 134.400 195.535 136.135 195.750 ;
        RECT 134.400 195.510 134.775 195.535 ;
        RECT 133.575 195.340 134.205 195.380 ;
        RECT 133.575 195.110 134.710 195.340 ;
        RECT 134.035 195.010 134.710 195.110 ;
        RECT 134.885 195.065 135.735 195.365 ;
        RECT 135.905 195.260 136.135 195.535 ;
        RECT 136.305 195.430 136.925 195.760 ;
        RECT 135.905 195.090 136.565 195.260 ;
        RECT 134.885 195.060 135.055 195.065 ;
        RECT 133.235 194.655 133.865 194.940 ;
        RECT 130.175 194.185 130.635 194.355 ;
        RECT 127.825 193.620 129.165 193.935 ;
        RECT 124.265 193.450 126.045 193.620 ;
        RECT 128.595 193.605 129.165 193.620 ;
        RECT 128.595 193.450 128.765 193.605 ;
        RECT 124.265 193.160 127.210 193.450 ;
        RECT 127.870 193.160 128.765 193.450 ;
        RECT 129.335 193.430 129.505 194.105 ;
        RECT 128.985 193.260 129.505 193.430 ;
        RECT 129.675 193.215 130.295 193.955 ;
        RECT 124.265 192.700 126.045 193.160 ;
        RECT 128.595 193.060 128.765 193.160 ;
        RECT 121.915 192.560 122.245 192.645 ;
        RECT 123.155 192.560 123.325 192.700 ;
        RECT 119.335 192.270 120.265 192.440 ;
        RECT 120.435 192.310 121.745 192.480 ;
        RECT 121.915 192.390 122.585 192.560 ;
        RECT 119.335 191.945 119.505 192.270 ;
        RECT 120.435 192.090 120.605 192.310 ;
        RECT 121.915 192.140 122.245 192.165 ;
        RECT 118.435 191.775 119.505 191.945 ;
        RECT 116.915 191.310 117.545 191.590 ;
        RECT 115.335 190.720 117.545 191.120 ;
        RECT 112.275 190.405 113.285 190.665 ;
        RECT 113.845 190.405 115.165 190.665 ;
        RECT 117.715 190.710 117.885 191.760 ;
        RECT 118.860 191.660 119.190 191.775 ;
        RECT 119.675 191.760 120.605 192.090 ;
        RECT 118.055 191.490 118.560 191.580 ;
        RECT 119.360 191.490 120.265 191.590 ;
        RECT 118.055 191.320 120.265 191.490 ;
        RECT 118.055 190.890 118.605 191.060 ;
        RECT 112.275 189.790 112.445 190.405 ;
        RECT 114.995 190.320 115.165 190.405 ;
        RECT 115.795 190.340 117.085 190.550 ;
        RECT 112.615 190.050 114.825 190.230 ;
        RECT 112.615 189.970 113.120 190.050 ;
        RECT 113.920 189.960 114.825 190.050 ;
        RECT 114.995 190.050 115.625 190.320 ;
        RECT 112.275 189.460 112.825 189.790 ;
        RECT 113.420 189.775 113.750 189.880 ;
        RECT 114.995 189.790 115.165 190.050 ;
        RECT 115.795 189.880 116.015 190.340 ;
        RECT 112.995 189.605 114.065 189.775 ;
        RECT 112.275 187.925 112.445 189.460 ;
        RECT 112.995 189.280 113.165 189.605 ;
        RECT 112.615 189.110 113.165 189.280 ;
        RECT 113.345 189.040 113.715 189.380 ;
        RECT 113.895 189.280 114.065 189.605 ;
        RECT 114.235 189.460 115.165 189.790 ;
        RECT 115.335 189.595 116.015 189.880 ;
        RECT 116.185 189.480 116.745 190.170 ;
        RECT 116.915 189.880 117.085 190.340 ;
        RECT 117.715 190.380 118.265 190.710 ;
        RECT 118.435 190.565 118.605 190.890 ;
        RECT 118.785 190.800 119.155 191.130 ;
        RECT 119.335 190.890 120.265 191.060 ;
        RECT 119.335 190.565 119.505 190.890 ;
        RECT 120.435 190.710 120.605 191.760 ;
        RECT 118.435 190.395 119.505 190.565 ;
        RECT 117.715 190.320 117.885 190.380 ;
        RECT 117.255 190.050 117.885 190.320 ;
        RECT 118.860 190.280 119.190 190.395 ;
        RECT 119.675 190.380 120.605 190.710 ;
        RECT 116.915 189.595 117.545 189.880 ;
        RECT 117.715 189.760 117.885 190.050 ;
        RECT 118.055 190.110 118.560 190.200 ;
        RECT 119.360 190.110 120.265 190.210 ;
        RECT 118.055 189.940 120.265 190.110 ;
        RECT 120.435 189.940 120.605 190.380 ;
        RECT 120.775 191.970 122.245 192.140 ;
        RECT 120.775 190.280 120.945 191.970 ;
        RECT 122.415 191.805 122.585 192.390 ;
        RECT 122.755 192.230 123.325 192.560 ;
        RECT 122.415 191.800 122.985 191.805 ;
        RECT 121.115 191.630 122.985 191.800 ;
        RECT 121.115 190.675 121.285 191.630 ;
        RECT 121.455 191.290 122.425 191.460 ;
        RECT 121.455 190.640 121.625 191.290 ;
        RECT 122.620 191.275 122.985 191.630 ;
        RECT 123.155 191.500 123.325 192.230 ;
        RECT 123.495 191.670 124.125 191.955 ;
        RECT 123.155 191.230 123.785 191.500 ;
        RECT 122.645 191.085 122.815 191.090 ;
        RECT 121.825 190.810 122.985 191.085 ;
        RECT 121.455 190.450 122.985 190.640 ;
        RECT 120.775 190.110 121.800 190.280 ;
        RECT 123.155 190.270 123.325 191.230 ;
        RECT 123.955 191.210 124.125 191.670 ;
        RECT 124.295 191.380 124.855 192.070 ;
        RECT 125.025 191.670 125.705 191.955 ;
        RECT 125.875 191.700 126.045 192.700 ;
        RECT 126.685 192.690 128.025 192.815 ;
        RECT 126.255 192.645 128.025 192.690 ;
        RECT 128.595 192.730 129.265 193.060 ;
        RECT 130.465 193.045 130.635 194.185 ;
        RECT 128.595 192.660 128.765 192.730 ;
        RECT 126.255 192.360 126.855 192.645 ;
        RECT 127.025 192.230 127.685 192.475 ;
        RECT 126.265 191.930 126.855 192.180 ;
        RECT 127.855 192.160 128.025 192.645 ;
        RECT 128.195 192.330 128.765 192.660 ;
        RECT 129.675 192.535 130.005 192.945 ;
        RECT 130.175 192.725 130.635 193.045 ;
        RECT 125.025 191.210 125.245 191.670 ;
        RECT 125.875 191.500 126.515 191.700 ;
        RECT 125.415 191.370 126.515 191.500 ;
        RECT 125.415 191.230 126.045 191.370 ;
        RECT 123.955 191.000 125.245 191.210 ;
        RECT 123.495 190.430 125.705 190.830 ;
        RECT 125.875 190.700 126.045 191.230 ;
        RECT 126.685 191.140 126.855 191.930 ;
        RECT 127.025 191.750 127.685 192.015 ;
        RECT 127.855 191.830 128.365 192.160 ;
        RECT 128.595 192.120 128.765 192.330 ;
        RECT 128.985 192.530 130.005 192.535 ;
        RECT 128.985 192.290 130.600 192.530 ;
        RECT 130.805 192.305 131.095 194.355 ;
        RECT 131.315 193.450 131.485 194.525 ;
        RECT 134.035 193.450 134.205 195.010 ;
        RECT 136.755 194.380 136.925 195.430 ;
        RECT 137.145 194.550 137.435 196.205 ;
        RECT 137.605 195.885 138.065 196.205 ;
        RECT 137.605 194.785 137.775 195.885 ;
        RECT 138.235 195.855 138.805 196.205 ;
        RECT 139.475 196.200 140.105 196.220 ;
        RECT 138.975 195.970 140.105 196.200 ;
        RECT 140.275 196.025 141.225 196.305 ;
        RECT 142.195 196.235 142.365 196.830 ;
        RECT 142.535 196.410 143.465 196.580 ;
        RECT 141.735 196.195 142.365 196.235 ;
        RECT 141.735 195.970 143.125 196.195 ;
        RECT 138.975 195.870 139.645 195.970 ;
        RECT 137.945 194.975 138.565 195.685 ;
        RECT 138.735 195.500 139.255 195.670 ;
        RECT 137.605 194.615 138.065 194.785 ;
        RECT 136.755 194.100 137.725 194.380 ;
        RECT 137.895 194.230 138.065 194.615 ;
        RECT 138.235 194.400 138.565 194.805 ;
        RECT 138.735 194.800 138.905 195.500 ;
        RECT 139.475 195.300 139.645 195.870 ;
        RECT 142.195 195.865 143.125 195.970 ;
        RECT 143.295 196.035 143.465 196.410 ;
        RECT 143.645 196.315 144.015 196.670 ;
        RECT 144.195 196.410 144.745 196.580 ;
        RECT 144.195 196.035 144.365 196.410 ;
        RECT 144.915 196.195 145.085 197.005 ;
        RECT 145.255 196.870 147.465 197.270 ;
        RECT 145.255 196.400 145.885 196.680 ;
        RECT 143.295 195.865 144.365 196.035 ;
        RECT 144.535 195.880 145.085 196.195 ;
        RECT 145.715 196.005 145.885 196.400 ;
        RECT 146.055 196.175 146.615 196.870 ;
        RECT 146.785 196.400 147.465 196.680 ;
        RECT 146.785 196.005 147.005 196.400 ;
        RECT 144.535 195.865 145.545 195.880 ;
        RECT 140.235 195.800 141.600 195.855 ;
        RECT 139.925 195.685 142.025 195.800 ;
        RECT 139.925 195.630 140.365 195.685 ;
        RECT 139.925 195.465 140.095 195.630 ;
        RECT 141.470 195.550 142.025 195.685 ;
        RECT 139.075 194.970 139.645 195.300 ;
        RECT 138.735 194.630 139.255 194.800 ;
        RECT 138.735 194.230 138.905 194.630 ;
        RECT 139.475 194.460 139.645 194.970 ;
        RECT 139.925 194.765 140.095 195.270 ;
        RECT 140.295 195.105 140.515 195.460 ;
        RECT 140.685 195.275 141.280 195.515 ;
        RECT 140.295 194.935 141.580 195.105 ;
        RECT 139.925 194.595 141.045 194.765 ;
        RECT 134.385 193.600 136.585 193.910 ;
        RECT 134.385 193.470 134.945 193.600 ;
        RECT 135.955 193.470 136.585 193.600 ;
        RECT 131.315 193.160 132.650 193.450 ;
        RECT 133.310 193.300 134.205 193.450 ;
        RECT 136.755 193.450 136.925 194.100 ;
        RECT 137.895 194.060 138.905 194.230 ;
        RECT 139.075 194.275 139.645 194.460 ;
        RECT 140.875 194.405 141.045 194.595 ;
        RECT 141.215 194.575 141.580 194.935 ;
        RECT 141.750 194.405 141.920 195.340 ;
        RECT 139.075 194.080 140.145 194.275 ;
        RECT 138.235 193.960 138.565 194.060 ;
        RECT 139.475 193.905 140.145 194.080 ;
        RECT 140.325 194.185 140.655 194.385 ;
        RECT 140.875 194.235 141.920 194.405 ;
        RECT 142.195 195.265 142.365 195.865 ;
        RECT 143.675 195.780 144.005 195.865 ;
        RECT 142.535 195.610 143.440 195.695 ;
        RECT 144.170 195.610 144.745 195.695 ;
        RECT 142.535 195.440 144.745 195.610 ;
        RECT 144.915 195.555 145.545 195.865 ;
        RECT 145.715 195.555 147.005 196.005 ;
        RECT 147.635 195.880 147.805 197.670 ;
        RECT 147.175 195.555 147.805 195.880 ;
        RECT 144.915 195.265 145.085 195.555 ;
        RECT 145.995 195.450 146.325 195.555 ;
        RECT 142.195 195.005 143.515 195.265 ;
        RECT 144.075 195.005 145.085 195.265 ;
        RECT 142.195 194.790 142.365 195.005 ;
        RECT 142.195 194.560 143.505 194.790 ;
        RECT 137.095 193.790 138.065 193.890 ;
        RECT 138.800 193.790 139.145 193.890 ;
        RECT 137.095 193.620 139.145 193.790 ;
        RECT 139.475 193.450 139.645 193.905 ;
        RECT 140.325 193.725 140.625 194.185 ;
        RECT 140.875 194.065 141.135 194.235 ;
        RECT 142.195 194.065 142.365 194.560 ;
        RECT 143.675 194.480 143.925 194.810 ;
        RECT 144.915 194.790 145.085 195.005 ;
        RECT 145.255 195.280 145.825 195.385 ;
        RECT 146.495 195.280 147.465 195.385 ;
        RECT 145.255 195.000 147.465 195.280 ;
        RECT 144.095 194.560 145.085 194.790 ;
        RECT 145.255 194.570 145.805 194.740 ;
        RECT 144.915 194.390 145.085 194.560 ;
        RECT 140.805 193.895 141.135 194.065 ;
        RECT 141.395 193.895 142.365 194.065 ;
        RECT 142.535 194.310 143.515 194.390 ;
        RECT 144.115 194.310 144.745 194.390 ;
        RECT 142.535 194.060 144.745 194.310 ;
        RECT 144.915 194.060 145.465 194.390 ;
        RECT 145.635 194.245 145.805 194.570 ;
        RECT 145.985 194.470 146.355 194.810 ;
        RECT 146.535 194.570 147.465 194.750 ;
        RECT 146.535 194.245 146.705 194.570 ;
        RECT 147.635 194.390 147.805 195.555 ;
        RECT 145.635 194.075 146.705 194.245 ;
        RECT 142.195 193.890 142.365 193.895 ;
        RECT 144.915 193.890 145.085 194.060 ;
        RECT 146.060 193.970 146.390 194.075 ;
        RECT 146.875 194.060 147.805 194.390 ;
        RECT 133.310 193.160 134.945 193.300 ;
        RECT 135.115 193.260 135.735 193.430 ;
        RECT 136.755 193.295 138.090 193.450 ;
        RECT 131.315 192.120 131.485 193.160 ;
        RECT 127.025 191.270 127.685 191.555 ;
        RECT 126.265 190.890 126.855 191.140 ;
        RECT 127.025 190.880 127.685 191.095 ;
        RECT 127.355 190.790 127.685 190.880 ;
        RECT 125.875 190.450 127.185 190.700 ;
        RECT 127.855 190.620 128.025 191.830 ;
        RECT 128.595 191.780 129.265 192.120 ;
        RECT 129.435 191.780 130.005 192.120 ;
        RECT 130.240 191.780 131.485 192.120 ;
        RECT 131.705 191.800 131.995 192.990 ;
        RECT 132.165 192.645 132.625 192.970 ;
        RECT 132.795 192.645 133.125 192.990 ;
        RECT 133.295 192.720 133.815 192.975 ;
        RECT 134.035 192.850 134.945 193.160 ;
        RECT 132.165 191.970 132.335 192.645 ;
        RECT 132.505 192.280 133.125 192.475 ;
        RECT 132.165 191.800 132.625 191.970 ;
        RECT 128.595 191.590 128.765 191.780 ;
        RECT 131.315 191.630 131.485 191.780 ;
        RECT 128.595 191.350 129.575 191.590 ;
        RECT 128.595 190.780 128.765 191.350 ;
        RECT 129.755 191.260 130.005 191.610 ;
        RECT 130.175 191.270 131.130 191.600 ;
        RECT 131.315 191.350 132.285 191.630 ;
        RECT 132.455 191.480 132.625 191.800 ;
        RECT 132.795 191.650 133.125 192.280 ;
        RECT 133.295 192.050 133.465 192.720 ;
        RECT 134.035 192.550 134.205 192.850 ;
        RECT 135.115 192.700 135.395 193.090 ;
        RECT 135.565 192.810 135.735 193.260 ;
        RECT 135.905 193.160 138.090 193.295 ;
        RECT 138.750 193.160 139.645 193.450 ;
        RECT 139.925 193.555 142.025 193.725 ;
        RECT 139.925 193.320 140.095 193.555 ;
        RECT 141.695 193.475 142.025 193.555 ;
        RECT 142.195 193.680 143.505 193.890 ;
        RECT 144.095 193.680 145.085 193.890 ;
        RECT 142.195 193.450 142.365 193.680 ;
        RECT 144.915 193.450 145.085 193.680 ;
        RECT 145.255 193.800 145.760 193.880 ;
        RECT 146.560 193.800 147.465 193.890 ;
        RECT 145.255 193.620 147.465 193.800 ;
        RECT 147.635 193.450 147.805 194.060 ;
        RECT 140.805 193.195 141.525 193.385 ;
        RECT 135.905 192.980 136.925 193.160 ;
        RECT 133.635 192.340 134.205 192.550 ;
        RECT 134.375 192.510 134.945 192.680 ;
        RECT 135.565 192.640 136.585 192.810 ;
        RECT 133.635 192.220 134.605 192.340 ;
        RECT 133.295 191.880 133.815 192.050 ;
        RECT 134.035 191.920 134.605 192.220 ;
        RECT 133.295 191.480 133.465 191.880 ;
        RECT 134.035 191.710 134.205 191.920 ;
        RECT 134.775 191.750 134.945 192.510 ;
        RECT 135.115 192.470 135.445 192.515 ;
        RECT 135.115 192.270 136.245 192.470 ;
        RECT 135.115 191.820 136.245 192.070 ;
        RECT 128.935 191.090 129.575 191.180 ;
        RECT 130.175 191.090 130.345 191.270 ;
        RECT 128.935 190.920 130.345 191.090 ;
        RECT 128.935 190.850 129.575 190.920 ;
        RECT 127.355 190.450 128.025 190.620 ;
        RECT 128.195 190.680 128.765 190.780 ;
        RECT 128.195 190.450 129.575 190.680 ;
        RECT 120.435 189.770 121.365 189.940 ;
        RECT 117.715 189.490 118.695 189.760 ;
        RECT 113.895 189.100 114.825 189.280 ;
        RECT 114.995 188.380 115.165 189.460 ;
        RECT 117.715 188.820 117.885 189.490 ;
        RECT 118.875 189.420 119.125 189.770 ;
        RECT 120.435 189.760 120.605 189.770 ;
        RECT 119.295 189.430 120.605 189.760 ;
        RECT 118.055 189.250 118.695 189.320 ;
        RECT 118.055 189.080 119.465 189.250 ;
        RECT 118.055 188.990 118.695 189.080 ;
        RECT 117.715 188.580 118.695 188.820 ;
        RECT 114.995 188.050 115.885 188.380 ;
        RECT 116.185 188.160 116.725 188.390 ;
        RECT 116.525 188.060 116.725 188.160 ;
        RECT 116.895 188.050 117.545 188.390 ;
        RECT 112.275 187.590 112.950 187.925 ;
        RECT 112.275 186.165 112.445 187.590 ;
        RECT 113.125 187.570 113.975 187.870 ;
        RECT 114.145 187.670 114.805 187.840 ;
        RECT 112.640 187.400 113.015 187.420 ;
        RECT 114.145 187.400 114.375 187.670 ;
        RECT 114.995 187.500 115.165 188.050 ;
        RECT 115.410 187.750 116.705 187.870 ;
        RECT 115.410 187.655 116.725 187.750 ;
        RECT 112.640 187.180 114.375 187.400 ;
        RECT 113.165 187.165 114.375 187.180 ;
        RECT 114.545 187.170 115.165 187.500 ;
        RECT 112.630 186.730 112.970 186.900 ;
        RECT 113.165 186.865 113.495 187.165 ;
        RECT 112.775 186.695 112.970 186.730 ;
        RECT 113.665 186.710 114.780 186.995 ;
        RECT 114.995 186.960 115.165 187.170 ;
        RECT 115.335 187.130 116.325 187.460 ;
        RECT 116.525 187.420 116.725 187.655 ;
        RECT 116.895 187.540 117.085 188.050 ;
        RECT 117.715 187.880 117.885 188.580 ;
        RECT 118.875 188.560 119.125 188.910 ;
        RECT 119.295 188.900 119.465 189.080 ;
        RECT 119.295 188.570 120.250 188.900 ;
        RECT 120.435 188.410 120.605 189.430 ;
        RECT 120.955 189.360 121.365 189.535 ;
        RECT 121.610 189.530 121.800 190.110 ;
        RECT 122.175 189.540 122.345 190.250 ;
        RECT 122.620 189.760 123.325 190.270 ;
        RECT 123.495 189.960 124.125 190.240 ;
        RECT 122.175 189.360 122.950 189.540 ;
        RECT 120.955 189.295 122.950 189.360 ;
        RECT 123.155 189.440 123.325 189.760 ;
        RECT 123.955 189.565 124.125 189.960 ;
        RECT 124.295 189.735 124.855 190.430 ;
        RECT 125.025 189.960 125.705 190.240 ;
        RECT 125.025 189.565 125.245 189.960 ;
        RECT 120.955 189.020 122.345 189.295 ;
        RECT 123.155 189.115 123.785 189.440 ;
        RECT 123.955 189.115 125.245 189.565 ;
        RECT 125.875 189.440 126.045 190.450 ;
        RECT 127.355 190.310 127.685 190.450 ;
        RECT 128.595 190.410 129.575 190.450 ;
        RECT 126.255 190.140 127.105 190.280 ;
        RECT 127.870 190.140 128.380 190.280 ;
        RECT 126.255 189.950 128.380 190.140 ;
        RECT 125.415 189.115 126.045 189.440 ;
        RECT 120.775 188.590 121.705 188.760 ;
        RECT 118.250 188.135 120.265 188.390 ;
        RECT 118.250 188.030 118.625 188.135 ;
        RECT 119.280 188.050 120.265 188.135 ;
        RECT 120.435 188.080 121.365 188.410 ;
        RECT 121.535 188.265 121.705 188.590 ;
        RECT 121.885 188.500 122.255 188.830 ;
        RECT 122.435 188.590 122.985 188.760 ;
        RECT 122.435 188.265 122.605 188.590 ;
        RECT 123.155 188.410 123.325 189.115 ;
        RECT 124.235 189.010 124.565 189.115 ;
        RECT 123.495 188.840 124.065 188.945 ;
        RECT 124.735 188.840 125.705 188.945 ;
        RECT 123.495 188.560 125.705 188.840 ;
        RECT 125.875 188.635 126.045 189.115 ;
        RECT 128.595 189.790 128.765 190.410 ;
        RECT 129.755 190.400 130.005 190.750 ;
        RECT 131.315 190.740 131.485 191.350 ;
        RECT 132.455 191.310 133.465 191.480 ;
        RECT 133.635 191.330 134.205 191.710 ;
        RECT 134.375 191.520 134.945 191.750 ;
        RECT 136.415 191.630 136.585 192.640 ;
        RECT 132.795 191.205 133.125 191.310 ;
        RECT 131.655 191.035 132.625 191.140 ;
        RECT 133.360 191.035 133.705 191.140 ;
        RECT 131.655 190.865 133.705 191.035 ;
        RECT 130.175 190.690 131.485 190.740 ;
        RECT 134.035 190.690 134.205 191.330 ;
        RECT 134.375 191.030 134.945 191.350 ;
        RECT 135.115 191.200 135.445 191.605 ;
        RECT 135.615 191.380 136.585 191.630 ;
        RECT 136.755 192.480 136.925 192.980 ;
        RECT 137.095 192.735 139.110 192.990 ;
        RECT 137.095 192.650 138.080 192.735 ;
        RECT 138.735 192.630 139.110 192.735 ;
        RECT 138.235 192.480 138.565 192.565 ;
        RECT 136.755 192.070 137.355 192.480 ;
        RECT 137.525 192.215 138.565 192.480 ;
        RECT 139.475 192.365 139.645 193.160 ;
        RECT 139.925 192.535 140.095 193.150 ;
        RECT 140.265 193.025 140.595 193.170 ;
        RECT 140.265 192.705 141.555 193.025 ;
        RECT 141.725 192.535 141.895 193.250 ;
        RECT 139.925 192.365 141.895 192.535 ;
        RECT 142.195 193.160 143.530 193.450 ;
        RECT 144.190 193.160 145.810 193.450 ;
        RECT 146.470 193.160 147.805 193.450 ;
        RECT 142.195 192.375 142.365 193.160 ;
        RECT 142.535 192.680 144.735 192.990 ;
        RECT 142.535 192.550 143.165 192.680 ;
        RECT 144.175 192.550 144.735 192.680 ;
        RECT 135.615 191.030 135.785 191.380 ;
        RECT 136.755 191.325 136.925 192.070 ;
        RECT 136.755 191.200 137.345 191.325 ;
        RECT 134.375 190.860 135.785 191.030 ;
        RECT 135.955 190.995 137.345 191.200 ;
        RECT 137.525 191.205 137.695 192.215 ;
        RECT 138.735 192.195 139.645 192.365 ;
        RECT 139.475 192.090 139.645 192.195 ;
        RECT 137.865 191.545 138.035 192.000 ;
        RECT 138.235 191.715 138.565 192.045 ;
        RECT 138.735 191.745 139.110 191.915 ;
        RECT 139.475 191.880 140.175 192.090 ;
        RECT 138.735 191.545 138.905 191.745 ;
        RECT 137.865 191.375 138.905 191.545 ;
        RECT 137.525 191.035 139.305 191.205 ;
        RECT 139.475 191.120 139.645 191.880 ;
        RECT 140.555 191.660 140.885 192.365 ;
        RECT 141.090 191.640 141.465 192.195 ;
        RECT 142.195 192.185 143.215 192.375 ;
        RECT 141.695 192.060 143.215 192.185 ;
        RECT 143.385 192.340 144.005 192.510 ;
        RECT 144.915 192.380 145.085 193.160 ;
        RECT 141.695 191.870 142.365 192.060 ;
        RECT 143.385 191.890 143.555 192.340 ;
        RECT 139.860 191.490 140.385 191.620 ;
        RECT 141.090 191.490 142.025 191.640 ;
        RECT 139.860 191.300 142.025 191.490 ;
        RECT 139.860 191.290 140.885 191.300 ;
        RECT 135.955 190.870 136.925 190.995 ;
        RECT 130.175 190.410 132.575 190.690 ;
        RECT 128.935 189.970 129.485 190.140 ;
        RECT 128.595 189.460 129.145 189.790 ;
        RECT 129.315 189.645 129.485 189.970 ;
        RECT 129.665 189.870 130.035 190.210 ;
        RECT 130.215 189.970 131.145 190.150 ;
        RECT 130.215 189.645 130.385 189.970 ;
        RECT 131.315 189.790 132.575 190.410 ;
        RECT 129.315 189.475 130.385 189.645 ;
        RECT 121.535 188.095 122.605 188.265 ;
        RECT 117.255 187.765 117.885 187.880 ;
        RECT 118.795 187.880 119.125 187.965 ;
        RECT 120.435 187.880 120.605 188.080 ;
        RECT 121.850 187.980 122.180 188.095 ;
        RECT 122.775 188.080 123.325 188.410 ;
        RECT 117.255 187.710 118.625 187.765 ;
        RECT 117.715 187.595 118.625 187.710 ;
        RECT 118.795 187.615 119.835 187.880 ;
        RECT 113.665 186.695 113.835 186.710 ;
        RECT 112.775 186.525 113.835 186.695 ;
        RECT 112.275 185.770 112.940 186.165 ;
        RECT 113.305 186.135 113.835 186.525 ;
        RECT 112.275 184.710 112.445 185.770 ;
        RECT 113.305 185.710 113.685 186.135 ;
        RECT 114.005 185.840 114.315 186.535 ;
        RECT 114.995 186.530 115.940 186.960 ;
        RECT 114.525 186.250 115.940 186.530 ;
        RECT 116.110 186.595 116.325 187.130 ;
        RECT 116.495 186.780 116.725 187.250 ;
        RECT 116.895 187.210 117.165 187.540 ;
        RECT 117.280 187.075 117.545 187.080 ;
        RECT 117.275 187.070 117.545 187.075 ;
        RECT 117.265 187.065 117.545 187.070 ;
        RECT 117.260 187.060 117.545 187.065 ;
        RECT 117.250 187.055 117.545 187.060 ;
        RECT 117.245 187.045 117.545 187.055 ;
        RECT 117.235 187.035 117.545 187.045 ;
        RECT 117.225 187.020 117.545 187.035 ;
        RECT 116.895 186.720 117.545 187.020 ;
        RECT 116.895 186.595 117.085 186.720 ;
        RECT 116.110 186.310 117.085 186.595 ;
        RECT 117.715 186.480 117.885 187.595 ;
        RECT 118.250 187.145 118.625 187.315 ;
        RECT 118.455 186.945 118.625 187.145 ;
        RECT 118.795 187.115 119.125 187.445 ;
        RECT 119.325 186.945 119.495 187.400 ;
        RECT 118.455 186.775 119.495 186.945 ;
        RECT 119.665 186.605 119.835 187.615 ;
        RECT 120.005 187.470 120.605 187.880 ;
        RECT 120.775 187.810 121.680 187.910 ;
        RECT 122.480 187.810 122.985 187.900 ;
        RECT 120.775 187.640 122.985 187.810 ;
        RECT 123.155 187.780 123.325 188.080 ;
        RECT 123.505 188.080 125.705 188.390 ;
        RECT 123.505 187.950 124.065 188.080 ;
        RECT 125.075 187.950 125.705 188.080 ;
        RECT 125.875 188.305 127.145 188.635 ;
        RECT 120.435 186.990 120.605 187.470 ;
        RECT 120.775 187.300 122.825 187.470 ;
        RECT 120.775 187.200 121.745 187.300 ;
        RECT 122.480 187.200 122.825 187.300 ;
        RECT 123.155 187.330 124.065 187.780 ;
        RECT 124.235 187.740 124.855 187.910 ;
        RECT 125.875 187.775 126.045 188.305 ;
        RECT 127.395 188.205 127.605 188.850 ;
        RECT 127.775 188.365 128.410 188.695 ;
        RECT 121.915 187.030 122.245 187.130 ;
        RECT 120.435 186.725 121.405 186.990 ;
        RECT 117.255 186.310 117.885 186.480 ;
        RECT 118.055 186.435 119.835 186.605 ;
        RECT 114.525 185.845 115.165 186.250 ;
        RECT 116.770 186.080 117.545 186.140 ;
        RECT 112.615 185.535 113.135 185.600 ;
        RECT 113.940 185.535 114.725 185.665 ;
        RECT 112.615 185.360 114.725 185.535 ;
        RECT 114.995 184.710 115.165 185.845 ;
        RECT 115.335 185.800 117.545 186.080 ;
        RECT 117.715 185.705 117.885 186.310 ;
        RECT 118.055 185.875 118.705 186.205 ;
        RECT 117.715 185.535 118.355 185.705 ;
        RECT 117.715 184.710 117.885 185.535 ;
        RECT 118.535 185.365 118.705 185.875 ;
        RECT 118.875 185.695 119.085 186.265 ;
        RECT 119.255 186.225 119.835 186.435 ;
        RECT 120.015 186.710 121.405 186.725 ;
        RECT 121.575 186.860 122.585 187.030 ;
        RECT 123.155 187.010 123.325 187.330 ;
        RECT 124.235 187.180 124.515 187.570 ;
        RECT 124.685 187.290 124.855 187.740 ;
        RECT 125.025 187.460 126.045 187.775 ;
        RECT 126.215 187.505 127.225 187.830 ;
        RECT 125.875 187.335 126.045 187.460 ;
        RECT 120.015 186.395 120.605 186.710 ;
        RECT 119.255 185.900 120.265 186.225 ;
        RECT 118.070 185.035 118.705 185.365 ;
        RECT 118.875 184.880 119.085 185.525 ;
        RECT 120.435 185.425 120.605 186.395 ;
        RECT 119.335 185.095 120.605 185.425 ;
        RECT 120.435 184.710 120.605 185.095 ;
        RECT 120.825 184.885 121.115 186.540 ;
        RECT 121.575 186.475 121.745 186.860 ;
        RECT 121.285 186.305 121.745 186.475 ;
        RECT 121.285 185.205 121.455 186.305 ;
        RECT 121.915 186.285 122.245 186.690 ;
        RECT 122.415 186.460 122.585 186.860 ;
        RECT 122.755 186.820 123.325 187.010 ;
        RECT 123.495 186.990 124.065 187.160 ;
        RECT 124.685 187.120 125.705 187.290 ;
        RECT 122.755 186.630 123.725 186.820 ;
        RECT 122.415 186.290 122.935 186.460 ;
        RECT 123.155 186.400 123.725 186.630 ;
        RECT 121.625 185.405 122.245 186.115 ;
        RECT 122.415 185.590 122.585 186.290 ;
        RECT 123.155 186.120 123.325 186.400 ;
        RECT 123.895 186.230 124.065 186.990 ;
        RECT 124.235 186.950 124.565 186.995 ;
        RECT 124.235 186.750 125.365 186.950 ;
        RECT 124.235 186.300 125.365 186.550 ;
        RECT 122.755 185.790 123.325 186.120 ;
        RECT 123.495 186.000 124.065 186.230 ;
        RECT 125.535 186.110 125.705 187.120 ;
        RECT 122.415 185.420 122.935 185.590 ;
        RECT 121.285 184.885 121.745 185.205 ;
        RECT 121.915 184.885 122.485 185.235 ;
        RECT 123.155 185.220 123.325 185.790 ;
        RECT 123.495 185.510 124.065 185.830 ;
        RECT 124.235 185.680 124.565 186.085 ;
        RECT 124.735 185.860 125.705 186.110 ;
        RECT 125.875 187.005 126.465 187.335 ;
        RECT 126.645 187.295 127.225 187.505 ;
        RECT 127.395 187.465 127.605 188.035 ;
        RECT 127.775 187.855 127.945 188.365 ;
        RECT 128.595 188.195 128.765 189.460 ;
        RECT 129.740 189.370 130.070 189.475 ;
        RECT 130.555 189.460 132.575 189.790 ;
        RECT 132.745 190.670 134.205 190.690 ;
        RECT 132.745 190.430 135.015 190.670 ;
        RECT 132.745 189.760 134.205 190.430 ;
        RECT 135.195 190.340 135.445 190.690 ;
        RECT 135.615 190.350 136.570 190.680 ;
        RECT 134.375 190.170 135.015 190.260 ;
        RECT 135.615 190.170 135.785 190.350 ;
        RECT 134.375 190.000 135.785 190.170 ;
        RECT 136.755 190.025 136.925 190.870 ;
        RECT 137.525 190.825 138.105 191.035 ;
        RECT 139.475 190.950 140.255 191.120 ;
        RECT 137.095 190.500 138.105 190.825 ;
        RECT 138.275 190.295 138.485 190.865 ;
        RECT 138.655 190.475 139.305 190.805 ;
        RECT 134.375 189.930 135.015 190.000 ;
        RECT 132.745 189.490 135.015 189.760 ;
        RECT 132.745 189.480 134.205 189.490 ;
        RECT 135.195 189.480 135.445 189.830 ;
        RECT 136.755 189.820 138.025 190.025 ;
        RECT 135.615 189.695 138.025 189.820 ;
        RECT 135.615 189.490 136.925 189.695 ;
        RECT 131.315 189.310 132.575 189.460 ;
        RECT 128.935 189.200 129.440 189.280 ;
        RECT 130.240 189.200 131.145 189.290 ;
        RECT 128.935 189.020 131.145 189.200 ;
        RECT 128.950 188.365 129.585 188.695 ;
        RECT 128.125 188.025 129.235 188.195 ;
        RECT 127.775 187.525 128.425 187.855 ;
        RECT 126.645 187.125 128.425 187.295 ;
        RECT 125.875 186.260 126.045 187.005 ;
        RECT 124.735 185.510 124.905 185.860 ;
        RECT 125.875 185.850 126.475 186.260 ;
        RECT 126.645 186.115 126.815 187.125 ;
        RECT 126.985 186.785 128.025 186.955 ;
        RECT 126.985 186.330 127.155 186.785 ;
        RECT 127.355 186.285 127.685 186.615 ;
        RECT 127.855 186.585 128.025 186.785 ;
        RECT 127.855 186.415 128.230 186.585 ;
        RECT 128.595 186.135 128.765 188.025 ;
        RECT 129.415 187.855 129.585 188.365 ;
        RECT 129.755 188.205 129.965 188.850 ;
        RECT 131.315 188.635 133.095 189.310 ;
        RECT 130.215 188.305 133.095 188.635 ;
        RECT 131.315 188.100 133.095 188.305 ;
        RECT 133.265 188.225 134.205 189.480 ;
        RECT 134.570 188.595 136.585 188.850 ;
        RECT 134.570 188.490 134.945 188.595 ;
        RECT 135.600 188.510 136.585 188.595 ;
        RECT 136.755 188.800 136.925 189.490 ;
        RECT 138.275 189.480 138.485 190.125 ;
        RECT 138.655 189.965 138.825 190.475 ;
        RECT 139.475 190.305 139.645 190.950 ;
        RECT 139.865 190.625 140.385 190.780 ;
        RECT 140.555 190.740 140.885 191.290 ;
        RECT 142.195 191.130 142.365 191.870 ;
        RECT 141.185 190.960 142.365 191.130 ;
        RECT 139.865 190.570 140.425 190.625 ;
        RECT 141.055 190.615 141.980 190.790 ;
        RECT 141.005 190.570 141.980 190.615 ;
        RECT 139.865 190.460 141.980 190.570 ;
        RECT 139.865 190.450 141.135 190.460 ;
        RECT 140.300 190.400 141.135 190.450 ;
        RECT 139.005 190.135 139.645 190.305 ;
        RECT 138.655 189.635 139.290 189.965 ;
        RECT 139.475 189.605 139.645 190.135 ;
        RECT 142.195 190.280 142.365 190.960 ;
        RECT 142.535 191.720 143.555 191.890 ;
        RECT 143.725 191.780 144.005 192.170 ;
        RECT 144.175 192.065 145.085 192.380 ;
        RECT 147.635 192.065 147.805 193.160 ;
        RECT 144.175 191.930 145.925 192.065 ;
        RECT 144.915 191.805 145.925 191.930 ;
        RECT 146.485 191.805 147.805 192.065 ;
        RECT 142.535 190.710 142.705 191.720 ;
        RECT 143.675 191.550 144.005 191.595 ;
        RECT 142.875 191.350 144.005 191.550 ;
        RECT 144.175 191.590 144.745 191.760 ;
        RECT 142.875 190.900 144.005 191.150 ;
        RECT 144.175 190.830 144.345 191.590 ;
        RECT 144.915 191.420 145.085 191.805 ;
        RECT 144.515 191.205 145.085 191.420 ;
        RECT 145.255 191.460 147.465 191.630 ;
        RECT 145.255 191.375 145.830 191.460 ;
        RECT 146.560 191.375 147.465 191.460 ;
        RECT 145.995 191.205 146.325 191.290 ;
        RECT 147.635 191.205 147.805 191.805 ;
        RECT 144.515 191.000 145.465 191.205 ;
        RECT 144.915 190.875 145.465 191.000 ;
        RECT 145.635 191.035 146.705 191.205 ;
        RECT 142.535 190.460 143.505 190.710 ;
        RECT 142.195 189.950 143.165 190.280 ;
        RECT 143.335 190.110 143.505 190.460 ;
        RECT 143.675 190.280 144.005 190.685 ;
        RECT 144.175 190.600 144.745 190.830 ;
        RECT 144.175 190.110 144.745 190.430 ;
        RECT 139.475 189.365 140.155 189.605 ;
        RECT 137.095 189.055 139.110 189.310 ;
        RECT 137.095 188.970 138.080 189.055 ;
        RECT 138.735 188.950 139.110 189.055 ;
        RECT 138.235 188.800 138.565 188.885 ;
        RECT 135.115 188.340 135.445 188.425 ;
        RECT 136.755 188.390 137.355 188.800 ;
        RECT 137.525 188.535 138.565 188.800 ;
        RECT 139.475 188.685 139.645 189.365 ;
        RECT 140.325 189.355 140.885 189.710 ;
        RECT 141.055 189.195 141.400 189.585 ;
        RECT 142.195 189.200 142.365 189.950 ;
        RECT 143.335 189.940 144.745 190.110 ;
        RECT 144.915 190.230 145.085 190.875 ;
        RECT 145.635 190.660 145.805 191.035 ;
        RECT 145.255 190.490 145.805 190.660 ;
        RECT 145.985 190.400 146.355 190.755 ;
        RECT 146.535 190.660 146.705 191.035 ;
        RECT 146.875 190.875 147.805 191.205 ;
        RECT 146.535 190.490 147.465 190.660 ;
        RECT 147.635 190.230 147.805 190.875 ;
        RECT 142.535 189.370 143.215 189.655 ;
        RECT 141.055 189.185 141.225 189.195 ;
        RECT 139.825 189.015 141.225 189.185 ;
        RECT 139.825 188.905 140.155 189.015 ;
        RECT 138.735 188.675 139.645 188.685 ;
        RECT 136.755 188.340 136.925 188.390 ;
        RECT 133.265 188.100 134.945 188.225 ;
        RECT 128.935 187.525 129.585 187.855 ;
        RECT 129.755 187.465 129.965 188.035 ;
        RECT 130.135 187.505 131.145 187.830 ;
        RECT 130.135 187.295 130.715 187.505 ;
        RECT 131.315 187.460 131.485 188.100 ;
        RECT 134.035 188.055 134.945 188.100 ;
        RECT 135.115 188.075 136.155 188.340 ;
        RECT 131.315 187.335 132.625 187.460 ;
        RECT 128.935 187.125 130.715 187.295 ;
        RECT 129.335 186.785 130.375 186.955 ;
        RECT 129.335 186.585 129.505 186.785 ;
        RECT 129.130 186.415 129.505 186.585 ;
        RECT 129.675 186.285 130.005 186.615 ;
        RECT 130.205 186.330 130.375 186.785 ;
        RECT 126.645 185.850 127.685 186.115 ;
        RECT 127.855 185.965 129.505 186.135 ;
        RECT 130.545 186.115 130.715 187.125 ;
        RECT 130.895 187.130 132.625 187.335 ;
        RECT 130.895 187.005 131.485 187.130 ;
        RECT 132.795 187.120 133.045 187.470 ;
        RECT 134.035 187.460 134.205 188.055 ;
        RECT 134.570 187.605 134.945 187.775 ;
        RECT 133.225 187.190 134.205 187.460 ;
        RECT 134.775 187.405 134.945 187.605 ;
        RECT 135.115 187.575 135.445 187.905 ;
        RECT 135.645 187.405 135.815 187.860 ;
        RECT 134.775 187.235 135.815 187.405 ;
        RECT 131.315 186.260 131.485 187.005 ;
        RECT 133.225 186.950 133.865 187.020 ;
        RECT 132.455 186.780 133.865 186.950 ;
        RECT 132.455 186.600 132.625 186.780 ;
        RECT 133.225 186.690 133.865 186.780 ;
        RECT 131.670 186.270 132.625 186.600 ;
        RECT 132.795 186.260 133.045 186.610 ;
        RECT 134.035 186.520 134.205 187.190 ;
        RECT 135.985 187.065 136.155 188.075 ;
        RECT 136.325 187.930 136.925 188.340 ;
        RECT 136.755 187.645 136.925 187.930 ;
        RECT 136.755 187.315 137.345 187.645 ;
        RECT 137.525 187.525 137.695 188.535 ;
        RECT 138.735 188.515 140.155 188.675 ;
        RECT 140.325 188.580 140.885 188.845 ;
        RECT 139.475 188.460 140.155 188.515 ;
        RECT 137.865 187.865 138.035 188.320 ;
        RECT 138.235 188.035 138.565 188.365 ;
        RECT 138.735 188.065 139.110 188.235 ;
        RECT 138.735 187.865 138.905 188.065 ;
        RECT 137.865 187.695 138.905 187.865 ;
        RECT 137.525 187.355 139.305 187.525 ;
        RECT 136.755 187.185 136.925 187.315 ;
        RECT 134.375 186.895 136.155 187.065 ;
        RECT 133.225 186.280 134.205 186.520 ;
        RECT 134.375 186.335 135.025 186.665 ;
        RECT 125.875 185.680 126.045 185.850 ;
        RECT 127.355 185.765 127.685 185.850 ;
        RECT 123.495 185.340 124.905 185.510 ;
        RECT 125.075 185.350 126.045 185.680 ;
        RECT 122.655 184.890 123.325 185.220 ;
        RECT 123.155 184.710 123.325 184.890 ;
        RECT 125.875 184.710 126.045 185.350 ;
        RECT 126.215 185.595 127.200 185.680 ;
        RECT 127.855 185.595 128.230 185.700 ;
        RECT 126.215 185.570 128.230 185.595 ;
        RECT 126.215 185.400 128.255 185.570 ;
        RECT 126.215 185.340 128.230 185.400 ;
        RECT 128.595 184.710 128.765 185.965 ;
        RECT 129.675 185.850 130.715 186.115 ;
        RECT 130.885 185.850 131.485 186.260 ;
        RECT 134.035 186.165 134.205 186.280 ;
        RECT 129.675 185.765 130.005 185.850 ;
        RECT 129.130 185.595 129.505 185.700 ;
        RECT 130.160 185.595 131.145 185.680 ;
        RECT 129.130 185.340 131.145 185.595 ;
        RECT 131.315 185.650 131.485 185.850 ;
        RECT 131.655 185.920 133.865 186.090 ;
        RECT 131.655 185.820 132.560 185.920 ;
        RECT 133.360 185.830 133.865 185.920 ;
        RECT 134.035 185.995 134.675 186.165 ;
        RECT 131.315 185.320 132.245 185.650 ;
        RECT 132.730 185.635 133.060 185.750 ;
        RECT 134.035 185.650 134.205 185.995 ;
        RECT 134.855 185.825 135.025 186.335 ;
        RECT 135.195 186.155 135.405 186.725 ;
        RECT 135.575 186.685 136.155 186.895 ;
        RECT 136.335 186.855 136.925 187.185 ;
        RECT 137.525 187.145 138.105 187.355 ;
        RECT 135.575 186.360 136.585 186.685 ;
        RECT 136.755 186.345 136.925 186.855 ;
        RECT 137.095 186.820 138.105 187.145 ;
        RECT 138.275 186.615 138.485 187.185 ;
        RECT 138.655 186.795 139.305 187.125 ;
        RECT 139.475 187.030 139.645 188.460 ;
        RECT 141.055 188.330 141.225 189.015 ;
        RECT 142.195 188.930 142.825 189.200 ;
        RECT 142.195 188.710 142.365 188.930 ;
        RECT 141.395 188.380 142.365 188.710 ;
        RECT 142.995 188.910 143.215 189.370 ;
        RECT 143.385 189.080 143.945 189.770 ;
        RECT 144.915 189.710 146.375 190.230 ;
        RECT 144.115 189.370 144.745 189.655 ;
        RECT 144.115 188.910 144.285 189.370 ;
        RECT 144.915 189.200 145.835 189.710 ;
        RECT 146.545 189.540 147.805 190.230 ;
        RECT 144.455 189.020 145.835 189.200 ;
        RECT 146.005 189.020 147.805 189.540 ;
        RECT 144.455 188.930 145.085 189.020 ;
        RECT 142.995 188.700 144.285 188.910 ;
        RECT 139.815 187.990 140.385 188.290 ;
        RECT 140.555 188.160 141.225 188.330 ;
        RECT 141.405 187.990 142.025 188.210 ;
        RECT 139.815 187.675 142.025 187.990 ;
        RECT 139.815 187.210 140.365 187.380 ;
        RECT 136.755 186.015 138.025 186.345 ;
        RECT 132.415 185.465 133.485 185.635 ;
        RECT 131.315 184.710 131.485 185.320 ;
        RECT 132.415 185.140 132.585 185.465 ;
        RECT 131.655 184.970 132.585 185.140 ;
        RECT 132.765 184.900 133.135 185.230 ;
        RECT 133.315 185.140 133.485 185.465 ;
        RECT 133.655 185.320 134.205 185.650 ;
        RECT 134.390 185.495 135.025 185.825 ;
        RECT 135.195 185.340 135.405 185.985 ;
        RECT 136.755 185.885 136.925 186.015 ;
        RECT 135.655 185.555 136.925 185.885 ;
        RECT 138.275 185.800 138.485 186.445 ;
        RECT 138.655 186.285 138.825 186.795 ;
        RECT 139.475 186.700 140.025 187.030 ;
        RECT 140.195 186.885 140.365 187.210 ;
        RECT 140.545 187.120 140.915 187.450 ;
        RECT 141.095 187.210 142.025 187.380 ;
        RECT 141.095 186.885 141.265 187.210 ;
        RECT 142.195 187.140 142.365 188.380 ;
        RECT 142.535 188.130 144.745 188.530 ;
        RECT 144.915 188.410 145.085 188.930 ;
        RECT 145.255 188.680 147.465 188.850 ;
        RECT 145.255 188.590 145.760 188.680 ;
        RECT 146.560 188.580 147.465 188.680 ;
        RECT 142.535 187.660 143.215 187.940 ;
        RECT 142.995 187.265 143.215 187.660 ;
        RECT 143.385 187.435 143.945 188.130 ;
        RECT 144.915 188.080 145.465 188.410 ;
        RECT 146.060 188.395 146.390 188.510 ;
        RECT 147.635 188.410 147.805 189.020 ;
        RECT 145.635 188.225 146.705 188.395 ;
        RECT 144.115 187.660 144.745 187.940 ;
        RECT 144.115 187.265 144.285 187.660 ;
        RECT 142.195 187.030 142.825 187.140 ;
        RECT 140.195 186.715 141.265 186.885 ;
        RECT 141.435 186.815 142.825 187.030 ;
        RECT 142.995 186.815 144.285 187.265 ;
        RECT 144.915 187.140 145.085 188.080 ;
        RECT 145.635 187.900 145.805 188.225 ;
        RECT 145.255 187.730 145.805 187.900 ;
        RECT 145.985 187.660 146.355 187.990 ;
        RECT 146.535 187.900 146.705 188.225 ;
        RECT 146.875 188.080 147.805 188.410 ;
        RECT 146.535 187.730 147.465 187.900 ;
        RECT 145.255 187.300 147.465 187.470 ;
        RECT 145.255 187.210 145.760 187.300 ;
        RECT 146.560 187.200 147.465 187.300 ;
        RECT 144.455 187.030 145.085 187.140 ;
        RECT 144.455 186.815 145.465 187.030 ;
        RECT 146.060 187.015 146.390 187.130 ;
        RECT 147.635 187.030 147.805 188.080 ;
        RECT 139.475 186.625 139.645 186.700 ;
        RECT 139.005 186.455 139.645 186.625 ;
        RECT 140.620 186.600 140.950 186.715 ;
        RECT 141.435 186.700 142.365 186.815 ;
        RECT 143.675 186.710 144.005 186.815 ;
        RECT 138.655 185.955 139.290 186.285 ;
        RECT 133.315 184.970 133.865 185.140 ;
        RECT 134.035 184.710 134.205 185.320 ;
        RECT 136.755 184.710 136.925 185.555 ;
        RECT 139.475 185.650 139.645 186.455 ;
        RECT 139.815 186.430 140.320 186.520 ;
        RECT 141.120 186.430 142.025 186.530 ;
        RECT 139.815 186.260 142.025 186.430 ;
        RECT 139.815 185.910 142.025 186.090 ;
        RECT 139.815 185.830 140.320 185.910 ;
        RECT 141.120 185.820 142.025 185.910 ;
        RECT 139.475 185.320 140.025 185.650 ;
        RECT 140.620 185.635 140.950 185.740 ;
        RECT 142.195 185.650 142.365 186.700 ;
        RECT 144.915 186.700 145.465 186.815 ;
        RECT 145.635 186.845 146.705 187.015 ;
        RECT 142.535 186.540 143.505 186.645 ;
        RECT 144.175 186.540 144.745 186.645 ;
        RECT 142.535 186.260 144.745 186.540 ;
        RECT 142.535 185.910 144.745 186.090 ;
        RECT 142.535 185.820 143.440 185.910 ;
        RECT 144.240 185.830 144.745 185.910 ;
        RECT 140.195 185.465 141.265 185.635 ;
        RECT 139.475 184.710 139.645 185.320 ;
        RECT 140.195 185.140 140.365 185.465 ;
        RECT 139.815 184.970 140.365 185.140 ;
        RECT 140.545 184.900 140.915 185.240 ;
        RECT 141.095 185.140 141.265 185.465 ;
        RECT 141.435 185.320 143.125 185.650 ;
        RECT 143.610 185.635 143.940 185.740 ;
        RECT 144.915 185.650 145.085 186.700 ;
        RECT 145.635 186.520 145.805 186.845 ;
        RECT 145.255 186.350 145.805 186.520 ;
        RECT 145.985 186.280 146.355 186.610 ;
        RECT 146.535 186.520 146.705 186.845 ;
        RECT 146.875 186.700 147.805 187.030 ;
        RECT 146.535 186.350 147.465 186.520 ;
        RECT 145.255 185.910 147.465 186.090 ;
        RECT 145.255 185.830 145.760 185.910 ;
        RECT 146.560 185.820 147.465 185.910 ;
        RECT 143.295 185.465 144.365 185.635 ;
        RECT 141.095 184.960 142.025 185.140 ;
        RECT 142.195 184.710 142.365 185.320 ;
        RECT 143.295 185.140 143.465 185.465 ;
        RECT 142.535 184.960 143.465 185.140 ;
        RECT 143.645 184.900 144.015 185.240 ;
        RECT 144.195 185.140 144.365 185.465 ;
        RECT 144.535 185.320 145.465 185.650 ;
        RECT 146.060 185.635 146.390 185.740 ;
        RECT 147.635 185.650 147.805 186.700 ;
        RECT 145.635 185.465 146.705 185.635 ;
        RECT 144.195 184.970 144.745 185.140 ;
        RECT 144.915 184.710 145.085 185.320 ;
        RECT 145.635 185.140 145.805 185.465 ;
        RECT 145.255 184.970 145.805 185.140 ;
        RECT 145.985 184.900 146.355 185.240 ;
        RECT 146.535 185.140 146.705 185.465 ;
        RECT 146.875 185.320 147.805 185.650 ;
        RECT 146.535 184.960 147.465 185.140 ;
        RECT 147.635 184.710 147.805 185.320 ;
        RECT 112.275 184.020 113.195 184.710 ;
        RECT 113.365 184.190 116.795 184.710 ;
        RECT 112.275 183.500 113.735 184.020 ;
        RECT 113.905 183.500 116.255 184.190 ;
        RECT 116.965 184.020 118.635 184.710 ;
        RECT 118.805 184.190 122.235 184.710 ;
        RECT 116.425 183.500 119.175 184.020 ;
        RECT 119.345 183.500 121.695 184.190 ;
        RECT 122.405 184.020 124.075 184.710 ;
        RECT 124.245 184.190 127.675 184.710 ;
        RECT 121.865 183.500 124.615 184.020 ;
        RECT 124.785 183.500 127.135 184.190 ;
        RECT 127.845 184.020 129.515 184.710 ;
        RECT 129.685 184.190 133.115 184.710 ;
        RECT 127.305 183.500 130.055 184.020 ;
        RECT 130.225 183.500 132.575 184.190 ;
        RECT 133.285 184.020 134.955 184.710 ;
        RECT 135.125 184.190 138.555 184.710 ;
        RECT 132.745 183.500 135.495 184.020 ;
        RECT 135.665 183.500 138.015 184.190 ;
        RECT 138.725 184.020 140.395 184.710 ;
        RECT 140.565 184.190 143.995 184.710 ;
        RECT 138.185 183.500 140.935 184.020 ;
        RECT 141.105 183.500 143.455 184.190 ;
        RECT 144.165 184.020 145.835 184.710 ;
        RECT 146.005 184.190 147.805 184.710 ;
        RECT 143.625 183.500 146.375 184.020 ;
        RECT 146.545 183.500 147.805 184.190 ;
        RECT 112.275 183.415 112.445 183.500 ;
        RECT 114.995 183.415 115.165 183.500 ;
        RECT 117.715 183.415 117.885 183.500 ;
        RECT 120.435 183.415 120.605 183.500 ;
        RECT 123.155 183.415 123.325 183.500 ;
        RECT 125.875 183.415 126.045 183.500 ;
        RECT 128.595 183.415 128.765 183.500 ;
        RECT 131.315 183.415 131.485 183.500 ;
        RECT 134.035 183.415 134.205 183.500 ;
        RECT 136.755 183.415 136.925 183.500 ;
        RECT 139.475 183.415 139.645 183.500 ;
        RECT 142.195 183.415 142.365 183.500 ;
        RECT 144.915 183.415 145.085 183.500 ;
        RECT 147.635 183.415 147.805 183.500 ;
        RECT 100.630 176.790 106.370 176.800 ;
        RECT 100.140 176.630 106.370 176.790 ;
        RECT 100.140 174.370 100.810 176.630 ;
        RECT 101.480 176.060 105.520 176.230 ;
        RECT 101.140 175.000 101.310 176.000 ;
        RECT 105.690 175.000 105.860 176.000 ;
        RECT 101.480 174.770 105.520 174.940 ;
        RECT 106.200 174.370 106.370 176.630 ;
        RECT 100.140 174.200 106.370 174.370 ;
        RECT 100.140 170.940 100.810 174.200 ;
        RECT 101.480 173.630 105.520 173.800 ;
        RECT 101.140 171.570 101.310 173.570 ;
        RECT 105.690 171.570 105.860 173.570 ;
        RECT 101.480 171.340 105.520 171.510 ;
        RECT 106.200 170.940 106.370 174.200 ;
        RECT 100.140 170.770 106.370 170.940 ;
        RECT 100.140 167.510 100.810 170.770 ;
        RECT 101.480 170.200 105.520 170.370 ;
        RECT 101.140 168.140 101.310 170.140 ;
        RECT 105.690 168.140 105.860 170.140 ;
        RECT 101.480 167.910 105.520 168.080 ;
        RECT 106.200 167.510 106.370 170.770 ;
        RECT 100.140 167.500 106.370 167.510 ;
        RECT 107.960 176.770 117.790 176.810 ;
        RECT 140.540 176.790 146.280 176.800 ;
        RECT 107.960 176.640 118.590 176.770 ;
        RECT 120.510 176.740 126.250 176.750 ;
        RECT 107.960 174.380 108.130 176.640 ;
        RECT 108.855 176.070 116.895 176.240 ;
        RECT 108.470 175.010 108.640 176.010 ;
        RECT 117.110 175.010 117.280 176.010 ;
        RECT 108.855 174.780 116.895 174.950 ;
        RECT 117.620 174.380 118.590 176.640 ;
        RECT 107.960 174.210 118.590 174.380 ;
        RECT 107.960 170.950 108.130 174.210 ;
        RECT 108.855 173.640 116.895 173.810 ;
        RECT 108.470 171.580 108.640 173.580 ;
        RECT 117.110 171.580 117.280 173.580 ;
        RECT 108.855 171.350 116.895 171.520 ;
        RECT 117.620 170.950 118.590 174.210 ;
        RECT 107.960 170.780 118.590 170.950 ;
        RECT 107.960 167.520 108.130 170.780 ;
        RECT 108.855 170.210 116.895 170.380 ;
        RECT 108.470 168.150 108.640 170.150 ;
        RECT 117.110 168.150 117.280 170.150 ;
        RECT 108.855 167.920 116.895 168.090 ;
        RECT 117.620 167.520 118.590 170.780 ;
        RECT 100.140 167.400 106.380 167.500 ;
        RECT 100.130 166.840 106.380 167.400 ;
        RECT 100.130 166.820 105.300 166.840 ;
        RECT 100.130 166.750 104.120 166.820 ;
        RECT 100.130 165.480 102.050 166.750 ;
        RECT 103.560 166.740 104.120 166.750 ;
        RECT 103.790 165.650 104.120 166.740 ;
        RECT 104.490 166.270 105.530 166.440 ;
        RECT 104.490 165.830 105.530 166.000 ;
        RECT 105.700 165.970 105.870 166.300 ;
        RECT 103.950 165.430 104.120 165.650 ;
        RECT 106.210 165.430 106.380 166.840 ;
        RECT 103.950 165.260 106.380 165.430 ;
        RECT 107.960 167.350 118.590 167.520 ;
        RECT 120.020 176.580 126.250 176.740 ;
        RECT 120.020 174.320 120.690 176.580 ;
        RECT 121.360 176.010 125.400 176.180 ;
        RECT 121.020 174.950 121.190 175.950 ;
        RECT 125.570 174.950 125.740 175.950 ;
        RECT 121.360 174.720 125.400 174.890 ;
        RECT 126.080 174.320 126.250 176.580 ;
        RECT 120.020 174.150 126.250 174.320 ;
        RECT 120.020 170.890 120.690 174.150 ;
        RECT 121.360 173.580 125.400 173.750 ;
        RECT 121.020 171.520 121.190 173.520 ;
        RECT 125.570 171.520 125.740 173.520 ;
        RECT 121.360 171.290 125.400 171.460 ;
        RECT 126.080 170.890 126.250 174.150 ;
        RECT 120.020 170.720 126.250 170.890 ;
        RECT 120.020 167.460 120.690 170.720 ;
        RECT 121.360 170.150 125.400 170.320 ;
        RECT 121.020 168.090 121.190 170.090 ;
        RECT 125.570 168.090 125.740 170.090 ;
        RECT 121.360 167.860 125.400 168.030 ;
        RECT 126.080 167.460 126.250 170.720 ;
        RECT 120.020 167.450 126.250 167.460 ;
        RECT 127.840 176.720 137.670 176.760 ;
        RECT 127.840 176.590 138.470 176.720 ;
        RECT 127.840 174.330 128.010 176.590 ;
        RECT 128.735 176.020 136.775 176.190 ;
        RECT 128.350 174.960 128.520 175.960 ;
        RECT 136.990 174.960 137.160 175.960 ;
        RECT 128.735 174.730 136.775 174.900 ;
        RECT 137.500 174.330 138.470 176.590 ;
        RECT 127.840 174.160 138.470 174.330 ;
        RECT 127.840 170.900 128.010 174.160 ;
        RECT 128.735 173.590 136.775 173.760 ;
        RECT 128.350 171.530 128.520 173.530 ;
        RECT 136.990 171.530 137.160 173.530 ;
        RECT 128.735 171.300 136.775 171.470 ;
        RECT 137.500 170.900 138.470 174.160 ;
        RECT 127.840 170.730 138.470 170.900 ;
        RECT 127.840 167.470 128.010 170.730 ;
        RECT 128.735 170.160 136.775 170.330 ;
        RECT 128.350 168.100 128.520 170.100 ;
        RECT 136.990 168.100 137.160 170.100 ;
        RECT 128.735 167.870 136.775 168.040 ;
        RECT 137.500 167.470 138.470 170.730 ;
        RECT 120.020 167.350 126.260 167.450 ;
        RECT 107.960 165.090 108.130 167.350 ;
        RECT 108.855 166.780 116.895 166.950 ;
        RECT 108.470 165.720 108.640 166.720 ;
        RECT 117.110 165.720 117.280 166.720 ;
        RECT 108.855 165.490 116.895 165.660 ;
        RECT 117.620 165.090 118.590 167.350 ;
        RECT 120.010 166.790 126.260 167.350 ;
        RECT 120.010 166.770 125.180 166.790 ;
        RECT 120.010 166.700 124.000 166.770 ;
        RECT 120.010 165.430 121.930 166.700 ;
        RECT 123.440 166.690 124.000 166.700 ;
        RECT 123.670 165.600 124.000 166.690 ;
        RECT 124.370 166.220 125.410 166.390 ;
        RECT 124.370 165.780 125.410 165.950 ;
        RECT 125.580 165.920 125.750 166.250 ;
        RECT 123.830 165.380 124.000 165.600 ;
        RECT 126.090 165.380 126.260 166.790 ;
        RECT 123.830 165.210 126.260 165.380 ;
        RECT 127.840 167.300 138.470 167.470 ;
        RECT 140.050 176.630 146.280 176.790 ;
        RECT 140.050 174.370 140.720 176.630 ;
        RECT 141.390 176.060 145.430 176.230 ;
        RECT 141.050 175.000 141.220 176.000 ;
        RECT 145.600 175.000 145.770 176.000 ;
        RECT 141.390 174.770 145.430 174.940 ;
        RECT 146.110 174.370 146.280 176.630 ;
        RECT 140.050 174.200 146.280 174.370 ;
        RECT 140.050 170.940 140.720 174.200 ;
        RECT 141.390 173.630 145.430 173.800 ;
        RECT 141.050 171.570 141.220 173.570 ;
        RECT 145.600 171.570 145.770 173.570 ;
        RECT 141.390 171.340 145.430 171.510 ;
        RECT 146.110 170.940 146.280 174.200 ;
        RECT 140.050 170.770 146.280 170.940 ;
        RECT 140.050 167.510 140.720 170.770 ;
        RECT 141.390 170.200 145.430 170.370 ;
        RECT 141.050 168.140 141.220 170.140 ;
        RECT 145.600 168.140 145.770 170.140 ;
        RECT 141.390 167.910 145.430 168.080 ;
        RECT 146.110 167.510 146.280 170.770 ;
        RECT 140.050 167.500 146.280 167.510 ;
        RECT 147.870 176.770 157.700 176.810 ;
        RECT 147.870 176.640 158.500 176.770 ;
        RECT 147.870 174.380 148.040 176.640 ;
        RECT 148.765 176.070 156.805 176.240 ;
        RECT 148.380 175.010 148.550 176.010 ;
        RECT 157.020 175.010 157.190 176.010 ;
        RECT 148.765 174.780 156.805 174.950 ;
        RECT 157.530 174.380 158.500 176.640 ;
        RECT 147.870 174.210 158.500 174.380 ;
        RECT 147.870 170.950 148.040 174.210 ;
        RECT 148.765 173.640 156.805 173.810 ;
        RECT 148.380 171.580 148.550 173.580 ;
        RECT 157.020 171.580 157.190 173.580 ;
        RECT 148.765 171.350 156.805 171.520 ;
        RECT 157.530 170.950 158.500 174.210 ;
        RECT 147.870 170.780 158.500 170.950 ;
        RECT 147.870 167.520 148.040 170.780 ;
        RECT 148.765 170.210 156.805 170.380 ;
        RECT 148.380 168.150 148.550 170.150 ;
        RECT 157.020 168.150 157.190 170.150 ;
        RECT 148.765 167.920 156.805 168.090 ;
        RECT 157.530 167.520 158.500 170.780 ;
        RECT 140.050 167.400 146.290 167.500 ;
        RECT 107.960 165.060 118.590 165.090 ;
        RECT 107.930 164.950 118.590 165.060 ;
        RECT 127.840 165.040 128.010 167.300 ;
        RECT 128.735 166.730 136.775 166.900 ;
        RECT 128.350 165.670 128.520 166.670 ;
        RECT 136.990 165.670 137.160 166.670 ;
        RECT 128.735 165.440 136.775 165.610 ;
        RECT 137.500 165.040 138.470 167.300 ;
        RECT 140.040 166.840 146.290 167.400 ;
        RECT 140.040 166.820 145.210 166.840 ;
        RECT 140.040 166.750 144.030 166.820 ;
        RECT 140.040 165.480 141.960 166.750 ;
        RECT 143.470 166.740 144.030 166.750 ;
        RECT 143.700 165.650 144.030 166.740 ;
        RECT 144.400 166.270 145.440 166.440 ;
        RECT 144.400 165.830 145.440 166.000 ;
        RECT 145.610 165.970 145.780 166.300 ;
        RECT 143.860 165.430 144.030 165.650 ;
        RECT 146.120 165.430 146.290 166.840 ;
        RECT 143.860 165.260 146.290 165.430 ;
        RECT 147.870 167.350 158.500 167.520 ;
        RECT 147.870 165.090 148.040 167.350 ;
        RECT 148.765 166.780 156.805 166.950 ;
        RECT 148.380 165.720 148.550 166.720 ;
        RECT 157.020 165.720 157.190 166.720 ;
        RECT 148.765 165.490 156.805 165.660 ;
        RECT 157.530 165.090 158.500 167.350 ;
        RECT 147.870 165.060 158.500 165.090 ;
        RECT 127.840 165.010 138.470 165.040 ;
        RECT 106.180 164.900 118.590 164.950 ;
        RECT 127.810 164.900 138.470 165.010 ;
        RECT 147.840 164.950 158.500 165.060 ;
        RECT 146.090 164.900 158.500 164.950 ;
        RECT 101.840 164.730 118.590 164.900 ;
        RECT 126.060 164.850 138.470 164.900 ;
        RECT 101.840 163.320 102.010 164.730 ;
        RECT 102.380 164.160 105.420 164.330 ;
        RECT 102.380 163.720 105.420 163.890 ;
        RECT 105.635 163.860 105.805 164.190 ;
        RECT 106.140 163.970 118.590 164.730 ;
        RECT 121.720 164.680 138.470 164.850 ;
        RECT 106.140 163.960 118.480 163.970 ;
        RECT 106.140 163.950 112.020 163.960 ;
        RECT 106.140 163.930 106.710 163.950 ;
        RECT 107.930 163.940 112.020 163.950 ;
        RECT 106.150 163.320 106.320 163.930 ;
        RECT 101.840 163.150 106.320 163.320 ;
        RECT 121.720 163.270 121.890 164.680 ;
        RECT 122.260 164.110 125.300 164.280 ;
        RECT 122.260 163.670 125.300 163.840 ;
        RECT 125.515 163.810 125.685 164.140 ;
        RECT 126.020 163.920 138.470 164.680 ;
        RECT 141.750 164.730 158.500 164.900 ;
        RECT 126.020 163.910 138.360 163.920 ;
        RECT 126.020 163.900 131.900 163.910 ;
        RECT 126.020 163.880 126.590 163.900 ;
        RECT 127.810 163.890 131.900 163.900 ;
        RECT 126.030 163.270 126.200 163.880 ;
        RECT 121.720 163.100 126.200 163.270 ;
        RECT 141.750 163.320 141.920 164.730 ;
        RECT 142.290 164.160 145.330 164.330 ;
        RECT 142.290 163.720 145.330 163.890 ;
        RECT 145.545 163.860 145.715 164.190 ;
        RECT 146.050 163.970 158.500 164.730 ;
        RECT 146.050 163.960 158.390 163.970 ;
        RECT 146.050 163.950 151.930 163.960 ;
        RECT 146.050 163.930 146.620 163.950 ;
        RECT 147.840 163.940 151.930 163.950 ;
        RECT 146.060 163.320 146.230 163.930 ;
        RECT 141.750 163.150 146.230 163.320 ;
        RECT 100.630 161.790 106.370 161.800 ;
        RECT 100.140 161.630 106.370 161.790 ;
        RECT 100.140 159.370 100.810 161.630 ;
        RECT 101.480 161.060 105.520 161.230 ;
        RECT 101.140 160.000 101.310 161.000 ;
        RECT 105.690 160.000 105.860 161.000 ;
        RECT 101.480 159.770 105.520 159.940 ;
        RECT 106.200 159.370 106.370 161.630 ;
        RECT 100.140 159.200 106.370 159.370 ;
        RECT 100.140 155.940 100.810 159.200 ;
        RECT 101.480 158.630 105.520 158.800 ;
        RECT 101.140 156.570 101.310 158.570 ;
        RECT 105.690 156.570 105.860 158.570 ;
        RECT 101.480 156.340 105.520 156.510 ;
        RECT 106.200 155.940 106.370 159.200 ;
        RECT 100.140 155.770 106.370 155.940 ;
        RECT 100.140 152.510 100.810 155.770 ;
        RECT 101.480 155.200 105.520 155.370 ;
        RECT 101.140 153.140 101.310 155.140 ;
        RECT 105.690 153.140 105.860 155.140 ;
        RECT 101.480 152.910 105.520 153.080 ;
        RECT 106.200 152.510 106.370 155.770 ;
        RECT 100.140 152.500 106.370 152.510 ;
        RECT 107.960 161.770 117.790 161.810 ;
        RECT 120.510 161.790 126.250 161.800 ;
        RECT 107.960 161.640 118.590 161.770 ;
        RECT 107.960 159.380 108.130 161.640 ;
        RECT 108.855 161.070 116.895 161.240 ;
        RECT 108.470 160.010 108.640 161.010 ;
        RECT 117.110 160.010 117.280 161.010 ;
        RECT 108.855 159.780 116.895 159.950 ;
        RECT 117.620 159.380 118.590 161.640 ;
        RECT 107.960 159.210 118.590 159.380 ;
        RECT 107.960 155.950 108.130 159.210 ;
        RECT 108.855 158.640 116.895 158.810 ;
        RECT 108.470 156.580 108.640 158.580 ;
        RECT 117.110 156.580 117.280 158.580 ;
        RECT 108.855 156.350 116.895 156.520 ;
        RECT 117.620 155.950 118.590 159.210 ;
        RECT 107.960 155.780 118.590 155.950 ;
        RECT 107.960 152.520 108.130 155.780 ;
        RECT 108.855 155.210 116.895 155.380 ;
        RECT 108.470 153.150 108.640 155.150 ;
        RECT 117.110 153.150 117.280 155.150 ;
        RECT 108.855 152.920 116.895 153.090 ;
        RECT 117.620 152.520 118.590 155.780 ;
        RECT 100.140 152.400 106.380 152.500 ;
        RECT 100.130 151.840 106.380 152.400 ;
        RECT 100.130 151.820 105.300 151.840 ;
        RECT 100.130 151.750 104.120 151.820 ;
        RECT 100.130 150.480 102.050 151.750 ;
        RECT 103.560 151.740 104.120 151.750 ;
        RECT 103.790 150.650 104.120 151.740 ;
        RECT 104.490 151.270 105.530 151.440 ;
        RECT 104.490 150.830 105.530 151.000 ;
        RECT 105.700 150.970 105.870 151.300 ;
        RECT 103.950 150.430 104.120 150.650 ;
        RECT 106.210 150.430 106.380 151.840 ;
        RECT 103.950 150.260 106.380 150.430 ;
        RECT 107.960 152.350 118.590 152.520 ;
        RECT 120.020 161.630 126.250 161.790 ;
        RECT 120.020 159.370 120.690 161.630 ;
        RECT 121.360 161.060 125.400 161.230 ;
        RECT 121.020 160.000 121.190 161.000 ;
        RECT 125.570 160.000 125.740 161.000 ;
        RECT 121.360 159.770 125.400 159.940 ;
        RECT 126.080 159.370 126.250 161.630 ;
        RECT 120.020 159.200 126.250 159.370 ;
        RECT 120.020 155.940 120.690 159.200 ;
        RECT 121.360 158.630 125.400 158.800 ;
        RECT 121.020 156.570 121.190 158.570 ;
        RECT 125.570 156.570 125.740 158.570 ;
        RECT 121.360 156.340 125.400 156.510 ;
        RECT 126.080 155.940 126.250 159.200 ;
        RECT 120.020 155.770 126.250 155.940 ;
        RECT 120.020 152.510 120.690 155.770 ;
        RECT 121.360 155.200 125.400 155.370 ;
        RECT 121.020 153.140 121.190 155.140 ;
        RECT 125.570 153.140 125.740 155.140 ;
        RECT 121.360 152.910 125.400 153.080 ;
        RECT 126.080 152.510 126.250 155.770 ;
        RECT 120.020 152.500 126.250 152.510 ;
        RECT 127.840 161.770 137.670 161.810 ;
        RECT 127.840 161.640 138.470 161.770 ;
        RECT 140.590 161.740 146.330 161.750 ;
        RECT 127.840 159.380 128.010 161.640 ;
        RECT 128.735 161.070 136.775 161.240 ;
        RECT 128.350 160.010 128.520 161.010 ;
        RECT 136.990 160.010 137.160 161.010 ;
        RECT 128.735 159.780 136.775 159.950 ;
        RECT 137.500 159.380 138.470 161.640 ;
        RECT 127.840 159.210 138.470 159.380 ;
        RECT 127.840 155.950 128.010 159.210 ;
        RECT 128.735 158.640 136.775 158.810 ;
        RECT 128.350 156.580 128.520 158.580 ;
        RECT 136.990 156.580 137.160 158.580 ;
        RECT 128.735 156.350 136.775 156.520 ;
        RECT 137.500 155.950 138.470 159.210 ;
        RECT 127.840 155.780 138.470 155.950 ;
        RECT 127.840 152.520 128.010 155.780 ;
        RECT 128.735 155.210 136.775 155.380 ;
        RECT 128.350 153.150 128.520 155.150 ;
        RECT 136.990 153.150 137.160 155.150 ;
        RECT 128.735 152.920 136.775 153.090 ;
        RECT 137.500 152.520 138.470 155.780 ;
        RECT 120.020 152.400 126.260 152.500 ;
        RECT 107.960 150.090 108.130 152.350 ;
        RECT 108.855 151.780 116.895 151.950 ;
        RECT 108.470 150.720 108.640 151.720 ;
        RECT 117.110 150.720 117.280 151.720 ;
        RECT 108.855 150.490 116.895 150.660 ;
        RECT 117.620 150.090 118.590 152.350 ;
        RECT 120.010 151.840 126.260 152.400 ;
        RECT 120.010 151.820 125.180 151.840 ;
        RECT 120.010 151.750 124.000 151.820 ;
        RECT 120.010 150.480 121.930 151.750 ;
        RECT 123.440 151.740 124.000 151.750 ;
        RECT 123.670 150.650 124.000 151.740 ;
        RECT 124.370 151.270 125.410 151.440 ;
        RECT 124.370 150.830 125.410 151.000 ;
        RECT 125.580 150.970 125.750 151.300 ;
        RECT 123.830 150.430 124.000 150.650 ;
        RECT 126.090 150.430 126.260 151.840 ;
        RECT 123.830 150.260 126.260 150.430 ;
        RECT 127.840 152.350 138.470 152.520 ;
        RECT 140.100 161.580 146.330 161.740 ;
        RECT 140.100 159.320 140.770 161.580 ;
        RECT 141.440 161.010 145.480 161.180 ;
        RECT 141.100 159.950 141.270 160.950 ;
        RECT 145.650 159.950 145.820 160.950 ;
        RECT 141.440 159.720 145.480 159.890 ;
        RECT 146.160 159.320 146.330 161.580 ;
        RECT 140.100 159.150 146.330 159.320 ;
        RECT 140.100 155.890 140.770 159.150 ;
        RECT 141.440 158.580 145.480 158.750 ;
        RECT 141.100 156.520 141.270 158.520 ;
        RECT 145.650 156.520 145.820 158.520 ;
        RECT 141.440 156.290 145.480 156.460 ;
        RECT 146.160 155.890 146.330 159.150 ;
        RECT 140.100 155.720 146.330 155.890 ;
        RECT 140.100 152.460 140.770 155.720 ;
        RECT 141.440 155.150 145.480 155.320 ;
        RECT 141.100 153.090 141.270 155.090 ;
        RECT 145.650 153.090 145.820 155.090 ;
        RECT 141.440 152.860 145.480 153.030 ;
        RECT 146.160 152.460 146.330 155.720 ;
        RECT 140.100 152.450 146.330 152.460 ;
        RECT 147.920 161.720 157.750 161.760 ;
        RECT 147.920 161.590 158.550 161.720 ;
        RECT 147.920 159.330 148.090 161.590 ;
        RECT 148.815 161.020 156.855 161.190 ;
        RECT 148.430 159.960 148.600 160.960 ;
        RECT 157.070 159.960 157.240 160.960 ;
        RECT 148.815 159.730 156.855 159.900 ;
        RECT 157.580 159.330 158.550 161.590 ;
        RECT 147.920 159.160 158.550 159.330 ;
        RECT 147.920 155.900 148.090 159.160 ;
        RECT 148.815 158.590 156.855 158.760 ;
        RECT 148.430 156.530 148.600 158.530 ;
        RECT 157.070 156.530 157.240 158.530 ;
        RECT 148.815 156.300 156.855 156.470 ;
        RECT 157.580 155.900 158.550 159.160 ;
        RECT 147.920 155.730 158.550 155.900 ;
        RECT 147.920 152.470 148.090 155.730 ;
        RECT 148.815 155.160 156.855 155.330 ;
        RECT 148.430 153.100 148.600 155.100 ;
        RECT 157.070 153.100 157.240 155.100 ;
        RECT 148.815 152.870 156.855 153.040 ;
        RECT 157.580 152.470 158.550 155.730 ;
        RECT 140.100 152.350 146.340 152.450 ;
        RECT 107.960 150.060 118.590 150.090 ;
        RECT 127.840 150.090 128.010 152.350 ;
        RECT 128.735 151.780 136.775 151.950 ;
        RECT 128.350 150.720 128.520 151.720 ;
        RECT 136.990 150.720 137.160 151.720 ;
        RECT 128.735 150.490 136.775 150.660 ;
        RECT 137.500 150.090 138.470 152.350 ;
        RECT 140.090 151.790 146.340 152.350 ;
        RECT 140.090 151.770 145.260 151.790 ;
        RECT 140.090 151.700 144.080 151.770 ;
        RECT 140.090 150.430 142.010 151.700 ;
        RECT 143.520 151.690 144.080 151.700 ;
        RECT 143.750 150.600 144.080 151.690 ;
        RECT 144.450 151.220 145.490 151.390 ;
        RECT 144.450 150.780 145.490 150.950 ;
        RECT 145.660 150.920 145.830 151.250 ;
        RECT 143.910 150.380 144.080 150.600 ;
        RECT 146.170 150.380 146.340 151.790 ;
        RECT 143.910 150.210 146.340 150.380 ;
        RECT 147.920 152.300 158.550 152.470 ;
        RECT 127.840 150.060 138.470 150.090 ;
        RECT 107.930 149.950 118.590 150.060 ;
        RECT 127.810 149.950 138.470 150.060 ;
        RECT 147.920 150.040 148.090 152.300 ;
        RECT 148.815 151.730 156.855 151.900 ;
        RECT 148.430 150.670 148.600 151.670 ;
        RECT 157.070 150.670 157.240 151.670 ;
        RECT 148.815 150.440 156.855 150.610 ;
        RECT 157.580 150.040 158.550 152.300 ;
        RECT 147.920 150.010 158.550 150.040 ;
        RECT 106.180 149.900 118.590 149.950 ;
        RECT 126.060 149.900 138.470 149.950 ;
        RECT 147.890 149.900 158.550 150.010 ;
        RECT 101.840 149.730 118.590 149.900 ;
        RECT 101.840 148.320 102.010 149.730 ;
        RECT 102.380 149.160 105.420 149.330 ;
        RECT 102.380 148.720 105.420 148.890 ;
        RECT 105.635 148.860 105.805 149.190 ;
        RECT 106.140 148.970 118.590 149.730 ;
        RECT 121.720 149.730 138.470 149.900 ;
        RECT 146.140 149.850 158.550 149.900 ;
        RECT 106.140 148.960 118.480 148.970 ;
        RECT 106.140 148.950 112.020 148.960 ;
        RECT 106.140 148.930 106.710 148.950 ;
        RECT 107.930 148.940 112.020 148.950 ;
        RECT 106.150 148.320 106.320 148.930 ;
        RECT 101.840 148.150 106.320 148.320 ;
        RECT 121.720 148.320 121.890 149.730 ;
        RECT 122.260 149.160 125.300 149.330 ;
        RECT 122.260 148.720 125.300 148.890 ;
        RECT 125.515 148.860 125.685 149.190 ;
        RECT 126.020 148.970 138.470 149.730 ;
        RECT 141.800 149.680 158.550 149.850 ;
        RECT 126.020 148.960 138.360 148.970 ;
        RECT 126.020 148.950 131.900 148.960 ;
        RECT 126.020 148.930 126.590 148.950 ;
        RECT 127.810 148.940 131.900 148.950 ;
        RECT 126.030 148.320 126.200 148.930 ;
        RECT 121.720 148.150 126.200 148.320 ;
        RECT 141.800 148.270 141.970 149.680 ;
        RECT 142.340 149.110 145.380 149.280 ;
        RECT 142.340 148.670 145.380 148.840 ;
        RECT 145.595 148.810 145.765 149.140 ;
        RECT 146.100 148.920 158.550 149.680 ;
        RECT 146.100 148.910 158.440 148.920 ;
        RECT 146.100 148.900 151.980 148.910 ;
        RECT 146.100 148.880 146.670 148.900 ;
        RECT 147.890 148.890 151.980 148.900 ;
        RECT 146.110 148.270 146.280 148.880 ;
        RECT 141.800 148.100 146.280 148.270 ;
        RECT 100.630 146.740 106.370 146.750 ;
        RECT 100.140 146.580 106.370 146.740 ;
        RECT 100.140 144.320 100.810 146.580 ;
        RECT 101.480 146.010 105.520 146.180 ;
        RECT 101.140 144.950 101.310 145.950 ;
        RECT 105.690 144.950 105.860 145.950 ;
        RECT 101.480 144.720 105.520 144.890 ;
        RECT 106.200 144.320 106.370 146.580 ;
        RECT 100.140 144.150 106.370 144.320 ;
        RECT 100.140 140.890 100.810 144.150 ;
        RECT 101.480 143.580 105.520 143.750 ;
        RECT 101.140 141.520 101.310 143.520 ;
        RECT 105.690 141.520 105.860 143.520 ;
        RECT 101.480 141.290 105.520 141.460 ;
        RECT 106.200 140.890 106.370 144.150 ;
        RECT 100.140 140.720 106.370 140.890 ;
        RECT 100.140 137.460 100.810 140.720 ;
        RECT 101.480 140.150 105.520 140.320 ;
        RECT 101.140 138.090 101.310 140.090 ;
        RECT 105.690 138.090 105.860 140.090 ;
        RECT 101.480 137.860 105.520 138.030 ;
        RECT 106.200 137.460 106.370 140.720 ;
        RECT 100.140 137.450 106.370 137.460 ;
        RECT 107.960 146.720 117.790 146.760 ;
        RECT 120.510 146.740 126.250 146.750 ;
        RECT 107.960 146.590 118.590 146.720 ;
        RECT 107.960 144.330 108.130 146.590 ;
        RECT 108.855 146.020 116.895 146.190 ;
        RECT 108.470 144.960 108.640 145.960 ;
        RECT 117.110 144.960 117.280 145.960 ;
        RECT 108.855 144.730 116.895 144.900 ;
        RECT 117.620 144.330 118.590 146.590 ;
        RECT 107.960 144.160 118.590 144.330 ;
        RECT 107.960 140.900 108.130 144.160 ;
        RECT 108.855 143.590 116.895 143.760 ;
        RECT 108.470 141.530 108.640 143.530 ;
        RECT 117.110 141.530 117.280 143.530 ;
        RECT 108.855 141.300 116.895 141.470 ;
        RECT 117.620 140.900 118.590 144.160 ;
        RECT 107.960 140.730 118.590 140.900 ;
        RECT 107.960 137.470 108.130 140.730 ;
        RECT 108.855 140.160 116.895 140.330 ;
        RECT 108.470 138.100 108.640 140.100 ;
        RECT 117.110 138.100 117.280 140.100 ;
        RECT 108.855 137.870 116.895 138.040 ;
        RECT 117.620 137.470 118.590 140.730 ;
        RECT 100.140 137.350 106.380 137.450 ;
        RECT 100.130 136.790 106.380 137.350 ;
        RECT 100.130 136.770 105.300 136.790 ;
        RECT 100.130 136.700 104.120 136.770 ;
        RECT 100.130 135.430 102.050 136.700 ;
        RECT 103.560 136.690 104.120 136.700 ;
        RECT 103.790 135.600 104.120 136.690 ;
        RECT 104.490 136.220 105.530 136.390 ;
        RECT 104.490 135.780 105.530 135.950 ;
        RECT 105.700 135.920 105.870 136.250 ;
        RECT 103.950 135.380 104.120 135.600 ;
        RECT 106.210 135.380 106.380 136.790 ;
        RECT 103.950 135.210 106.380 135.380 ;
        RECT 107.960 137.300 118.590 137.470 ;
        RECT 120.020 146.580 126.250 146.740 ;
        RECT 120.020 144.320 120.690 146.580 ;
        RECT 121.360 146.010 125.400 146.180 ;
        RECT 121.020 144.950 121.190 145.950 ;
        RECT 125.570 144.950 125.740 145.950 ;
        RECT 121.360 144.720 125.400 144.890 ;
        RECT 126.080 144.320 126.250 146.580 ;
        RECT 120.020 144.150 126.250 144.320 ;
        RECT 120.020 140.890 120.690 144.150 ;
        RECT 121.360 143.580 125.400 143.750 ;
        RECT 121.020 141.520 121.190 143.520 ;
        RECT 125.570 141.520 125.740 143.520 ;
        RECT 121.360 141.290 125.400 141.460 ;
        RECT 126.080 140.890 126.250 144.150 ;
        RECT 120.020 140.720 126.250 140.890 ;
        RECT 120.020 137.460 120.690 140.720 ;
        RECT 121.360 140.150 125.400 140.320 ;
        RECT 121.020 138.090 121.190 140.090 ;
        RECT 125.570 138.090 125.740 140.090 ;
        RECT 121.360 137.860 125.400 138.030 ;
        RECT 126.080 137.460 126.250 140.720 ;
        RECT 120.020 137.450 126.250 137.460 ;
        RECT 127.840 146.720 137.670 146.760 ;
        RECT 140.540 146.740 146.280 146.750 ;
        RECT 127.840 146.590 138.470 146.720 ;
        RECT 127.840 144.330 128.010 146.590 ;
        RECT 128.735 146.020 136.775 146.190 ;
        RECT 128.350 144.960 128.520 145.960 ;
        RECT 136.990 144.960 137.160 145.960 ;
        RECT 128.735 144.730 136.775 144.900 ;
        RECT 137.500 144.330 138.470 146.590 ;
        RECT 127.840 144.160 138.470 144.330 ;
        RECT 127.840 140.900 128.010 144.160 ;
        RECT 128.735 143.590 136.775 143.760 ;
        RECT 128.350 141.530 128.520 143.530 ;
        RECT 136.990 141.530 137.160 143.530 ;
        RECT 128.735 141.300 136.775 141.470 ;
        RECT 137.500 140.900 138.470 144.160 ;
        RECT 127.840 140.730 138.470 140.900 ;
        RECT 127.840 137.470 128.010 140.730 ;
        RECT 128.735 140.160 136.775 140.330 ;
        RECT 128.350 138.100 128.520 140.100 ;
        RECT 136.990 138.100 137.160 140.100 ;
        RECT 128.735 137.870 136.775 138.040 ;
        RECT 137.500 137.470 138.470 140.730 ;
        RECT 120.020 137.350 126.260 137.450 ;
        RECT 107.960 135.040 108.130 137.300 ;
        RECT 108.855 136.730 116.895 136.900 ;
        RECT 108.470 135.670 108.640 136.670 ;
        RECT 117.110 135.670 117.280 136.670 ;
        RECT 108.855 135.440 116.895 135.610 ;
        RECT 117.620 135.040 118.590 137.300 ;
        RECT 120.010 136.790 126.260 137.350 ;
        RECT 120.010 136.770 125.180 136.790 ;
        RECT 120.010 136.700 124.000 136.770 ;
        RECT 120.010 135.430 121.930 136.700 ;
        RECT 123.440 136.690 124.000 136.700 ;
        RECT 123.670 135.600 124.000 136.690 ;
        RECT 124.370 136.220 125.410 136.390 ;
        RECT 124.370 135.780 125.410 135.950 ;
        RECT 125.580 135.920 125.750 136.250 ;
        RECT 123.830 135.380 124.000 135.600 ;
        RECT 126.090 135.380 126.260 136.790 ;
        RECT 123.830 135.210 126.260 135.380 ;
        RECT 127.840 137.300 138.470 137.470 ;
        RECT 140.050 146.580 146.280 146.740 ;
        RECT 140.050 144.320 140.720 146.580 ;
        RECT 141.390 146.010 145.430 146.180 ;
        RECT 141.050 144.950 141.220 145.950 ;
        RECT 145.600 144.950 145.770 145.950 ;
        RECT 141.390 144.720 145.430 144.890 ;
        RECT 146.110 144.320 146.280 146.580 ;
        RECT 140.050 144.150 146.280 144.320 ;
        RECT 140.050 140.890 140.720 144.150 ;
        RECT 141.390 143.580 145.430 143.750 ;
        RECT 141.050 141.520 141.220 143.520 ;
        RECT 145.600 141.520 145.770 143.520 ;
        RECT 141.390 141.290 145.430 141.460 ;
        RECT 146.110 140.890 146.280 144.150 ;
        RECT 140.050 140.720 146.280 140.890 ;
        RECT 140.050 137.460 140.720 140.720 ;
        RECT 141.390 140.150 145.430 140.320 ;
        RECT 141.050 138.090 141.220 140.090 ;
        RECT 145.600 138.090 145.770 140.090 ;
        RECT 141.390 137.860 145.430 138.030 ;
        RECT 146.110 137.460 146.280 140.720 ;
        RECT 140.050 137.450 146.280 137.460 ;
        RECT 147.870 146.720 157.700 146.760 ;
        RECT 147.870 146.590 158.500 146.720 ;
        RECT 147.870 144.330 148.040 146.590 ;
        RECT 148.765 146.020 156.805 146.190 ;
        RECT 148.380 144.960 148.550 145.960 ;
        RECT 157.020 144.960 157.190 145.960 ;
        RECT 148.765 144.730 156.805 144.900 ;
        RECT 157.530 144.330 158.500 146.590 ;
        RECT 147.870 144.160 158.500 144.330 ;
        RECT 147.870 140.900 148.040 144.160 ;
        RECT 148.765 143.590 156.805 143.760 ;
        RECT 148.380 141.530 148.550 143.530 ;
        RECT 157.020 141.530 157.190 143.530 ;
        RECT 148.765 141.300 156.805 141.470 ;
        RECT 157.530 140.900 158.500 144.160 ;
        RECT 147.870 140.730 158.500 140.900 ;
        RECT 147.870 137.470 148.040 140.730 ;
        RECT 148.765 140.160 156.805 140.330 ;
        RECT 148.380 138.100 148.550 140.100 ;
        RECT 157.020 138.100 157.190 140.100 ;
        RECT 148.765 137.870 156.805 138.040 ;
        RECT 157.530 137.470 158.500 140.730 ;
        RECT 140.050 137.350 146.290 137.450 ;
        RECT 107.960 135.010 118.590 135.040 ;
        RECT 127.840 135.040 128.010 137.300 ;
        RECT 128.735 136.730 136.775 136.900 ;
        RECT 128.350 135.670 128.520 136.670 ;
        RECT 136.990 135.670 137.160 136.670 ;
        RECT 128.735 135.440 136.775 135.610 ;
        RECT 137.500 135.040 138.470 137.300 ;
        RECT 140.040 136.790 146.290 137.350 ;
        RECT 140.040 136.770 145.210 136.790 ;
        RECT 140.040 136.700 144.030 136.770 ;
        RECT 140.040 135.430 141.960 136.700 ;
        RECT 143.470 136.690 144.030 136.700 ;
        RECT 143.700 135.600 144.030 136.690 ;
        RECT 144.400 136.220 145.440 136.390 ;
        RECT 144.400 135.780 145.440 135.950 ;
        RECT 145.610 135.920 145.780 136.250 ;
        RECT 143.860 135.380 144.030 135.600 ;
        RECT 146.120 135.380 146.290 136.790 ;
        RECT 143.860 135.210 146.290 135.380 ;
        RECT 147.870 137.300 158.500 137.470 ;
        RECT 127.840 135.010 138.470 135.040 ;
        RECT 147.870 135.040 148.040 137.300 ;
        RECT 148.765 136.730 156.805 136.900 ;
        RECT 148.380 135.670 148.550 136.670 ;
        RECT 157.020 135.670 157.190 136.670 ;
        RECT 148.765 135.440 156.805 135.610 ;
        RECT 157.530 135.040 158.500 137.300 ;
        RECT 147.870 135.010 158.500 135.040 ;
        RECT 107.930 134.900 118.590 135.010 ;
        RECT 127.810 134.900 138.470 135.010 ;
        RECT 147.840 134.900 158.500 135.010 ;
        RECT 106.180 134.850 118.590 134.900 ;
        RECT 126.060 134.850 138.470 134.900 ;
        RECT 146.090 134.850 158.500 134.900 ;
        RECT 101.840 134.680 118.590 134.850 ;
        RECT 101.840 133.270 102.010 134.680 ;
        RECT 102.380 134.110 105.420 134.280 ;
        RECT 102.380 133.670 105.420 133.840 ;
        RECT 105.635 133.810 105.805 134.140 ;
        RECT 106.140 133.920 118.590 134.680 ;
        RECT 121.720 134.680 138.470 134.850 ;
        RECT 106.140 133.910 118.480 133.920 ;
        RECT 106.140 133.900 112.020 133.910 ;
        RECT 106.140 133.880 106.710 133.900 ;
        RECT 107.930 133.890 112.020 133.900 ;
        RECT 106.150 133.270 106.320 133.880 ;
        RECT 101.840 133.100 106.320 133.270 ;
        RECT 121.720 133.270 121.890 134.680 ;
        RECT 122.260 134.110 125.300 134.280 ;
        RECT 122.260 133.670 125.300 133.840 ;
        RECT 125.515 133.810 125.685 134.140 ;
        RECT 126.020 133.920 138.470 134.680 ;
        RECT 141.750 134.680 158.500 134.850 ;
        RECT 126.020 133.910 138.360 133.920 ;
        RECT 126.020 133.900 131.900 133.910 ;
        RECT 126.020 133.880 126.590 133.900 ;
        RECT 127.810 133.890 131.900 133.900 ;
        RECT 126.030 133.270 126.200 133.880 ;
        RECT 121.720 133.100 126.200 133.270 ;
        RECT 141.750 133.270 141.920 134.680 ;
        RECT 142.290 134.110 145.330 134.280 ;
        RECT 142.290 133.670 145.330 133.840 ;
        RECT 145.545 133.810 145.715 134.140 ;
        RECT 146.050 133.920 158.500 134.680 ;
        RECT 146.050 133.910 158.390 133.920 ;
        RECT 146.050 133.900 151.930 133.910 ;
        RECT 146.050 133.880 146.620 133.900 ;
        RECT 147.840 133.890 151.930 133.900 ;
        RECT 146.060 133.270 146.230 133.880 ;
        RECT 141.750 133.100 146.230 133.270 ;
        RECT 120.510 131.800 126.250 131.810 ;
        RECT 100.630 131.740 106.370 131.750 ;
        RECT 100.140 131.580 106.370 131.740 ;
        RECT 100.140 129.320 100.810 131.580 ;
        RECT 101.480 131.010 105.520 131.180 ;
        RECT 101.140 129.950 101.310 130.950 ;
        RECT 105.690 129.950 105.860 130.950 ;
        RECT 101.480 129.720 105.520 129.890 ;
        RECT 106.200 129.320 106.370 131.580 ;
        RECT 100.140 129.150 106.370 129.320 ;
        RECT 100.140 125.890 100.810 129.150 ;
        RECT 101.480 128.580 105.520 128.750 ;
        RECT 101.140 126.520 101.310 128.520 ;
        RECT 105.690 126.520 105.860 128.520 ;
        RECT 101.480 126.290 105.520 126.460 ;
        RECT 106.200 125.890 106.370 129.150 ;
        RECT 100.140 125.720 106.370 125.890 ;
        RECT 100.140 122.460 100.810 125.720 ;
        RECT 101.480 125.150 105.520 125.320 ;
        RECT 101.140 123.090 101.310 125.090 ;
        RECT 105.690 123.090 105.860 125.090 ;
        RECT 101.480 122.860 105.520 123.030 ;
        RECT 106.200 122.460 106.370 125.720 ;
        RECT 100.140 122.450 106.370 122.460 ;
        RECT 107.960 131.720 117.790 131.760 ;
        RECT 107.960 131.590 118.590 131.720 ;
        RECT 107.960 129.330 108.130 131.590 ;
        RECT 108.855 131.020 116.895 131.190 ;
        RECT 108.470 129.960 108.640 130.960 ;
        RECT 117.110 129.960 117.280 130.960 ;
        RECT 108.855 129.730 116.895 129.900 ;
        RECT 117.620 129.330 118.590 131.590 ;
        RECT 107.960 129.160 118.590 129.330 ;
        RECT 107.960 125.900 108.130 129.160 ;
        RECT 108.855 128.590 116.895 128.760 ;
        RECT 108.470 126.530 108.640 128.530 ;
        RECT 117.110 126.530 117.280 128.530 ;
        RECT 108.855 126.300 116.895 126.470 ;
        RECT 117.620 125.900 118.590 129.160 ;
        RECT 107.960 125.730 118.590 125.900 ;
        RECT 107.960 122.470 108.130 125.730 ;
        RECT 108.855 125.160 116.895 125.330 ;
        RECT 108.470 123.100 108.640 125.100 ;
        RECT 117.110 123.100 117.280 125.100 ;
        RECT 108.855 122.870 116.895 123.040 ;
        RECT 117.620 122.470 118.590 125.730 ;
        RECT 100.140 122.350 106.380 122.450 ;
        RECT 100.130 121.790 106.380 122.350 ;
        RECT 100.130 121.770 105.300 121.790 ;
        RECT 100.130 121.700 104.120 121.770 ;
        RECT 100.130 120.430 102.050 121.700 ;
        RECT 103.560 121.690 104.120 121.700 ;
        RECT 103.790 120.600 104.120 121.690 ;
        RECT 104.490 121.220 105.530 121.390 ;
        RECT 104.490 120.780 105.530 120.950 ;
        RECT 105.700 120.920 105.870 121.250 ;
        RECT 103.950 120.380 104.120 120.600 ;
        RECT 106.210 120.380 106.380 121.790 ;
        RECT 103.950 120.210 106.380 120.380 ;
        RECT 107.960 122.300 118.590 122.470 ;
        RECT 120.020 131.640 126.250 131.800 ;
        RECT 120.020 129.380 120.690 131.640 ;
        RECT 121.360 131.070 125.400 131.240 ;
        RECT 121.020 130.010 121.190 131.010 ;
        RECT 125.570 130.010 125.740 131.010 ;
        RECT 121.360 129.780 125.400 129.950 ;
        RECT 126.080 129.380 126.250 131.640 ;
        RECT 120.020 129.210 126.250 129.380 ;
        RECT 120.020 125.950 120.690 129.210 ;
        RECT 121.360 128.640 125.400 128.810 ;
        RECT 121.020 126.580 121.190 128.580 ;
        RECT 125.570 126.580 125.740 128.580 ;
        RECT 121.360 126.350 125.400 126.520 ;
        RECT 126.080 125.950 126.250 129.210 ;
        RECT 120.020 125.780 126.250 125.950 ;
        RECT 120.020 122.520 120.690 125.780 ;
        RECT 121.360 125.210 125.400 125.380 ;
        RECT 121.020 123.150 121.190 125.150 ;
        RECT 125.570 123.150 125.740 125.150 ;
        RECT 121.360 122.920 125.400 123.090 ;
        RECT 126.080 122.520 126.250 125.780 ;
        RECT 120.020 122.510 126.250 122.520 ;
        RECT 127.840 131.780 137.670 131.820 ;
        RECT 140.540 131.800 146.280 131.810 ;
        RECT 127.840 131.650 138.470 131.780 ;
        RECT 127.840 129.390 128.010 131.650 ;
        RECT 128.735 131.080 136.775 131.250 ;
        RECT 128.350 130.020 128.520 131.020 ;
        RECT 136.990 130.020 137.160 131.020 ;
        RECT 128.735 129.790 136.775 129.960 ;
        RECT 137.500 129.390 138.470 131.650 ;
        RECT 127.840 129.220 138.470 129.390 ;
        RECT 127.840 125.960 128.010 129.220 ;
        RECT 128.735 128.650 136.775 128.820 ;
        RECT 128.350 126.590 128.520 128.590 ;
        RECT 136.990 126.590 137.160 128.590 ;
        RECT 128.735 126.360 136.775 126.530 ;
        RECT 137.500 125.960 138.470 129.220 ;
        RECT 127.840 125.790 138.470 125.960 ;
        RECT 127.840 122.530 128.010 125.790 ;
        RECT 128.735 125.220 136.775 125.390 ;
        RECT 128.350 123.160 128.520 125.160 ;
        RECT 136.990 123.160 137.160 125.160 ;
        RECT 128.735 122.930 136.775 123.100 ;
        RECT 137.500 122.530 138.470 125.790 ;
        RECT 120.020 122.410 126.260 122.510 ;
        RECT 107.960 120.040 108.130 122.300 ;
        RECT 108.855 121.730 116.895 121.900 ;
        RECT 108.470 120.670 108.640 121.670 ;
        RECT 117.110 120.670 117.280 121.670 ;
        RECT 108.855 120.440 116.895 120.610 ;
        RECT 117.620 120.040 118.590 122.300 ;
        RECT 120.010 121.850 126.260 122.410 ;
        RECT 120.010 121.830 125.180 121.850 ;
        RECT 120.010 121.760 124.000 121.830 ;
        RECT 120.010 120.490 121.930 121.760 ;
        RECT 123.440 121.750 124.000 121.760 ;
        RECT 123.670 120.660 124.000 121.750 ;
        RECT 124.370 121.280 125.410 121.450 ;
        RECT 124.370 120.840 125.410 121.010 ;
        RECT 125.580 120.980 125.750 121.310 ;
        RECT 123.830 120.440 124.000 120.660 ;
        RECT 126.090 120.440 126.260 121.850 ;
        RECT 123.830 120.270 126.260 120.440 ;
        RECT 127.840 122.360 138.470 122.530 ;
        RECT 140.050 131.640 146.280 131.800 ;
        RECT 140.050 129.380 140.720 131.640 ;
        RECT 141.390 131.070 145.430 131.240 ;
        RECT 141.050 130.010 141.220 131.010 ;
        RECT 145.600 130.010 145.770 131.010 ;
        RECT 141.390 129.780 145.430 129.950 ;
        RECT 146.110 129.380 146.280 131.640 ;
        RECT 140.050 129.210 146.280 129.380 ;
        RECT 140.050 125.950 140.720 129.210 ;
        RECT 141.390 128.640 145.430 128.810 ;
        RECT 141.050 126.580 141.220 128.580 ;
        RECT 145.600 126.580 145.770 128.580 ;
        RECT 141.390 126.350 145.430 126.520 ;
        RECT 146.110 125.950 146.280 129.210 ;
        RECT 140.050 125.780 146.280 125.950 ;
        RECT 140.050 122.520 140.720 125.780 ;
        RECT 141.390 125.210 145.430 125.380 ;
        RECT 141.050 123.150 141.220 125.150 ;
        RECT 145.600 123.150 145.770 125.150 ;
        RECT 141.390 122.920 145.430 123.090 ;
        RECT 146.110 122.520 146.280 125.780 ;
        RECT 140.050 122.510 146.280 122.520 ;
        RECT 147.870 131.780 157.700 131.820 ;
        RECT 147.870 131.650 158.500 131.780 ;
        RECT 147.870 129.390 148.040 131.650 ;
        RECT 148.765 131.080 156.805 131.250 ;
        RECT 148.380 130.020 148.550 131.020 ;
        RECT 157.020 130.020 157.190 131.020 ;
        RECT 148.765 129.790 156.805 129.960 ;
        RECT 157.530 129.390 158.500 131.650 ;
        RECT 147.870 129.220 158.500 129.390 ;
        RECT 147.870 125.960 148.040 129.220 ;
        RECT 148.765 128.650 156.805 128.820 ;
        RECT 148.380 126.590 148.550 128.590 ;
        RECT 157.020 126.590 157.190 128.590 ;
        RECT 148.765 126.360 156.805 126.530 ;
        RECT 157.530 125.960 158.500 129.220 ;
        RECT 147.870 125.790 158.500 125.960 ;
        RECT 147.870 122.530 148.040 125.790 ;
        RECT 148.765 125.220 156.805 125.390 ;
        RECT 148.380 123.160 148.550 125.160 ;
        RECT 157.020 123.160 157.190 125.160 ;
        RECT 148.765 122.930 156.805 123.100 ;
        RECT 157.530 122.530 158.500 125.790 ;
        RECT 140.050 122.410 146.290 122.510 ;
        RECT 127.840 120.100 128.010 122.360 ;
        RECT 128.735 121.790 136.775 121.960 ;
        RECT 128.350 120.730 128.520 121.730 ;
        RECT 136.990 120.730 137.160 121.730 ;
        RECT 128.735 120.500 136.775 120.670 ;
        RECT 137.500 120.100 138.470 122.360 ;
        RECT 140.040 121.850 146.290 122.410 ;
        RECT 140.040 121.830 145.210 121.850 ;
        RECT 140.040 121.760 144.030 121.830 ;
        RECT 140.040 120.490 141.960 121.760 ;
        RECT 143.470 121.750 144.030 121.760 ;
        RECT 143.700 120.660 144.030 121.750 ;
        RECT 144.400 121.280 145.440 121.450 ;
        RECT 144.400 120.840 145.440 121.010 ;
        RECT 145.610 120.980 145.780 121.310 ;
        RECT 143.860 120.440 144.030 120.660 ;
        RECT 146.120 120.440 146.290 121.850 ;
        RECT 143.860 120.270 146.290 120.440 ;
        RECT 147.870 122.360 158.500 122.530 ;
        RECT 127.840 120.070 138.470 120.100 ;
        RECT 147.870 120.100 148.040 122.360 ;
        RECT 148.765 121.790 156.805 121.960 ;
        RECT 148.380 120.730 148.550 121.730 ;
        RECT 157.020 120.730 157.190 121.730 ;
        RECT 148.765 120.500 156.805 120.670 ;
        RECT 157.530 120.100 158.500 122.360 ;
        RECT 147.870 120.070 158.500 120.100 ;
        RECT 107.960 120.010 118.590 120.040 ;
        RECT 107.930 119.900 118.590 120.010 ;
        RECT 127.810 119.960 138.470 120.070 ;
        RECT 147.840 119.960 158.500 120.070 ;
        RECT 126.060 119.910 138.470 119.960 ;
        RECT 146.090 119.910 158.500 119.960 ;
        RECT 106.180 119.850 118.590 119.900 ;
        RECT 101.840 119.680 118.590 119.850 ;
        RECT 101.840 118.270 102.010 119.680 ;
        RECT 102.380 119.110 105.420 119.280 ;
        RECT 102.380 118.670 105.420 118.840 ;
        RECT 105.635 118.810 105.805 119.140 ;
        RECT 106.140 118.920 118.590 119.680 ;
        RECT 121.720 119.740 138.470 119.910 ;
        RECT 106.140 118.910 118.480 118.920 ;
        RECT 106.140 118.900 112.020 118.910 ;
        RECT 106.140 118.880 106.710 118.900 ;
        RECT 107.930 118.890 112.020 118.900 ;
        RECT 106.150 118.270 106.320 118.880 ;
        RECT 101.840 118.100 106.320 118.270 ;
        RECT 121.720 118.330 121.890 119.740 ;
        RECT 122.260 119.170 125.300 119.340 ;
        RECT 122.260 118.730 125.300 118.900 ;
        RECT 125.515 118.870 125.685 119.200 ;
        RECT 126.020 118.980 138.470 119.740 ;
        RECT 141.750 119.740 158.500 119.910 ;
        RECT 126.020 118.970 138.360 118.980 ;
        RECT 126.020 118.960 131.900 118.970 ;
        RECT 126.020 118.940 126.590 118.960 ;
        RECT 127.810 118.950 131.900 118.960 ;
        RECT 126.030 118.330 126.200 118.940 ;
        RECT 121.720 118.160 126.200 118.330 ;
        RECT 141.750 118.330 141.920 119.740 ;
        RECT 142.290 119.170 145.330 119.340 ;
        RECT 142.290 118.730 145.330 118.900 ;
        RECT 145.545 118.870 145.715 119.200 ;
        RECT 146.050 118.980 158.500 119.740 ;
        RECT 146.050 118.970 158.390 118.980 ;
        RECT 146.050 118.960 151.930 118.970 ;
        RECT 146.050 118.940 146.620 118.960 ;
        RECT 147.840 118.950 151.930 118.960 ;
        RECT 146.060 118.330 146.230 118.940 ;
        RECT 141.750 118.160 146.230 118.330 ;
        RECT 100.580 116.800 106.320 116.810 ;
        RECT 100.090 116.640 106.320 116.800 ;
        RECT 100.090 114.380 100.760 116.640 ;
        RECT 101.430 116.070 105.470 116.240 ;
        RECT 101.090 115.010 101.260 116.010 ;
        RECT 105.640 115.010 105.810 116.010 ;
        RECT 101.430 114.780 105.470 114.950 ;
        RECT 106.150 114.380 106.320 116.640 ;
        RECT 100.090 114.210 106.320 114.380 ;
        RECT 100.090 110.950 100.760 114.210 ;
        RECT 101.430 113.640 105.470 113.810 ;
        RECT 101.090 111.580 101.260 113.580 ;
        RECT 105.640 111.580 105.810 113.580 ;
        RECT 101.430 111.350 105.470 111.520 ;
        RECT 106.150 110.950 106.320 114.210 ;
        RECT 100.090 110.780 106.320 110.950 ;
        RECT 100.090 107.520 100.760 110.780 ;
        RECT 101.430 110.210 105.470 110.380 ;
        RECT 101.090 108.150 101.260 110.150 ;
        RECT 105.640 108.150 105.810 110.150 ;
        RECT 101.430 107.920 105.470 108.090 ;
        RECT 106.150 107.520 106.320 110.780 ;
        RECT 100.090 107.510 106.320 107.520 ;
        RECT 107.910 116.780 117.740 116.820 ;
        RECT 120.510 116.800 126.250 116.810 ;
        RECT 107.910 116.650 118.540 116.780 ;
        RECT 107.910 114.390 108.080 116.650 ;
        RECT 108.805 116.080 116.845 116.250 ;
        RECT 108.420 115.020 108.590 116.020 ;
        RECT 117.060 115.020 117.230 116.020 ;
        RECT 108.805 114.790 116.845 114.960 ;
        RECT 117.570 114.390 118.540 116.650 ;
        RECT 107.910 114.220 118.540 114.390 ;
        RECT 107.910 110.960 108.080 114.220 ;
        RECT 108.805 113.650 116.845 113.820 ;
        RECT 108.420 111.590 108.590 113.590 ;
        RECT 117.060 111.590 117.230 113.590 ;
        RECT 108.805 111.360 116.845 111.530 ;
        RECT 117.570 110.960 118.540 114.220 ;
        RECT 107.910 110.790 118.540 110.960 ;
        RECT 107.910 107.530 108.080 110.790 ;
        RECT 108.805 110.220 116.845 110.390 ;
        RECT 108.420 108.160 108.590 110.160 ;
        RECT 117.060 108.160 117.230 110.160 ;
        RECT 108.805 107.930 116.845 108.100 ;
        RECT 117.570 107.530 118.540 110.790 ;
        RECT 100.090 107.410 106.330 107.510 ;
        RECT 100.080 106.850 106.330 107.410 ;
        RECT 100.080 106.830 105.250 106.850 ;
        RECT 100.080 106.760 104.070 106.830 ;
        RECT 100.080 105.490 102.000 106.760 ;
        RECT 103.510 106.750 104.070 106.760 ;
        RECT 103.740 105.660 104.070 106.750 ;
        RECT 104.440 106.280 105.480 106.450 ;
        RECT 104.440 105.840 105.480 106.010 ;
        RECT 105.650 105.980 105.820 106.310 ;
        RECT 103.900 105.440 104.070 105.660 ;
        RECT 106.160 105.440 106.330 106.850 ;
        RECT 103.900 105.270 106.330 105.440 ;
        RECT 107.910 107.360 118.540 107.530 ;
        RECT 120.020 116.640 126.250 116.800 ;
        RECT 120.020 114.380 120.690 116.640 ;
        RECT 121.360 116.070 125.400 116.240 ;
        RECT 121.020 115.010 121.190 116.010 ;
        RECT 125.570 115.010 125.740 116.010 ;
        RECT 121.360 114.780 125.400 114.950 ;
        RECT 126.080 114.380 126.250 116.640 ;
        RECT 120.020 114.210 126.250 114.380 ;
        RECT 120.020 110.950 120.690 114.210 ;
        RECT 121.360 113.640 125.400 113.810 ;
        RECT 121.020 111.580 121.190 113.580 ;
        RECT 125.570 111.580 125.740 113.580 ;
        RECT 121.360 111.350 125.400 111.520 ;
        RECT 126.080 110.950 126.250 114.210 ;
        RECT 120.020 110.780 126.250 110.950 ;
        RECT 120.020 107.520 120.690 110.780 ;
        RECT 121.360 110.210 125.400 110.380 ;
        RECT 121.020 108.150 121.190 110.150 ;
        RECT 125.570 108.150 125.740 110.150 ;
        RECT 121.360 107.920 125.400 108.090 ;
        RECT 126.080 107.520 126.250 110.780 ;
        RECT 120.020 107.510 126.250 107.520 ;
        RECT 127.840 116.780 137.670 116.820 ;
        RECT 140.540 116.800 146.280 116.810 ;
        RECT 127.840 116.650 138.470 116.780 ;
        RECT 127.840 114.390 128.010 116.650 ;
        RECT 128.735 116.080 136.775 116.250 ;
        RECT 128.350 115.020 128.520 116.020 ;
        RECT 136.990 115.020 137.160 116.020 ;
        RECT 128.735 114.790 136.775 114.960 ;
        RECT 137.500 114.390 138.470 116.650 ;
        RECT 127.840 114.220 138.470 114.390 ;
        RECT 127.840 110.960 128.010 114.220 ;
        RECT 128.735 113.650 136.775 113.820 ;
        RECT 128.350 111.590 128.520 113.590 ;
        RECT 136.990 111.590 137.160 113.590 ;
        RECT 128.735 111.360 136.775 111.530 ;
        RECT 137.500 110.960 138.470 114.220 ;
        RECT 127.840 110.790 138.470 110.960 ;
        RECT 127.840 107.530 128.010 110.790 ;
        RECT 128.735 110.220 136.775 110.390 ;
        RECT 128.350 108.160 128.520 110.160 ;
        RECT 136.990 108.160 137.160 110.160 ;
        RECT 128.735 107.930 136.775 108.100 ;
        RECT 137.500 107.530 138.470 110.790 ;
        RECT 120.020 107.410 126.260 107.510 ;
        RECT 107.910 105.100 108.080 107.360 ;
        RECT 108.805 106.790 116.845 106.960 ;
        RECT 108.420 105.730 108.590 106.730 ;
        RECT 117.060 105.730 117.230 106.730 ;
        RECT 108.805 105.500 116.845 105.670 ;
        RECT 117.570 105.100 118.540 107.360 ;
        RECT 120.010 106.850 126.260 107.410 ;
        RECT 120.010 106.830 125.180 106.850 ;
        RECT 120.010 106.760 124.000 106.830 ;
        RECT 120.010 105.490 121.930 106.760 ;
        RECT 123.440 106.750 124.000 106.760 ;
        RECT 123.670 105.660 124.000 106.750 ;
        RECT 124.370 106.280 125.410 106.450 ;
        RECT 124.370 105.840 125.410 106.010 ;
        RECT 125.580 105.980 125.750 106.310 ;
        RECT 123.830 105.440 124.000 105.660 ;
        RECT 126.090 105.440 126.260 106.850 ;
        RECT 123.830 105.270 126.260 105.440 ;
        RECT 127.840 107.360 138.470 107.530 ;
        RECT 140.050 116.640 146.280 116.800 ;
        RECT 140.050 114.380 140.720 116.640 ;
        RECT 141.390 116.070 145.430 116.240 ;
        RECT 141.050 115.010 141.220 116.010 ;
        RECT 145.600 115.010 145.770 116.010 ;
        RECT 141.390 114.780 145.430 114.950 ;
        RECT 146.110 114.380 146.280 116.640 ;
        RECT 140.050 114.210 146.280 114.380 ;
        RECT 140.050 110.950 140.720 114.210 ;
        RECT 141.390 113.640 145.430 113.810 ;
        RECT 141.050 111.580 141.220 113.580 ;
        RECT 145.600 111.580 145.770 113.580 ;
        RECT 141.390 111.350 145.430 111.520 ;
        RECT 146.110 110.950 146.280 114.210 ;
        RECT 140.050 110.780 146.280 110.950 ;
        RECT 140.050 107.520 140.720 110.780 ;
        RECT 141.390 110.210 145.430 110.380 ;
        RECT 141.050 108.150 141.220 110.150 ;
        RECT 145.600 108.150 145.770 110.150 ;
        RECT 141.390 107.920 145.430 108.090 ;
        RECT 146.110 107.520 146.280 110.780 ;
        RECT 140.050 107.510 146.280 107.520 ;
        RECT 147.870 116.780 157.700 116.820 ;
        RECT 147.870 116.650 158.500 116.780 ;
        RECT 147.870 114.390 148.040 116.650 ;
        RECT 148.765 116.080 156.805 116.250 ;
        RECT 148.380 115.020 148.550 116.020 ;
        RECT 157.020 115.020 157.190 116.020 ;
        RECT 148.765 114.790 156.805 114.960 ;
        RECT 157.530 114.390 158.500 116.650 ;
        RECT 147.870 114.220 158.500 114.390 ;
        RECT 147.870 110.960 148.040 114.220 ;
        RECT 148.765 113.650 156.805 113.820 ;
        RECT 148.380 111.590 148.550 113.590 ;
        RECT 157.020 111.590 157.190 113.590 ;
        RECT 148.765 111.360 156.805 111.530 ;
        RECT 157.530 110.960 158.500 114.220 ;
        RECT 147.870 110.790 158.500 110.960 ;
        RECT 147.870 107.530 148.040 110.790 ;
        RECT 148.765 110.220 156.805 110.390 ;
        RECT 148.380 108.160 148.550 110.160 ;
        RECT 157.020 108.160 157.190 110.160 ;
        RECT 148.765 107.930 156.805 108.100 ;
        RECT 157.530 107.530 158.500 110.790 ;
        RECT 140.050 107.410 146.290 107.510 ;
        RECT 107.910 105.070 118.540 105.100 ;
        RECT 127.840 105.100 128.010 107.360 ;
        RECT 128.735 106.790 136.775 106.960 ;
        RECT 128.350 105.730 128.520 106.730 ;
        RECT 136.990 105.730 137.160 106.730 ;
        RECT 128.735 105.500 136.775 105.670 ;
        RECT 137.500 105.100 138.470 107.360 ;
        RECT 140.040 106.850 146.290 107.410 ;
        RECT 140.040 106.830 145.210 106.850 ;
        RECT 140.040 106.760 144.030 106.830 ;
        RECT 140.040 105.490 141.960 106.760 ;
        RECT 143.470 106.750 144.030 106.760 ;
        RECT 143.700 105.660 144.030 106.750 ;
        RECT 144.400 106.280 145.440 106.450 ;
        RECT 144.400 105.840 145.440 106.010 ;
        RECT 145.610 105.980 145.780 106.310 ;
        RECT 143.860 105.440 144.030 105.660 ;
        RECT 146.120 105.440 146.290 106.850 ;
        RECT 143.860 105.270 146.290 105.440 ;
        RECT 147.870 107.360 158.500 107.530 ;
        RECT 127.840 105.070 138.470 105.100 ;
        RECT 147.870 105.100 148.040 107.360 ;
        RECT 148.765 106.790 156.805 106.960 ;
        RECT 148.380 105.730 148.550 106.730 ;
        RECT 157.020 105.730 157.190 106.730 ;
        RECT 148.765 105.500 156.805 105.670 ;
        RECT 157.530 105.100 158.500 107.360 ;
        RECT 147.870 105.070 158.500 105.100 ;
        RECT 107.880 104.960 118.540 105.070 ;
        RECT 127.810 104.960 138.470 105.070 ;
        RECT 147.840 104.960 158.500 105.070 ;
        RECT 106.130 104.910 118.540 104.960 ;
        RECT 126.060 104.910 138.470 104.960 ;
        RECT 146.090 104.910 158.500 104.960 ;
        RECT 101.790 104.740 118.540 104.910 ;
        RECT 101.790 103.330 101.960 104.740 ;
        RECT 102.330 104.170 105.370 104.340 ;
        RECT 102.330 103.730 105.370 103.900 ;
        RECT 105.585 103.870 105.755 104.200 ;
        RECT 106.090 103.980 118.540 104.740 ;
        RECT 121.720 104.740 138.470 104.910 ;
        RECT 106.090 103.970 118.430 103.980 ;
        RECT 106.090 103.960 111.970 103.970 ;
        RECT 106.090 103.940 106.660 103.960 ;
        RECT 107.880 103.950 111.970 103.960 ;
        RECT 106.100 103.330 106.270 103.940 ;
        RECT 101.790 103.160 106.270 103.330 ;
        RECT 121.720 103.330 121.890 104.740 ;
        RECT 122.260 104.170 125.300 104.340 ;
        RECT 122.260 103.730 125.300 103.900 ;
        RECT 125.515 103.870 125.685 104.200 ;
        RECT 126.020 103.980 138.470 104.740 ;
        RECT 141.750 104.740 158.500 104.910 ;
        RECT 126.020 103.970 138.360 103.980 ;
        RECT 126.020 103.960 131.900 103.970 ;
        RECT 126.020 103.940 126.590 103.960 ;
        RECT 127.810 103.950 131.900 103.960 ;
        RECT 126.030 103.330 126.200 103.940 ;
        RECT 121.720 103.160 126.200 103.330 ;
        RECT 141.750 103.330 141.920 104.740 ;
        RECT 142.290 104.170 145.330 104.340 ;
        RECT 142.290 103.730 145.330 103.900 ;
        RECT 145.545 103.870 145.715 104.200 ;
        RECT 146.050 103.980 158.500 104.740 ;
        RECT 146.050 103.970 158.390 103.980 ;
        RECT 146.050 103.960 151.930 103.970 ;
        RECT 146.050 103.940 146.620 103.960 ;
        RECT 147.840 103.950 151.930 103.960 ;
        RECT 146.060 103.330 146.230 103.940 ;
        RECT 141.750 103.160 146.230 103.330 ;
      LAYER met1 ;
        RECT 115.800 220.285 116.060 220.605 ;
        RECT 112.120 183.415 112.600 219.295 ;
        RECT 113.420 207.865 113.680 208.185 ;
        RECT 112.755 206.960 112.985 207.250 ;
        RECT 112.800 205.425 112.940 206.960 ;
        RECT 112.740 205.105 113.000 205.425 ;
        RECT 112.755 204.660 112.985 204.950 ;
        RECT 112.800 202.665 112.940 204.660 ;
        RECT 113.435 203.955 113.665 204.030 ;
        RECT 113.435 203.815 114.640 203.955 ;
        RECT 113.435 203.740 113.665 203.815 ;
        RECT 113.435 203.280 113.665 203.570 ;
        RECT 113.480 203.125 113.620 203.280 ;
        RECT 113.420 202.805 113.680 203.125 ;
        RECT 114.115 202.795 114.345 203.085 ;
        RECT 112.740 202.345 113.000 202.665 ;
        RECT 113.775 202.400 114.005 202.690 ;
        RECT 113.095 201.945 113.325 202.235 ;
        RECT 113.140 200.825 113.280 201.945 ;
        RECT 113.820 201.500 113.960 202.400 ;
        RECT 113.775 201.210 114.005 201.500 ;
        RECT 113.080 200.505 113.340 200.825 ;
        RECT 113.820 198.980 113.960 201.210 ;
        RECT 114.160 200.985 114.300 202.795 ;
        RECT 114.115 200.695 114.345 200.985 ;
        RECT 114.160 199.415 114.300 200.695 ;
        RECT 114.115 199.125 114.345 199.415 ;
        RECT 113.775 198.690 114.005 198.980 ;
        RECT 112.740 198.435 113.000 198.525 ;
        RECT 112.740 198.295 113.280 198.435 ;
        RECT 112.740 198.205 113.000 198.295 ;
        RECT 112.755 195.675 112.985 195.750 ;
        RECT 113.140 195.675 113.280 198.295 ;
        RECT 114.500 198.065 114.640 203.815 ;
        RECT 114.440 197.745 114.700 198.065 ;
        RECT 114.115 196.380 114.345 196.670 ;
        RECT 112.755 195.535 113.280 195.675 ;
        RECT 112.755 195.460 112.985 195.535 ;
        RECT 114.160 194.845 114.300 196.380 ;
        RECT 113.420 194.525 113.680 194.845 ;
        RECT 114.100 194.525 114.360 194.845 ;
        RECT 112.740 192.225 113.000 192.545 ;
        RECT 112.800 191.150 112.940 192.225 ;
        RECT 113.420 191.765 113.680 192.085 ;
        RECT 112.755 190.860 112.985 191.150 ;
        RECT 114.455 189.940 114.685 190.230 ;
        RECT 113.760 189.465 114.020 189.785 ;
        RECT 113.420 189.005 113.680 189.325 ;
        RECT 113.820 187.930 113.960 189.465 ;
        RECT 114.100 188.545 114.360 188.865 ;
        RECT 113.775 187.640 114.005 187.930 ;
        RECT 114.160 186.550 114.300 188.545 ;
        RECT 114.500 188.405 114.640 189.940 ;
        RECT 114.440 188.085 114.700 188.405 ;
        RECT 114.115 186.260 114.345 186.550 ;
        RECT 114.440 185.785 114.700 186.105 ;
        RECT 114.500 185.630 114.640 185.785 ;
        RECT 114.455 185.340 114.685 185.630 ;
        RECT 114.840 183.415 115.320 219.295 ;
        RECT 115.860 217.370 116.000 220.285 ;
        RECT 116.480 217.525 116.740 217.845 ;
        RECT 115.815 217.080 116.045 217.370 ;
        RECT 116.540 216.450 116.680 217.525 ;
        RECT 116.495 216.160 116.725 216.450 ;
        RECT 117.160 214.765 117.420 215.085 ;
        RECT 117.160 212.925 117.420 213.245 ;
        RECT 117.160 212.465 117.420 212.785 ;
        RECT 116.155 211.560 116.385 211.850 ;
        RECT 116.200 206.345 116.340 211.560 ;
        RECT 117.160 210.165 117.420 210.485 ;
        RECT 117.220 208.185 117.360 210.165 ;
        RECT 117.160 207.865 117.420 208.185 ;
        RECT 116.140 206.025 116.400 206.345 ;
        RECT 117.220 205.870 117.360 207.865 ;
        RECT 117.175 205.580 117.405 205.870 ;
        RECT 116.155 203.270 116.385 203.560 ;
        RECT 115.815 202.835 116.045 203.125 ;
        RECT 115.860 201.555 116.000 202.835 ;
        RECT 115.815 201.265 116.045 201.555 ;
        RECT 115.460 200.505 115.720 200.825 ;
        RECT 115.520 198.510 115.660 200.505 ;
        RECT 115.860 199.455 116.000 201.265 ;
        RECT 116.200 201.040 116.340 203.270 ;
        RECT 117.160 201.655 117.420 201.745 ;
        RECT 116.540 201.515 117.420 201.655 ;
        RECT 116.155 200.750 116.385 201.040 ;
        RECT 116.200 199.850 116.340 200.750 ;
        RECT 116.540 200.305 116.680 201.515 ;
        RECT 117.160 201.425 117.420 201.515 ;
        RECT 116.820 200.505 117.080 200.825 ;
        RECT 116.495 200.015 116.725 200.305 ;
        RECT 116.155 199.560 116.385 199.850 ;
        RECT 115.815 199.165 116.045 199.455 ;
        RECT 116.495 198.895 116.725 198.970 ;
        RECT 116.880 198.895 117.020 200.505 ;
        RECT 116.495 198.755 117.020 198.895 ;
        RECT 116.495 198.680 116.725 198.755 ;
        RECT 115.475 198.220 115.705 198.510 ;
        RECT 116.495 196.380 116.725 196.670 ;
        RECT 116.140 194.985 116.400 195.305 ;
        RECT 116.140 194.525 116.400 194.845 ;
        RECT 116.200 190.230 116.340 194.525 ;
        RECT 116.540 192.990 116.680 196.380 ;
        RECT 117.160 195.905 117.420 196.225 ;
        RECT 116.495 192.700 116.725 192.990 ;
        RECT 116.155 189.940 116.385 190.230 ;
        RECT 116.140 189.465 116.400 189.785 ;
        RECT 116.200 188.390 116.340 189.465 ;
        RECT 116.480 189.005 116.740 189.325 ;
        RECT 116.155 188.100 116.385 188.390 ;
        RECT 116.155 187.640 116.385 187.930 ;
        RECT 116.200 185.185 116.340 187.640 ;
        RECT 116.540 187.010 116.680 189.005 ;
        RECT 116.495 186.720 116.725 187.010 ;
        RECT 117.160 186.245 117.420 186.565 ;
        RECT 117.220 186.090 117.360 186.245 ;
        RECT 117.175 185.800 117.405 186.090 ;
        RECT 116.140 184.865 116.400 185.185 ;
        RECT 117.560 183.415 118.040 219.295 ;
        RECT 119.880 217.525 120.140 217.845 ;
        RECT 119.215 215.230 119.445 215.520 ;
        RECT 118.520 214.765 118.780 215.085 ;
        RECT 118.580 212.265 118.720 214.765 ;
        RECT 119.260 213.000 119.400 215.230 ;
        RECT 119.555 214.795 119.785 215.085 ;
        RECT 119.600 213.515 119.740 214.795 ;
        RECT 119.555 213.225 119.785 213.515 ;
        RECT 119.215 212.710 119.445 213.000 ;
        RECT 118.535 211.975 118.765 212.265 ;
        RECT 119.260 211.810 119.400 212.710 ;
        RECT 119.215 211.520 119.445 211.810 ;
        RECT 119.600 211.415 119.740 213.225 ;
        RECT 119.555 211.125 119.785 211.415 ;
        RECT 119.200 210.625 119.460 210.945 ;
        RECT 118.875 205.580 119.105 205.870 ;
        RECT 118.920 201.285 119.060 205.580 ;
        RECT 118.860 200.965 119.120 201.285 ;
        RECT 119.880 200.505 120.140 200.825 ;
        RECT 119.940 199.430 120.080 200.505 ;
        RECT 119.895 199.140 120.125 199.430 ;
        RECT 118.875 195.215 119.105 195.290 ;
        RECT 118.875 195.075 119.400 195.215 ;
        RECT 118.875 195.000 119.105 195.075 ;
        RECT 118.860 193.605 119.120 193.925 ;
        RECT 118.195 192.915 118.425 192.990 ;
        RECT 118.195 192.775 118.720 192.915 ;
        RECT 118.195 192.700 118.425 192.775 ;
        RECT 118.195 189.940 118.425 190.230 ;
        RECT 118.240 189.785 118.380 189.940 ;
        RECT 118.180 189.465 118.440 189.785 ;
        RECT 118.580 189.695 118.720 192.775 ;
        RECT 118.860 192.225 119.120 192.545 ;
        RECT 118.860 190.845 119.120 191.165 ;
        RECT 118.875 189.695 119.105 189.770 ;
        RECT 118.580 189.555 119.105 189.695 ;
        RECT 118.180 189.005 118.440 189.325 ;
        RECT 118.580 187.395 118.720 189.555 ;
        RECT 118.875 189.480 119.105 189.555 ;
        RECT 118.875 188.560 119.105 188.850 ;
        RECT 118.920 188.405 119.060 188.560 ;
        RECT 118.860 188.085 119.120 188.405 ;
        RECT 118.860 187.395 119.120 187.485 ;
        RECT 118.580 187.255 119.120 187.395 ;
        RECT 118.860 187.165 119.120 187.255 ;
        RECT 118.860 185.785 119.120 186.105 ;
        RECT 119.260 185.645 119.400 195.075 ;
        RECT 119.555 194.080 119.785 194.370 ;
        RECT 119.600 188.865 119.740 194.080 ;
        RECT 119.895 191.320 120.125 191.610 ;
        RECT 119.940 189.325 120.080 191.320 ;
        RECT 119.880 189.005 120.140 189.325 ;
        RECT 119.540 188.545 119.800 188.865 ;
        RECT 119.895 188.100 120.125 188.390 ;
        RECT 119.940 187.945 120.080 188.100 ;
        RECT 119.880 187.625 120.140 187.945 ;
        RECT 119.200 185.325 119.460 185.645 ;
        RECT 118.860 184.865 119.120 185.185 ;
        RECT 120.280 183.415 120.760 219.295 ;
        RECT 121.240 217.985 121.500 218.305 ;
        RECT 121.300 217.370 121.440 217.985 ;
        RECT 121.580 217.525 121.840 217.845 ;
        RECT 121.255 217.080 121.485 217.370 ;
        RECT 121.640 215.070 121.780 217.525 ;
        RECT 121.935 216.160 122.165 216.450 ;
        RECT 121.595 214.780 121.825 215.070 ;
        RECT 120.900 212.925 121.160 213.245 ;
        RECT 120.960 211.850 121.100 212.925 ;
        RECT 121.240 212.465 121.500 212.785 ;
        RECT 120.915 211.560 121.145 211.850 ;
        RECT 120.915 202.820 121.145 203.110 ;
        RECT 120.960 201.745 121.100 202.820 ;
        RECT 120.900 201.425 121.160 201.745 ;
        RECT 121.300 200.735 121.440 212.465 ;
        RECT 121.580 210.165 121.840 210.485 ;
        RECT 121.980 210.025 122.120 216.160 ;
        RECT 121.920 209.705 122.180 210.025 ;
        RECT 121.935 206.960 122.165 207.250 ;
        RECT 121.580 206.025 121.840 206.345 ;
        RECT 121.595 205.120 121.825 205.410 ;
        RECT 121.640 201.195 121.780 205.120 ;
        RECT 121.980 204.950 122.120 206.960 ;
        RECT 121.935 204.660 122.165 204.950 ;
        RECT 121.640 201.055 122.460 201.195 ;
        RECT 120.960 200.595 121.440 200.735 ;
        RECT 120.960 194.385 121.100 200.595 ;
        RECT 121.920 200.505 122.180 200.825 ;
        RECT 121.255 200.035 121.485 200.325 ;
        RECT 121.300 198.225 121.440 200.035 ;
        RECT 121.595 199.640 121.825 199.930 ;
        RECT 121.640 198.740 121.780 199.640 ;
        RECT 121.935 199.185 122.165 199.475 ;
        RECT 121.595 198.450 121.825 198.740 ;
        RECT 121.255 197.935 121.485 198.225 ;
        RECT 121.300 196.655 121.440 197.935 ;
        RECT 121.255 196.365 121.485 196.655 ;
        RECT 121.640 196.220 121.780 198.450 ;
        RECT 121.595 195.930 121.825 196.220 ;
        RECT 121.980 195.675 122.120 199.185 ;
        RECT 122.320 196.225 122.460 201.055 ;
        RECT 122.260 195.905 122.520 196.225 ;
        RECT 121.300 195.535 122.120 195.675 ;
        RECT 120.900 194.065 121.160 194.385 ;
        RECT 120.915 193.620 121.145 193.910 ;
        RECT 120.960 192.085 121.100 193.620 ;
        RECT 121.300 192.990 121.440 195.535 ;
        RECT 121.920 194.985 122.180 195.305 ;
        RECT 121.580 194.065 121.840 194.385 ;
        RECT 121.255 192.700 121.485 192.990 ;
        RECT 120.900 191.765 121.160 192.085 ;
        RECT 121.640 190.690 121.780 194.065 ;
        RECT 121.595 190.400 121.825 190.690 ;
        RECT 121.595 190.155 121.825 190.230 ;
        RECT 121.980 190.155 122.120 194.985 ;
        RECT 122.600 190.845 122.860 191.165 ;
        RECT 121.595 190.015 122.120 190.155 ;
        RECT 121.595 189.940 121.825 190.015 ;
        RECT 121.580 189.005 121.840 189.325 ;
        RECT 120.900 188.085 121.160 188.405 ;
        RECT 120.960 186.550 121.100 188.085 ;
        RECT 121.255 187.640 121.485 187.930 ;
        RECT 120.915 186.260 121.145 186.550 ;
        RECT 121.300 185.185 121.440 187.640 ;
        RECT 121.640 186.105 121.780 189.005 ;
        RECT 121.920 188.545 122.180 188.865 ;
        RECT 121.920 187.165 122.180 187.485 ;
        RECT 122.600 187.165 122.860 187.485 ;
        RECT 121.980 186.550 122.120 187.165 ;
        RECT 122.260 186.705 122.520 187.025 ;
        RECT 121.935 186.260 122.165 186.550 ;
        RECT 121.580 185.785 121.840 186.105 ;
        RECT 121.240 184.865 121.500 185.185 ;
        RECT 122.320 185.170 122.460 186.705 ;
        RECT 122.275 184.880 122.505 185.170 ;
        RECT 123.000 183.415 123.480 219.295 ;
        RECT 124.640 217.755 124.900 217.845 ;
        RECT 124.360 217.615 124.900 217.755 ;
        RECT 123.975 216.205 124.205 216.495 ;
        RECT 124.020 215.545 124.160 216.205 ;
        RECT 123.960 215.225 124.220 215.545 ;
        RECT 124.360 210.945 124.500 217.615 ;
        RECT 124.640 217.525 124.900 217.615 ;
        RECT 124.995 217.055 125.225 217.345 ;
        RECT 124.655 216.660 124.885 216.950 ;
        RECT 124.700 215.760 124.840 216.660 ;
        RECT 124.655 215.470 124.885 215.760 ;
        RECT 124.700 213.240 124.840 215.470 ;
        RECT 125.040 215.245 125.180 217.055 ;
        RECT 124.995 214.955 125.225 215.245 ;
        RECT 125.040 213.675 125.180 214.955 ;
        RECT 124.995 213.385 125.225 213.675 ;
        RECT 124.655 212.950 124.885 213.240 ;
        RECT 124.300 210.625 124.560 210.945 ;
        RECT 125.335 210.640 125.565 210.930 ;
        RECT 124.360 205.870 124.500 210.625 ;
        RECT 125.380 210.025 125.520 210.640 ;
        RECT 125.320 209.705 125.580 210.025 ;
        RECT 124.315 205.795 124.545 205.870 ;
        RECT 123.680 205.655 124.545 205.795 ;
        RECT 123.680 200.825 123.820 205.655 ;
        RECT 124.315 205.580 124.545 205.655 ;
        RECT 124.995 205.095 125.225 205.385 ;
        RECT 123.960 204.645 124.220 204.965 ;
        RECT 124.655 204.700 124.885 204.990 ;
        RECT 124.020 204.415 124.160 204.645 ;
        RECT 124.315 204.415 124.545 204.535 ;
        RECT 124.020 204.275 124.545 204.415 ;
        RECT 124.315 204.245 124.545 204.275 ;
        RECT 124.700 203.800 124.840 204.700 ;
        RECT 124.655 203.510 124.885 203.800 ;
        RECT 124.700 201.280 124.840 203.510 ;
        RECT 125.040 203.285 125.180 205.095 ;
        RECT 124.995 202.995 125.225 203.285 ;
        RECT 125.040 201.715 125.180 202.995 ;
        RECT 124.995 201.425 125.225 201.715 ;
        RECT 124.655 200.990 124.885 201.280 ;
        RECT 123.620 200.505 123.880 200.825 ;
        RECT 123.635 198.680 123.865 198.970 ;
        RECT 123.680 198.065 123.820 198.680 ;
        RECT 124.655 198.220 124.885 198.510 ;
        RECT 123.620 197.745 123.880 198.065 ;
        RECT 124.700 197.605 124.840 198.220 ;
        RECT 124.640 197.285 124.900 197.605 ;
        RECT 124.980 196.365 125.240 196.685 ;
        RECT 125.335 195.920 125.565 196.210 ;
        RECT 125.380 195.305 125.520 195.920 ;
        RECT 125.320 194.985 125.580 195.305 ;
        RECT 124.300 191.765 124.560 192.085 ;
        RECT 123.620 190.845 123.880 191.165 ;
        RECT 123.680 188.850 123.820 190.845 ;
        RECT 124.640 189.465 124.900 189.785 ;
        RECT 124.300 189.005 124.560 189.325 ;
        RECT 123.635 188.560 123.865 188.850 ;
        RECT 124.360 187.470 124.500 189.005 ;
        RECT 124.315 187.180 124.545 187.470 ;
        RECT 124.300 186.705 124.560 187.025 ;
        RECT 124.300 186.245 124.560 186.565 ;
        RECT 124.315 186.015 124.545 186.090 ;
        RECT 124.700 186.015 124.840 189.465 ;
        RECT 125.320 189.005 125.580 189.325 ;
        RECT 125.380 188.390 125.520 189.005 ;
        RECT 125.335 188.100 125.565 188.390 ;
        RECT 124.315 185.875 124.840 186.015 ;
        RECT 124.315 185.800 124.545 185.875 ;
        RECT 125.720 183.415 126.200 219.295 ;
        RECT 128.040 217.985 128.300 218.305 ;
        RECT 126.680 217.525 126.940 217.845 ;
        RECT 127.360 217.525 127.620 217.845 ;
        RECT 126.340 215.225 126.600 215.545 ;
        RECT 126.740 211.315 126.880 217.525 ;
        RECT 127.420 216.450 127.560 217.525 ;
        RECT 128.100 217.370 128.240 217.985 ;
        RECT 128.055 217.080 128.285 217.370 ;
        RECT 127.375 216.160 127.605 216.450 ;
        RECT 128.055 213.400 128.285 213.690 ;
        RECT 127.035 212.940 127.265 213.230 ;
        RECT 127.080 212.785 127.220 212.940 ;
        RECT 128.100 212.785 128.240 213.400 ;
        RECT 127.020 212.465 127.280 212.785 ;
        RECT 128.040 212.465 128.300 212.785 ;
        RECT 127.020 212.005 127.280 212.325 ;
        RECT 127.035 211.315 127.265 211.390 ;
        RECT 126.740 211.175 127.265 211.315 ;
        RECT 127.035 211.100 127.265 211.175 ;
        RECT 126.695 210.615 126.925 210.905 ;
        RECT 126.740 208.805 126.880 210.615 ;
        RECT 127.035 210.220 127.265 210.510 ;
        RECT 127.080 209.320 127.220 210.220 ;
        RECT 127.715 209.765 127.945 210.055 ;
        RECT 127.035 209.030 127.265 209.320 ;
        RECT 126.695 208.515 126.925 208.805 ;
        RECT 126.740 207.235 126.880 208.515 ;
        RECT 126.695 206.945 126.925 207.235 ;
        RECT 127.080 206.800 127.220 209.030 ;
        RECT 127.035 206.510 127.265 206.800 ;
        RECT 127.760 206.345 127.900 209.765 ;
        RECT 127.700 206.025 127.960 206.345 ;
        RECT 127.760 204.965 127.900 206.025 ;
        RECT 126.680 204.645 126.940 204.965 ;
        RECT 127.700 204.645 127.960 204.965 ;
        RECT 126.740 204.030 126.880 204.645 ;
        RECT 128.040 204.185 128.300 204.505 ;
        RECT 126.695 203.740 126.925 204.030 ;
        RECT 127.375 201.900 127.605 202.190 ;
        RECT 127.035 201.655 127.265 201.730 ;
        RECT 126.740 201.515 127.265 201.655 ;
        RECT 126.740 196.225 126.880 201.515 ;
        RECT 127.035 201.440 127.265 201.515 ;
        RECT 127.035 200.520 127.265 200.810 ;
        RECT 127.080 198.525 127.220 200.520 ;
        RECT 127.420 199.890 127.560 201.900 ;
        RECT 127.375 199.600 127.605 199.890 ;
        RECT 127.020 198.205 127.280 198.525 ;
        RECT 127.020 197.745 127.280 198.065 ;
        RECT 127.080 197.130 127.220 197.745 ;
        RECT 128.100 197.605 128.240 204.185 ;
        RECT 128.040 197.285 128.300 197.605 ;
        RECT 127.035 196.840 127.265 197.130 ;
        RECT 126.680 195.905 126.940 196.225 ;
        RECT 126.740 190.230 126.880 195.905 ;
        RECT 127.360 193.605 127.620 193.925 ;
        RECT 127.420 192.530 127.560 193.605 ;
        RECT 127.375 192.240 127.605 192.530 ;
        RECT 127.375 191.995 127.605 192.070 ;
        RECT 127.375 191.855 127.900 191.995 ;
        RECT 127.375 191.780 127.605 191.855 ;
        RECT 127.360 191.305 127.620 191.625 ;
        RECT 127.035 190.860 127.265 191.150 ;
        RECT 126.695 189.940 126.925 190.230 ;
        RECT 127.080 187.485 127.220 190.860 ;
        RECT 127.760 189.785 127.900 191.855 ;
        RECT 127.700 189.465 127.960 189.785 ;
        RECT 127.375 188.560 127.605 188.850 ;
        RECT 127.420 188.405 127.560 188.560 ;
        RECT 127.360 188.085 127.620 188.405 ;
        RECT 127.360 187.625 127.620 187.945 ;
        RECT 128.040 187.625 128.300 187.945 ;
        RECT 127.020 187.165 127.280 187.485 ;
        RECT 127.375 186.260 127.605 186.550 ;
        RECT 127.420 186.105 127.560 186.260 ;
        RECT 127.360 185.785 127.620 186.105 ;
        RECT 128.100 185.630 128.240 187.625 ;
        RECT 128.055 185.340 128.285 185.630 ;
        RECT 128.440 183.415 128.920 219.295 ;
        RECT 130.080 217.525 130.340 217.845 ;
        RECT 130.140 216.450 130.280 217.525 ;
        RECT 130.095 216.160 130.325 216.450 ;
        RECT 130.760 212.925 131.020 213.245 ;
        RECT 129.060 212.465 129.320 212.785 ;
        RECT 129.740 209.705 130.000 210.025 ;
        RECT 129.755 205.795 129.985 205.870 ;
        RECT 129.460 205.655 129.985 205.795 ;
        RECT 129.460 200.350 129.600 205.655 ;
        RECT 129.755 205.580 129.985 205.655 ;
        RECT 129.755 204.875 129.985 204.950 ;
        RECT 129.755 204.735 130.280 204.875 ;
        RECT 129.755 204.660 129.985 204.735 ;
        RECT 129.740 204.185 130.000 204.505 ;
        RECT 130.140 203.495 130.280 204.735 ;
        RECT 130.760 204.645 131.020 204.965 ;
        RECT 130.760 204.185 131.020 204.505 ;
        RECT 130.435 203.495 130.665 203.570 ;
        RECT 130.140 203.355 130.665 203.495 ;
        RECT 130.435 203.280 130.665 203.355 ;
        RECT 130.095 202.820 130.325 203.110 ;
        RECT 129.755 201.900 129.985 202.190 ;
        RECT 129.800 201.745 129.940 201.900 ;
        RECT 129.740 201.425 130.000 201.745 ;
        RECT 129.740 200.505 130.000 200.825 ;
        RECT 129.415 200.060 129.645 200.350 ;
        RECT 130.140 197.515 130.280 202.820 ;
        RECT 130.480 200.365 130.620 203.280 ;
        RECT 130.820 202.650 130.960 204.185 ;
        RECT 130.775 202.360 131.005 202.650 ;
        RECT 130.420 200.045 130.680 200.365 ;
        RECT 130.140 197.375 130.620 197.515 ;
        RECT 130.080 196.825 130.340 197.145 ;
        RECT 130.480 196.225 130.620 197.375 ;
        RECT 130.420 195.905 130.680 196.225 ;
        RECT 129.075 195.000 129.305 195.290 ;
        RECT 129.120 194.385 129.260 195.000 ;
        RECT 129.060 194.065 129.320 194.385 ;
        RECT 129.755 194.295 129.985 194.370 ;
        RECT 129.755 194.155 130.280 194.295 ;
        RECT 129.755 194.080 129.985 194.155 ;
        RECT 129.755 193.160 129.985 193.450 ;
        RECT 129.415 191.780 129.645 192.070 ;
        RECT 129.060 191.305 129.320 191.625 ;
        RECT 129.120 191.150 129.260 191.305 ;
        RECT 129.075 190.860 129.305 191.150 ;
        RECT 129.460 189.785 129.600 191.780 ;
        RECT 129.800 191.610 129.940 193.160 ;
        RECT 129.755 191.320 129.985 191.610 ;
        RECT 129.800 191.165 129.940 191.320 ;
        RECT 129.740 190.845 130.000 191.165 ;
        RECT 129.755 190.615 129.985 190.690 ;
        RECT 130.140 190.615 130.280 194.155 ;
        RECT 130.760 193.605 131.020 193.925 ;
        RECT 129.755 190.475 130.280 190.615 ;
        RECT 129.755 190.400 129.985 190.475 ;
        RECT 129.740 189.925 130.000 190.245 ;
        RECT 129.400 189.465 129.660 189.785 ;
        RECT 129.075 189.235 129.305 189.310 ;
        RECT 129.075 189.095 129.600 189.235 ;
        RECT 129.075 189.020 129.305 189.095 ;
        RECT 129.460 188.775 129.600 189.095 ;
        RECT 129.755 188.775 129.985 188.850 ;
        RECT 129.460 188.635 129.985 188.775 ;
        RECT 129.460 187.025 129.600 188.635 ;
        RECT 129.755 188.560 129.985 188.635 ;
        RECT 129.740 187.625 130.000 187.945 ;
        RECT 130.140 187.855 130.280 190.475 ;
        RECT 130.420 187.855 130.680 187.945 ;
        RECT 130.140 187.715 130.680 187.855 ;
        RECT 130.420 187.625 130.680 187.715 ;
        RECT 129.740 187.165 130.000 187.485 ;
        RECT 129.400 186.705 129.660 187.025 ;
        RECT 129.800 186.550 129.940 187.165 ;
        RECT 129.755 186.260 129.985 186.550 ;
        RECT 130.760 186.245 131.020 186.565 ;
        RECT 130.820 185.630 130.960 186.245 ;
        RECT 130.775 185.340 131.005 185.630 ;
        RECT 131.160 183.415 131.640 219.295 ;
        RECT 131.780 217.525 132.040 217.845 ;
        RECT 133.140 217.525 133.400 217.845 ;
        RECT 132.475 215.230 132.705 215.520 ;
        RECT 132.135 214.795 132.365 215.085 ;
        RECT 132.180 213.515 132.320 214.795 ;
        RECT 132.135 213.225 132.365 213.515 ;
        RECT 132.180 211.415 132.320 213.225 ;
        RECT 132.520 213.000 132.660 215.230 ;
        RECT 132.475 212.710 132.705 213.000 ;
        RECT 132.520 211.810 132.660 212.710 ;
        RECT 133.200 212.265 133.340 217.525 ;
        RECT 133.155 211.975 133.385 212.265 ;
        RECT 132.475 211.520 132.705 211.810 ;
        RECT 132.135 211.125 132.365 211.415 ;
        RECT 132.800 210.625 133.060 210.945 ;
        RECT 133.140 206.945 133.400 207.265 ;
        RECT 131.780 200.965 132.040 201.285 ;
        RECT 131.840 200.810 131.980 200.965 ;
        RECT 131.795 200.520 132.025 200.810 ;
        RECT 132.460 200.505 132.720 200.825 ;
        RECT 131.780 195.905 132.040 196.225 ;
        RECT 131.840 192.990 131.980 195.905 ;
        RECT 132.520 195.290 132.660 200.505 ;
        RECT 133.480 197.745 133.740 198.065 ;
        RECT 133.480 195.445 133.740 195.765 ;
        RECT 132.475 195.000 132.705 195.290 ;
        RECT 131.795 192.700 132.025 192.990 ;
        RECT 132.800 192.685 133.060 193.005 ;
        RECT 132.800 191.765 133.060 192.085 ;
        RECT 133.540 191.150 133.680 195.445 ;
        RECT 133.495 190.860 133.725 191.150 ;
        RECT 131.780 189.465 132.040 189.785 ;
        RECT 131.840 186.550 131.980 189.465 ;
        RECT 132.800 187.395 133.060 187.485 ;
        RECT 132.800 187.255 133.340 187.395 ;
        RECT 132.800 187.165 133.060 187.255 ;
        RECT 131.795 186.260 132.025 186.550 ;
        RECT 132.815 186.260 133.045 186.550 ;
        RECT 132.860 186.105 133.000 186.260 ;
        RECT 132.800 185.785 133.060 186.105 ;
        RECT 133.200 186.015 133.340 187.255 ;
        RECT 133.495 186.015 133.725 186.090 ;
        RECT 133.200 185.875 133.725 186.015 ;
        RECT 133.495 185.800 133.725 185.875 ;
        RECT 132.800 184.865 133.060 185.185 ;
        RECT 133.880 183.415 134.360 219.295 ;
        RECT 134.500 217.525 134.760 217.845 ;
        RECT 134.515 215.700 134.745 215.990 ;
        RECT 134.560 213.245 134.700 215.700 ;
        RECT 135.520 215.225 135.780 215.545 ;
        RECT 135.535 214.320 135.765 214.610 ;
        RECT 135.195 213.400 135.425 213.690 ;
        RECT 135.580 213.615 135.720 214.320 ;
        RECT 135.580 213.475 136.400 213.615 ;
        RECT 134.500 212.925 134.760 213.245 ;
        RECT 134.900 212.355 135.040 212.760 ;
        RECT 134.855 212.325 135.085 212.355 ;
        RECT 134.840 212.005 135.100 212.325 ;
        RECT 134.900 204.875 135.040 212.005 ;
        RECT 135.240 210.945 135.380 213.400 ;
        RECT 135.875 212.915 136.105 213.205 ;
        RECT 135.535 212.520 135.765 212.810 ;
        RECT 135.580 211.620 135.720 212.520 ;
        RECT 135.535 211.330 135.765 211.620 ;
        RECT 135.180 210.625 135.440 210.945 ;
        RECT 135.240 208.185 135.380 210.625 ;
        RECT 135.580 209.100 135.720 211.330 ;
        RECT 135.920 211.105 136.060 212.915 ;
        RECT 135.875 210.815 136.105 211.105 ;
        RECT 135.920 209.535 136.060 210.815 ;
        RECT 135.875 209.245 136.105 209.535 ;
        RECT 135.535 208.810 135.765 209.100 ;
        RECT 135.180 207.865 135.440 208.185 ;
        RECT 135.875 206.715 136.105 206.790 ;
        RECT 134.560 204.735 135.040 204.875 ;
        RECT 135.240 206.575 136.105 206.715 ;
        RECT 134.560 198.525 134.700 204.735 ;
        RECT 134.855 204.245 135.085 204.535 ;
        RECT 134.500 198.205 134.760 198.525 ;
        RECT 134.560 197.590 134.700 198.205 ;
        RECT 134.900 198.065 135.040 204.245 ;
        RECT 134.840 197.745 135.100 198.065 ;
        RECT 135.240 197.605 135.380 206.575 ;
        RECT 135.875 206.500 136.105 206.575 ;
        RECT 135.520 205.565 135.780 205.885 ;
        RECT 135.875 205.095 136.105 205.385 ;
        RECT 135.535 204.700 135.765 204.990 ;
        RECT 135.580 203.800 135.720 204.700 ;
        RECT 135.535 203.510 135.765 203.800 ;
        RECT 135.580 201.280 135.720 203.510 ;
        RECT 135.920 203.285 136.060 205.095 ;
        RECT 136.260 204.965 136.400 213.475 ;
        RECT 136.200 204.645 136.460 204.965 ;
        RECT 135.875 202.995 136.105 203.285 ;
        RECT 135.920 201.715 136.060 202.995 ;
        RECT 135.875 201.425 136.105 201.715 ;
        RECT 135.535 200.990 135.765 201.280 ;
        RECT 136.215 198.680 136.445 198.970 ;
        RECT 136.260 198.525 136.400 198.680 ;
        RECT 136.200 198.205 136.460 198.525 ;
        RECT 134.515 197.300 134.745 197.590 ;
        RECT 135.180 197.285 135.440 197.605 ;
        RECT 134.840 196.595 135.100 196.685 ;
        RECT 135.240 196.595 135.380 197.285 ;
        RECT 135.860 196.825 136.120 197.145 ;
        RECT 134.840 196.455 135.380 196.595 ;
        RECT 134.840 196.365 135.100 196.455 ;
        RECT 134.900 195.290 135.040 196.365 ;
        RECT 134.855 195.000 135.085 195.290 ;
        RECT 134.515 193.620 134.745 193.910 ;
        RECT 134.560 193.005 134.700 193.620 ;
        RECT 134.500 192.685 134.760 193.005 ;
        RECT 135.195 192.915 135.425 192.990 ;
        RECT 134.900 192.775 135.425 192.915 ;
        RECT 134.900 192.455 135.040 192.775 ;
        RECT 135.195 192.700 135.425 192.775 ;
        RECT 134.560 192.315 135.040 192.455 ;
        RECT 135.535 192.455 135.765 192.530 ;
        RECT 135.535 192.315 136.060 192.455 ;
        RECT 134.560 187.855 134.700 192.315 ;
        RECT 135.535 192.240 135.765 192.315 ;
        RECT 135.535 191.780 135.765 192.070 ;
        RECT 135.195 191.535 135.425 191.610 ;
        RECT 134.900 191.395 135.425 191.535 ;
        RECT 134.900 190.230 135.040 191.395 ;
        RECT 135.195 191.320 135.425 191.395 ;
        RECT 135.180 190.845 135.440 191.165 ;
        RECT 135.240 190.690 135.380 190.845 ;
        RECT 135.195 190.400 135.425 190.690 ;
        RECT 134.855 189.940 135.085 190.230 ;
        RECT 135.195 189.480 135.425 189.770 ;
        RECT 135.240 188.405 135.380 189.480 ;
        RECT 135.580 189.325 135.720 191.780 ;
        RECT 135.920 190.245 136.060 192.315 ;
        RECT 135.860 189.925 136.120 190.245 ;
        RECT 135.520 189.005 135.780 189.325 ;
        RECT 135.180 188.085 135.440 188.405 ;
        RECT 135.180 187.855 135.440 187.945 ;
        RECT 134.560 187.715 135.440 187.855 ;
        RECT 135.180 187.625 135.440 187.715 ;
        RECT 135.180 186.245 135.440 186.565 ;
        RECT 135.180 185.785 135.440 186.105 ;
        RECT 135.240 185.630 135.380 185.785 ;
        RECT 135.920 185.645 136.060 189.925 ;
        RECT 136.215 188.560 136.445 188.850 ;
        RECT 136.260 187.025 136.400 188.560 ;
        RECT 136.200 186.705 136.460 187.025 ;
        RECT 135.195 185.340 135.425 185.630 ;
        RECT 135.860 185.325 136.120 185.645 ;
        RECT 136.600 183.415 137.080 219.295 ;
        RECT 138.920 217.985 139.180 218.305 ;
        RECT 138.980 217.370 139.120 217.985 ;
        RECT 138.935 217.080 139.165 217.370 ;
        RECT 138.255 216.160 138.485 216.450 ;
        RECT 137.560 215.225 137.820 215.545 ;
        RECT 137.620 213.615 137.760 215.225 ;
        RECT 137.915 213.615 138.145 213.690 ;
        RECT 137.620 213.475 138.145 213.615 ;
        RECT 137.235 200.980 137.465 201.270 ;
        RECT 137.280 200.825 137.420 200.980 ;
        RECT 137.220 200.505 137.480 200.825 ;
        RECT 137.620 195.765 137.760 213.475 ;
        RECT 137.915 213.400 138.145 213.475 ;
        RECT 137.915 212.480 138.145 212.770 ;
        RECT 137.960 212.325 138.100 212.480 ;
        RECT 137.900 212.005 138.160 212.325 ;
        RECT 138.300 210.945 138.440 216.160 ;
        RECT 138.920 215.685 139.180 216.005 ;
        RECT 138.935 213.860 139.165 214.150 ;
        RECT 138.240 210.625 138.500 210.945 ;
        RECT 138.980 210.485 139.120 213.860 ;
        RECT 138.920 210.165 139.180 210.485 ;
        RECT 138.920 207.865 139.180 208.185 ;
        RECT 138.980 205.885 139.120 207.865 ;
        RECT 138.920 205.565 139.180 205.885 ;
        RECT 138.920 204.645 139.180 204.965 ;
        RECT 138.255 201.440 138.485 201.730 ;
        RECT 138.300 201.285 138.440 201.440 ;
        RECT 138.980 201.285 139.120 204.645 ;
        RECT 138.240 200.965 138.500 201.285 ;
        RECT 138.920 200.965 139.180 201.285 ;
        RECT 137.915 197.760 138.145 198.050 ;
        RECT 137.960 197.605 138.100 197.760 ;
        RECT 137.900 197.285 138.160 197.605 ;
        RECT 138.580 195.905 138.840 196.225 ;
        RECT 137.560 195.445 137.820 195.765 ;
        RECT 137.915 195.000 138.145 195.290 ;
        RECT 137.235 194.755 137.465 194.830 ;
        RECT 137.235 194.615 137.760 194.755 ;
        RECT 137.235 194.540 137.465 194.615 ;
        RECT 137.220 193.605 137.480 193.925 ;
        RECT 137.620 191.165 137.760 194.615 ;
        RECT 137.960 191.995 138.100 195.000 ;
        RECT 138.255 194.755 138.485 194.830 ;
        RECT 138.255 194.615 139.120 194.755 ;
        RECT 138.255 194.540 138.485 194.615 ;
        RECT 138.595 192.700 138.825 192.990 ;
        RECT 138.240 191.995 138.500 192.085 ;
        RECT 137.960 191.855 138.500 191.995 ;
        RECT 138.240 191.765 138.500 191.855 ;
        RECT 138.640 191.625 138.780 192.700 ;
        RECT 138.580 191.305 138.840 191.625 ;
        RECT 137.560 190.845 137.820 191.165 ;
        RECT 138.580 190.845 138.840 191.165 ;
        RECT 138.255 190.615 138.485 190.690 ;
        RECT 137.960 190.475 138.485 190.615 ;
        RECT 137.960 189.310 138.100 190.475 ;
        RECT 138.255 190.400 138.485 190.475 ;
        RECT 138.255 189.695 138.485 189.770 ;
        RECT 138.640 189.695 138.780 190.845 ;
        RECT 138.255 189.555 138.780 189.695 ;
        RECT 138.255 189.480 138.485 189.555 ;
        RECT 137.915 189.020 138.145 189.310 ;
        RECT 138.240 188.085 138.500 188.405 ;
        RECT 138.240 186.705 138.500 187.025 ;
        RECT 138.255 185.800 138.485 186.090 ;
        RECT 138.640 186.015 138.780 189.555 ;
        RECT 138.980 188.405 139.120 194.615 ;
        RECT 138.920 188.085 139.180 188.405 ;
        RECT 138.920 186.015 139.180 186.105 ;
        RECT 138.640 185.875 139.180 186.015 ;
        RECT 138.300 185.645 138.440 185.800 ;
        RECT 138.920 185.785 139.180 185.875 ;
        RECT 138.240 185.325 138.500 185.645 ;
        RECT 139.320 183.415 139.800 219.295 ;
        RECT 140.635 217.540 140.865 217.830 ;
        RECT 140.295 216.205 140.525 216.495 ;
        RECT 140.340 216.005 140.480 216.205 ;
        RECT 140.280 215.685 140.540 216.005 ;
        RECT 139.940 210.855 140.200 210.945 ;
        RECT 139.940 210.715 140.480 210.855 ;
        RECT 139.940 210.625 140.200 210.715 ;
        RECT 139.940 210.165 140.200 210.485 ;
        RECT 140.340 207.635 140.480 210.715 ;
        RECT 140.680 208.185 140.820 217.540 ;
        RECT 141.315 217.055 141.545 217.345 ;
        RECT 140.975 216.660 141.205 216.950 ;
        RECT 141.020 215.760 141.160 216.660 ;
        RECT 140.975 215.470 141.205 215.760 ;
        RECT 141.020 213.240 141.160 215.470 ;
        RECT 141.360 215.245 141.500 217.055 ;
        RECT 141.315 214.955 141.545 215.245 ;
        RECT 141.360 213.675 141.500 214.955 ;
        RECT 141.315 213.385 141.545 213.675 ;
        RECT 140.975 212.950 141.205 213.240 ;
        RECT 140.620 207.865 140.880 208.185 ;
        RECT 140.635 207.635 140.865 207.710 ;
        RECT 140.340 207.495 140.865 207.635 ;
        RECT 140.635 207.420 140.865 207.495 ;
        RECT 141.640 205.565 141.900 205.885 ;
        RECT 140.635 203.740 140.865 204.030 ;
        RECT 140.295 203.280 140.525 203.570 ;
        RECT 139.940 201.425 140.200 201.745 ;
        RECT 140.000 199.430 140.140 201.425 ;
        RECT 139.955 199.140 140.185 199.430 ;
        RECT 140.340 195.765 140.480 203.280 ;
        RECT 140.680 201.745 140.820 203.740 ;
        RECT 140.975 202.575 141.205 202.650 ;
        RECT 140.975 202.435 141.500 202.575 ;
        RECT 140.975 202.360 141.205 202.435 ;
        RECT 140.620 201.425 140.880 201.745 ;
        RECT 140.620 200.965 140.880 201.285 ;
        RECT 140.620 200.045 140.880 200.365 ;
        RECT 140.680 198.525 140.820 200.045 ;
        RECT 140.620 198.205 140.880 198.525 ;
        RECT 140.620 197.745 140.880 198.065 ;
        RECT 140.680 197.145 140.820 197.745 ;
        RECT 140.960 197.285 141.220 197.605 ;
        RECT 141.360 197.515 141.500 202.435 ;
        RECT 141.640 200.505 141.900 200.825 ;
        RECT 141.700 198.510 141.840 200.505 ;
        RECT 141.655 198.220 141.885 198.510 ;
        RECT 141.360 197.375 141.840 197.515 ;
        RECT 140.620 196.825 140.880 197.145 ;
        RECT 141.315 196.815 141.545 197.105 ;
        RECT 140.975 196.420 141.205 196.710 ;
        RECT 140.635 195.965 140.865 196.255 ;
        RECT 140.280 195.445 140.540 195.765 ;
        RECT 140.680 194.845 140.820 195.965 ;
        RECT 141.020 195.520 141.160 196.420 ;
        RECT 140.975 195.230 141.205 195.520 ;
        RECT 140.620 194.525 140.880 194.845 ;
        RECT 141.020 193.000 141.160 195.230 ;
        RECT 141.360 195.005 141.500 196.815 ;
        RECT 141.700 195.765 141.840 197.375 ;
        RECT 141.640 195.445 141.900 195.765 ;
        RECT 141.315 194.715 141.545 195.005 ;
        RECT 141.360 193.435 141.500 194.715 ;
        RECT 141.315 193.145 141.545 193.435 ;
        RECT 140.975 192.710 141.205 193.000 ;
        RECT 141.700 192.455 141.840 195.445 ;
        RECT 140.680 192.315 141.840 192.455 ;
        RECT 140.680 189.770 140.820 192.315 ;
        RECT 141.640 190.385 141.900 190.705 ;
        RECT 140.635 189.480 140.865 189.770 ;
        RECT 140.620 188.545 140.880 188.865 ;
        RECT 141.640 187.625 141.900 187.945 ;
        RECT 140.620 187.165 140.880 187.485 ;
        RECT 139.940 186.245 140.200 186.565 ;
        RECT 139.940 185.785 140.200 186.105 ;
        RECT 140.620 184.865 140.880 185.185 ;
        RECT 142.040 183.415 142.520 219.295 ;
        RECT 144.360 213.385 144.620 213.705 ;
        RECT 143.355 211.090 143.585 211.380 ;
        RECT 143.015 210.655 143.245 210.945 ;
        RECT 143.060 209.375 143.200 210.655 ;
        RECT 143.015 209.085 143.245 209.375 ;
        RECT 142.660 207.865 142.920 208.185 ;
        RECT 142.720 206.255 142.860 207.865 ;
        RECT 143.060 207.275 143.200 209.085 ;
        RECT 143.400 208.860 143.540 211.090 ;
        RECT 143.355 208.570 143.585 208.860 ;
        RECT 144.360 208.785 144.620 209.105 ;
        RECT 143.400 207.670 143.540 208.570 ;
        RECT 143.695 207.780 143.925 208.070 ;
        RECT 143.355 207.380 143.585 207.670 ;
        RECT 143.015 206.985 143.245 207.275 ;
        RECT 143.355 206.500 143.585 206.790 ;
        RECT 143.400 206.330 143.540 206.500 ;
        RECT 143.355 206.255 143.585 206.330 ;
        RECT 142.720 206.115 143.585 206.255 ;
        RECT 142.720 197.605 142.860 206.115 ;
        RECT 143.355 206.040 143.585 206.115 ;
        RECT 143.740 205.885 143.880 207.780 ;
        RECT 144.020 206.485 144.280 206.805 ;
        RECT 143.015 205.555 143.245 205.845 ;
        RECT 143.680 205.565 143.940 205.885 ;
        RECT 143.060 203.745 143.200 205.555 ;
        RECT 143.355 205.160 143.585 205.450 ;
        RECT 143.400 204.260 143.540 205.160 ;
        RECT 144.080 205.105 144.220 206.485 ;
        RECT 144.035 204.815 144.265 205.105 ;
        RECT 143.355 203.970 143.585 204.260 ;
        RECT 143.015 203.455 143.245 203.745 ;
        RECT 143.060 202.175 143.200 203.455 ;
        RECT 143.015 201.885 143.245 202.175 ;
        RECT 143.400 201.740 143.540 203.970 ;
        RECT 144.420 203.955 144.560 208.785 ;
        RECT 144.080 203.815 144.560 203.955 ;
        RECT 143.355 201.450 143.585 201.740 ;
        RECT 143.000 200.965 143.260 201.285 ;
        RECT 142.660 197.285 142.920 197.605 ;
        RECT 143.060 195.750 143.200 200.965 ;
        RECT 143.340 200.045 143.600 200.365 ;
        RECT 143.400 196.595 143.540 200.045 ;
        RECT 144.080 198.970 144.220 203.815 ;
        RECT 144.375 199.140 144.605 199.430 ;
        RECT 144.035 198.680 144.265 198.970 ;
        RECT 144.420 198.525 144.560 199.140 ;
        RECT 144.360 198.205 144.620 198.525 ;
        RECT 144.020 197.745 144.280 198.065 ;
        RECT 143.680 196.825 143.940 197.145 ;
        RECT 143.695 196.595 143.925 196.670 ;
        RECT 143.400 196.455 143.925 196.595 ;
        RECT 143.695 196.380 143.925 196.455 ;
        RECT 143.340 195.905 143.600 196.225 ;
        RECT 143.015 195.460 143.245 195.750 ;
        RECT 142.660 194.525 142.920 194.845 ;
        RECT 142.720 192.990 142.860 194.525 ;
        RECT 143.015 194.080 143.245 194.370 ;
        RECT 142.675 192.700 142.905 192.990 ;
        RECT 143.060 191.610 143.200 194.080 ;
        RECT 143.400 193.835 143.540 195.905 ;
        RECT 143.680 195.445 143.940 195.765 ;
        RECT 143.740 194.830 143.880 195.445 ;
        RECT 143.695 194.540 143.925 194.830 ;
        RECT 143.680 193.835 143.940 193.925 ;
        RECT 143.400 193.695 143.940 193.835 ;
        RECT 143.680 193.605 143.940 193.695 ;
        RECT 143.740 192.070 143.880 193.605 ;
        RECT 143.695 191.780 143.925 192.070 ;
        RECT 143.015 191.320 143.245 191.610 ;
        RECT 143.680 190.845 143.940 191.165 ;
        RECT 143.000 190.385 143.260 190.705 ;
        RECT 143.695 190.400 143.925 190.690 ;
        RECT 143.060 189.695 143.200 190.385 ;
        RECT 143.355 189.695 143.585 189.770 ;
        RECT 143.060 189.555 143.585 189.695 ;
        RECT 143.355 189.480 143.585 189.555 ;
        RECT 142.660 188.545 142.920 188.865 ;
        RECT 142.720 186.550 142.860 188.545 ;
        RECT 143.740 187.945 143.880 190.400 ;
        RECT 143.680 187.625 143.940 187.945 ;
        RECT 143.000 187.165 143.260 187.485 ;
        RECT 142.675 186.260 142.905 186.550 ;
        RECT 143.060 186.090 143.200 187.165 ;
        RECT 143.015 185.800 143.245 186.090 ;
        RECT 143.680 184.865 143.940 185.185 ;
        RECT 144.760 183.415 145.240 219.295 ;
        RECT 146.060 213.385 146.320 213.705 ;
        RECT 146.120 211.390 146.260 213.385 ;
        RECT 146.075 211.315 146.305 211.390 ;
        RECT 146.075 211.175 146.600 211.315 ;
        RECT 146.075 211.100 146.305 211.175 ;
        RECT 146.060 208.785 146.320 209.105 ;
        RECT 146.060 208.325 146.320 208.645 ;
        RECT 146.075 207.420 146.305 207.710 ;
        RECT 145.380 206.485 145.640 206.805 ;
        RECT 145.380 201.425 145.640 201.745 ;
        RECT 146.120 199.355 146.260 207.420 ;
        RECT 146.460 204.950 146.600 211.175 ;
        RECT 147.095 210.180 147.325 210.470 ;
        RECT 146.755 207.880 146.985 208.170 ;
        RECT 146.415 204.660 146.645 204.950 ;
        RECT 146.800 200.825 146.940 207.880 ;
        RECT 147.140 205.425 147.280 210.180 ;
        RECT 147.080 205.105 147.340 205.425 ;
        RECT 146.740 200.505 147.000 200.825 ;
        RECT 147.095 199.600 147.325 199.890 ;
        RECT 146.120 199.215 146.940 199.355 ;
        RECT 146.075 198.680 146.305 198.970 ;
        RECT 146.120 198.525 146.260 198.680 ;
        RECT 146.060 198.205 146.320 198.525 ;
        RECT 145.380 197.745 145.640 198.065 ;
        RECT 145.440 195.290 145.580 197.745 ;
        RECT 146.060 195.445 146.320 195.765 ;
        RECT 145.395 195.000 145.625 195.290 ;
        RECT 146.120 194.830 146.260 195.445 ;
        RECT 146.075 194.540 146.305 194.830 ;
        RECT 146.800 193.925 146.940 199.215 ;
        RECT 147.140 198.985 147.280 199.600 ;
        RECT 147.080 198.665 147.340 198.985 ;
        RECT 146.740 193.605 147.000 193.925 ;
        RECT 147.080 192.225 147.340 192.545 ;
        RECT 145.380 191.765 145.640 192.085 ;
        RECT 145.440 188.850 145.580 191.765 ;
        RECT 147.140 191.610 147.280 192.225 ;
        RECT 147.095 191.320 147.325 191.610 ;
        RECT 146.060 190.385 146.320 190.705 ;
        RECT 145.395 188.560 145.625 188.850 ;
        RECT 145.380 188.085 145.640 188.405 ;
        RECT 145.440 187.470 145.580 188.085 ;
        RECT 146.060 187.625 146.320 187.945 ;
        RECT 145.395 187.180 145.625 187.470 ;
        RECT 146.060 186.245 146.320 186.565 ;
        RECT 145.395 185.800 145.625 186.090 ;
        RECT 145.440 185.645 145.580 185.800 ;
        RECT 145.380 185.325 145.640 185.645 ;
        RECT 146.060 184.865 146.320 185.185 ;
        RECT 147.480 183.415 147.960 219.295 ;
        RECT 100.050 176.770 100.310 176.800 ;
        RECT 100.050 174.670 100.880 176.770 ;
        RECT 106.550 176.380 107.800 176.820 ;
        RECT 104.490 176.370 109.730 176.380 ;
        RECT 101.540 176.270 116.840 176.370 ;
        RECT 101.540 176.260 116.875 176.270 ;
        RECT 101.500 176.140 116.875 176.260 ;
        RECT 101.500 176.030 105.500 176.140 ;
        RECT 106.550 176.060 108.290 176.140 ;
        RECT 108.870 176.060 116.875 176.140 ;
        RECT 106.550 175.980 107.800 176.060 ;
        RECT 108.875 176.040 116.875 176.060 ;
        RECT 101.110 175.730 101.340 175.980 ;
        RECT 105.660 175.840 105.890 175.980 ;
        RECT 108.440 175.840 108.670 175.990 ;
        RECT 105.660 175.730 108.670 175.840 ;
        RECT 117.080 175.730 117.310 175.990 ;
        RECT 101.110 175.290 117.310 175.730 ;
        RECT 101.110 175.020 101.340 175.290 ;
        RECT 105.660 175.260 117.310 175.290 ;
        RECT 105.660 175.170 108.670 175.260 ;
        RECT 105.660 175.020 105.890 175.170 ;
        RECT 108.440 175.030 108.670 175.170 ;
        RECT 117.080 175.030 117.310 175.260 ;
        RECT 101.500 174.740 105.500 174.970 ;
        RECT 108.875 174.760 116.875 174.980 ;
        RECT 117.640 174.760 118.600 176.800 ;
        RECT 139.960 176.770 140.220 176.800 ;
        RECT 108.875 174.750 118.600 174.760 ;
        RECT 101.500 174.670 105.490 174.740 ;
        RECT 100.050 174.560 105.490 174.670 ;
        RECT 108.930 174.590 118.600 174.750 ;
        RECT 100.050 174.470 103.180 174.560 ;
        RECT 116.670 174.540 118.600 174.590 ;
        RECT 100.050 171.200 100.880 174.470 ;
        RECT 104.530 174.010 109.780 174.020 ;
        RECT 104.530 173.900 116.840 174.010 ;
        RECT 101.560 173.840 116.840 173.900 ;
        RECT 101.560 173.830 116.875 173.840 ;
        RECT 101.500 173.700 116.875 173.830 ;
        RECT 101.500 173.690 106.660 173.700 ;
        RECT 101.500 173.600 105.500 173.690 ;
        RECT 108.875 173.610 116.875 173.700 ;
        RECT 108.960 173.600 116.850 173.610 ;
        RECT 101.110 173.240 101.340 173.550 ;
        RECT 101.560 173.240 105.460 173.600 ;
        RECT 105.660 173.240 105.890 173.550 ;
        RECT 101.110 171.900 105.890 173.240 ;
        RECT 101.110 171.590 101.340 171.900 ;
        RECT 105.660 171.590 105.890 171.900 ;
        RECT 108.440 173.020 108.670 173.560 ;
        RECT 109.480 173.020 110.490 173.050 ;
        RECT 117.080 173.020 117.310 173.560 ;
        RECT 108.440 172.120 117.310 173.020 ;
        RECT 108.440 171.600 108.670 172.120 ;
        RECT 109.480 172.050 110.490 172.120 ;
        RECT 117.080 171.600 117.310 172.120 ;
        RECT 101.500 171.310 105.500 171.540 ;
        RECT 108.875 171.320 116.875 171.550 ;
        RECT 100.050 171.160 101.180 171.200 ;
        RECT 100.050 171.080 101.420 171.160 ;
        RECT 101.790 171.090 105.450 171.310 ;
        RECT 101.790 171.080 103.230 171.090 ;
        RECT 100.050 171.040 103.230 171.080 ;
        RECT 100.050 170.950 102.740 171.040 ;
        RECT 108.940 171.030 116.830 171.320 ;
        RECT 100.050 170.890 102.070 170.950 ;
        RECT 100.050 170.840 101.820 170.890 ;
        RECT 100.050 167.500 100.880 170.840 ;
        RECT 108.930 170.540 116.850 170.550 ;
        RECT 105.160 170.530 116.850 170.540 ;
        RECT 101.540 170.410 116.850 170.530 ;
        RECT 101.540 170.400 116.875 170.410 ;
        RECT 101.500 170.280 116.875 170.400 ;
        RECT 101.500 170.170 105.500 170.280 ;
        RECT 101.110 169.830 101.340 170.120 ;
        RECT 101.560 169.830 105.450 170.170 ;
        RECT 105.660 169.830 105.890 170.120 ;
        RECT 101.110 168.460 105.890 169.830 ;
        RECT 101.110 168.160 101.340 168.460 ;
        RECT 105.660 168.160 105.890 168.460 ;
        RECT 101.500 167.880 105.500 168.110 ;
        RECT 101.750 167.650 105.320 167.880 ;
        RECT 101.750 167.500 105.440 167.650 ;
        RECT 100.050 167.220 105.440 167.500 ;
        RECT 106.690 167.330 107.310 170.280 ;
        RECT 108.875 170.180 116.875 170.280 ;
        RECT 108.930 170.170 116.850 170.180 ;
        RECT 108.440 169.470 108.670 170.130 ;
        RECT 109.450 169.470 110.450 169.560 ;
        RECT 117.080 169.470 117.310 170.130 ;
        RECT 108.440 168.650 117.310 169.470 ;
        RECT 108.440 168.170 108.670 168.650 ;
        RECT 109.450 168.560 110.450 168.650 ;
        RECT 117.080 168.170 117.310 168.650 ;
        RECT 108.875 167.890 116.875 168.120 ;
        RECT 100.050 166.760 105.450 167.220 ;
        RECT 100.050 165.420 102.050 166.760 ;
        RECT 103.800 166.750 105.450 166.760 ;
        RECT 102.490 165.480 103.490 166.200 ;
        RECT 103.800 165.940 104.110 166.750 ;
        RECT 104.570 166.470 105.450 166.750 ;
        RECT 105.690 166.930 107.310 167.330 ;
        RECT 108.960 166.980 116.830 167.890 ;
        RECT 104.510 166.240 105.510 166.470 ;
        RECT 105.690 166.280 106.040 166.930 ;
        RECT 106.690 166.920 107.310 166.930 ;
        RECT 108.875 166.750 116.875 166.980 ;
        RECT 108.960 166.740 116.830 166.750 ;
        RECT 104.570 166.030 105.450 166.050 ;
        RECT 103.840 165.650 104.110 165.940 ;
        RECT 104.510 165.800 105.510 166.030 ;
        RECT 105.670 165.990 106.040 166.280 ;
        RECT 105.700 165.930 106.040 165.990 ;
        RECT 106.800 166.600 107.560 166.650 ;
        RECT 108.440 166.600 108.670 166.700 ;
        RECT 106.800 166.390 108.670 166.600 ;
        RECT 117.080 166.390 117.310 166.700 ;
        RECT 106.800 165.970 109.340 166.390 ;
        RECT 116.710 165.970 117.310 166.390 ;
        RECT 104.570 165.650 105.450 165.800 ;
        RECT 104.580 165.480 105.310 165.650 ;
        RECT 100.130 165.410 102.050 165.420 ;
        RECT 102.460 164.360 105.310 165.480 ;
        RECT 105.700 165.180 106.050 165.930 ;
        RECT 106.800 165.810 108.670 165.970 ;
        RECT 106.800 165.760 107.560 165.810 ;
        RECT 108.440 165.740 108.670 165.810 ;
        RECT 117.080 165.740 117.310 165.970 ;
        RECT 108.875 165.460 116.875 165.690 ;
        RECT 105.700 165.120 105.990 165.180 ;
        RECT 105.610 165.000 105.990 165.120 ;
        RECT 108.970 165.060 116.830 165.460 ;
        RECT 117.640 165.060 118.600 174.540 ;
        RECT 119.930 176.720 120.190 176.750 ;
        RECT 119.930 174.620 120.760 176.720 ;
        RECT 126.430 176.330 127.680 176.770 ;
        RECT 124.370 176.320 129.610 176.330 ;
        RECT 121.420 176.220 136.720 176.320 ;
        RECT 121.420 176.210 136.755 176.220 ;
        RECT 121.380 176.090 136.755 176.210 ;
        RECT 121.380 175.980 125.380 176.090 ;
        RECT 126.430 176.010 128.170 176.090 ;
        RECT 128.750 176.010 136.755 176.090 ;
        RECT 126.430 175.930 127.680 176.010 ;
        RECT 128.755 175.990 136.755 176.010 ;
        RECT 120.990 175.680 121.220 175.930 ;
        RECT 125.540 175.790 125.770 175.930 ;
        RECT 128.320 175.790 128.550 175.940 ;
        RECT 125.540 175.680 128.550 175.790 ;
        RECT 136.960 175.680 137.190 175.940 ;
        RECT 120.990 175.240 137.190 175.680 ;
        RECT 120.990 174.970 121.220 175.240 ;
        RECT 125.540 175.210 137.190 175.240 ;
        RECT 125.540 175.120 128.550 175.210 ;
        RECT 125.540 174.970 125.770 175.120 ;
        RECT 128.320 174.980 128.550 175.120 ;
        RECT 136.960 174.980 137.190 175.210 ;
        RECT 121.380 174.690 125.380 174.920 ;
        RECT 128.755 174.710 136.755 174.930 ;
        RECT 137.520 174.710 138.480 176.750 ;
        RECT 128.755 174.700 138.480 174.710 ;
        RECT 121.380 174.620 125.370 174.690 ;
        RECT 119.930 174.510 125.370 174.620 ;
        RECT 128.810 174.540 138.480 174.700 ;
        RECT 119.930 174.420 123.060 174.510 ;
        RECT 136.550 174.490 138.480 174.540 ;
        RECT 119.930 171.150 120.760 174.420 ;
        RECT 124.410 173.960 129.660 173.970 ;
        RECT 124.410 173.850 136.720 173.960 ;
        RECT 121.440 173.790 136.720 173.850 ;
        RECT 121.440 173.780 136.755 173.790 ;
        RECT 121.380 173.650 136.755 173.780 ;
        RECT 121.380 173.640 126.540 173.650 ;
        RECT 121.380 173.550 125.380 173.640 ;
        RECT 128.755 173.560 136.755 173.650 ;
        RECT 128.840 173.550 136.730 173.560 ;
        RECT 120.990 173.190 121.220 173.500 ;
        RECT 121.440 173.190 125.340 173.550 ;
        RECT 125.540 173.190 125.770 173.500 ;
        RECT 120.990 171.850 125.770 173.190 ;
        RECT 120.990 171.540 121.220 171.850 ;
        RECT 125.540 171.540 125.770 171.850 ;
        RECT 128.320 172.970 128.550 173.510 ;
        RECT 129.360 172.970 130.370 173.000 ;
        RECT 136.960 172.970 137.190 173.510 ;
        RECT 128.320 172.070 137.190 172.970 ;
        RECT 128.320 171.550 128.550 172.070 ;
        RECT 129.360 172.000 130.370 172.070 ;
        RECT 136.960 171.550 137.190 172.070 ;
        RECT 121.380 171.260 125.380 171.490 ;
        RECT 128.755 171.270 136.755 171.500 ;
        RECT 119.930 171.110 121.060 171.150 ;
        RECT 119.930 171.030 121.300 171.110 ;
        RECT 121.670 171.040 125.330 171.260 ;
        RECT 121.670 171.030 123.110 171.040 ;
        RECT 119.930 170.990 123.110 171.030 ;
        RECT 119.930 170.900 122.620 170.990 ;
        RECT 128.820 170.980 136.710 171.270 ;
        RECT 119.930 170.840 121.950 170.900 ;
        RECT 119.930 170.790 121.700 170.840 ;
        RECT 119.930 167.450 120.760 170.790 ;
        RECT 128.810 170.490 136.730 170.500 ;
        RECT 125.040 170.480 136.730 170.490 ;
        RECT 121.420 170.360 136.730 170.480 ;
        RECT 121.420 170.350 136.755 170.360 ;
        RECT 121.380 170.230 136.755 170.350 ;
        RECT 121.380 170.120 125.380 170.230 ;
        RECT 120.990 169.780 121.220 170.070 ;
        RECT 121.440 169.780 125.330 170.120 ;
        RECT 125.540 169.780 125.770 170.070 ;
        RECT 120.990 168.410 125.770 169.780 ;
        RECT 120.990 168.110 121.220 168.410 ;
        RECT 125.540 168.110 125.770 168.410 ;
        RECT 121.380 167.830 125.380 168.060 ;
        RECT 121.630 167.600 125.200 167.830 ;
        RECT 121.630 167.450 125.320 167.600 ;
        RECT 119.930 167.170 125.320 167.450 ;
        RECT 126.570 167.280 127.190 170.230 ;
        RECT 128.755 170.130 136.755 170.230 ;
        RECT 128.810 170.120 136.730 170.130 ;
        RECT 128.320 169.420 128.550 170.080 ;
        RECT 129.330 169.420 130.330 169.510 ;
        RECT 136.960 169.420 137.190 170.080 ;
        RECT 128.320 168.600 137.190 169.420 ;
        RECT 128.320 168.120 128.550 168.600 ;
        RECT 129.330 168.510 130.330 168.600 ;
        RECT 136.960 168.120 137.190 168.600 ;
        RECT 128.755 167.840 136.755 168.070 ;
        RECT 119.930 166.710 125.330 167.170 ;
        RECT 119.930 165.370 121.930 166.710 ;
        RECT 123.680 166.700 125.330 166.710 ;
        RECT 122.370 165.430 123.370 166.150 ;
        RECT 123.680 165.890 123.990 166.700 ;
        RECT 124.450 166.420 125.330 166.700 ;
        RECT 125.570 166.880 127.190 167.280 ;
        RECT 128.840 166.930 136.710 167.840 ;
        RECT 124.390 166.190 125.390 166.420 ;
        RECT 125.570 166.230 125.920 166.880 ;
        RECT 126.570 166.870 127.190 166.880 ;
        RECT 128.755 166.700 136.755 166.930 ;
        RECT 128.840 166.690 136.710 166.700 ;
        RECT 124.450 165.980 125.330 166.000 ;
        RECT 123.720 165.600 123.990 165.890 ;
        RECT 124.390 165.750 125.390 165.980 ;
        RECT 125.550 165.940 125.920 166.230 ;
        RECT 125.580 165.880 125.920 165.940 ;
        RECT 126.680 166.550 127.440 166.600 ;
        RECT 128.320 166.550 128.550 166.650 ;
        RECT 126.680 166.340 128.550 166.550 ;
        RECT 136.960 166.340 137.190 166.650 ;
        RECT 126.680 165.920 129.220 166.340 ;
        RECT 136.590 165.920 137.190 166.340 ;
        RECT 124.450 165.600 125.330 165.750 ;
        RECT 124.460 165.430 125.190 165.600 ;
        RECT 120.010 165.360 121.930 165.370 ;
        RECT 102.400 164.130 105.400 164.360 ;
        RECT 105.610 164.170 105.950 165.000 ;
        RECT 107.960 164.990 118.600 165.060 ;
        RECT 102.450 164.100 105.310 164.130 ;
        RECT 102.450 164.080 103.620 164.100 ;
        RECT 104.580 164.090 105.310 164.100 ;
        RECT 102.400 163.690 105.400 163.920 ;
        RECT 105.605 163.880 105.950 164.170 ;
        RECT 106.140 163.950 118.600 164.990 ;
        RECT 122.340 164.310 125.190 165.430 ;
        RECT 125.580 165.130 125.930 165.880 ;
        RECT 126.680 165.760 128.550 165.920 ;
        RECT 126.680 165.710 127.440 165.760 ;
        RECT 128.320 165.690 128.550 165.760 ;
        RECT 136.960 165.690 137.190 165.920 ;
        RECT 128.755 165.410 136.755 165.640 ;
        RECT 125.580 165.070 125.870 165.130 ;
        RECT 125.490 164.950 125.870 165.070 ;
        RECT 128.850 165.010 136.710 165.410 ;
        RECT 137.520 165.010 138.480 174.490 ;
        RECT 139.960 174.670 140.790 176.770 ;
        RECT 146.460 176.380 147.710 176.820 ;
        RECT 144.400 176.370 149.640 176.380 ;
        RECT 141.450 176.270 156.750 176.370 ;
        RECT 141.450 176.260 156.785 176.270 ;
        RECT 141.410 176.140 156.785 176.260 ;
        RECT 141.410 176.030 145.410 176.140 ;
        RECT 146.460 176.060 148.200 176.140 ;
        RECT 148.780 176.060 156.785 176.140 ;
        RECT 146.460 175.980 147.710 176.060 ;
        RECT 148.785 176.040 156.785 176.060 ;
        RECT 141.020 175.730 141.250 175.980 ;
        RECT 145.570 175.840 145.800 175.980 ;
        RECT 148.350 175.840 148.580 175.990 ;
        RECT 145.570 175.730 148.580 175.840 ;
        RECT 156.990 175.730 157.220 175.990 ;
        RECT 141.020 175.290 157.220 175.730 ;
        RECT 141.020 175.020 141.250 175.290 ;
        RECT 145.570 175.260 157.220 175.290 ;
        RECT 145.570 175.170 148.580 175.260 ;
        RECT 145.570 175.020 145.800 175.170 ;
        RECT 148.350 175.030 148.580 175.170 ;
        RECT 156.990 175.030 157.220 175.260 ;
        RECT 141.410 174.740 145.410 174.970 ;
        RECT 148.785 174.760 156.785 174.980 ;
        RECT 157.550 174.760 158.510 176.800 ;
        RECT 148.785 174.750 158.510 174.760 ;
        RECT 141.410 174.670 145.400 174.740 ;
        RECT 139.960 174.560 145.400 174.670 ;
        RECT 148.840 174.590 158.510 174.750 ;
        RECT 139.960 174.470 143.090 174.560 ;
        RECT 156.580 174.540 158.510 174.590 ;
        RECT 139.960 171.200 140.790 174.470 ;
        RECT 144.440 174.010 149.690 174.020 ;
        RECT 144.440 173.900 156.750 174.010 ;
        RECT 141.470 173.840 156.750 173.900 ;
        RECT 141.470 173.830 156.785 173.840 ;
        RECT 141.410 173.700 156.785 173.830 ;
        RECT 141.410 173.690 146.570 173.700 ;
        RECT 141.410 173.600 145.410 173.690 ;
        RECT 148.785 173.610 156.785 173.700 ;
        RECT 148.870 173.600 156.760 173.610 ;
        RECT 141.020 173.240 141.250 173.550 ;
        RECT 141.470 173.240 145.370 173.600 ;
        RECT 145.570 173.240 145.800 173.550 ;
        RECT 141.020 171.900 145.800 173.240 ;
        RECT 141.020 171.590 141.250 171.900 ;
        RECT 145.570 171.590 145.800 171.900 ;
        RECT 148.350 173.020 148.580 173.560 ;
        RECT 149.390 173.020 150.400 173.050 ;
        RECT 156.990 173.020 157.220 173.560 ;
        RECT 148.350 172.120 157.220 173.020 ;
        RECT 148.350 171.600 148.580 172.120 ;
        RECT 149.390 172.050 150.400 172.120 ;
        RECT 156.990 171.600 157.220 172.120 ;
        RECT 141.410 171.310 145.410 171.540 ;
        RECT 148.785 171.320 156.785 171.550 ;
        RECT 139.960 171.160 141.090 171.200 ;
        RECT 139.960 171.080 141.330 171.160 ;
        RECT 141.700 171.090 145.360 171.310 ;
        RECT 141.700 171.080 143.140 171.090 ;
        RECT 139.960 171.040 143.140 171.080 ;
        RECT 139.960 170.950 142.650 171.040 ;
        RECT 148.850 171.030 156.740 171.320 ;
        RECT 139.960 170.890 141.980 170.950 ;
        RECT 139.960 170.840 141.730 170.890 ;
        RECT 139.960 167.500 140.790 170.840 ;
        RECT 148.840 170.540 156.760 170.550 ;
        RECT 145.070 170.530 156.760 170.540 ;
        RECT 141.450 170.410 156.760 170.530 ;
        RECT 141.450 170.400 156.785 170.410 ;
        RECT 141.410 170.280 156.785 170.400 ;
        RECT 141.410 170.170 145.410 170.280 ;
        RECT 141.020 169.830 141.250 170.120 ;
        RECT 141.470 169.830 145.360 170.170 ;
        RECT 145.570 169.830 145.800 170.120 ;
        RECT 141.020 168.460 145.800 169.830 ;
        RECT 141.020 168.160 141.250 168.460 ;
        RECT 145.570 168.160 145.800 168.460 ;
        RECT 141.410 167.880 145.410 168.110 ;
        RECT 141.660 167.650 145.230 167.880 ;
        RECT 141.660 167.500 145.350 167.650 ;
        RECT 139.960 167.220 145.350 167.500 ;
        RECT 146.600 167.330 147.220 170.280 ;
        RECT 148.785 170.180 156.785 170.280 ;
        RECT 148.840 170.170 156.760 170.180 ;
        RECT 148.350 169.470 148.580 170.130 ;
        RECT 149.360 169.470 150.360 169.560 ;
        RECT 156.990 169.470 157.220 170.130 ;
        RECT 148.350 168.650 157.220 169.470 ;
        RECT 148.350 168.170 148.580 168.650 ;
        RECT 149.360 168.560 150.360 168.650 ;
        RECT 156.990 168.170 157.220 168.650 ;
        RECT 148.785 167.890 156.785 168.120 ;
        RECT 139.960 166.760 145.360 167.220 ;
        RECT 139.960 165.420 141.960 166.760 ;
        RECT 143.710 166.750 145.360 166.760 ;
        RECT 142.400 165.480 143.400 166.200 ;
        RECT 143.710 165.940 144.020 166.750 ;
        RECT 144.480 166.470 145.360 166.750 ;
        RECT 145.600 166.930 147.220 167.330 ;
        RECT 148.870 166.980 156.740 167.890 ;
        RECT 144.420 166.240 145.420 166.470 ;
        RECT 145.600 166.280 145.950 166.930 ;
        RECT 146.600 166.920 147.220 166.930 ;
        RECT 148.785 166.750 156.785 166.980 ;
        RECT 148.870 166.740 156.740 166.750 ;
        RECT 144.480 166.030 145.360 166.050 ;
        RECT 143.750 165.650 144.020 165.940 ;
        RECT 144.420 165.800 145.420 166.030 ;
        RECT 145.580 165.990 145.950 166.280 ;
        RECT 145.610 165.930 145.950 165.990 ;
        RECT 146.710 166.600 147.470 166.650 ;
        RECT 148.350 166.600 148.580 166.700 ;
        RECT 146.710 166.390 148.580 166.600 ;
        RECT 156.990 166.390 157.220 166.700 ;
        RECT 146.710 165.970 149.250 166.390 ;
        RECT 156.620 165.970 157.220 166.390 ;
        RECT 144.480 165.650 145.360 165.800 ;
        RECT 144.490 165.480 145.220 165.650 ;
        RECT 140.040 165.410 141.960 165.420 ;
        RECT 122.280 164.080 125.280 164.310 ;
        RECT 125.490 164.120 125.830 164.950 ;
        RECT 127.840 164.940 138.480 165.010 ;
        RECT 122.330 164.050 125.190 164.080 ;
        RECT 122.330 164.030 123.500 164.050 ;
        RECT 124.460 164.040 125.190 164.050 ;
        RECT 106.140 163.930 118.470 163.950 ;
        RECT 106.410 163.920 111.850 163.930 ;
        RECT 112.850 163.920 118.470 163.930 ;
        RECT 105.610 163.770 105.950 163.880 ;
        RECT 122.280 163.640 125.280 163.870 ;
        RECT 125.485 163.830 125.830 164.120 ;
        RECT 126.020 163.900 138.480 164.940 ;
        RECT 142.370 164.360 145.220 165.480 ;
        RECT 145.610 165.180 145.960 165.930 ;
        RECT 146.710 165.810 148.580 165.970 ;
        RECT 146.710 165.760 147.470 165.810 ;
        RECT 148.350 165.740 148.580 165.810 ;
        RECT 156.990 165.740 157.220 165.970 ;
        RECT 148.785 165.460 156.785 165.690 ;
        RECT 145.610 165.120 145.900 165.180 ;
        RECT 145.520 165.000 145.900 165.120 ;
        RECT 148.880 165.060 156.740 165.460 ;
        RECT 157.550 165.060 158.510 174.540 ;
        RECT 142.310 164.130 145.310 164.360 ;
        RECT 145.520 164.170 145.860 165.000 ;
        RECT 147.870 164.990 158.510 165.060 ;
        RECT 142.360 164.100 145.220 164.130 ;
        RECT 142.360 164.080 143.530 164.100 ;
        RECT 144.490 164.090 145.220 164.100 ;
        RECT 126.020 163.880 138.350 163.900 ;
        RECT 126.290 163.870 131.730 163.880 ;
        RECT 132.730 163.870 138.350 163.880 ;
        RECT 125.490 163.720 125.830 163.830 ;
        RECT 142.310 163.690 145.310 163.920 ;
        RECT 145.515 163.880 145.860 164.170 ;
        RECT 146.050 163.950 158.510 164.990 ;
        RECT 146.050 163.930 158.380 163.950 ;
        RECT 146.320 163.920 151.760 163.930 ;
        RECT 152.760 163.920 158.380 163.930 ;
        RECT 145.520 163.770 145.860 163.880 ;
        RECT 100.050 161.770 100.310 161.800 ;
        RECT 100.050 159.670 100.880 161.770 ;
        RECT 106.550 161.380 107.800 161.820 ;
        RECT 104.490 161.370 109.730 161.380 ;
        RECT 101.540 161.270 116.840 161.370 ;
        RECT 101.540 161.260 116.875 161.270 ;
        RECT 101.500 161.140 116.875 161.260 ;
        RECT 101.500 161.030 105.500 161.140 ;
        RECT 106.550 161.060 108.290 161.140 ;
        RECT 108.870 161.060 116.875 161.140 ;
        RECT 106.550 160.980 107.800 161.060 ;
        RECT 108.875 161.040 116.875 161.060 ;
        RECT 101.110 160.730 101.340 160.980 ;
        RECT 105.660 160.840 105.890 160.980 ;
        RECT 108.440 160.840 108.670 160.990 ;
        RECT 105.660 160.730 108.670 160.840 ;
        RECT 117.080 160.730 117.310 160.990 ;
        RECT 101.110 160.290 117.310 160.730 ;
        RECT 101.110 160.020 101.340 160.290 ;
        RECT 105.660 160.260 117.310 160.290 ;
        RECT 105.660 160.170 108.670 160.260 ;
        RECT 105.660 160.020 105.890 160.170 ;
        RECT 108.440 160.030 108.670 160.170 ;
        RECT 117.080 160.030 117.310 160.260 ;
        RECT 101.500 159.740 105.500 159.970 ;
        RECT 108.875 159.760 116.875 159.980 ;
        RECT 117.640 159.760 118.600 161.800 ;
        RECT 108.875 159.750 118.600 159.760 ;
        RECT 101.500 159.670 105.490 159.740 ;
        RECT 100.050 159.560 105.490 159.670 ;
        RECT 108.930 159.590 118.600 159.750 ;
        RECT 100.050 159.470 103.180 159.560 ;
        RECT 116.670 159.540 118.600 159.590 ;
        RECT 100.050 156.200 100.880 159.470 ;
        RECT 104.530 159.010 109.780 159.020 ;
        RECT 104.530 158.900 116.840 159.010 ;
        RECT 101.560 158.840 116.840 158.900 ;
        RECT 101.560 158.830 116.875 158.840 ;
        RECT 101.500 158.700 116.875 158.830 ;
        RECT 101.500 158.690 106.660 158.700 ;
        RECT 101.500 158.600 105.500 158.690 ;
        RECT 108.875 158.610 116.875 158.700 ;
        RECT 108.960 158.600 116.850 158.610 ;
        RECT 101.110 158.240 101.340 158.550 ;
        RECT 101.560 158.240 105.460 158.600 ;
        RECT 105.660 158.240 105.890 158.550 ;
        RECT 101.110 156.900 105.890 158.240 ;
        RECT 101.110 156.590 101.340 156.900 ;
        RECT 105.660 156.590 105.890 156.900 ;
        RECT 108.440 158.020 108.670 158.560 ;
        RECT 109.480 158.020 110.490 158.050 ;
        RECT 117.080 158.020 117.310 158.560 ;
        RECT 108.440 157.120 117.310 158.020 ;
        RECT 108.440 156.600 108.670 157.120 ;
        RECT 109.480 157.050 110.490 157.120 ;
        RECT 117.080 156.600 117.310 157.120 ;
        RECT 101.500 156.310 105.500 156.540 ;
        RECT 108.875 156.320 116.875 156.550 ;
        RECT 100.050 156.160 101.180 156.200 ;
        RECT 100.050 156.080 101.420 156.160 ;
        RECT 101.790 156.090 105.450 156.310 ;
        RECT 101.790 156.080 103.230 156.090 ;
        RECT 100.050 156.040 103.230 156.080 ;
        RECT 100.050 155.950 102.740 156.040 ;
        RECT 108.940 156.030 116.830 156.320 ;
        RECT 100.050 155.890 102.070 155.950 ;
        RECT 100.050 155.840 101.820 155.890 ;
        RECT 100.050 152.500 100.880 155.840 ;
        RECT 108.930 155.540 116.850 155.550 ;
        RECT 105.160 155.530 116.850 155.540 ;
        RECT 101.540 155.410 116.850 155.530 ;
        RECT 101.540 155.400 116.875 155.410 ;
        RECT 101.500 155.280 116.875 155.400 ;
        RECT 101.500 155.170 105.500 155.280 ;
        RECT 101.110 154.830 101.340 155.120 ;
        RECT 101.560 154.830 105.450 155.170 ;
        RECT 105.660 154.830 105.890 155.120 ;
        RECT 101.110 153.460 105.890 154.830 ;
        RECT 101.110 153.160 101.340 153.460 ;
        RECT 105.660 153.160 105.890 153.460 ;
        RECT 101.500 152.880 105.500 153.110 ;
        RECT 101.750 152.650 105.320 152.880 ;
        RECT 101.750 152.500 105.440 152.650 ;
        RECT 100.050 152.220 105.440 152.500 ;
        RECT 106.690 152.330 107.310 155.280 ;
        RECT 108.875 155.180 116.875 155.280 ;
        RECT 108.930 155.170 116.850 155.180 ;
        RECT 108.440 154.470 108.670 155.130 ;
        RECT 109.450 154.470 110.450 154.560 ;
        RECT 117.080 154.470 117.310 155.130 ;
        RECT 108.440 153.650 117.310 154.470 ;
        RECT 108.440 153.170 108.670 153.650 ;
        RECT 109.450 153.560 110.450 153.650 ;
        RECT 117.080 153.170 117.310 153.650 ;
        RECT 108.875 152.890 116.875 153.120 ;
        RECT 100.050 151.760 105.450 152.220 ;
        RECT 100.050 150.420 102.050 151.760 ;
        RECT 103.800 151.750 105.450 151.760 ;
        RECT 102.490 150.480 103.490 151.200 ;
        RECT 103.800 150.940 104.110 151.750 ;
        RECT 104.570 151.470 105.450 151.750 ;
        RECT 105.690 151.930 107.310 152.330 ;
        RECT 108.960 151.980 116.830 152.890 ;
        RECT 104.510 151.240 105.510 151.470 ;
        RECT 105.690 151.280 106.040 151.930 ;
        RECT 106.690 151.920 107.310 151.930 ;
        RECT 108.875 151.750 116.875 151.980 ;
        RECT 108.960 151.740 116.830 151.750 ;
        RECT 104.570 151.030 105.450 151.050 ;
        RECT 103.840 150.650 104.110 150.940 ;
        RECT 104.510 150.800 105.510 151.030 ;
        RECT 105.670 150.990 106.040 151.280 ;
        RECT 105.700 150.930 106.040 150.990 ;
        RECT 106.800 151.600 107.560 151.650 ;
        RECT 108.440 151.600 108.670 151.700 ;
        RECT 106.800 151.390 108.670 151.600 ;
        RECT 117.080 151.390 117.310 151.700 ;
        RECT 106.800 150.970 109.340 151.390 ;
        RECT 116.710 150.970 117.310 151.390 ;
        RECT 104.570 150.650 105.450 150.800 ;
        RECT 104.580 150.480 105.310 150.650 ;
        RECT 100.130 150.410 102.050 150.420 ;
        RECT 102.460 149.360 105.310 150.480 ;
        RECT 105.700 150.180 106.050 150.930 ;
        RECT 106.800 150.810 108.670 150.970 ;
        RECT 106.800 150.760 107.560 150.810 ;
        RECT 108.440 150.740 108.670 150.810 ;
        RECT 117.080 150.740 117.310 150.970 ;
        RECT 108.875 150.460 116.875 150.690 ;
        RECT 105.700 150.120 105.990 150.180 ;
        RECT 105.610 150.000 105.990 150.120 ;
        RECT 108.970 150.060 116.830 150.460 ;
        RECT 117.640 150.060 118.600 159.540 ;
        RECT 119.930 161.770 120.190 161.800 ;
        RECT 119.930 159.670 120.760 161.770 ;
        RECT 126.430 161.380 127.680 161.820 ;
        RECT 124.370 161.370 129.610 161.380 ;
        RECT 121.420 161.270 136.720 161.370 ;
        RECT 121.420 161.260 136.755 161.270 ;
        RECT 121.380 161.140 136.755 161.260 ;
        RECT 121.380 161.030 125.380 161.140 ;
        RECT 126.430 161.060 128.170 161.140 ;
        RECT 128.750 161.060 136.755 161.140 ;
        RECT 126.430 160.980 127.680 161.060 ;
        RECT 128.755 161.040 136.755 161.060 ;
        RECT 120.990 160.730 121.220 160.980 ;
        RECT 125.540 160.840 125.770 160.980 ;
        RECT 128.320 160.840 128.550 160.990 ;
        RECT 125.540 160.730 128.550 160.840 ;
        RECT 136.960 160.730 137.190 160.990 ;
        RECT 120.990 160.290 137.190 160.730 ;
        RECT 120.990 160.020 121.220 160.290 ;
        RECT 125.540 160.260 137.190 160.290 ;
        RECT 125.540 160.170 128.550 160.260 ;
        RECT 125.540 160.020 125.770 160.170 ;
        RECT 128.320 160.030 128.550 160.170 ;
        RECT 136.960 160.030 137.190 160.260 ;
        RECT 121.380 159.740 125.380 159.970 ;
        RECT 128.755 159.760 136.755 159.980 ;
        RECT 137.520 159.760 138.480 161.800 ;
        RECT 128.755 159.750 138.480 159.760 ;
        RECT 121.380 159.670 125.370 159.740 ;
        RECT 119.930 159.560 125.370 159.670 ;
        RECT 128.810 159.590 138.480 159.750 ;
        RECT 119.930 159.470 123.060 159.560 ;
        RECT 136.550 159.540 138.480 159.590 ;
        RECT 119.930 156.200 120.760 159.470 ;
        RECT 124.410 159.010 129.660 159.020 ;
        RECT 124.410 158.900 136.720 159.010 ;
        RECT 121.440 158.840 136.720 158.900 ;
        RECT 121.440 158.830 136.755 158.840 ;
        RECT 121.380 158.700 136.755 158.830 ;
        RECT 121.380 158.690 126.540 158.700 ;
        RECT 121.380 158.600 125.380 158.690 ;
        RECT 128.755 158.610 136.755 158.700 ;
        RECT 128.840 158.600 136.730 158.610 ;
        RECT 120.990 158.240 121.220 158.550 ;
        RECT 121.440 158.240 125.340 158.600 ;
        RECT 125.540 158.240 125.770 158.550 ;
        RECT 120.990 156.900 125.770 158.240 ;
        RECT 120.990 156.590 121.220 156.900 ;
        RECT 125.540 156.590 125.770 156.900 ;
        RECT 128.320 158.020 128.550 158.560 ;
        RECT 129.360 158.020 130.370 158.050 ;
        RECT 136.960 158.020 137.190 158.560 ;
        RECT 128.320 157.120 137.190 158.020 ;
        RECT 128.320 156.600 128.550 157.120 ;
        RECT 129.360 157.050 130.370 157.120 ;
        RECT 136.960 156.600 137.190 157.120 ;
        RECT 121.380 156.310 125.380 156.540 ;
        RECT 128.755 156.320 136.755 156.550 ;
        RECT 119.930 156.160 121.060 156.200 ;
        RECT 119.930 156.080 121.300 156.160 ;
        RECT 121.670 156.090 125.330 156.310 ;
        RECT 121.670 156.080 123.110 156.090 ;
        RECT 119.930 156.040 123.110 156.080 ;
        RECT 119.930 155.950 122.620 156.040 ;
        RECT 128.820 156.030 136.710 156.320 ;
        RECT 119.930 155.890 121.950 155.950 ;
        RECT 119.930 155.840 121.700 155.890 ;
        RECT 119.930 152.500 120.760 155.840 ;
        RECT 128.810 155.540 136.730 155.550 ;
        RECT 125.040 155.530 136.730 155.540 ;
        RECT 121.420 155.410 136.730 155.530 ;
        RECT 121.420 155.400 136.755 155.410 ;
        RECT 121.380 155.280 136.755 155.400 ;
        RECT 121.380 155.170 125.380 155.280 ;
        RECT 120.990 154.830 121.220 155.120 ;
        RECT 121.440 154.830 125.330 155.170 ;
        RECT 125.540 154.830 125.770 155.120 ;
        RECT 120.990 153.460 125.770 154.830 ;
        RECT 120.990 153.160 121.220 153.460 ;
        RECT 125.540 153.160 125.770 153.460 ;
        RECT 121.380 152.880 125.380 153.110 ;
        RECT 121.630 152.650 125.200 152.880 ;
        RECT 121.630 152.500 125.320 152.650 ;
        RECT 119.930 152.220 125.320 152.500 ;
        RECT 126.570 152.330 127.190 155.280 ;
        RECT 128.755 155.180 136.755 155.280 ;
        RECT 128.810 155.170 136.730 155.180 ;
        RECT 128.320 154.470 128.550 155.130 ;
        RECT 129.330 154.470 130.330 154.560 ;
        RECT 136.960 154.470 137.190 155.130 ;
        RECT 128.320 153.650 137.190 154.470 ;
        RECT 128.320 153.170 128.550 153.650 ;
        RECT 129.330 153.560 130.330 153.650 ;
        RECT 136.960 153.170 137.190 153.650 ;
        RECT 128.755 152.890 136.755 153.120 ;
        RECT 119.930 151.760 125.330 152.220 ;
        RECT 119.930 150.420 121.930 151.760 ;
        RECT 123.680 151.750 125.330 151.760 ;
        RECT 122.370 150.480 123.370 151.200 ;
        RECT 123.680 150.940 123.990 151.750 ;
        RECT 124.450 151.470 125.330 151.750 ;
        RECT 125.570 151.930 127.190 152.330 ;
        RECT 128.840 151.980 136.710 152.890 ;
        RECT 124.390 151.240 125.390 151.470 ;
        RECT 125.570 151.280 125.920 151.930 ;
        RECT 126.570 151.920 127.190 151.930 ;
        RECT 128.755 151.750 136.755 151.980 ;
        RECT 128.840 151.740 136.710 151.750 ;
        RECT 124.450 151.030 125.330 151.050 ;
        RECT 123.720 150.650 123.990 150.940 ;
        RECT 124.390 150.800 125.390 151.030 ;
        RECT 125.550 150.990 125.920 151.280 ;
        RECT 125.580 150.930 125.920 150.990 ;
        RECT 126.680 151.600 127.440 151.650 ;
        RECT 128.320 151.600 128.550 151.700 ;
        RECT 126.680 151.390 128.550 151.600 ;
        RECT 136.960 151.390 137.190 151.700 ;
        RECT 126.680 150.970 129.220 151.390 ;
        RECT 136.590 150.970 137.190 151.390 ;
        RECT 124.450 150.650 125.330 150.800 ;
        RECT 124.460 150.480 125.190 150.650 ;
        RECT 120.010 150.410 121.930 150.420 ;
        RECT 102.400 149.130 105.400 149.360 ;
        RECT 105.610 149.170 105.950 150.000 ;
        RECT 107.960 149.990 118.600 150.060 ;
        RECT 102.450 149.100 105.310 149.130 ;
        RECT 102.450 149.080 103.620 149.100 ;
        RECT 104.580 149.090 105.310 149.100 ;
        RECT 102.400 148.690 105.400 148.920 ;
        RECT 105.605 148.880 105.950 149.170 ;
        RECT 106.140 148.950 118.600 149.990 ;
        RECT 122.340 149.360 125.190 150.480 ;
        RECT 125.580 150.180 125.930 150.930 ;
        RECT 126.680 150.810 128.550 150.970 ;
        RECT 126.680 150.760 127.440 150.810 ;
        RECT 128.320 150.740 128.550 150.810 ;
        RECT 136.960 150.740 137.190 150.970 ;
        RECT 128.755 150.460 136.755 150.690 ;
        RECT 125.580 150.120 125.870 150.180 ;
        RECT 125.490 150.000 125.870 150.120 ;
        RECT 128.850 150.060 136.710 150.460 ;
        RECT 137.520 150.060 138.480 159.540 ;
        RECT 140.010 161.720 140.270 161.750 ;
        RECT 140.010 159.620 140.840 161.720 ;
        RECT 146.510 161.330 147.760 161.770 ;
        RECT 144.450 161.320 149.690 161.330 ;
        RECT 141.500 161.220 156.800 161.320 ;
        RECT 141.500 161.210 156.835 161.220 ;
        RECT 141.460 161.090 156.835 161.210 ;
        RECT 141.460 160.980 145.460 161.090 ;
        RECT 146.510 161.010 148.250 161.090 ;
        RECT 148.830 161.010 156.835 161.090 ;
        RECT 146.510 160.930 147.760 161.010 ;
        RECT 148.835 160.990 156.835 161.010 ;
        RECT 141.070 160.680 141.300 160.930 ;
        RECT 145.620 160.790 145.850 160.930 ;
        RECT 148.400 160.790 148.630 160.940 ;
        RECT 145.620 160.680 148.630 160.790 ;
        RECT 157.040 160.680 157.270 160.940 ;
        RECT 141.070 160.240 157.270 160.680 ;
        RECT 141.070 159.970 141.300 160.240 ;
        RECT 145.620 160.210 157.270 160.240 ;
        RECT 145.620 160.120 148.630 160.210 ;
        RECT 145.620 159.970 145.850 160.120 ;
        RECT 148.400 159.980 148.630 160.120 ;
        RECT 157.040 159.980 157.270 160.210 ;
        RECT 141.460 159.690 145.460 159.920 ;
        RECT 148.835 159.710 156.835 159.930 ;
        RECT 157.600 159.710 158.560 161.750 ;
        RECT 148.835 159.700 158.560 159.710 ;
        RECT 141.460 159.620 145.450 159.690 ;
        RECT 140.010 159.510 145.450 159.620 ;
        RECT 148.890 159.540 158.560 159.700 ;
        RECT 140.010 159.420 143.140 159.510 ;
        RECT 156.630 159.490 158.560 159.540 ;
        RECT 140.010 156.150 140.840 159.420 ;
        RECT 144.490 158.960 149.740 158.970 ;
        RECT 144.490 158.850 156.800 158.960 ;
        RECT 141.520 158.790 156.800 158.850 ;
        RECT 141.520 158.780 156.835 158.790 ;
        RECT 141.460 158.650 156.835 158.780 ;
        RECT 141.460 158.640 146.620 158.650 ;
        RECT 141.460 158.550 145.460 158.640 ;
        RECT 148.835 158.560 156.835 158.650 ;
        RECT 148.920 158.550 156.810 158.560 ;
        RECT 141.070 158.190 141.300 158.500 ;
        RECT 141.520 158.190 145.420 158.550 ;
        RECT 145.620 158.190 145.850 158.500 ;
        RECT 141.070 156.850 145.850 158.190 ;
        RECT 141.070 156.540 141.300 156.850 ;
        RECT 145.620 156.540 145.850 156.850 ;
        RECT 148.400 157.970 148.630 158.510 ;
        RECT 149.440 157.970 150.450 158.000 ;
        RECT 157.040 157.970 157.270 158.510 ;
        RECT 148.400 157.070 157.270 157.970 ;
        RECT 148.400 156.550 148.630 157.070 ;
        RECT 149.440 157.000 150.450 157.070 ;
        RECT 157.040 156.550 157.270 157.070 ;
        RECT 141.460 156.260 145.460 156.490 ;
        RECT 148.835 156.270 156.835 156.500 ;
        RECT 140.010 156.110 141.140 156.150 ;
        RECT 140.010 156.030 141.380 156.110 ;
        RECT 141.750 156.040 145.410 156.260 ;
        RECT 141.750 156.030 143.190 156.040 ;
        RECT 140.010 155.990 143.190 156.030 ;
        RECT 140.010 155.900 142.700 155.990 ;
        RECT 148.900 155.980 156.790 156.270 ;
        RECT 140.010 155.840 142.030 155.900 ;
        RECT 140.010 155.790 141.780 155.840 ;
        RECT 140.010 152.450 140.840 155.790 ;
        RECT 148.890 155.490 156.810 155.500 ;
        RECT 145.120 155.480 156.810 155.490 ;
        RECT 141.500 155.360 156.810 155.480 ;
        RECT 141.500 155.350 156.835 155.360 ;
        RECT 141.460 155.230 156.835 155.350 ;
        RECT 141.460 155.120 145.460 155.230 ;
        RECT 141.070 154.780 141.300 155.070 ;
        RECT 141.520 154.780 145.410 155.120 ;
        RECT 145.620 154.780 145.850 155.070 ;
        RECT 141.070 153.410 145.850 154.780 ;
        RECT 141.070 153.110 141.300 153.410 ;
        RECT 145.620 153.110 145.850 153.410 ;
        RECT 141.460 152.830 145.460 153.060 ;
        RECT 141.710 152.600 145.280 152.830 ;
        RECT 141.710 152.450 145.400 152.600 ;
        RECT 140.010 152.170 145.400 152.450 ;
        RECT 146.650 152.280 147.270 155.230 ;
        RECT 148.835 155.130 156.835 155.230 ;
        RECT 148.890 155.120 156.810 155.130 ;
        RECT 148.400 154.420 148.630 155.080 ;
        RECT 149.410 154.420 150.410 154.510 ;
        RECT 157.040 154.420 157.270 155.080 ;
        RECT 148.400 153.600 157.270 154.420 ;
        RECT 148.400 153.120 148.630 153.600 ;
        RECT 149.410 153.510 150.410 153.600 ;
        RECT 157.040 153.120 157.270 153.600 ;
        RECT 148.835 152.840 156.835 153.070 ;
        RECT 140.010 151.710 145.410 152.170 ;
        RECT 140.010 150.370 142.010 151.710 ;
        RECT 143.760 151.700 145.410 151.710 ;
        RECT 142.450 150.430 143.450 151.150 ;
        RECT 143.760 150.890 144.070 151.700 ;
        RECT 144.530 151.420 145.410 151.700 ;
        RECT 145.650 151.880 147.270 152.280 ;
        RECT 148.920 151.930 156.790 152.840 ;
        RECT 144.470 151.190 145.470 151.420 ;
        RECT 145.650 151.230 146.000 151.880 ;
        RECT 146.650 151.870 147.270 151.880 ;
        RECT 148.835 151.700 156.835 151.930 ;
        RECT 148.920 151.690 156.790 151.700 ;
        RECT 144.530 150.980 145.410 151.000 ;
        RECT 143.800 150.600 144.070 150.890 ;
        RECT 144.470 150.750 145.470 150.980 ;
        RECT 145.630 150.940 146.000 151.230 ;
        RECT 145.660 150.880 146.000 150.940 ;
        RECT 146.760 151.550 147.520 151.600 ;
        RECT 148.400 151.550 148.630 151.650 ;
        RECT 146.760 151.340 148.630 151.550 ;
        RECT 157.040 151.340 157.270 151.650 ;
        RECT 146.760 150.920 149.300 151.340 ;
        RECT 156.670 150.920 157.270 151.340 ;
        RECT 144.530 150.600 145.410 150.750 ;
        RECT 144.540 150.430 145.270 150.600 ;
        RECT 140.090 150.360 142.010 150.370 ;
        RECT 122.280 149.130 125.280 149.360 ;
        RECT 125.490 149.170 125.830 150.000 ;
        RECT 127.840 149.990 138.480 150.060 ;
        RECT 122.330 149.100 125.190 149.130 ;
        RECT 122.330 149.080 123.500 149.100 ;
        RECT 124.460 149.090 125.190 149.100 ;
        RECT 106.140 148.930 118.470 148.950 ;
        RECT 106.410 148.920 111.850 148.930 ;
        RECT 112.850 148.920 118.470 148.930 ;
        RECT 105.610 148.770 105.950 148.880 ;
        RECT 122.280 148.690 125.280 148.920 ;
        RECT 125.485 148.880 125.830 149.170 ;
        RECT 126.020 148.950 138.480 149.990 ;
        RECT 142.420 149.310 145.270 150.430 ;
        RECT 145.660 150.130 146.010 150.880 ;
        RECT 146.760 150.760 148.630 150.920 ;
        RECT 146.760 150.710 147.520 150.760 ;
        RECT 148.400 150.690 148.630 150.760 ;
        RECT 157.040 150.690 157.270 150.920 ;
        RECT 148.835 150.410 156.835 150.640 ;
        RECT 145.660 150.070 145.950 150.130 ;
        RECT 145.570 149.950 145.950 150.070 ;
        RECT 148.930 150.010 156.790 150.410 ;
        RECT 157.600 150.010 158.560 159.490 ;
        RECT 142.360 149.080 145.360 149.310 ;
        RECT 145.570 149.120 145.910 149.950 ;
        RECT 147.920 149.940 158.560 150.010 ;
        RECT 142.410 149.050 145.270 149.080 ;
        RECT 142.410 149.030 143.580 149.050 ;
        RECT 144.540 149.040 145.270 149.050 ;
        RECT 126.020 148.930 138.350 148.950 ;
        RECT 126.290 148.920 131.730 148.930 ;
        RECT 132.730 148.920 138.350 148.930 ;
        RECT 125.490 148.770 125.830 148.880 ;
        RECT 142.360 148.640 145.360 148.870 ;
        RECT 145.565 148.830 145.910 149.120 ;
        RECT 146.100 148.900 158.560 149.940 ;
        RECT 146.100 148.880 158.430 148.900 ;
        RECT 146.370 148.870 151.810 148.880 ;
        RECT 152.810 148.870 158.430 148.880 ;
        RECT 145.570 148.720 145.910 148.830 ;
        RECT 100.050 146.720 100.310 146.750 ;
        RECT 100.050 144.620 100.880 146.720 ;
        RECT 106.550 146.330 107.800 146.770 ;
        RECT 104.490 146.320 109.730 146.330 ;
        RECT 101.540 146.220 116.840 146.320 ;
        RECT 101.540 146.210 116.875 146.220 ;
        RECT 101.500 146.090 116.875 146.210 ;
        RECT 101.500 145.980 105.500 146.090 ;
        RECT 106.550 146.010 108.290 146.090 ;
        RECT 108.870 146.010 116.875 146.090 ;
        RECT 106.550 145.930 107.800 146.010 ;
        RECT 108.875 145.990 116.875 146.010 ;
        RECT 101.110 145.680 101.340 145.930 ;
        RECT 105.660 145.790 105.890 145.930 ;
        RECT 108.440 145.790 108.670 145.940 ;
        RECT 105.660 145.680 108.670 145.790 ;
        RECT 117.080 145.680 117.310 145.940 ;
        RECT 101.110 145.240 117.310 145.680 ;
        RECT 101.110 144.970 101.340 145.240 ;
        RECT 105.660 145.210 117.310 145.240 ;
        RECT 105.660 145.120 108.670 145.210 ;
        RECT 105.660 144.970 105.890 145.120 ;
        RECT 108.440 144.980 108.670 145.120 ;
        RECT 117.080 144.980 117.310 145.210 ;
        RECT 101.500 144.690 105.500 144.920 ;
        RECT 108.875 144.710 116.875 144.930 ;
        RECT 117.640 144.710 118.600 146.750 ;
        RECT 108.875 144.700 118.600 144.710 ;
        RECT 101.500 144.620 105.490 144.690 ;
        RECT 100.050 144.510 105.490 144.620 ;
        RECT 108.930 144.540 118.600 144.700 ;
        RECT 100.050 144.420 103.180 144.510 ;
        RECT 116.670 144.490 118.600 144.540 ;
        RECT 100.050 141.150 100.880 144.420 ;
        RECT 104.530 143.960 109.780 143.970 ;
        RECT 104.530 143.850 116.840 143.960 ;
        RECT 101.560 143.790 116.840 143.850 ;
        RECT 101.560 143.780 116.875 143.790 ;
        RECT 101.500 143.650 116.875 143.780 ;
        RECT 101.500 143.640 106.660 143.650 ;
        RECT 101.500 143.550 105.500 143.640 ;
        RECT 108.875 143.560 116.875 143.650 ;
        RECT 108.960 143.550 116.850 143.560 ;
        RECT 101.110 143.190 101.340 143.500 ;
        RECT 101.560 143.190 105.460 143.550 ;
        RECT 105.660 143.190 105.890 143.500 ;
        RECT 101.110 141.850 105.890 143.190 ;
        RECT 101.110 141.540 101.340 141.850 ;
        RECT 105.660 141.540 105.890 141.850 ;
        RECT 108.440 142.970 108.670 143.510 ;
        RECT 109.480 142.970 110.490 143.000 ;
        RECT 117.080 142.970 117.310 143.510 ;
        RECT 108.440 142.070 117.310 142.970 ;
        RECT 108.440 141.550 108.670 142.070 ;
        RECT 109.480 142.000 110.490 142.070 ;
        RECT 117.080 141.550 117.310 142.070 ;
        RECT 101.500 141.260 105.500 141.490 ;
        RECT 108.875 141.270 116.875 141.500 ;
        RECT 100.050 141.110 101.180 141.150 ;
        RECT 100.050 141.030 101.420 141.110 ;
        RECT 101.790 141.040 105.450 141.260 ;
        RECT 101.790 141.030 103.230 141.040 ;
        RECT 100.050 140.990 103.230 141.030 ;
        RECT 100.050 140.900 102.740 140.990 ;
        RECT 108.940 140.980 116.830 141.270 ;
        RECT 100.050 140.840 102.070 140.900 ;
        RECT 100.050 140.790 101.820 140.840 ;
        RECT 100.050 137.450 100.880 140.790 ;
        RECT 108.930 140.490 116.850 140.500 ;
        RECT 105.160 140.480 116.850 140.490 ;
        RECT 101.540 140.360 116.850 140.480 ;
        RECT 101.540 140.350 116.875 140.360 ;
        RECT 101.500 140.230 116.875 140.350 ;
        RECT 101.500 140.120 105.500 140.230 ;
        RECT 101.110 139.780 101.340 140.070 ;
        RECT 101.560 139.780 105.450 140.120 ;
        RECT 105.660 139.780 105.890 140.070 ;
        RECT 101.110 138.410 105.890 139.780 ;
        RECT 101.110 138.110 101.340 138.410 ;
        RECT 105.660 138.110 105.890 138.410 ;
        RECT 101.500 137.830 105.500 138.060 ;
        RECT 101.750 137.600 105.320 137.830 ;
        RECT 101.750 137.450 105.440 137.600 ;
        RECT 100.050 137.170 105.440 137.450 ;
        RECT 106.690 137.280 107.310 140.230 ;
        RECT 108.875 140.130 116.875 140.230 ;
        RECT 108.930 140.120 116.850 140.130 ;
        RECT 108.440 139.420 108.670 140.080 ;
        RECT 109.450 139.420 110.450 139.510 ;
        RECT 117.080 139.420 117.310 140.080 ;
        RECT 108.440 138.600 117.310 139.420 ;
        RECT 108.440 138.120 108.670 138.600 ;
        RECT 109.450 138.510 110.450 138.600 ;
        RECT 117.080 138.120 117.310 138.600 ;
        RECT 108.875 137.840 116.875 138.070 ;
        RECT 100.050 136.710 105.450 137.170 ;
        RECT 100.050 135.370 102.050 136.710 ;
        RECT 103.800 136.700 105.450 136.710 ;
        RECT 102.490 135.430 103.490 136.150 ;
        RECT 103.800 135.890 104.110 136.700 ;
        RECT 104.570 136.420 105.450 136.700 ;
        RECT 105.690 136.880 107.310 137.280 ;
        RECT 108.960 136.930 116.830 137.840 ;
        RECT 104.510 136.190 105.510 136.420 ;
        RECT 105.690 136.230 106.040 136.880 ;
        RECT 106.690 136.870 107.310 136.880 ;
        RECT 108.875 136.700 116.875 136.930 ;
        RECT 108.960 136.690 116.830 136.700 ;
        RECT 104.570 135.980 105.450 136.000 ;
        RECT 103.840 135.600 104.110 135.890 ;
        RECT 104.510 135.750 105.510 135.980 ;
        RECT 105.670 135.940 106.040 136.230 ;
        RECT 105.700 135.880 106.040 135.940 ;
        RECT 106.800 136.550 107.560 136.600 ;
        RECT 108.440 136.550 108.670 136.650 ;
        RECT 106.800 136.340 108.670 136.550 ;
        RECT 117.080 136.340 117.310 136.650 ;
        RECT 106.800 135.920 109.340 136.340 ;
        RECT 116.710 135.920 117.310 136.340 ;
        RECT 104.570 135.600 105.450 135.750 ;
        RECT 104.580 135.430 105.310 135.600 ;
        RECT 100.130 135.360 102.050 135.370 ;
        RECT 102.460 134.310 105.310 135.430 ;
        RECT 105.700 135.130 106.050 135.880 ;
        RECT 106.800 135.760 108.670 135.920 ;
        RECT 106.800 135.710 107.560 135.760 ;
        RECT 108.440 135.690 108.670 135.760 ;
        RECT 117.080 135.690 117.310 135.920 ;
        RECT 108.875 135.410 116.875 135.640 ;
        RECT 105.700 135.070 105.990 135.130 ;
        RECT 105.610 134.950 105.990 135.070 ;
        RECT 108.970 135.010 116.830 135.410 ;
        RECT 117.640 135.010 118.600 144.490 ;
        RECT 119.930 146.720 120.190 146.750 ;
        RECT 119.930 144.620 120.760 146.720 ;
        RECT 126.430 146.330 127.680 146.770 ;
        RECT 124.370 146.320 129.610 146.330 ;
        RECT 121.420 146.220 136.720 146.320 ;
        RECT 121.420 146.210 136.755 146.220 ;
        RECT 121.380 146.090 136.755 146.210 ;
        RECT 121.380 145.980 125.380 146.090 ;
        RECT 126.430 146.010 128.170 146.090 ;
        RECT 128.750 146.010 136.755 146.090 ;
        RECT 126.430 145.930 127.680 146.010 ;
        RECT 128.755 145.990 136.755 146.010 ;
        RECT 120.990 145.680 121.220 145.930 ;
        RECT 125.540 145.790 125.770 145.930 ;
        RECT 128.320 145.790 128.550 145.940 ;
        RECT 125.540 145.680 128.550 145.790 ;
        RECT 136.960 145.680 137.190 145.940 ;
        RECT 120.990 145.240 137.190 145.680 ;
        RECT 120.990 144.970 121.220 145.240 ;
        RECT 125.540 145.210 137.190 145.240 ;
        RECT 125.540 145.120 128.550 145.210 ;
        RECT 125.540 144.970 125.770 145.120 ;
        RECT 128.320 144.980 128.550 145.120 ;
        RECT 136.960 144.980 137.190 145.210 ;
        RECT 121.380 144.690 125.380 144.920 ;
        RECT 128.755 144.710 136.755 144.930 ;
        RECT 137.520 144.710 138.480 146.750 ;
        RECT 128.755 144.700 138.480 144.710 ;
        RECT 121.380 144.620 125.370 144.690 ;
        RECT 119.930 144.510 125.370 144.620 ;
        RECT 128.810 144.540 138.480 144.700 ;
        RECT 119.930 144.420 123.060 144.510 ;
        RECT 136.550 144.490 138.480 144.540 ;
        RECT 119.930 141.150 120.760 144.420 ;
        RECT 124.410 143.960 129.660 143.970 ;
        RECT 124.410 143.850 136.720 143.960 ;
        RECT 121.440 143.790 136.720 143.850 ;
        RECT 121.440 143.780 136.755 143.790 ;
        RECT 121.380 143.650 136.755 143.780 ;
        RECT 121.380 143.640 126.540 143.650 ;
        RECT 121.380 143.550 125.380 143.640 ;
        RECT 128.755 143.560 136.755 143.650 ;
        RECT 128.840 143.550 136.730 143.560 ;
        RECT 120.990 143.190 121.220 143.500 ;
        RECT 121.440 143.190 125.340 143.550 ;
        RECT 125.540 143.190 125.770 143.500 ;
        RECT 120.990 141.850 125.770 143.190 ;
        RECT 120.990 141.540 121.220 141.850 ;
        RECT 125.540 141.540 125.770 141.850 ;
        RECT 128.320 142.970 128.550 143.510 ;
        RECT 129.360 142.970 130.370 143.000 ;
        RECT 136.960 142.970 137.190 143.510 ;
        RECT 128.320 142.070 137.190 142.970 ;
        RECT 128.320 141.550 128.550 142.070 ;
        RECT 129.360 142.000 130.370 142.070 ;
        RECT 136.960 141.550 137.190 142.070 ;
        RECT 121.380 141.260 125.380 141.490 ;
        RECT 128.755 141.270 136.755 141.500 ;
        RECT 119.930 141.110 121.060 141.150 ;
        RECT 119.930 141.030 121.300 141.110 ;
        RECT 121.670 141.040 125.330 141.260 ;
        RECT 121.670 141.030 123.110 141.040 ;
        RECT 119.930 140.990 123.110 141.030 ;
        RECT 119.930 140.900 122.620 140.990 ;
        RECT 128.820 140.980 136.710 141.270 ;
        RECT 119.930 140.840 121.950 140.900 ;
        RECT 119.930 140.790 121.700 140.840 ;
        RECT 119.930 137.450 120.760 140.790 ;
        RECT 128.810 140.490 136.730 140.500 ;
        RECT 125.040 140.480 136.730 140.490 ;
        RECT 121.420 140.360 136.730 140.480 ;
        RECT 121.420 140.350 136.755 140.360 ;
        RECT 121.380 140.230 136.755 140.350 ;
        RECT 121.380 140.120 125.380 140.230 ;
        RECT 120.990 139.780 121.220 140.070 ;
        RECT 121.440 139.780 125.330 140.120 ;
        RECT 125.540 139.780 125.770 140.070 ;
        RECT 120.990 138.410 125.770 139.780 ;
        RECT 120.990 138.110 121.220 138.410 ;
        RECT 125.540 138.110 125.770 138.410 ;
        RECT 121.380 137.830 125.380 138.060 ;
        RECT 121.630 137.600 125.200 137.830 ;
        RECT 121.630 137.450 125.320 137.600 ;
        RECT 119.930 137.170 125.320 137.450 ;
        RECT 126.570 137.280 127.190 140.230 ;
        RECT 128.755 140.130 136.755 140.230 ;
        RECT 128.810 140.120 136.730 140.130 ;
        RECT 128.320 139.420 128.550 140.080 ;
        RECT 129.330 139.420 130.330 139.510 ;
        RECT 136.960 139.420 137.190 140.080 ;
        RECT 128.320 138.600 137.190 139.420 ;
        RECT 128.320 138.120 128.550 138.600 ;
        RECT 129.330 138.510 130.330 138.600 ;
        RECT 136.960 138.120 137.190 138.600 ;
        RECT 128.755 137.840 136.755 138.070 ;
        RECT 119.930 136.710 125.330 137.170 ;
        RECT 119.930 135.370 121.930 136.710 ;
        RECT 123.680 136.700 125.330 136.710 ;
        RECT 122.370 135.430 123.370 136.150 ;
        RECT 123.680 135.890 123.990 136.700 ;
        RECT 124.450 136.420 125.330 136.700 ;
        RECT 125.570 136.880 127.190 137.280 ;
        RECT 128.840 136.930 136.710 137.840 ;
        RECT 124.390 136.190 125.390 136.420 ;
        RECT 125.570 136.230 125.920 136.880 ;
        RECT 126.570 136.870 127.190 136.880 ;
        RECT 128.755 136.700 136.755 136.930 ;
        RECT 128.840 136.690 136.710 136.700 ;
        RECT 124.450 135.980 125.330 136.000 ;
        RECT 123.720 135.600 123.990 135.890 ;
        RECT 124.390 135.750 125.390 135.980 ;
        RECT 125.550 135.940 125.920 136.230 ;
        RECT 125.580 135.880 125.920 135.940 ;
        RECT 126.680 136.550 127.440 136.600 ;
        RECT 128.320 136.550 128.550 136.650 ;
        RECT 126.680 136.340 128.550 136.550 ;
        RECT 136.960 136.340 137.190 136.650 ;
        RECT 126.680 135.920 129.220 136.340 ;
        RECT 136.590 135.920 137.190 136.340 ;
        RECT 124.450 135.600 125.330 135.750 ;
        RECT 124.460 135.430 125.190 135.600 ;
        RECT 120.010 135.360 121.930 135.370 ;
        RECT 102.400 134.080 105.400 134.310 ;
        RECT 105.610 134.120 105.950 134.950 ;
        RECT 107.960 134.940 118.600 135.010 ;
        RECT 102.450 134.050 105.310 134.080 ;
        RECT 102.450 134.030 103.620 134.050 ;
        RECT 104.580 134.040 105.310 134.050 ;
        RECT 102.400 133.640 105.400 133.870 ;
        RECT 105.605 133.830 105.950 134.120 ;
        RECT 106.140 133.900 118.600 134.940 ;
        RECT 122.340 134.310 125.190 135.430 ;
        RECT 125.580 135.130 125.930 135.880 ;
        RECT 126.680 135.760 128.550 135.920 ;
        RECT 126.680 135.710 127.440 135.760 ;
        RECT 128.320 135.690 128.550 135.760 ;
        RECT 136.960 135.690 137.190 135.920 ;
        RECT 128.755 135.410 136.755 135.640 ;
        RECT 125.580 135.070 125.870 135.130 ;
        RECT 125.490 134.950 125.870 135.070 ;
        RECT 128.850 135.010 136.710 135.410 ;
        RECT 137.520 135.010 138.480 144.490 ;
        RECT 139.960 146.720 140.220 146.750 ;
        RECT 139.960 144.620 140.790 146.720 ;
        RECT 146.460 146.330 147.710 146.770 ;
        RECT 144.400 146.320 149.640 146.330 ;
        RECT 141.450 146.220 156.750 146.320 ;
        RECT 141.450 146.210 156.785 146.220 ;
        RECT 141.410 146.090 156.785 146.210 ;
        RECT 141.410 145.980 145.410 146.090 ;
        RECT 146.460 146.010 148.200 146.090 ;
        RECT 148.780 146.010 156.785 146.090 ;
        RECT 146.460 145.930 147.710 146.010 ;
        RECT 148.785 145.990 156.785 146.010 ;
        RECT 141.020 145.680 141.250 145.930 ;
        RECT 145.570 145.790 145.800 145.930 ;
        RECT 148.350 145.790 148.580 145.940 ;
        RECT 145.570 145.680 148.580 145.790 ;
        RECT 156.990 145.680 157.220 145.940 ;
        RECT 141.020 145.240 157.220 145.680 ;
        RECT 141.020 144.970 141.250 145.240 ;
        RECT 145.570 145.210 157.220 145.240 ;
        RECT 145.570 145.120 148.580 145.210 ;
        RECT 145.570 144.970 145.800 145.120 ;
        RECT 148.350 144.980 148.580 145.120 ;
        RECT 156.990 144.980 157.220 145.210 ;
        RECT 141.410 144.690 145.410 144.920 ;
        RECT 148.785 144.710 156.785 144.930 ;
        RECT 157.550 144.710 158.510 146.750 ;
        RECT 148.785 144.700 158.510 144.710 ;
        RECT 141.410 144.620 145.400 144.690 ;
        RECT 139.960 144.510 145.400 144.620 ;
        RECT 148.840 144.540 158.510 144.700 ;
        RECT 139.960 144.420 143.090 144.510 ;
        RECT 156.580 144.490 158.510 144.540 ;
        RECT 139.960 141.150 140.790 144.420 ;
        RECT 144.440 143.960 149.690 143.970 ;
        RECT 144.440 143.850 156.750 143.960 ;
        RECT 141.470 143.790 156.750 143.850 ;
        RECT 141.470 143.780 156.785 143.790 ;
        RECT 141.410 143.650 156.785 143.780 ;
        RECT 141.410 143.640 146.570 143.650 ;
        RECT 141.410 143.550 145.410 143.640 ;
        RECT 148.785 143.560 156.785 143.650 ;
        RECT 148.870 143.550 156.760 143.560 ;
        RECT 141.020 143.190 141.250 143.500 ;
        RECT 141.470 143.190 145.370 143.550 ;
        RECT 145.570 143.190 145.800 143.500 ;
        RECT 141.020 141.850 145.800 143.190 ;
        RECT 141.020 141.540 141.250 141.850 ;
        RECT 145.570 141.540 145.800 141.850 ;
        RECT 148.350 142.970 148.580 143.510 ;
        RECT 149.390 142.970 150.400 143.000 ;
        RECT 156.990 142.970 157.220 143.510 ;
        RECT 148.350 142.070 157.220 142.970 ;
        RECT 148.350 141.550 148.580 142.070 ;
        RECT 149.390 142.000 150.400 142.070 ;
        RECT 156.990 141.550 157.220 142.070 ;
        RECT 141.410 141.260 145.410 141.490 ;
        RECT 148.785 141.270 156.785 141.500 ;
        RECT 139.960 141.110 141.090 141.150 ;
        RECT 139.960 141.030 141.330 141.110 ;
        RECT 141.700 141.040 145.360 141.260 ;
        RECT 141.700 141.030 143.140 141.040 ;
        RECT 139.960 140.990 143.140 141.030 ;
        RECT 139.960 140.900 142.650 140.990 ;
        RECT 148.850 140.980 156.740 141.270 ;
        RECT 139.960 140.840 141.980 140.900 ;
        RECT 139.960 140.790 141.730 140.840 ;
        RECT 139.960 137.450 140.790 140.790 ;
        RECT 148.840 140.490 156.760 140.500 ;
        RECT 145.070 140.480 156.760 140.490 ;
        RECT 141.450 140.360 156.760 140.480 ;
        RECT 141.450 140.350 156.785 140.360 ;
        RECT 141.410 140.230 156.785 140.350 ;
        RECT 141.410 140.120 145.410 140.230 ;
        RECT 141.020 139.780 141.250 140.070 ;
        RECT 141.470 139.780 145.360 140.120 ;
        RECT 145.570 139.780 145.800 140.070 ;
        RECT 141.020 138.410 145.800 139.780 ;
        RECT 141.020 138.110 141.250 138.410 ;
        RECT 145.570 138.110 145.800 138.410 ;
        RECT 141.410 137.830 145.410 138.060 ;
        RECT 141.660 137.600 145.230 137.830 ;
        RECT 141.660 137.450 145.350 137.600 ;
        RECT 139.960 137.170 145.350 137.450 ;
        RECT 146.600 137.280 147.220 140.230 ;
        RECT 148.785 140.130 156.785 140.230 ;
        RECT 148.840 140.120 156.760 140.130 ;
        RECT 148.350 139.420 148.580 140.080 ;
        RECT 149.360 139.420 150.360 139.510 ;
        RECT 156.990 139.420 157.220 140.080 ;
        RECT 148.350 138.600 157.220 139.420 ;
        RECT 148.350 138.120 148.580 138.600 ;
        RECT 149.360 138.510 150.360 138.600 ;
        RECT 156.990 138.120 157.220 138.600 ;
        RECT 148.785 137.840 156.785 138.070 ;
        RECT 139.960 136.710 145.360 137.170 ;
        RECT 139.960 135.370 141.960 136.710 ;
        RECT 143.710 136.700 145.360 136.710 ;
        RECT 142.400 135.430 143.400 136.150 ;
        RECT 143.710 135.890 144.020 136.700 ;
        RECT 144.480 136.420 145.360 136.700 ;
        RECT 145.600 136.880 147.220 137.280 ;
        RECT 148.870 136.930 156.740 137.840 ;
        RECT 144.420 136.190 145.420 136.420 ;
        RECT 145.600 136.230 145.950 136.880 ;
        RECT 146.600 136.870 147.220 136.880 ;
        RECT 148.785 136.700 156.785 136.930 ;
        RECT 148.870 136.690 156.740 136.700 ;
        RECT 144.480 135.980 145.360 136.000 ;
        RECT 143.750 135.600 144.020 135.890 ;
        RECT 144.420 135.750 145.420 135.980 ;
        RECT 145.580 135.940 145.950 136.230 ;
        RECT 145.610 135.880 145.950 135.940 ;
        RECT 146.710 136.550 147.470 136.600 ;
        RECT 148.350 136.550 148.580 136.650 ;
        RECT 146.710 136.340 148.580 136.550 ;
        RECT 156.990 136.340 157.220 136.650 ;
        RECT 146.710 135.920 149.250 136.340 ;
        RECT 156.620 135.920 157.220 136.340 ;
        RECT 144.480 135.600 145.360 135.750 ;
        RECT 144.490 135.430 145.220 135.600 ;
        RECT 140.040 135.360 141.960 135.370 ;
        RECT 122.280 134.080 125.280 134.310 ;
        RECT 125.490 134.120 125.830 134.950 ;
        RECT 127.840 134.940 138.480 135.010 ;
        RECT 122.330 134.050 125.190 134.080 ;
        RECT 122.330 134.030 123.500 134.050 ;
        RECT 124.460 134.040 125.190 134.050 ;
        RECT 106.140 133.880 118.470 133.900 ;
        RECT 106.410 133.870 111.850 133.880 ;
        RECT 112.850 133.870 118.470 133.880 ;
        RECT 105.610 133.720 105.950 133.830 ;
        RECT 122.280 133.640 125.280 133.870 ;
        RECT 125.485 133.830 125.830 134.120 ;
        RECT 126.020 133.900 138.480 134.940 ;
        RECT 142.370 134.310 145.220 135.430 ;
        RECT 145.610 135.130 145.960 135.880 ;
        RECT 146.710 135.760 148.580 135.920 ;
        RECT 146.710 135.710 147.470 135.760 ;
        RECT 148.350 135.690 148.580 135.760 ;
        RECT 156.990 135.690 157.220 135.920 ;
        RECT 148.785 135.410 156.785 135.640 ;
        RECT 145.610 135.070 145.900 135.130 ;
        RECT 145.520 134.950 145.900 135.070 ;
        RECT 148.880 135.010 156.740 135.410 ;
        RECT 157.550 135.010 158.510 144.490 ;
        RECT 142.310 134.080 145.310 134.310 ;
        RECT 145.520 134.120 145.860 134.950 ;
        RECT 147.870 134.940 158.510 135.010 ;
        RECT 142.360 134.050 145.220 134.080 ;
        RECT 142.360 134.030 143.530 134.050 ;
        RECT 144.490 134.040 145.220 134.050 ;
        RECT 126.020 133.880 138.350 133.900 ;
        RECT 126.290 133.870 131.730 133.880 ;
        RECT 132.730 133.870 138.350 133.880 ;
        RECT 125.490 133.720 125.830 133.830 ;
        RECT 142.310 133.640 145.310 133.870 ;
        RECT 145.515 133.830 145.860 134.120 ;
        RECT 146.050 133.900 158.510 134.940 ;
        RECT 146.050 133.880 158.380 133.900 ;
        RECT 146.320 133.870 151.760 133.880 ;
        RECT 152.760 133.870 158.380 133.880 ;
        RECT 145.520 133.720 145.860 133.830 ;
        RECT 119.930 131.780 120.190 131.810 ;
        RECT 100.050 131.720 100.310 131.750 ;
        RECT 100.050 129.620 100.880 131.720 ;
        RECT 106.550 131.330 107.800 131.770 ;
        RECT 104.490 131.320 109.730 131.330 ;
        RECT 101.540 131.220 116.840 131.320 ;
        RECT 101.540 131.210 116.875 131.220 ;
        RECT 101.500 131.090 116.875 131.210 ;
        RECT 101.500 130.980 105.500 131.090 ;
        RECT 106.550 131.010 108.290 131.090 ;
        RECT 108.870 131.010 116.875 131.090 ;
        RECT 106.550 130.930 107.800 131.010 ;
        RECT 108.875 130.990 116.875 131.010 ;
        RECT 101.110 130.680 101.340 130.930 ;
        RECT 105.660 130.790 105.890 130.930 ;
        RECT 108.440 130.790 108.670 130.940 ;
        RECT 105.660 130.680 108.670 130.790 ;
        RECT 117.080 130.680 117.310 130.940 ;
        RECT 101.110 130.240 117.310 130.680 ;
        RECT 101.110 129.970 101.340 130.240 ;
        RECT 105.660 130.210 117.310 130.240 ;
        RECT 105.660 130.120 108.670 130.210 ;
        RECT 105.660 129.970 105.890 130.120 ;
        RECT 108.440 129.980 108.670 130.120 ;
        RECT 117.080 129.980 117.310 130.210 ;
        RECT 101.500 129.690 105.500 129.920 ;
        RECT 108.875 129.710 116.875 129.930 ;
        RECT 117.640 129.710 118.600 131.750 ;
        RECT 108.875 129.700 118.600 129.710 ;
        RECT 101.500 129.620 105.490 129.690 ;
        RECT 100.050 129.510 105.490 129.620 ;
        RECT 108.930 129.540 118.600 129.700 ;
        RECT 100.050 129.420 103.180 129.510 ;
        RECT 116.670 129.490 118.600 129.540 ;
        RECT 100.050 126.150 100.880 129.420 ;
        RECT 104.530 128.960 109.780 128.970 ;
        RECT 104.530 128.850 116.840 128.960 ;
        RECT 101.560 128.790 116.840 128.850 ;
        RECT 101.560 128.780 116.875 128.790 ;
        RECT 101.500 128.650 116.875 128.780 ;
        RECT 101.500 128.640 106.660 128.650 ;
        RECT 101.500 128.550 105.500 128.640 ;
        RECT 108.875 128.560 116.875 128.650 ;
        RECT 108.960 128.550 116.850 128.560 ;
        RECT 101.110 128.190 101.340 128.500 ;
        RECT 101.560 128.190 105.460 128.550 ;
        RECT 105.660 128.190 105.890 128.500 ;
        RECT 101.110 126.850 105.890 128.190 ;
        RECT 101.110 126.540 101.340 126.850 ;
        RECT 105.660 126.540 105.890 126.850 ;
        RECT 108.440 127.970 108.670 128.510 ;
        RECT 109.480 127.970 110.490 128.000 ;
        RECT 117.080 127.970 117.310 128.510 ;
        RECT 108.440 127.070 117.310 127.970 ;
        RECT 108.440 126.550 108.670 127.070 ;
        RECT 109.480 127.000 110.490 127.070 ;
        RECT 117.080 126.550 117.310 127.070 ;
        RECT 101.500 126.260 105.500 126.490 ;
        RECT 108.875 126.270 116.875 126.500 ;
        RECT 100.050 126.110 101.180 126.150 ;
        RECT 100.050 126.030 101.420 126.110 ;
        RECT 101.790 126.040 105.450 126.260 ;
        RECT 101.790 126.030 103.230 126.040 ;
        RECT 100.050 125.990 103.230 126.030 ;
        RECT 100.050 125.900 102.740 125.990 ;
        RECT 108.940 125.980 116.830 126.270 ;
        RECT 100.050 125.840 102.070 125.900 ;
        RECT 100.050 125.790 101.820 125.840 ;
        RECT 100.050 122.450 100.880 125.790 ;
        RECT 108.930 125.490 116.850 125.500 ;
        RECT 105.160 125.480 116.850 125.490 ;
        RECT 101.540 125.360 116.850 125.480 ;
        RECT 101.540 125.350 116.875 125.360 ;
        RECT 101.500 125.230 116.875 125.350 ;
        RECT 101.500 125.120 105.500 125.230 ;
        RECT 101.110 124.780 101.340 125.070 ;
        RECT 101.560 124.780 105.450 125.120 ;
        RECT 105.660 124.780 105.890 125.070 ;
        RECT 101.110 123.410 105.890 124.780 ;
        RECT 101.110 123.110 101.340 123.410 ;
        RECT 105.660 123.110 105.890 123.410 ;
        RECT 101.500 122.830 105.500 123.060 ;
        RECT 101.750 122.600 105.320 122.830 ;
        RECT 101.750 122.450 105.440 122.600 ;
        RECT 100.050 122.170 105.440 122.450 ;
        RECT 106.690 122.280 107.310 125.230 ;
        RECT 108.875 125.130 116.875 125.230 ;
        RECT 108.930 125.120 116.850 125.130 ;
        RECT 108.440 124.420 108.670 125.080 ;
        RECT 109.450 124.420 110.450 124.510 ;
        RECT 117.080 124.420 117.310 125.080 ;
        RECT 108.440 123.600 117.310 124.420 ;
        RECT 108.440 123.120 108.670 123.600 ;
        RECT 109.450 123.510 110.450 123.600 ;
        RECT 117.080 123.120 117.310 123.600 ;
        RECT 108.875 122.840 116.875 123.070 ;
        RECT 100.050 121.710 105.450 122.170 ;
        RECT 100.050 120.370 102.050 121.710 ;
        RECT 103.800 121.700 105.450 121.710 ;
        RECT 102.490 120.430 103.490 121.150 ;
        RECT 103.800 120.890 104.110 121.700 ;
        RECT 104.570 121.420 105.450 121.700 ;
        RECT 105.690 121.880 107.310 122.280 ;
        RECT 108.960 121.930 116.830 122.840 ;
        RECT 104.510 121.190 105.510 121.420 ;
        RECT 105.690 121.230 106.040 121.880 ;
        RECT 106.690 121.870 107.310 121.880 ;
        RECT 108.875 121.700 116.875 121.930 ;
        RECT 108.960 121.690 116.830 121.700 ;
        RECT 104.570 120.980 105.450 121.000 ;
        RECT 103.840 120.600 104.110 120.890 ;
        RECT 104.510 120.750 105.510 120.980 ;
        RECT 105.670 120.940 106.040 121.230 ;
        RECT 105.700 120.880 106.040 120.940 ;
        RECT 106.800 121.550 107.560 121.600 ;
        RECT 108.440 121.550 108.670 121.650 ;
        RECT 106.800 121.340 108.670 121.550 ;
        RECT 117.080 121.340 117.310 121.650 ;
        RECT 106.800 120.920 109.340 121.340 ;
        RECT 116.710 120.920 117.310 121.340 ;
        RECT 104.570 120.600 105.450 120.750 ;
        RECT 104.580 120.430 105.310 120.600 ;
        RECT 100.130 120.360 102.050 120.370 ;
        RECT 102.460 119.310 105.310 120.430 ;
        RECT 105.700 120.130 106.050 120.880 ;
        RECT 106.800 120.760 108.670 120.920 ;
        RECT 106.800 120.710 107.560 120.760 ;
        RECT 108.440 120.690 108.670 120.760 ;
        RECT 117.080 120.690 117.310 120.920 ;
        RECT 108.875 120.410 116.875 120.640 ;
        RECT 105.700 120.070 105.990 120.130 ;
        RECT 105.610 119.950 105.990 120.070 ;
        RECT 108.970 120.010 116.830 120.410 ;
        RECT 117.640 120.010 118.600 129.490 ;
        RECT 119.930 129.680 120.760 131.780 ;
        RECT 126.430 131.390 127.680 131.830 ;
        RECT 124.370 131.380 129.610 131.390 ;
        RECT 121.420 131.280 136.720 131.380 ;
        RECT 121.420 131.270 136.755 131.280 ;
        RECT 121.380 131.150 136.755 131.270 ;
        RECT 121.380 131.040 125.380 131.150 ;
        RECT 126.430 131.070 128.170 131.150 ;
        RECT 128.750 131.070 136.755 131.150 ;
        RECT 126.430 130.990 127.680 131.070 ;
        RECT 128.755 131.050 136.755 131.070 ;
        RECT 120.990 130.740 121.220 130.990 ;
        RECT 125.540 130.850 125.770 130.990 ;
        RECT 128.320 130.850 128.550 131.000 ;
        RECT 125.540 130.740 128.550 130.850 ;
        RECT 136.960 130.740 137.190 131.000 ;
        RECT 120.990 130.300 137.190 130.740 ;
        RECT 120.990 130.030 121.220 130.300 ;
        RECT 125.540 130.270 137.190 130.300 ;
        RECT 125.540 130.180 128.550 130.270 ;
        RECT 125.540 130.030 125.770 130.180 ;
        RECT 128.320 130.040 128.550 130.180 ;
        RECT 136.960 130.040 137.190 130.270 ;
        RECT 121.380 129.750 125.380 129.980 ;
        RECT 128.755 129.770 136.755 129.990 ;
        RECT 137.520 129.770 138.480 131.810 ;
        RECT 128.755 129.760 138.480 129.770 ;
        RECT 121.380 129.680 125.370 129.750 ;
        RECT 119.930 129.570 125.370 129.680 ;
        RECT 128.810 129.600 138.480 129.760 ;
        RECT 119.930 129.480 123.060 129.570 ;
        RECT 136.550 129.550 138.480 129.600 ;
        RECT 119.930 126.210 120.760 129.480 ;
        RECT 124.410 129.020 129.660 129.030 ;
        RECT 124.410 128.910 136.720 129.020 ;
        RECT 121.440 128.850 136.720 128.910 ;
        RECT 121.440 128.840 136.755 128.850 ;
        RECT 121.380 128.710 136.755 128.840 ;
        RECT 121.380 128.700 126.540 128.710 ;
        RECT 121.380 128.610 125.380 128.700 ;
        RECT 128.755 128.620 136.755 128.710 ;
        RECT 128.840 128.610 136.730 128.620 ;
        RECT 120.990 128.250 121.220 128.560 ;
        RECT 121.440 128.250 125.340 128.610 ;
        RECT 125.540 128.250 125.770 128.560 ;
        RECT 120.990 126.910 125.770 128.250 ;
        RECT 120.990 126.600 121.220 126.910 ;
        RECT 125.540 126.600 125.770 126.910 ;
        RECT 128.320 128.030 128.550 128.570 ;
        RECT 129.360 128.030 130.370 128.060 ;
        RECT 136.960 128.030 137.190 128.570 ;
        RECT 128.320 127.130 137.190 128.030 ;
        RECT 128.320 126.610 128.550 127.130 ;
        RECT 129.360 127.060 130.370 127.130 ;
        RECT 136.960 126.610 137.190 127.130 ;
        RECT 121.380 126.320 125.380 126.550 ;
        RECT 128.755 126.330 136.755 126.560 ;
        RECT 119.930 126.170 121.060 126.210 ;
        RECT 119.930 126.090 121.300 126.170 ;
        RECT 121.670 126.100 125.330 126.320 ;
        RECT 121.670 126.090 123.110 126.100 ;
        RECT 119.930 126.050 123.110 126.090 ;
        RECT 119.930 125.960 122.620 126.050 ;
        RECT 128.820 126.040 136.710 126.330 ;
        RECT 119.930 125.900 121.950 125.960 ;
        RECT 119.930 125.850 121.700 125.900 ;
        RECT 119.930 122.510 120.760 125.850 ;
        RECT 128.810 125.550 136.730 125.560 ;
        RECT 125.040 125.540 136.730 125.550 ;
        RECT 121.420 125.420 136.730 125.540 ;
        RECT 121.420 125.410 136.755 125.420 ;
        RECT 121.380 125.290 136.755 125.410 ;
        RECT 121.380 125.180 125.380 125.290 ;
        RECT 120.990 124.840 121.220 125.130 ;
        RECT 121.440 124.840 125.330 125.180 ;
        RECT 125.540 124.840 125.770 125.130 ;
        RECT 120.990 123.470 125.770 124.840 ;
        RECT 120.990 123.170 121.220 123.470 ;
        RECT 125.540 123.170 125.770 123.470 ;
        RECT 121.380 122.890 125.380 123.120 ;
        RECT 121.630 122.660 125.200 122.890 ;
        RECT 121.630 122.510 125.320 122.660 ;
        RECT 119.930 122.230 125.320 122.510 ;
        RECT 126.570 122.340 127.190 125.290 ;
        RECT 128.755 125.190 136.755 125.290 ;
        RECT 128.810 125.180 136.730 125.190 ;
        RECT 128.320 124.480 128.550 125.140 ;
        RECT 129.330 124.480 130.330 124.570 ;
        RECT 136.960 124.480 137.190 125.140 ;
        RECT 128.320 123.660 137.190 124.480 ;
        RECT 128.320 123.180 128.550 123.660 ;
        RECT 129.330 123.570 130.330 123.660 ;
        RECT 136.960 123.180 137.190 123.660 ;
        RECT 128.755 122.900 136.755 123.130 ;
        RECT 119.930 121.770 125.330 122.230 ;
        RECT 119.930 120.430 121.930 121.770 ;
        RECT 123.680 121.760 125.330 121.770 ;
        RECT 122.370 120.490 123.370 121.210 ;
        RECT 123.680 120.950 123.990 121.760 ;
        RECT 124.450 121.480 125.330 121.760 ;
        RECT 125.570 121.940 127.190 122.340 ;
        RECT 128.840 121.990 136.710 122.900 ;
        RECT 124.390 121.250 125.390 121.480 ;
        RECT 125.570 121.290 125.920 121.940 ;
        RECT 126.570 121.930 127.190 121.940 ;
        RECT 128.755 121.760 136.755 121.990 ;
        RECT 128.840 121.750 136.710 121.760 ;
        RECT 124.450 121.040 125.330 121.060 ;
        RECT 123.720 120.660 123.990 120.950 ;
        RECT 124.390 120.810 125.390 121.040 ;
        RECT 125.550 121.000 125.920 121.290 ;
        RECT 125.580 120.940 125.920 121.000 ;
        RECT 126.680 121.610 127.440 121.660 ;
        RECT 128.320 121.610 128.550 121.710 ;
        RECT 126.680 121.400 128.550 121.610 ;
        RECT 136.960 121.400 137.190 121.710 ;
        RECT 126.680 120.980 129.220 121.400 ;
        RECT 136.590 120.980 137.190 121.400 ;
        RECT 124.450 120.660 125.330 120.810 ;
        RECT 124.460 120.490 125.190 120.660 ;
        RECT 120.010 120.420 121.930 120.430 ;
        RECT 102.400 119.080 105.400 119.310 ;
        RECT 105.610 119.120 105.950 119.950 ;
        RECT 107.960 119.940 118.600 120.010 ;
        RECT 102.450 119.050 105.310 119.080 ;
        RECT 102.450 119.030 103.620 119.050 ;
        RECT 104.580 119.040 105.310 119.050 ;
        RECT 102.400 118.640 105.400 118.870 ;
        RECT 105.605 118.830 105.950 119.120 ;
        RECT 106.140 118.900 118.600 119.940 ;
        RECT 122.340 119.370 125.190 120.490 ;
        RECT 125.580 120.190 125.930 120.940 ;
        RECT 126.680 120.820 128.550 120.980 ;
        RECT 126.680 120.770 127.440 120.820 ;
        RECT 128.320 120.750 128.550 120.820 ;
        RECT 136.960 120.750 137.190 120.980 ;
        RECT 128.755 120.470 136.755 120.700 ;
        RECT 125.580 120.130 125.870 120.190 ;
        RECT 125.490 120.010 125.870 120.130 ;
        RECT 128.850 120.070 136.710 120.470 ;
        RECT 137.520 120.070 138.480 129.550 ;
        RECT 139.960 131.780 140.220 131.810 ;
        RECT 139.960 129.680 140.790 131.780 ;
        RECT 146.460 131.390 147.710 131.830 ;
        RECT 144.400 131.380 149.640 131.390 ;
        RECT 141.450 131.280 156.750 131.380 ;
        RECT 141.450 131.270 156.785 131.280 ;
        RECT 141.410 131.150 156.785 131.270 ;
        RECT 141.410 131.040 145.410 131.150 ;
        RECT 146.460 131.070 148.200 131.150 ;
        RECT 148.780 131.070 156.785 131.150 ;
        RECT 146.460 130.990 147.710 131.070 ;
        RECT 148.785 131.050 156.785 131.070 ;
        RECT 141.020 130.740 141.250 130.990 ;
        RECT 145.570 130.850 145.800 130.990 ;
        RECT 148.350 130.850 148.580 131.000 ;
        RECT 145.570 130.740 148.580 130.850 ;
        RECT 156.990 130.740 157.220 131.000 ;
        RECT 141.020 130.300 157.220 130.740 ;
        RECT 141.020 130.030 141.250 130.300 ;
        RECT 145.570 130.270 157.220 130.300 ;
        RECT 145.570 130.180 148.580 130.270 ;
        RECT 145.570 130.030 145.800 130.180 ;
        RECT 148.350 130.040 148.580 130.180 ;
        RECT 156.990 130.040 157.220 130.270 ;
        RECT 141.410 129.750 145.410 129.980 ;
        RECT 148.785 129.770 156.785 129.990 ;
        RECT 157.550 129.770 158.510 131.810 ;
        RECT 148.785 129.760 158.510 129.770 ;
        RECT 141.410 129.680 145.400 129.750 ;
        RECT 139.960 129.570 145.400 129.680 ;
        RECT 148.840 129.600 158.510 129.760 ;
        RECT 139.960 129.480 143.090 129.570 ;
        RECT 156.580 129.550 158.510 129.600 ;
        RECT 139.960 126.210 140.790 129.480 ;
        RECT 144.440 129.020 149.690 129.030 ;
        RECT 144.440 128.910 156.750 129.020 ;
        RECT 141.470 128.850 156.750 128.910 ;
        RECT 141.470 128.840 156.785 128.850 ;
        RECT 141.410 128.710 156.785 128.840 ;
        RECT 141.410 128.700 146.570 128.710 ;
        RECT 141.410 128.610 145.410 128.700 ;
        RECT 148.785 128.620 156.785 128.710 ;
        RECT 148.870 128.610 156.760 128.620 ;
        RECT 141.020 128.250 141.250 128.560 ;
        RECT 141.470 128.250 145.370 128.610 ;
        RECT 145.570 128.250 145.800 128.560 ;
        RECT 141.020 126.910 145.800 128.250 ;
        RECT 141.020 126.600 141.250 126.910 ;
        RECT 145.570 126.600 145.800 126.910 ;
        RECT 148.350 128.030 148.580 128.570 ;
        RECT 149.390 128.030 150.400 128.060 ;
        RECT 156.990 128.030 157.220 128.570 ;
        RECT 148.350 127.130 157.220 128.030 ;
        RECT 148.350 126.610 148.580 127.130 ;
        RECT 149.390 127.060 150.400 127.130 ;
        RECT 156.990 126.610 157.220 127.130 ;
        RECT 141.410 126.320 145.410 126.550 ;
        RECT 148.785 126.330 156.785 126.560 ;
        RECT 139.960 126.170 141.090 126.210 ;
        RECT 139.960 126.090 141.330 126.170 ;
        RECT 141.700 126.100 145.360 126.320 ;
        RECT 141.700 126.090 143.140 126.100 ;
        RECT 139.960 126.050 143.140 126.090 ;
        RECT 139.960 125.960 142.650 126.050 ;
        RECT 148.850 126.040 156.740 126.330 ;
        RECT 139.960 125.900 141.980 125.960 ;
        RECT 139.960 125.850 141.730 125.900 ;
        RECT 139.960 122.510 140.790 125.850 ;
        RECT 148.840 125.550 156.760 125.560 ;
        RECT 145.070 125.540 156.760 125.550 ;
        RECT 141.450 125.420 156.760 125.540 ;
        RECT 141.450 125.410 156.785 125.420 ;
        RECT 141.410 125.290 156.785 125.410 ;
        RECT 141.410 125.180 145.410 125.290 ;
        RECT 141.020 124.840 141.250 125.130 ;
        RECT 141.470 124.840 145.360 125.180 ;
        RECT 145.570 124.840 145.800 125.130 ;
        RECT 141.020 123.470 145.800 124.840 ;
        RECT 141.020 123.170 141.250 123.470 ;
        RECT 145.570 123.170 145.800 123.470 ;
        RECT 141.410 122.890 145.410 123.120 ;
        RECT 141.660 122.660 145.230 122.890 ;
        RECT 141.660 122.510 145.350 122.660 ;
        RECT 139.960 122.230 145.350 122.510 ;
        RECT 146.600 122.340 147.220 125.290 ;
        RECT 148.785 125.190 156.785 125.290 ;
        RECT 148.840 125.180 156.760 125.190 ;
        RECT 148.350 124.480 148.580 125.140 ;
        RECT 149.360 124.480 150.360 124.570 ;
        RECT 156.990 124.480 157.220 125.140 ;
        RECT 148.350 123.660 157.220 124.480 ;
        RECT 148.350 123.180 148.580 123.660 ;
        RECT 149.360 123.570 150.360 123.660 ;
        RECT 156.990 123.180 157.220 123.660 ;
        RECT 148.785 122.900 156.785 123.130 ;
        RECT 139.960 121.770 145.360 122.230 ;
        RECT 139.960 120.430 141.960 121.770 ;
        RECT 143.710 121.760 145.360 121.770 ;
        RECT 142.400 120.490 143.400 121.210 ;
        RECT 143.710 120.950 144.020 121.760 ;
        RECT 144.480 121.480 145.360 121.760 ;
        RECT 145.600 121.940 147.220 122.340 ;
        RECT 148.870 121.990 156.740 122.900 ;
        RECT 144.420 121.250 145.420 121.480 ;
        RECT 145.600 121.290 145.950 121.940 ;
        RECT 146.600 121.930 147.220 121.940 ;
        RECT 148.785 121.760 156.785 121.990 ;
        RECT 148.870 121.750 156.740 121.760 ;
        RECT 144.480 121.040 145.360 121.060 ;
        RECT 143.750 120.660 144.020 120.950 ;
        RECT 144.420 120.810 145.420 121.040 ;
        RECT 145.580 121.000 145.950 121.290 ;
        RECT 145.610 120.940 145.950 121.000 ;
        RECT 146.710 121.610 147.470 121.660 ;
        RECT 148.350 121.610 148.580 121.710 ;
        RECT 146.710 121.400 148.580 121.610 ;
        RECT 156.990 121.400 157.220 121.710 ;
        RECT 146.710 120.980 149.250 121.400 ;
        RECT 156.620 120.980 157.220 121.400 ;
        RECT 144.480 120.660 145.360 120.810 ;
        RECT 144.490 120.490 145.220 120.660 ;
        RECT 140.040 120.420 141.960 120.430 ;
        RECT 122.280 119.140 125.280 119.370 ;
        RECT 125.490 119.180 125.830 120.010 ;
        RECT 127.840 120.000 138.480 120.070 ;
        RECT 122.330 119.110 125.190 119.140 ;
        RECT 122.330 119.090 123.500 119.110 ;
        RECT 124.460 119.100 125.190 119.110 ;
        RECT 106.140 118.880 118.470 118.900 ;
        RECT 106.410 118.870 111.850 118.880 ;
        RECT 112.850 118.870 118.470 118.880 ;
        RECT 105.610 118.720 105.950 118.830 ;
        RECT 122.280 118.700 125.280 118.930 ;
        RECT 125.485 118.890 125.830 119.180 ;
        RECT 126.020 118.960 138.480 120.000 ;
        RECT 142.370 119.370 145.220 120.490 ;
        RECT 145.610 120.190 145.960 120.940 ;
        RECT 146.710 120.820 148.580 120.980 ;
        RECT 146.710 120.770 147.470 120.820 ;
        RECT 148.350 120.750 148.580 120.820 ;
        RECT 156.990 120.750 157.220 120.980 ;
        RECT 148.785 120.470 156.785 120.700 ;
        RECT 145.610 120.130 145.900 120.190 ;
        RECT 145.520 120.010 145.900 120.130 ;
        RECT 148.880 120.070 156.740 120.470 ;
        RECT 157.550 120.070 158.510 129.550 ;
        RECT 142.310 119.140 145.310 119.370 ;
        RECT 145.520 119.180 145.860 120.010 ;
        RECT 147.870 120.000 158.510 120.070 ;
        RECT 142.360 119.110 145.220 119.140 ;
        RECT 142.360 119.090 143.530 119.110 ;
        RECT 144.490 119.100 145.220 119.110 ;
        RECT 126.020 118.940 138.350 118.960 ;
        RECT 126.290 118.930 131.730 118.940 ;
        RECT 132.730 118.930 138.350 118.940 ;
        RECT 125.490 118.780 125.830 118.890 ;
        RECT 142.310 118.700 145.310 118.930 ;
        RECT 145.515 118.890 145.860 119.180 ;
        RECT 146.050 118.960 158.510 120.000 ;
        RECT 146.050 118.940 158.380 118.960 ;
        RECT 146.320 118.930 151.760 118.940 ;
        RECT 152.760 118.930 158.380 118.940 ;
        RECT 145.520 118.780 145.860 118.890 ;
        RECT 100.000 116.780 100.260 116.810 ;
        RECT 100.000 114.680 100.830 116.780 ;
        RECT 106.500 116.390 107.750 116.830 ;
        RECT 104.440 116.380 109.680 116.390 ;
        RECT 101.490 116.280 116.790 116.380 ;
        RECT 101.490 116.270 116.825 116.280 ;
        RECT 101.450 116.150 116.825 116.270 ;
        RECT 101.450 116.040 105.450 116.150 ;
        RECT 106.500 116.070 108.240 116.150 ;
        RECT 108.820 116.070 116.825 116.150 ;
        RECT 106.500 115.990 107.750 116.070 ;
        RECT 108.825 116.050 116.825 116.070 ;
        RECT 101.060 115.740 101.290 115.990 ;
        RECT 105.610 115.850 105.840 115.990 ;
        RECT 108.390 115.850 108.620 116.000 ;
        RECT 105.610 115.740 108.620 115.850 ;
        RECT 117.030 115.740 117.260 116.000 ;
        RECT 101.060 115.300 117.260 115.740 ;
        RECT 101.060 115.030 101.290 115.300 ;
        RECT 105.610 115.270 117.260 115.300 ;
        RECT 105.610 115.180 108.620 115.270 ;
        RECT 105.610 115.030 105.840 115.180 ;
        RECT 108.390 115.040 108.620 115.180 ;
        RECT 117.030 115.040 117.260 115.270 ;
        RECT 101.450 114.750 105.450 114.980 ;
        RECT 108.825 114.770 116.825 114.990 ;
        RECT 117.590 114.770 118.550 116.810 ;
        RECT 108.825 114.760 118.550 114.770 ;
        RECT 101.450 114.680 105.440 114.750 ;
        RECT 100.000 114.570 105.440 114.680 ;
        RECT 108.880 114.600 118.550 114.760 ;
        RECT 100.000 114.480 103.130 114.570 ;
        RECT 116.620 114.550 118.550 114.600 ;
        RECT 100.000 111.210 100.830 114.480 ;
        RECT 104.480 114.020 109.730 114.030 ;
        RECT 104.480 113.910 116.790 114.020 ;
        RECT 101.510 113.850 116.790 113.910 ;
        RECT 101.510 113.840 116.825 113.850 ;
        RECT 101.450 113.710 116.825 113.840 ;
        RECT 101.450 113.700 106.610 113.710 ;
        RECT 101.450 113.610 105.450 113.700 ;
        RECT 108.825 113.620 116.825 113.710 ;
        RECT 108.910 113.610 116.800 113.620 ;
        RECT 101.060 113.250 101.290 113.560 ;
        RECT 101.510 113.250 105.410 113.610 ;
        RECT 105.610 113.250 105.840 113.560 ;
        RECT 101.060 111.910 105.840 113.250 ;
        RECT 101.060 111.600 101.290 111.910 ;
        RECT 105.610 111.600 105.840 111.910 ;
        RECT 108.390 113.030 108.620 113.570 ;
        RECT 109.430 113.030 110.440 113.060 ;
        RECT 117.030 113.030 117.260 113.570 ;
        RECT 108.390 112.130 117.260 113.030 ;
        RECT 108.390 111.610 108.620 112.130 ;
        RECT 109.430 112.060 110.440 112.130 ;
        RECT 117.030 111.610 117.260 112.130 ;
        RECT 101.450 111.320 105.450 111.550 ;
        RECT 108.825 111.330 116.825 111.560 ;
        RECT 100.000 111.170 101.130 111.210 ;
        RECT 100.000 111.090 101.370 111.170 ;
        RECT 101.740 111.100 105.400 111.320 ;
        RECT 101.740 111.090 103.180 111.100 ;
        RECT 100.000 111.050 103.180 111.090 ;
        RECT 100.000 110.960 102.690 111.050 ;
        RECT 108.890 111.040 116.780 111.330 ;
        RECT 100.000 110.900 102.020 110.960 ;
        RECT 100.000 110.850 101.770 110.900 ;
        RECT 100.000 107.510 100.830 110.850 ;
        RECT 108.880 110.550 116.800 110.560 ;
        RECT 105.110 110.540 116.800 110.550 ;
        RECT 101.490 110.420 116.800 110.540 ;
        RECT 101.490 110.410 116.825 110.420 ;
        RECT 101.450 110.290 116.825 110.410 ;
        RECT 101.450 110.180 105.450 110.290 ;
        RECT 101.060 109.840 101.290 110.130 ;
        RECT 101.510 109.840 105.400 110.180 ;
        RECT 105.610 109.840 105.840 110.130 ;
        RECT 101.060 108.470 105.840 109.840 ;
        RECT 101.060 108.170 101.290 108.470 ;
        RECT 105.610 108.170 105.840 108.470 ;
        RECT 101.450 107.890 105.450 108.120 ;
        RECT 101.700 107.660 105.270 107.890 ;
        RECT 101.700 107.510 105.390 107.660 ;
        RECT 100.000 107.230 105.390 107.510 ;
        RECT 106.640 107.340 107.260 110.290 ;
        RECT 108.825 110.190 116.825 110.290 ;
        RECT 108.880 110.180 116.800 110.190 ;
        RECT 108.390 109.480 108.620 110.140 ;
        RECT 109.400 109.480 110.400 109.570 ;
        RECT 117.030 109.480 117.260 110.140 ;
        RECT 108.390 108.660 117.260 109.480 ;
        RECT 108.390 108.180 108.620 108.660 ;
        RECT 109.400 108.570 110.400 108.660 ;
        RECT 117.030 108.180 117.260 108.660 ;
        RECT 108.825 107.900 116.825 108.130 ;
        RECT 100.000 106.770 105.400 107.230 ;
        RECT 100.000 105.430 102.000 106.770 ;
        RECT 103.750 106.760 105.400 106.770 ;
        RECT 102.440 105.490 103.440 106.210 ;
        RECT 103.750 105.950 104.060 106.760 ;
        RECT 104.520 106.480 105.400 106.760 ;
        RECT 105.640 106.940 107.260 107.340 ;
        RECT 108.910 106.990 116.780 107.900 ;
        RECT 104.460 106.250 105.460 106.480 ;
        RECT 105.640 106.290 105.990 106.940 ;
        RECT 106.640 106.930 107.260 106.940 ;
        RECT 108.825 106.760 116.825 106.990 ;
        RECT 108.910 106.750 116.780 106.760 ;
        RECT 104.520 106.040 105.400 106.060 ;
        RECT 103.790 105.660 104.060 105.950 ;
        RECT 104.460 105.810 105.460 106.040 ;
        RECT 105.620 106.000 105.990 106.290 ;
        RECT 105.650 105.940 105.990 106.000 ;
        RECT 106.750 106.610 107.510 106.660 ;
        RECT 108.390 106.610 108.620 106.710 ;
        RECT 106.750 106.400 108.620 106.610 ;
        RECT 117.030 106.400 117.260 106.710 ;
        RECT 106.750 105.980 109.290 106.400 ;
        RECT 116.660 105.980 117.260 106.400 ;
        RECT 104.520 105.660 105.400 105.810 ;
        RECT 104.530 105.490 105.260 105.660 ;
        RECT 100.080 105.420 102.000 105.430 ;
        RECT 102.410 104.370 105.260 105.490 ;
        RECT 105.650 105.190 106.000 105.940 ;
        RECT 106.750 105.820 108.620 105.980 ;
        RECT 106.750 105.770 107.510 105.820 ;
        RECT 108.390 105.750 108.620 105.820 ;
        RECT 117.030 105.750 117.260 105.980 ;
        RECT 108.825 105.470 116.825 105.700 ;
        RECT 105.650 105.130 105.940 105.190 ;
        RECT 105.560 105.010 105.940 105.130 ;
        RECT 108.920 105.070 116.780 105.470 ;
        RECT 117.590 105.070 118.550 114.550 ;
        RECT 119.930 116.780 120.190 116.810 ;
        RECT 119.930 114.680 120.760 116.780 ;
        RECT 126.430 116.390 127.680 116.830 ;
        RECT 124.370 116.380 129.610 116.390 ;
        RECT 121.420 116.280 136.720 116.380 ;
        RECT 121.420 116.270 136.755 116.280 ;
        RECT 121.380 116.150 136.755 116.270 ;
        RECT 121.380 116.040 125.380 116.150 ;
        RECT 126.430 116.070 128.170 116.150 ;
        RECT 128.750 116.070 136.755 116.150 ;
        RECT 126.430 115.990 127.680 116.070 ;
        RECT 128.755 116.050 136.755 116.070 ;
        RECT 120.990 115.740 121.220 115.990 ;
        RECT 125.540 115.850 125.770 115.990 ;
        RECT 128.320 115.850 128.550 116.000 ;
        RECT 125.540 115.740 128.550 115.850 ;
        RECT 136.960 115.740 137.190 116.000 ;
        RECT 120.990 115.300 137.190 115.740 ;
        RECT 120.990 115.030 121.220 115.300 ;
        RECT 125.540 115.270 137.190 115.300 ;
        RECT 125.540 115.180 128.550 115.270 ;
        RECT 125.540 115.030 125.770 115.180 ;
        RECT 128.320 115.040 128.550 115.180 ;
        RECT 136.960 115.040 137.190 115.270 ;
        RECT 121.380 114.750 125.380 114.980 ;
        RECT 128.755 114.770 136.755 114.990 ;
        RECT 137.520 114.770 138.480 116.810 ;
        RECT 128.755 114.760 138.480 114.770 ;
        RECT 121.380 114.680 125.370 114.750 ;
        RECT 119.930 114.570 125.370 114.680 ;
        RECT 128.810 114.600 138.480 114.760 ;
        RECT 119.930 114.480 123.060 114.570 ;
        RECT 136.550 114.550 138.480 114.600 ;
        RECT 119.930 111.210 120.760 114.480 ;
        RECT 124.410 114.020 129.660 114.030 ;
        RECT 124.410 113.910 136.720 114.020 ;
        RECT 121.440 113.850 136.720 113.910 ;
        RECT 121.440 113.840 136.755 113.850 ;
        RECT 121.380 113.710 136.755 113.840 ;
        RECT 121.380 113.700 126.540 113.710 ;
        RECT 121.380 113.610 125.380 113.700 ;
        RECT 128.755 113.620 136.755 113.710 ;
        RECT 128.840 113.610 136.730 113.620 ;
        RECT 120.990 113.250 121.220 113.560 ;
        RECT 121.440 113.250 125.340 113.610 ;
        RECT 125.540 113.250 125.770 113.560 ;
        RECT 120.990 111.910 125.770 113.250 ;
        RECT 120.990 111.600 121.220 111.910 ;
        RECT 125.540 111.600 125.770 111.910 ;
        RECT 128.320 113.030 128.550 113.570 ;
        RECT 129.360 113.030 130.370 113.060 ;
        RECT 136.960 113.030 137.190 113.570 ;
        RECT 128.320 112.130 137.190 113.030 ;
        RECT 128.320 111.610 128.550 112.130 ;
        RECT 129.360 112.060 130.370 112.130 ;
        RECT 136.960 111.610 137.190 112.130 ;
        RECT 121.380 111.320 125.380 111.550 ;
        RECT 128.755 111.330 136.755 111.560 ;
        RECT 119.930 111.170 121.060 111.210 ;
        RECT 119.930 111.090 121.300 111.170 ;
        RECT 121.670 111.100 125.330 111.320 ;
        RECT 121.670 111.090 123.110 111.100 ;
        RECT 119.930 111.050 123.110 111.090 ;
        RECT 119.930 110.960 122.620 111.050 ;
        RECT 128.820 111.040 136.710 111.330 ;
        RECT 119.930 110.900 121.950 110.960 ;
        RECT 119.930 110.850 121.700 110.900 ;
        RECT 119.930 107.510 120.760 110.850 ;
        RECT 128.810 110.550 136.730 110.560 ;
        RECT 125.040 110.540 136.730 110.550 ;
        RECT 121.420 110.420 136.730 110.540 ;
        RECT 121.420 110.410 136.755 110.420 ;
        RECT 121.380 110.290 136.755 110.410 ;
        RECT 121.380 110.180 125.380 110.290 ;
        RECT 120.990 109.840 121.220 110.130 ;
        RECT 121.440 109.840 125.330 110.180 ;
        RECT 125.540 109.840 125.770 110.130 ;
        RECT 120.990 108.470 125.770 109.840 ;
        RECT 120.990 108.170 121.220 108.470 ;
        RECT 125.540 108.170 125.770 108.470 ;
        RECT 121.380 107.890 125.380 108.120 ;
        RECT 121.630 107.660 125.200 107.890 ;
        RECT 121.630 107.510 125.320 107.660 ;
        RECT 119.930 107.230 125.320 107.510 ;
        RECT 126.570 107.340 127.190 110.290 ;
        RECT 128.755 110.190 136.755 110.290 ;
        RECT 128.810 110.180 136.730 110.190 ;
        RECT 128.320 109.480 128.550 110.140 ;
        RECT 129.330 109.480 130.330 109.570 ;
        RECT 136.960 109.480 137.190 110.140 ;
        RECT 128.320 108.660 137.190 109.480 ;
        RECT 128.320 108.180 128.550 108.660 ;
        RECT 129.330 108.570 130.330 108.660 ;
        RECT 136.960 108.180 137.190 108.660 ;
        RECT 128.755 107.900 136.755 108.130 ;
        RECT 119.930 106.770 125.330 107.230 ;
        RECT 119.930 105.430 121.930 106.770 ;
        RECT 123.680 106.760 125.330 106.770 ;
        RECT 122.370 105.490 123.370 106.210 ;
        RECT 123.680 105.950 123.990 106.760 ;
        RECT 124.450 106.480 125.330 106.760 ;
        RECT 125.570 106.940 127.190 107.340 ;
        RECT 128.840 106.990 136.710 107.900 ;
        RECT 124.390 106.250 125.390 106.480 ;
        RECT 125.570 106.290 125.920 106.940 ;
        RECT 126.570 106.930 127.190 106.940 ;
        RECT 128.755 106.760 136.755 106.990 ;
        RECT 128.840 106.750 136.710 106.760 ;
        RECT 124.450 106.040 125.330 106.060 ;
        RECT 123.720 105.660 123.990 105.950 ;
        RECT 124.390 105.810 125.390 106.040 ;
        RECT 125.550 106.000 125.920 106.290 ;
        RECT 125.580 105.940 125.920 106.000 ;
        RECT 126.680 106.610 127.440 106.660 ;
        RECT 128.320 106.610 128.550 106.710 ;
        RECT 126.680 106.400 128.550 106.610 ;
        RECT 136.960 106.400 137.190 106.710 ;
        RECT 126.680 105.980 129.220 106.400 ;
        RECT 136.590 105.980 137.190 106.400 ;
        RECT 124.450 105.660 125.330 105.810 ;
        RECT 124.460 105.490 125.190 105.660 ;
        RECT 120.010 105.420 121.930 105.430 ;
        RECT 102.350 104.140 105.350 104.370 ;
        RECT 105.560 104.180 105.900 105.010 ;
        RECT 107.910 105.000 118.550 105.070 ;
        RECT 102.400 104.110 105.260 104.140 ;
        RECT 102.400 104.090 103.570 104.110 ;
        RECT 104.530 104.100 105.260 104.110 ;
        RECT 102.350 103.700 105.350 103.930 ;
        RECT 105.555 103.890 105.900 104.180 ;
        RECT 106.090 103.960 118.550 105.000 ;
        RECT 122.340 104.370 125.190 105.490 ;
        RECT 125.580 105.190 125.930 105.940 ;
        RECT 126.680 105.820 128.550 105.980 ;
        RECT 126.680 105.770 127.440 105.820 ;
        RECT 128.320 105.750 128.550 105.820 ;
        RECT 136.960 105.750 137.190 105.980 ;
        RECT 128.755 105.470 136.755 105.700 ;
        RECT 125.580 105.130 125.870 105.190 ;
        RECT 125.490 105.010 125.870 105.130 ;
        RECT 128.850 105.070 136.710 105.470 ;
        RECT 137.520 105.070 138.480 114.550 ;
        RECT 139.960 116.780 140.220 116.810 ;
        RECT 139.960 114.680 140.790 116.780 ;
        RECT 146.460 116.390 147.710 116.830 ;
        RECT 144.400 116.380 149.640 116.390 ;
        RECT 141.450 116.280 156.750 116.380 ;
        RECT 141.450 116.270 156.785 116.280 ;
        RECT 141.410 116.150 156.785 116.270 ;
        RECT 141.410 116.040 145.410 116.150 ;
        RECT 146.460 116.070 148.200 116.150 ;
        RECT 148.780 116.070 156.785 116.150 ;
        RECT 146.460 115.990 147.710 116.070 ;
        RECT 148.785 116.050 156.785 116.070 ;
        RECT 141.020 115.740 141.250 115.990 ;
        RECT 145.570 115.850 145.800 115.990 ;
        RECT 148.350 115.850 148.580 116.000 ;
        RECT 145.570 115.740 148.580 115.850 ;
        RECT 156.990 115.740 157.220 116.000 ;
        RECT 141.020 115.300 157.220 115.740 ;
        RECT 141.020 115.030 141.250 115.300 ;
        RECT 145.570 115.270 157.220 115.300 ;
        RECT 145.570 115.180 148.580 115.270 ;
        RECT 145.570 115.030 145.800 115.180 ;
        RECT 148.350 115.040 148.580 115.180 ;
        RECT 156.990 115.040 157.220 115.270 ;
        RECT 141.410 114.750 145.410 114.980 ;
        RECT 148.785 114.770 156.785 114.990 ;
        RECT 157.550 114.770 158.510 116.810 ;
        RECT 148.785 114.760 158.510 114.770 ;
        RECT 141.410 114.680 145.400 114.750 ;
        RECT 139.960 114.570 145.400 114.680 ;
        RECT 148.840 114.600 158.510 114.760 ;
        RECT 139.960 114.480 143.090 114.570 ;
        RECT 156.580 114.550 158.510 114.600 ;
        RECT 139.960 111.210 140.790 114.480 ;
        RECT 144.440 114.020 149.690 114.030 ;
        RECT 144.440 113.910 156.750 114.020 ;
        RECT 141.470 113.850 156.750 113.910 ;
        RECT 141.470 113.840 156.785 113.850 ;
        RECT 141.410 113.710 156.785 113.840 ;
        RECT 141.410 113.700 146.570 113.710 ;
        RECT 141.410 113.610 145.410 113.700 ;
        RECT 148.785 113.620 156.785 113.710 ;
        RECT 148.870 113.610 156.760 113.620 ;
        RECT 141.020 113.250 141.250 113.560 ;
        RECT 141.470 113.250 145.370 113.610 ;
        RECT 145.570 113.250 145.800 113.560 ;
        RECT 141.020 111.910 145.800 113.250 ;
        RECT 141.020 111.600 141.250 111.910 ;
        RECT 145.570 111.600 145.800 111.910 ;
        RECT 148.350 113.030 148.580 113.570 ;
        RECT 149.390 113.030 150.400 113.060 ;
        RECT 156.990 113.030 157.220 113.570 ;
        RECT 148.350 112.130 157.220 113.030 ;
        RECT 148.350 111.610 148.580 112.130 ;
        RECT 149.390 112.060 150.400 112.130 ;
        RECT 156.990 111.610 157.220 112.130 ;
        RECT 141.410 111.320 145.410 111.550 ;
        RECT 148.785 111.330 156.785 111.560 ;
        RECT 139.960 111.170 141.090 111.210 ;
        RECT 139.960 111.090 141.330 111.170 ;
        RECT 141.700 111.100 145.360 111.320 ;
        RECT 141.700 111.090 143.140 111.100 ;
        RECT 139.960 111.050 143.140 111.090 ;
        RECT 139.960 110.960 142.650 111.050 ;
        RECT 148.850 111.040 156.740 111.330 ;
        RECT 139.960 110.900 141.980 110.960 ;
        RECT 139.960 110.850 141.730 110.900 ;
        RECT 139.960 107.510 140.790 110.850 ;
        RECT 148.840 110.550 156.760 110.560 ;
        RECT 145.070 110.540 156.760 110.550 ;
        RECT 141.450 110.420 156.760 110.540 ;
        RECT 141.450 110.410 156.785 110.420 ;
        RECT 141.410 110.290 156.785 110.410 ;
        RECT 141.410 110.180 145.410 110.290 ;
        RECT 141.020 109.840 141.250 110.130 ;
        RECT 141.470 109.840 145.360 110.180 ;
        RECT 145.570 109.840 145.800 110.130 ;
        RECT 141.020 108.470 145.800 109.840 ;
        RECT 141.020 108.170 141.250 108.470 ;
        RECT 145.570 108.170 145.800 108.470 ;
        RECT 141.410 107.890 145.410 108.120 ;
        RECT 141.660 107.660 145.230 107.890 ;
        RECT 141.660 107.510 145.350 107.660 ;
        RECT 139.960 107.230 145.350 107.510 ;
        RECT 146.600 107.340 147.220 110.290 ;
        RECT 148.785 110.190 156.785 110.290 ;
        RECT 148.840 110.180 156.760 110.190 ;
        RECT 148.350 109.480 148.580 110.140 ;
        RECT 149.360 109.480 150.360 109.570 ;
        RECT 156.990 109.480 157.220 110.140 ;
        RECT 148.350 108.660 157.220 109.480 ;
        RECT 148.350 108.180 148.580 108.660 ;
        RECT 149.360 108.570 150.360 108.660 ;
        RECT 156.990 108.180 157.220 108.660 ;
        RECT 148.785 107.900 156.785 108.130 ;
        RECT 139.960 106.770 145.360 107.230 ;
        RECT 139.960 105.430 141.960 106.770 ;
        RECT 143.710 106.760 145.360 106.770 ;
        RECT 142.400 105.490 143.400 106.210 ;
        RECT 143.710 105.950 144.020 106.760 ;
        RECT 144.480 106.480 145.360 106.760 ;
        RECT 145.600 106.940 147.220 107.340 ;
        RECT 148.870 106.990 156.740 107.900 ;
        RECT 144.420 106.250 145.420 106.480 ;
        RECT 145.600 106.290 145.950 106.940 ;
        RECT 146.600 106.930 147.220 106.940 ;
        RECT 148.785 106.760 156.785 106.990 ;
        RECT 148.870 106.750 156.740 106.760 ;
        RECT 144.480 106.040 145.360 106.060 ;
        RECT 143.750 105.660 144.020 105.950 ;
        RECT 144.420 105.810 145.420 106.040 ;
        RECT 145.580 106.000 145.950 106.290 ;
        RECT 145.610 105.940 145.950 106.000 ;
        RECT 146.710 106.610 147.470 106.660 ;
        RECT 148.350 106.610 148.580 106.710 ;
        RECT 146.710 106.400 148.580 106.610 ;
        RECT 156.990 106.400 157.220 106.710 ;
        RECT 146.710 105.980 149.250 106.400 ;
        RECT 156.620 105.980 157.220 106.400 ;
        RECT 144.480 105.660 145.360 105.810 ;
        RECT 144.490 105.490 145.220 105.660 ;
        RECT 140.040 105.420 141.960 105.430 ;
        RECT 122.280 104.140 125.280 104.370 ;
        RECT 125.490 104.180 125.830 105.010 ;
        RECT 127.840 105.000 138.480 105.070 ;
        RECT 122.330 104.110 125.190 104.140 ;
        RECT 122.330 104.090 123.500 104.110 ;
        RECT 124.460 104.100 125.190 104.110 ;
        RECT 106.090 103.940 118.420 103.960 ;
        RECT 106.360 103.930 111.800 103.940 ;
        RECT 112.800 103.930 118.420 103.940 ;
        RECT 105.560 103.780 105.900 103.890 ;
        RECT 122.280 103.700 125.280 103.930 ;
        RECT 125.485 103.890 125.830 104.180 ;
        RECT 126.020 103.960 138.480 105.000 ;
        RECT 142.370 104.370 145.220 105.490 ;
        RECT 145.610 105.190 145.960 105.940 ;
        RECT 146.710 105.820 148.580 105.980 ;
        RECT 146.710 105.770 147.470 105.820 ;
        RECT 148.350 105.750 148.580 105.820 ;
        RECT 156.990 105.750 157.220 105.980 ;
        RECT 148.785 105.470 156.785 105.700 ;
        RECT 145.610 105.130 145.900 105.190 ;
        RECT 145.520 105.010 145.900 105.130 ;
        RECT 148.880 105.070 156.740 105.470 ;
        RECT 157.550 105.070 158.510 114.550 ;
        RECT 142.310 104.140 145.310 104.370 ;
        RECT 145.520 104.180 145.860 105.010 ;
        RECT 147.870 105.000 158.510 105.070 ;
        RECT 142.360 104.110 145.220 104.140 ;
        RECT 142.360 104.090 143.530 104.110 ;
        RECT 144.490 104.100 145.220 104.110 ;
        RECT 126.020 103.940 138.350 103.960 ;
        RECT 126.290 103.930 131.730 103.940 ;
        RECT 132.730 103.930 138.350 103.940 ;
        RECT 125.490 103.780 125.830 103.890 ;
        RECT 142.310 103.700 145.310 103.930 ;
        RECT 145.515 103.890 145.860 104.180 ;
        RECT 146.050 103.960 158.510 105.000 ;
        RECT 146.050 103.940 158.380 103.960 ;
        RECT 146.320 103.930 151.760 103.940 ;
        RECT 152.760 103.930 158.380 103.940 ;
        RECT 145.520 103.780 145.860 103.890 ;
      LAYER met2 ;
        RECT 115.915 220.575 116.285 220.585 ;
        RECT 115.770 220.315 116.285 220.575 ;
        RECT 115.915 220.305 116.285 220.315 ;
        RECT 121.210 218.215 121.530 218.275 ;
        RECT 125.435 218.215 125.805 218.285 ;
        RECT 121.210 218.075 125.805 218.215 ;
        RECT 121.210 218.015 121.530 218.075 ;
        RECT 125.435 218.005 125.805 218.075 ;
        RECT 128.010 218.215 128.330 218.275 ;
        RECT 132.235 218.215 132.605 218.285 ;
        RECT 139.035 218.275 139.405 218.285 ;
        RECT 128.010 218.075 132.605 218.215 ;
        RECT 128.010 218.015 128.330 218.075 ;
        RECT 132.235 218.005 132.605 218.075 ;
        RECT 138.890 218.015 139.405 218.275 ;
        RECT 139.035 218.005 139.405 218.015 ;
        RECT 116.450 217.755 116.770 217.815 ;
        RECT 119.850 217.755 120.170 217.815 ;
        RECT 121.550 217.755 121.870 217.815 ;
        RECT 116.450 217.615 121.870 217.755 ;
        RECT 116.450 217.555 116.770 217.615 ;
        RECT 119.850 217.555 120.170 217.615 ;
        RECT 121.550 217.555 121.870 217.615 ;
        RECT 124.610 217.755 124.930 217.815 ;
        RECT 126.650 217.755 126.970 217.815 ;
        RECT 124.610 217.615 126.970 217.755 ;
        RECT 124.610 217.555 124.930 217.615 ;
        RECT 126.650 217.555 126.970 217.615 ;
        RECT 127.330 217.755 127.650 217.815 ;
        RECT 130.050 217.755 130.370 217.815 ;
        RECT 131.750 217.755 132.070 217.815 ;
        RECT 127.330 217.615 132.070 217.755 ;
        RECT 127.330 217.555 127.650 217.615 ;
        RECT 130.050 217.555 130.370 217.615 ;
        RECT 131.750 217.555 132.070 217.615 ;
        RECT 133.110 217.755 133.430 217.815 ;
        RECT 134.470 217.755 134.790 217.815 ;
        RECT 133.110 217.615 134.790 217.755 ;
        RECT 133.110 217.555 133.430 217.615 ;
        RECT 134.470 217.555 134.790 217.615 ;
        RECT 138.890 215.915 139.210 215.975 ;
        RECT 140.250 215.915 140.570 215.975 ;
        RECT 138.890 215.775 140.570 215.915 ;
        RECT 138.890 215.715 139.210 215.775 ;
        RECT 140.250 215.715 140.570 215.775 ;
        RECT 123.930 215.455 124.250 215.515 ;
        RECT 126.310 215.455 126.630 215.515 ;
        RECT 123.930 215.315 126.630 215.455 ;
        RECT 123.930 215.255 124.250 215.315 ;
        RECT 126.310 215.255 126.630 215.315 ;
        RECT 135.490 215.455 135.810 215.515 ;
        RECT 137.530 215.455 137.850 215.515 ;
        RECT 135.490 215.315 137.850 215.455 ;
        RECT 135.490 215.255 135.810 215.315 ;
        RECT 137.530 215.255 137.850 215.315 ;
        RECT 117.130 214.995 117.450 215.055 ;
        RECT 118.490 214.995 118.810 215.055 ;
        RECT 117.130 214.855 118.810 214.995 ;
        RECT 117.130 214.795 117.450 214.855 ;
        RECT 118.490 214.795 118.810 214.855 ;
        RECT 144.330 213.615 144.650 213.675 ;
        RECT 146.030 213.615 146.350 213.675 ;
        RECT 144.330 213.475 146.350 213.615 ;
        RECT 144.330 213.415 144.650 213.475 ;
        RECT 146.030 213.415 146.350 213.475 ;
        RECT 117.130 213.155 117.450 213.215 ;
        RECT 120.870 213.155 121.190 213.215 ;
        RECT 117.130 213.015 121.190 213.155 ;
        RECT 117.130 212.955 117.450 213.015 ;
        RECT 120.870 212.955 121.190 213.015 ;
        RECT 130.730 213.155 131.050 213.215 ;
        RECT 134.470 213.155 134.790 213.215 ;
        RECT 130.730 213.015 134.790 213.155 ;
        RECT 130.730 212.955 131.050 213.015 ;
        RECT 134.470 212.955 134.790 213.015 ;
        RECT 117.130 212.695 117.450 212.755 ;
        RECT 121.210 212.695 121.530 212.755 ;
        RECT 126.990 212.695 127.310 212.755 ;
        RECT 117.130 212.555 127.310 212.695 ;
        RECT 117.130 212.495 117.450 212.555 ;
        RECT 121.210 212.495 121.530 212.555 ;
        RECT 126.990 212.495 127.310 212.555 ;
        RECT 128.010 212.695 128.330 212.755 ;
        RECT 129.030 212.695 129.350 212.755 ;
        RECT 128.010 212.555 129.350 212.695 ;
        RECT 128.010 212.495 128.330 212.555 ;
        RECT 129.030 212.495 129.350 212.555 ;
        RECT 126.990 212.235 127.310 212.295 ;
        RECT 134.810 212.235 135.130 212.295 ;
        RECT 137.870 212.235 138.190 212.295 ;
        RECT 126.990 212.095 138.190 212.235 ;
        RECT 126.990 212.035 127.310 212.095 ;
        RECT 134.810 212.035 135.130 212.095 ;
        RECT 137.870 212.035 138.190 212.095 ;
        RECT 119.170 210.855 119.490 210.915 ;
        RECT 124.270 210.855 124.590 210.915 ;
        RECT 119.170 210.715 124.590 210.855 ;
        RECT 119.170 210.655 119.490 210.715 ;
        RECT 124.270 210.655 124.590 210.715 ;
        RECT 132.770 210.855 133.090 210.915 ;
        RECT 135.150 210.855 135.470 210.915 ;
        RECT 132.770 210.715 135.470 210.855 ;
        RECT 132.770 210.655 133.090 210.715 ;
        RECT 135.150 210.655 135.470 210.715 ;
        RECT 138.210 210.855 138.530 210.915 ;
        RECT 139.910 210.855 140.230 210.915 ;
        RECT 138.210 210.715 140.230 210.855 ;
        RECT 138.210 210.655 138.530 210.715 ;
        RECT 139.910 210.655 140.230 210.715 ;
        RECT 117.130 210.395 117.450 210.455 ;
        RECT 121.550 210.395 121.870 210.455 ;
        RECT 117.130 210.255 121.870 210.395 ;
        RECT 117.130 210.195 117.450 210.255 ;
        RECT 121.550 210.195 121.870 210.255 ;
        RECT 138.890 210.395 139.210 210.455 ;
        RECT 139.910 210.395 140.230 210.455 ;
        RECT 138.890 210.255 140.230 210.395 ;
        RECT 138.890 210.195 139.210 210.255 ;
        RECT 139.910 210.195 140.230 210.255 ;
        RECT 121.890 209.935 122.210 209.995 ;
        RECT 125.290 209.935 125.610 209.995 ;
        RECT 129.710 209.935 130.030 209.995 ;
        RECT 121.890 209.795 130.030 209.935 ;
        RECT 121.890 209.735 122.210 209.795 ;
        RECT 125.290 209.735 125.610 209.795 ;
        RECT 129.710 209.735 130.030 209.795 ;
        RECT 144.330 209.015 144.650 209.075 ;
        RECT 146.030 209.015 146.350 209.075 ;
        RECT 144.330 208.875 146.350 209.015 ;
        RECT 144.330 208.815 144.650 208.875 ;
        RECT 146.030 208.815 146.350 208.875 ;
        RECT 143.795 208.555 144.165 208.625 ;
        RECT 146.030 208.555 146.350 208.615 ;
        RECT 143.795 208.415 146.350 208.555 ;
        RECT 143.795 208.345 144.165 208.415 ;
        RECT 146.030 208.355 146.350 208.415 ;
        RECT 113.390 208.095 113.710 208.155 ;
        RECT 117.130 208.095 117.450 208.155 ;
        RECT 113.390 207.955 117.450 208.095 ;
        RECT 113.390 207.895 113.710 207.955 ;
        RECT 117.130 207.895 117.450 207.955 ;
        RECT 135.150 208.095 135.470 208.155 ;
        RECT 138.890 208.095 139.210 208.155 ;
        RECT 140.590 208.095 140.910 208.155 ;
        RECT 142.630 208.095 142.950 208.155 ;
        RECT 135.150 207.955 142.950 208.095 ;
        RECT 135.150 207.895 135.470 207.955 ;
        RECT 138.890 207.895 139.210 207.955 ;
        RECT 140.590 207.895 140.910 207.955 ;
        RECT 142.630 207.895 142.950 207.955 ;
        RECT 133.110 207.175 133.430 207.235 ;
        RECT 142.435 207.175 142.805 207.245 ;
        RECT 133.110 207.035 142.805 207.175 ;
        RECT 133.110 206.975 133.430 207.035 ;
        RECT 142.435 206.965 142.805 207.035 ;
        RECT 143.990 206.715 144.310 206.775 ;
        RECT 145.350 206.715 145.670 206.775 ;
        RECT 143.990 206.575 145.670 206.715 ;
        RECT 143.990 206.515 144.310 206.575 ;
        RECT 145.350 206.515 145.670 206.575 ;
        RECT 116.110 206.255 116.430 206.315 ;
        RECT 121.550 206.255 121.870 206.315 ;
        RECT 127.670 206.255 127.990 206.315 ;
        RECT 116.110 206.115 127.990 206.255 ;
        RECT 116.110 206.055 116.430 206.115 ;
        RECT 121.550 206.055 121.870 206.115 ;
        RECT 127.670 206.055 127.990 206.115 ;
        RECT 135.490 205.795 135.810 205.855 ;
        RECT 138.890 205.795 139.210 205.855 ;
        RECT 135.490 205.655 139.210 205.795 ;
        RECT 135.490 205.595 135.810 205.655 ;
        RECT 138.890 205.595 139.210 205.655 ;
        RECT 141.610 205.795 141.930 205.855 ;
        RECT 143.650 205.795 143.970 205.855 ;
        RECT 141.610 205.655 143.970 205.795 ;
        RECT 141.610 205.595 141.930 205.655 ;
        RECT 143.650 205.595 143.970 205.655 ;
        RECT 101.480 205.335 105.480 205.405 ;
        RECT 112.710 205.335 113.030 205.395 ;
        RECT 101.480 205.195 113.030 205.335 ;
        RECT 101.480 205.125 105.480 205.195 ;
        RECT 112.710 205.135 113.030 205.195 ;
        RECT 147.050 205.335 147.370 205.395 ;
        RECT 155.245 205.335 159.245 205.405 ;
        RECT 147.050 205.195 159.245 205.335 ;
        RECT 147.050 205.135 147.370 205.195 ;
        RECT 155.245 205.125 159.245 205.195 ;
        RECT 123.930 204.875 124.250 204.935 ;
        RECT 126.650 204.875 126.970 204.935 ;
        RECT 123.930 204.735 126.970 204.875 ;
        RECT 123.930 204.675 124.250 204.735 ;
        RECT 126.650 204.675 126.970 204.735 ;
        RECT 127.670 204.875 127.990 204.935 ;
        RECT 130.730 204.875 131.050 204.935 ;
        RECT 136.170 204.875 136.490 204.935 ;
        RECT 138.890 204.875 139.210 204.935 ;
        RECT 127.670 204.735 139.210 204.875 ;
        RECT 127.670 204.675 127.990 204.735 ;
        RECT 130.730 204.675 131.050 204.735 ;
        RECT 136.170 204.675 136.490 204.735 ;
        RECT 138.890 204.675 139.210 204.735 ;
        RECT 128.010 204.415 128.330 204.475 ;
        RECT 129.710 204.415 130.030 204.475 ;
        RECT 128.010 204.275 130.030 204.415 ;
        RECT 128.010 204.215 128.330 204.275 ;
        RECT 129.710 204.215 130.030 204.275 ;
        RECT 130.730 204.415 131.050 204.475 ;
        RECT 143.795 204.415 144.165 204.485 ;
        RECT 130.730 204.275 144.165 204.415 ;
        RECT 130.730 204.215 131.050 204.275 ;
        RECT 143.795 204.205 144.165 204.275 ;
        RECT 113.390 202.835 113.710 203.095 ;
        RECT 112.710 202.575 113.030 202.635 ;
        RECT 107.190 202.435 113.030 202.575 ;
        RECT 101.480 202.115 105.480 202.185 ;
        RECT 107.190 202.115 107.330 202.435 ;
        RECT 112.710 202.375 113.030 202.435 ;
        RECT 101.480 201.975 107.330 202.115 ;
        RECT 101.480 201.905 105.480 201.975 ;
        RECT 113.480 201.655 113.620 202.835 ;
        RECT 114.895 202.205 115.265 203.745 ;
        RECT 120.335 202.205 120.705 203.745 ;
        RECT 125.775 202.205 126.145 203.745 ;
        RECT 131.215 202.205 131.585 203.745 ;
        RECT 136.655 202.205 137.025 203.745 ;
        RECT 142.095 202.205 142.465 203.745 ;
        RECT 147.535 202.205 147.905 203.745 ;
        RECT 155.245 202.115 159.245 202.185 ;
        RECT 148.670 201.975 159.245 202.115 ;
        RECT 117.130 201.655 117.450 201.715 ;
        RECT 120.870 201.655 121.190 201.715 ;
        RECT 113.480 201.515 116.850 201.655 ;
        RECT 116.710 200.795 116.850 201.515 ;
        RECT 117.130 201.515 121.190 201.655 ;
        RECT 117.130 201.455 117.450 201.515 ;
        RECT 120.870 201.455 121.190 201.515 ;
        RECT 129.710 201.655 130.030 201.715 ;
        RECT 139.910 201.655 140.230 201.715 ;
        RECT 129.710 201.515 140.230 201.655 ;
        RECT 129.710 201.455 130.030 201.515 ;
        RECT 139.910 201.455 140.230 201.515 ;
        RECT 140.590 201.655 140.910 201.715 ;
        RECT 145.350 201.655 145.670 201.715 ;
        RECT 140.590 201.515 145.670 201.655 ;
        RECT 140.590 201.455 140.910 201.515 ;
        RECT 145.350 201.455 145.670 201.515 ;
        RECT 118.830 201.195 119.150 201.255 ;
        RECT 131.750 201.195 132.070 201.255 ;
        RECT 138.210 201.195 138.530 201.255 ;
        RECT 118.830 201.055 138.530 201.195 ;
        RECT 118.830 200.995 119.150 201.055 ;
        RECT 131.750 200.995 132.070 201.055 ;
        RECT 138.210 200.995 138.530 201.055 ;
        RECT 138.890 201.195 139.210 201.255 ;
        RECT 140.590 201.195 140.910 201.255 ;
        RECT 138.890 201.055 140.910 201.195 ;
        RECT 138.890 200.995 139.210 201.055 ;
        RECT 140.590 200.995 140.910 201.055 ;
        RECT 142.970 201.195 143.290 201.255 ;
        RECT 148.670 201.195 148.810 201.975 ;
        RECT 155.245 201.905 159.245 201.975 ;
        RECT 142.970 201.055 148.810 201.195 ;
        RECT 142.970 200.995 143.290 201.055 ;
        RECT 113.050 200.735 113.370 200.795 ;
        RECT 115.430 200.735 115.750 200.795 ;
        RECT 113.050 200.595 115.750 200.735 ;
        RECT 116.710 200.735 117.110 200.795 ;
        RECT 119.850 200.735 120.170 200.795 ;
        RECT 121.890 200.735 122.210 200.795 ;
        RECT 123.590 200.735 123.910 200.795 ;
        RECT 116.710 200.595 123.910 200.735 ;
        RECT 113.050 200.535 113.370 200.595 ;
        RECT 115.430 200.535 115.750 200.595 ;
        RECT 116.790 200.535 117.110 200.595 ;
        RECT 119.850 200.535 120.170 200.595 ;
        RECT 121.890 200.535 122.210 200.595 ;
        RECT 123.590 200.535 123.910 200.595 ;
        RECT 129.710 200.735 130.030 200.795 ;
        RECT 132.430 200.735 132.750 200.795 ;
        RECT 137.190 200.735 137.510 200.795 ;
        RECT 129.710 200.595 132.750 200.735 ;
        RECT 129.710 200.535 130.030 200.595 ;
        RECT 132.430 200.535 132.750 200.595 ;
        RECT 133.030 200.595 137.510 200.735 ;
        RECT 101.480 198.895 105.480 198.965 ;
        RECT 112.175 198.905 112.545 200.445 ;
        RECT 117.615 198.905 117.985 200.445 ;
        RECT 123.055 198.905 123.425 200.445 ;
        RECT 128.495 198.905 128.865 200.445 ;
        RECT 130.390 200.275 130.710 200.335 ;
        RECT 133.030 200.275 133.170 200.595 ;
        RECT 137.190 200.535 137.510 200.595 ;
        RECT 141.610 200.735 141.930 200.795 ;
        RECT 146.710 200.735 147.030 200.795 ;
        RECT 141.610 200.595 147.030 200.735 ;
        RECT 141.610 200.535 141.930 200.595 ;
        RECT 146.710 200.535 147.030 200.595 ;
        RECT 130.390 200.135 133.170 200.275 ;
        RECT 130.390 200.075 130.710 200.135 ;
        RECT 133.935 198.905 134.305 200.445 ;
        RECT 139.375 198.905 139.745 200.445 ;
        RECT 140.590 200.275 140.910 200.335 ;
        RECT 143.310 200.275 143.630 200.335 ;
        RECT 140.590 200.135 143.630 200.275 ;
        RECT 140.590 200.075 140.910 200.135 ;
        RECT 143.310 200.075 143.630 200.135 ;
        RECT 144.815 198.905 145.185 200.445 ;
        RECT 147.050 198.895 147.370 198.955 ;
        RECT 155.245 198.895 159.245 198.965 ;
        RECT 101.480 198.755 107.330 198.895 ;
        RECT 101.480 198.685 105.480 198.755 ;
        RECT 107.190 198.435 107.330 198.755 ;
        RECT 147.050 198.755 159.245 198.895 ;
        RECT 147.050 198.695 147.370 198.755 ;
        RECT 155.245 198.685 159.245 198.755 ;
        RECT 112.710 198.435 113.030 198.495 ;
        RECT 107.190 198.295 113.030 198.435 ;
        RECT 112.710 198.235 113.030 198.295 ;
        RECT 126.990 198.435 127.310 198.495 ;
        RECT 134.470 198.435 134.790 198.495 ;
        RECT 136.170 198.435 136.490 198.495 ;
        RECT 140.590 198.435 140.910 198.495 ;
        RECT 126.990 198.295 135.890 198.435 ;
        RECT 126.990 198.235 127.310 198.295 ;
        RECT 134.470 198.235 134.790 198.295 ;
        RECT 114.410 197.975 114.730 198.035 ;
        RECT 123.590 197.975 123.910 198.035 ;
        RECT 126.990 197.975 127.310 198.035 ;
        RECT 114.410 197.835 127.310 197.975 ;
        RECT 114.410 197.775 114.730 197.835 ;
        RECT 123.590 197.775 123.910 197.835 ;
        RECT 126.990 197.775 127.310 197.835 ;
        RECT 133.450 197.975 133.770 198.035 ;
        RECT 134.810 197.975 135.130 198.035 ;
        RECT 133.450 197.835 135.130 197.975 ;
        RECT 135.750 197.975 135.890 198.295 ;
        RECT 136.170 198.295 140.910 198.435 ;
        RECT 136.170 198.235 136.490 198.295 ;
        RECT 140.590 198.235 140.910 198.295 ;
        RECT 144.330 198.435 144.650 198.495 ;
        RECT 146.030 198.435 146.350 198.495 ;
        RECT 144.330 198.295 146.350 198.435 ;
        RECT 144.330 198.235 144.650 198.295 ;
        RECT 146.030 198.235 146.350 198.295 ;
        RECT 140.590 197.975 140.910 198.035 ;
        RECT 135.750 197.835 140.910 197.975 ;
        RECT 133.450 197.775 133.770 197.835 ;
        RECT 134.810 197.775 135.130 197.835 ;
        RECT 140.590 197.775 140.910 197.835 ;
        RECT 143.990 197.975 144.310 198.035 ;
        RECT 145.350 197.975 145.670 198.035 ;
        RECT 143.990 197.835 145.670 197.975 ;
        RECT 143.990 197.775 144.310 197.835 ;
        RECT 145.350 197.775 145.670 197.835 ;
        RECT 124.610 197.515 124.930 197.575 ;
        RECT 124.610 197.315 125.010 197.515 ;
        RECT 128.010 197.315 128.330 197.575 ;
        RECT 135.150 197.515 135.470 197.575 ;
        RECT 137.870 197.515 138.190 197.575 ;
        RECT 135.150 197.375 138.190 197.515 ;
        RECT 135.150 197.315 135.470 197.375 ;
        RECT 137.870 197.315 138.190 197.375 ;
        RECT 140.930 197.515 141.250 197.575 ;
        RECT 142.630 197.515 142.950 197.575 ;
        RECT 140.930 197.375 142.950 197.515 ;
        RECT 140.930 197.315 141.250 197.375 ;
        RECT 142.630 197.315 142.950 197.375 ;
        RECT 124.870 197.055 125.010 197.315 ;
        RECT 128.100 197.055 128.240 197.315 ;
        RECT 130.050 197.055 130.370 197.115 ;
        RECT 135.830 197.055 136.150 197.115 ;
        RECT 124.870 196.915 136.150 197.055 ;
        RECT 130.050 196.855 130.370 196.915 ;
        RECT 135.830 196.855 136.150 196.915 ;
        RECT 140.590 197.055 140.910 197.115 ;
        RECT 143.650 197.055 143.970 197.115 ;
        RECT 140.590 196.915 143.970 197.055 ;
        RECT 140.590 196.855 140.910 196.915 ;
        RECT 143.650 196.855 143.970 196.915 ;
        RECT 124.950 196.595 125.270 196.655 ;
        RECT 134.810 196.595 135.130 196.655 ;
        RECT 124.950 196.455 135.130 196.595 ;
        RECT 124.950 196.395 125.270 196.455 ;
        RECT 134.810 196.395 135.130 196.455 ;
        RECT 117.130 196.135 117.450 196.195 ;
        RECT 122.230 196.135 122.550 196.195 ;
        RECT 126.650 196.135 126.970 196.195 ;
        RECT 117.130 195.995 126.970 196.135 ;
        RECT 117.130 195.935 117.450 195.995 ;
        RECT 122.230 195.935 122.550 195.995 ;
        RECT 126.650 195.935 126.970 195.995 ;
        RECT 130.390 196.135 130.710 196.195 ;
        RECT 131.750 196.135 132.070 196.195 ;
        RECT 138.550 196.135 138.870 196.195 ;
        RECT 143.310 196.135 143.630 196.195 ;
        RECT 130.390 195.995 143.630 196.135 ;
        RECT 130.390 195.935 130.710 195.995 ;
        RECT 131.750 195.935 132.070 195.995 ;
        RECT 138.550 195.935 138.870 195.995 ;
        RECT 143.310 195.935 143.630 195.995 ;
        RECT 133.450 195.675 133.770 195.735 ;
        RECT 137.530 195.675 137.850 195.735 ;
        RECT 140.250 195.675 140.570 195.735 ;
        RECT 141.610 195.675 141.930 195.735 ;
        RECT 143.650 195.675 143.970 195.735 ;
        RECT 133.450 195.535 140.570 195.675 ;
        RECT 133.450 195.475 133.770 195.535 ;
        RECT 137.530 195.475 137.850 195.535 ;
        RECT 140.250 195.475 140.570 195.535 ;
        RECT 141.190 195.535 143.970 195.675 ;
        RECT 116.110 195.215 116.430 195.275 ;
        RECT 121.890 195.215 122.210 195.275 ;
        RECT 125.290 195.215 125.610 195.275 ;
        RECT 141.190 195.215 141.330 195.535 ;
        RECT 141.610 195.475 141.930 195.535 ;
        RECT 143.650 195.475 143.970 195.535 ;
        RECT 146.030 195.675 146.350 195.735 ;
        RECT 155.245 195.675 159.245 195.745 ;
        RECT 146.030 195.535 159.245 195.675 ;
        RECT 146.030 195.475 146.350 195.535 ;
        RECT 155.245 195.465 159.245 195.535 ;
        RECT 116.110 195.075 141.330 195.215 ;
        RECT 116.110 195.015 116.430 195.075 ;
        RECT 121.890 195.015 122.210 195.075 ;
        RECT 125.290 195.015 125.610 195.075 ;
        RECT 113.390 194.755 113.710 194.815 ;
        RECT 114.070 194.755 114.390 194.815 ;
        RECT 116.110 194.755 116.430 194.815 ;
        RECT 113.390 194.615 116.430 194.755 ;
        RECT 113.390 194.555 113.710 194.615 ;
        RECT 114.070 194.555 114.390 194.615 ;
        RECT 116.110 194.555 116.430 194.615 ;
        RECT 140.590 194.755 140.910 194.815 ;
        RECT 142.630 194.755 142.950 194.815 ;
        RECT 140.590 194.615 142.950 194.755 ;
        RECT 140.590 194.555 140.910 194.615 ;
        RECT 142.630 194.555 142.950 194.615 ;
        RECT 120.870 194.295 121.190 194.355 ;
        RECT 121.550 194.295 121.870 194.355 ;
        RECT 129.030 194.295 129.350 194.355 ;
        RECT 120.870 194.155 129.350 194.295 ;
        RECT 120.870 194.095 121.190 194.155 ;
        RECT 121.550 194.095 121.870 194.155 ;
        RECT 129.030 194.095 129.350 194.155 ;
        RECT 115.235 193.835 115.605 193.905 ;
        RECT 118.830 193.835 119.150 193.895 ;
        RECT 115.235 193.695 119.150 193.835 ;
        RECT 115.235 193.625 115.605 193.695 ;
        RECT 118.830 193.635 119.150 193.695 ;
        RECT 127.330 193.835 127.650 193.895 ;
        RECT 130.730 193.835 131.050 193.895 ;
        RECT 137.190 193.835 137.510 193.895 ;
        RECT 127.330 193.695 137.510 193.835 ;
        RECT 127.330 193.635 127.650 193.695 ;
        RECT 130.730 193.635 131.050 193.695 ;
        RECT 137.190 193.635 137.510 193.695 ;
        RECT 143.650 193.835 143.970 193.895 ;
        RECT 146.710 193.835 147.030 193.895 ;
        RECT 143.650 193.695 147.030 193.835 ;
        RECT 143.650 193.635 143.970 193.695 ;
        RECT 146.710 193.635 147.030 193.695 ;
        RECT 132.770 192.915 133.090 192.975 ;
        RECT 134.470 192.915 134.790 192.975 ;
        RECT 132.770 192.775 134.790 192.915 ;
        RECT 132.770 192.715 133.090 192.775 ;
        RECT 134.470 192.715 134.790 192.775 ;
        RECT 101.480 192.455 105.480 192.525 ;
        RECT 112.710 192.455 113.030 192.515 ;
        RECT 101.480 192.315 113.030 192.455 ;
        RECT 101.480 192.245 105.480 192.315 ;
        RECT 112.710 192.255 113.030 192.315 ;
        RECT 118.830 192.455 119.150 192.515 ;
        RECT 125.435 192.455 125.805 192.525 ;
        RECT 118.830 192.315 125.805 192.455 ;
        RECT 118.830 192.255 119.150 192.315 ;
        RECT 125.435 192.245 125.805 192.315 ;
        RECT 147.050 192.455 147.370 192.515 ;
        RECT 155.245 192.455 159.245 192.525 ;
        RECT 147.050 192.315 159.245 192.455 ;
        RECT 147.050 192.255 147.370 192.315 ;
        RECT 155.245 192.245 159.245 192.315 ;
        RECT 113.390 191.995 113.710 192.055 ;
        RECT 120.870 191.995 121.190 192.055 ;
        RECT 124.270 191.995 124.590 192.055 ;
        RECT 113.390 191.855 124.590 191.995 ;
        RECT 113.390 191.795 113.710 191.855 ;
        RECT 120.870 191.795 121.190 191.855 ;
        RECT 124.270 191.795 124.590 191.855 ;
        RECT 132.770 191.995 133.090 192.055 ;
        RECT 138.210 191.995 138.530 192.055 ;
        RECT 145.350 191.995 145.670 192.055 ;
        RECT 132.770 191.855 145.670 191.995 ;
        RECT 132.770 191.795 133.090 191.855 ;
        RECT 138.210 191.795 138.530 191.855 ;
        RECT 145.350 191.795 145.670 191.855 ;
        RECT 127.330 191.535 127.650 191.595 ;
        RECT 129.030 191.535 129.350 191.595 ;
        RECT 127.330 191.395 129.350 191.535 ;
        RECT 127.330 191.335 127.650 191.395 ;
        RECT 129.030 191.335 129.350 191.395 ;
        RECT 138.550 191.535 138.870 191.595 ;
        RECT 138.550 191.395 143.880 191.535 ;
        RECT 138.550 191.335 138.870 191.395 ;
        RECT 143.740 191.145 143.880 191.395 ;
        RECT 118.635 191.135 119.005 191.145 ;
        RECT 143.740 191.135 144.165 191.145 ;
        RECT 118.635 190.875 119.150 191.135 ;
        RECT 122.570 191.075 122.890 191.135 ;
        RECT 123.590 191.075 123.910 191.135 ;
        RECT 122.570 190.935 123.910 191.075 ;
        RECT 122.570 190.875 122.890 190.935 ;
        RECT 123.590 190.875 123.910 190.935 ;
        RECT 129.710 191.075 130.030 191.135 ;
        RECT 135.150 191.075 135.470 191.135 ;
        RECT 137.530 191.075 137.850 191.135 ;
        RECT 138.550 191.075 138.870 191.135 ;
        RECT 129.710 190.935 130.450 191.075 ;
        RECT 129.710 190.875 130.030 190.935 ;
        RECT 118.635 190.865 119.005 190.875 ;
        RECT 128.835 190.155 129.205 190.225 ;
        RECT 129.710 190.155 130.030 190.215 ;
        RECT 128.835 190.015 130.030 190.155 ;
        RECT 130.310 190.155 130.450 190.935 ;
        RECT 135.150 190.935 138.870 191.075 ;
        RECT 135.150 190.875 135.470 190.935 ;
        RECT 137.530 190.875 137.850 190.935 ;
        RECT 138.550 190.875 138.870 190.935 ;
        RECT 143.650 190.875 144.165 191.135 ;
        RECT 143.795 190.865 144.165 190.875 ;
        RECT 141.610 190.615 141.930 190.675 ;
        RECT 142.970 190.615 143.290 190.675 ;
        RECT 146.030 190.615 146.350 190.675 ;
        RECT 141.610 190.475 146.350 190.615 ;
        RECT 141.610 190.415 141.930 190.475 ;
        RECT 142.970 190.415 143.290 190.475 ;
        RECT 146.030 190.415 146.350 190.475 ;
        RECT 135.830 190.155 136.150 190.215 ;
        RECT 130.310 190.015 136.150 190.155 ;
        RECT 128.835 189.945 129.205 190.015 ;
        RECT 129.710 189.955 130.030 190.015 ;
        RECT 135.830 189.955 136.150 190.015 ;
        RECT 113.730 189.695 114.050 189.755 ;
        RECT 116.110 189.695 116.430 189.755 ;
        RECT 118.150 189.695 118.470 189.755 ;
        RECT 113.730 189.555 118.470 189.695 ;
        RECT 113.730 189.495 114.050 189.555 ;
        RECT 116.110 189.495 116.430 189.555 ;
        RECT 118.150 189.495 118.470 189.555 ;
        RECT 124.610 189.695 124.930 189.755 ;
        RECT 127.670 189.695 127.990 189.755 ;
        RECT 129.370 189.695 129.690 189.755 ;
        RECT 131.750 189.695 132.070 189.755 ;
        RECT 124.610 189.555 132.070 189.695 ;
        RECT 124.610 189.495 124.930 189.555 ;
        RECT 127.670 189.495 127.990 189.555 ;
        RECT 129.370 189.495 129.690 189.555 ;
        RECT 131.750 189.495 132.070 189.555 ;
        RECT 111.835 189.235 112.205 189.305 ;
        RECT 113.390 189.235 113.710 189.295 ;
        RECT 111.835 189.095 113.710 189.235 ;
        RECT 111.835 189.025 112.205 189.095 ;
        RECT 113.390 189.035 113.710 189.095 ;
        RECT 116.450 189.235 116.770 189.295 ;
        RECT 118.150 189.235 118.470 189.295 ;
        RECT 116.450 189.095 118.470 189.235 ;
        RECT 116.450 189.035 116.770 189.095 ;
        RECT 118.150 189.035 118.470 189.095 ;
        RECT 119.850 189.235 120.170 189.295 ;
        RECT 121.550 189.235 121.870 189.295 ;
        RECT 124.270 189.235 124.590 189.295 ;
        RECT 119.850 189.095 124.590 189.235 ;
        RECT 119.850 189.035 120.170 189.095 ;
        RECT 121.550 189.035 121.870 189.095 ;
        RECT 124.270 189.035 124.590 189.095 ;
        RECT 125.290 189.235 125.610 189.295 ;
        RECT 135.490 189.235 135.810 189.295 ;
        RECT 125.290 189.095 135.810 189.235 ;
        RECT 125.290 189.035 125.610 189.095 ;
        RECT 135.490 189.035 135.810 189.095 ;
        RECT 122.035 188.835 122.405 188.845 ;
        RECT 114.070 188.775 114.390 188.835 ;
        RECT 119.510 188.775 119.830 188.835 ;
        RECT 114.070 188.635 119.830 188.775 ;
        RECT 114.070 188.575 114.390 188.635 ;
        RECT 119.510 188.575 119.830 188.635 ;
        RECT 121.890 188.575 122.405 188.835 ;
        RECT 140.590 188.775 140.910 188.835 ;
        RECT 142.630 188.775 142.950 188.835 ;
        RECT 140.590 188.635 142.950 188.775 ;
        RECT 140.590 188.575 140.910 188.635 ;
        RECT 142.630 188.575 142.950 188.635 ;
        RECT 122.035 188.565 122.405 188.575 ;
        RECT 114.410 188.315 114.730 188.375 ;
        RECT 118.830 188.315 119.150 188.375 ;
        RECT 120.870 188.315 121.190 188.375 ;
        RECT 127.330 188.315 127.650 188.375 ;
        RECT 114.410 188.175 127.650 188.315 ;
        RECT 114.410 188.115 114.730 188.175 ;
        RECT 118.830 188.115 119.150 188.175 ;
        RECT 120.870 188.115 121.190 188.175 ;
        RECT 127.330 188.115 127.650 188.175 ;
        RECT 135.150 188.315 135.470 188.375 ;
        RECT 138.210 188.315 138.530 188.375 ;
        RECT 138.890 188.315 139.210 188.375 ;
        RECT 145.350 188.315 145.670 188.375 ;
        RECT 135.150 188.175 145.670 188.315 ;
        RECT 135.150 188.115 135.470 188.175 ;
        RECT 138.210 188.115 138.530 188.175 ;
        RECT 138.890 188.115 139.210 188.175 ;
        RECT 145.350 188.115 145.670 188.175 ;
        RECT 119.850 187.855 120.170 187.915 ;
        RECT 127.330 187.855 127.650 187.915 ;
        RECT 119.850 187.715 127.650 187.855 ;
        RECT 119.850 187.655 120.170 187.715 ;
        RECT 127.330 187.655 127.650 187.715 ;
        RECT 128.010 187.855 128.330 187.915 ;
        RECT 129.710 187.855 130.030 187.915 ;
        RECT 128.010 187.715 130.030 187.855 ;
        RECT 128.010 187.655 128.330 187.715 ;
        RECT 129.710 187.655 130.030 187.715 ;
        RECT 130.390 187.855 130.710 187.915 ;
        RECT 135.150 187.855 135.470 187.915 ;
        RECT 141.610 187.855 141.930 187.915 ;
        RECT 143.650 187.855 143.970 187.915 ;
        RECT 130.390 187.715 141.330 187.855 ;
        RECT 130.390 187.655 130.710 187.715 ;
        RECT 135.150 187.655 135.470 187.715 ;
        RECT 118.830 187.395 119.150 187.455 ;
        RECT 121.890 187.395 122.210 187.455 ;
        RECT 118.830 187.255 122.210 187.395 ;
        RECT 118.830 187.195 119.150 187.255 ;
        RECT 121.890 187.195 122.210 187.255 ;
        RECT 122.570 187.395 122.890 187.455 ;
        RECT 126.990 187.395 127.310 187.455 ;
        RECT 122.570 187.255 127.310 187.395 ;
        RECT 122.570 187.195 122.890 187.255 ;
        RECT 126.990 187.195 127.310 187.255 ;
        RECT 129.710 187.395 130.030 187.455 ;
        RECT 132.770 187.395 133.090 187.455 ;
        RECT 129.710 187.255 133.090 187.395 ;
        RECT 129.710 187.195 130.030 187.255 ;
        RECT 132.770 187.195 133.090 187.255 ;
        RECT 135.635 187.395 136.005 187.465 ;
        RECT 140.590 187.395 140.910 187.455 ;
        RECT 135.635 187.255 140.910 187.395 ;
        RECT 141.190 187.395 141.330 187.715 ;
        RECT 141.610 187.715 143.970 187.855 ;
        RECT 141.610 187.655 141.930 187.715 ;
        RECT 143.650 187.655 143.970 187.715 ;
        RECT 146.030 187.855 146.350 187.915 ;
        RECT 149.235 187.855 149.605 187.925 ;
        RECT 146.030 187.715 149.605 187.855 ;
        RECT 146.030 187.655 146.350 187.715 ;
        RECT 149.235 187.645 149.605 187.715 ;
        RECT 142.970 187.395 143.290 187.455 ;
        RECT 141.190 187.255 143.290 187.395 ;
        RECT 135.635 187.185 136.005 187.255 ;
        RECT 140.590 187.195 140.910 187.255 ;
        RECT 142.970 187.195 143.290 187.255 ;
        RECT 122.230 186.935 122.550 186.995 ;
        RECT 124.270 186.935 124.590 186.995 ;
        RECT 129.370 186.935 129.690 186.995 ;
        RECT 122.230 186.795 129.690 186.935 ;
        RECT 122.230 186.735 122.550 186.795 ;
        RECT 124.270 186.735 124.590 186.795 ;
        RECT 129.370 186.735 129.690 186.795 ;
        RECT 136.170 186.935 136.490 186.995 ;
        RECT 138.210 186.935 138.530 186.995 ;
        RECT 136.170 186.795 138.530 186.935 ;
        RECT 136.170 186.735 136.490 186.795 ;
        RECT 138.210 186.735 138.530 186.795 ;
        RECT 145.835 186.535 146.205 186.545 ;
        RECT 117.130 186.475 117.450 186.535 ;
        RECT 124.270 186.475 124.590 186.535 ;
        RECT 117.130 186.335 124.590 186.475 ;
        RECT 117.130 186.275 117.450 186.335 ;
        RECT 124.270 186.275 124.590 186.335 ;
        RECT 130.730 186.475 131.050 186.535 ;
        RECT 135.150 186.475 135.470 186.535 ;
        RECT 139.910 186.475 140.230 186.535 ;
        RECT 130.730 186.335 135.470 186.475 ;
        RECT 130.730 186.275 131.050 186.335 ;
        RECT 135.150 186.275 135.470 186.335 ;
        RECT 135.750 186.335 140.230 186.475 ;
        RECT 114.410 186.015 114.730 186.075 ;
        RECT 118.830 186.015 119.150 186.075 ;
        RECT 114.410 185.875 119.150 186.015 ;
        RECT 114.410 185.815 114.730 185.875 ;
        RECT 118.830 185.815 119.150 185.875 ;
        RECT 121.550 186.015 121.870 186.075 ;
        RECT 127.330 186.015 127.650 186.075 ;
        RECT 121.550 185.875 127.650 186.015 ;
        RECT 121.550 185.815 121.870 185.875 ;
        RECT 127.330 185.815 127.650 185.875 ;
        RECT 132.770 186.015 133.090 186.075 ;
        RECT 135.150 186.015 135.470 186.075 ;
        RECT 135.750 186.015 135.890 186.335 ;
        RECT 139.910 186.275 140.230 186.335 ;
        RECT 145.835 186.275 146.350 186.535 ;
        RECT 145.835 186.265 146.205 186.275 ;
        RECT 132.770 185.875 135.890 186.015 ;
        RECT 138.890 186.015 139.210 186.075 ;
        RECT 139.910 186.015 140.230 186.075 ;
        RECT 138.890 185.875 140.230 186.015 ;
        RECT 132.770 185.815 133.090 185.875 ;
        RECT 135.150 185.815 135.470 185.875 ;
        RECT 138.890 185.815 139.210 185.875 ;
        RECT 139.910 185.815 140.230 185.875 ;
        RECT 108.435 185.555 108.805 185.625 ;
        RECT 119.170 185.555 119.490 185.615 ;
        RECT 108.435 185.415 119.490 185.555 ;
        RECT 108.435 185.345 108.805 185.415 ;
        RECT 119.170 185.355 119.490 185.415 ;
        RECT 135.830 185.555 136.150 185.615 ;
        RECT 138.210 185.555 138.530 185.615 ;
        RECT 145.350 185.555 145.670 185.615 ;
        RECT 135.830 185.415 145.670 185.555 ;
        RECT 135.830 185.355 136.150 185.415 ;
        RECT 138.210 185.355 138.530 185.415 ;
        RECT 145.350 185.355 145.670 185.415 ;
        RECT 116.110 185.095 116.430 185.155 ;
        RECT 118.830 185.095 119.150 185.155 ;
        RECT 121.210 185.095 121.530 185.155 ;
        RECT 116.110 184.955 121.530 185.095 ;
        RECT 116.110 184.895 116.430 184.955 ;
        RECT 118.830 184.895 119.150 184.955 ;
        RECT 121.210 184.895 121.530 184.955 ;
        RECT 132.235 185.095 132.605 185.165 ;
        RECT 132.770 185.095 133.090 185.155 ;
        RECT 132.235 184.955 133.090 185.095 ;
        RECT 132.235 184.885 132.605 184.955 ;
        RECT 132.770 184.895 133.090 184.955 ;
        RECT 139.035 185.095 139.405 185.165 ;
        RECT 140.590 185.095 140.910 185.155 ;
        RECT 139.035 184.955 140.910 185.095 ;
        RECT 139.035 184.885 139.405 184.955 ;
        RECT 140.590 184.895 140.910 184.955 ;
        RECT 142.435 185.095 142.805 185.165 ;
        RECT 143.650 185.095 143.970 185.155 ;
        RECT 142.435 184.955 143.970 185.095 ;
        RECT 142.435 184.885 142.805 184.955 ;
        RECT 143.650 184.895 143.970 184.955 ;
        RECT 146.030 185.095 146.350 185.155 ;
        RECT 152.635 185.095 153.005 185.165 ;
        RECT 146.030 184.955 153.005 185.095 ;
        RECT 146.030 184.895 146.350 184.955 ;
        RECT 152.635 184.885 153.005 184.955 ;
        RECT 106.840 176.770 107.540 176.780 ;
        RECT 146.750 176.770 147.450 176.780 ;
        RECT 106.500 176.030 107.850 176.770 ;
        RECT 126.720 176.720 127.420 176.730 ;
        RECT 106.840 166.600 107.540 176.030 ;
        RECT 126.380 175.980 127.730 176.720 ;
        RECT 146.410 176.030 147.760 176.770 ;
        RECT 108.890 171.080 116.880 171.470 ;
        RECT 111.430 168.020 114.090 171.080 ;
        RECT 108.930 167.570 116.870 168.020 ;
        RECT 106.750 165.810 107.610 166.600 ;
        RECT 126.720 166.550 127.420 175.980 ;
        RECT 128.770 171.030 136.760 171.420 ;
        RECT 131.310 167.970 133.970 171.030 ;
        RECT 128.810 167.520 136.750 167.970 ;
        RECT 146.750 166.600 147.450 176.030 ;
        RECT 148.800 171.080 156.790 171.470 ;
        RECT 151.340 168.020 154.000 171.080 ;
        RECT 148.840 167.570 156.780 168.020 ;
        RECT 126.630 165.760 127.490 166.550 ;
        RECT 146.660 165.810 147.520 166.600 ;
        RECT 106.840 161.770 107.540 161.780 ;
        RECT 126.720 161.770 127.420 161.780 ;
        RECT 106.500 161.030 107.850 161.770 ;
        RECT 126.380 161.030 127.730 161.770 ;
        RECT 146.800 161.720 147.500 161.730 ;
        RECT 106.840 151.600 107.540 161.030 ;
        RECT 108.890 156.080 116.880 156.470 ;
        RECT 111.430 153.020 114.090 156.080 ;
        RECT 108.930 152.570 116.870 153.020 ;
        RECT 126.720 151.600 127.420 161.030 ;
        RECT 146.460 160.980 147.810 161.720 ;
        RECT 128.770 156.080 136.760 156.470 ;
        RECT 131.310 153.020 133.970 156.080 ;
        RECT 128.810 152.570 136.750 153.020 ;
        RECT 106.750 150.810 107.610 151.600 ;
        RECT 126.630 150.810 127.490 151.600 ;
        RECT 146.800 151.550 147.500 160.980 ;
        RECT 148.850 156.030 156.840 156.420 ;
        RECT 151.390 152.970 154.050 156.030 ;
        RECT 148.890 152.520 156.830 152.970 ;
        RECT 146.710 150.760 147.570 151.550 ;
        RECT 106.840 146.720 107.540 146.730 ;
        RECT 126.720 146.720 127.420 146.730 ;
        RECT 146.750 146.720 147.450 146.730 ;
        RECT 106.500 145.980 107.850 146.720 ;
        RECT 126.380 145.980 127.730 146.720 ;
        RECT 146.410 145.980 147.760 146.720 ;
        RECT 106.840 136.550 107.540 145.980 ;
        RECT 108.890 141.030 116.880 141.420 ;
        RECT 111.430 137.970 114.090 141.030 ;
        RECT 108.930 137.520 116.870 137.970 ;
        RECT 126.720 136.550 127.420 145.980 ;
        RECT 128.770 141.030 136.760 141.420 ;
        RECT 131.310 137.970 133.970 141.030 ;
        RECT 128.810 137.520 136.750 137.970 ;
        RECT 146.750 136.550 147.450 145.980 ;
        RECT 148.800 141.030 156.790 141.420 ;
        RECT 151.340 137.970 154.000 141.030 ;
        RECT 148.840 137.520 156.780 137.970 ;
        RECT 106.750 135.760 107.610 136.550 ;
        RECT 126.630 135.760 127.490 136.550 ;
        RECT 146.660 135.760 147.520 136.550 ;
        RECT 126.720 131.780 127.420 131.790 ;
        RECT 146.750 131.780 147.450 131.790 ;
        RECT 106.840 131.720 107.540 131.730 ;
        RECT 106.500 130.980 107.850 131.720 ;
        RECT 126.380 131.040 127.730 131.780 ;
        RECT 146.410 131.040 147.760 131.780 ;
        RECT 106.840 121.550 107.540 130.980 ;
        RECT 108.890 126.030 116.880 126.420 ;
        RECT 111.430 122.970 114.090 126.030 ;
        RECT 108.930 122.520 116.870 122.970 ;
        RECT 126.720 121.610 127.420 131.040 ;
        RECT 128.770 126.090 136.760 126.480 ;
        RECT 131.310 123.030 133.970 126.090 ;
        RECT 128.810 122.580 136.750 123.030 ;
        RECT 146.750 121.610 147.450 131.040 ;
        RECT 148.800 126.090 156.790 126.480 ;
        RECT 151.340 123.030 154.000 126.090 ;
        RECT 148.840 122.580 156.780 123.030 ;
        RECT 106.750 120.760 107.610 121.550 ;
        RECT 126.630 120.820 127.490 121.610 ;
        RECT 146.660 120.820 147.520 121.610 ;
        RECT 106.790 116.780 107.490 116.790 ;
        RECT 126.720 116.780 127.420 116.790 ;
        RECT 146.750 116.780 147.450 116.790 ;
        RECT 106.450 116.040 107.800 116.780 ;
        RECT 126.380 116.040 127.730 116.780 ;
        RECT 146.410 116.040 147.760 116.780 ;
        RECT 106.790 106.610 107.490 116.040 ;
        RECT 108.840 111.090 116.830 111.480 ;
        RECT 111.380 108.030 114.040 111.090 ;
        RECT 108.880 107.580 116.820 108.030 ;
        RECT 126.720 106.610 127.420 116.040 ;
        RECT 128.770 111.090 136.760 111.480 ;
        RECT 131.310 108.030 133.970 111.090 ;
        RECT 128.810 107.580 136.750 108.030 ;
        RECT 146.750 106.610 147.450 116.040 ;
        RECT 148.800 111.090 156.790 111.480 ;
        RECT 151.340 108.030 154.000 111.090 ;
        RECT 148.840 107.580 156.780 108.030 ;
        RECT 106.700 105.820 107.560 106.610 ;
        RECT 126.630 105.820 127.490 106.610 ;
        RECT 146.660 105.820 147.520 106.610 ;
      LAYER met3 ;
        RECT 115.120 220.825 115.720 224.815 ;
        RECT 115.120 220.815 116.250 220.825 ;
        RECT 125.320 220.815 125.920 224.815 ;
        RECT 132.120 220.815 132.720 224.815 ;
        RECT 138.920 220.815 139.520 224.815 ;
        RECT 142.320 220.815 142.920 224.815 ;
        RECT 115.270 220.610 116.250 220.815 ;
        RECT 115.270 220.525 116.265 220.610 ;
        RECT 115.935 220.280 116.265 220.525 ;
        RECT 125.470 218.310 125.770 220.815 ;
        RECT 132.270 218.310 132.570 220.815 ;
        RECT 139.070 218.310 139.370 220.815 ;
        RECT 125.455 217.980 125.785 218.310 ;
        RECT 132.255 217.980 132.585 218.310 ;
        RECT 139.055 217.980 139.385 218.310 ;
        RECT 142.470 207.270 142.770 220.815 ;
        RECT 143.815 208.320 144.145 208.650 ;
        RECT 142.455 206.940 142.785 207.270 ;
        RECT 143.830 204.510 144.130 208.320 ;
        RECT 143.815 204.180 144.145 204.510 ;
        RECT 114.915 202.185 115.245 203.765 ;
        RECT 120.355 202.185 120.685 203.765 ;
        RECT 125.795 202.185 126.125 203.765 ;
        RECT 131.235 202.185 131.565 203.765 ;
        RECT 136.675 202.185 137.005 203.765 ;
        RECT 142.115 202.185 142.445 203.765 ;
        RECT 112.195 198.885 112.525 200.465 ;
        RECT 117.635 198.885 117.965 200.465 ;
        RECT 123.075 198.885 123.405 200.465 ;
        RECT 128.515 198.885 128.845 200.465 ;
        RECT 133.955 198.885 134.285 200.465 ;
        RECT 139.395 198.885 139.725 200.465 ;
        RECT 115.255 193.600 115.585 193.930 ;
        RECT 111.855 189.000 112.185 189.330 ;
        RECT 108.455 185.320 108.785 185.650 ;
        RECT 108.470 181.770 108.770 185.320 ;
        RECT 111.870 181.770 112.170 189.000 ;
        RECT 115.270 181.770 115.570 193.600 ;
        RECT 125.455 192.220 125.785 192.550 ;
        RECT 118.655 190.840 118.985 191.170 ;
        RECT 118.670 181.770 118.970 190.840 ;
        RECT 122.055 188.540 122.385 188.870 ;
        RECT 122.070 181.770 122.370 188.540 ;
        RECT 125.470 181.770 125.770 192.220 ;
        RECT 143.830 191.170 144.130 204.180 ;
        RECT 147.555 202.185 147.885 203.765 ;
        RECT 144.835 198.885 145.165 200.465 ;
        RECT 143.815 190.840 144.145 191.170 ;
        RECT 128.855 189.920 129.185 190.250 ;
        RECT 128.870 181.770 129.170 189.920 ;
        RECT 149.255 187.620 149.585 187.950 ;
        RECT 135.655 187.160 135.985 187.490 ;
        RECT 132.255 184.860 132.585 185.190 ;
        RECT 132.270 181.770 132.570 184.860 ;
        RECT 135.670 181.770 135.970 187.160 ;
        RECT 145.855 186.240 146.185 186.570 ;
        RECT 139.055 184.860 139.385 185.190 ;
        RECT 142.455 184.860 142.785 185.190 ;
        RECT 139.070 181.770 139.370 184.860 ;
        RECT 142.470 181.770 142.770 184.860 ;
        RECT 145.870 181.770 146.170 186.240 ;
        RECT 149.270 181.770 149.570 187.620 ;
        RECT 152.655 184.860 152.985 185.190 ;
        RECT 152.670 181.770 152.970 184.860 ;
        RECT 108.320 177.770 108.920 181.770 ;
        RECT 111.720 177.770 112.320 181.770 ;
        RECT 115.120 177.770 115.720 181.770 ;
        RECT 118.520 177.770 119.120 181.770 ;
        RECT 121.920 177.770 122.520 181.770 ;
        RECT 125.320 177.770 125.920 181.770 ;
        RECT 128.720 177.770 129.320 181.770 ;
        RECT 132.120 177.770 132.720 181.770 ;
        RECT 135.520 177.770 136.120 181.770 ;
        RECT 138.920 177.770 139.520 181.770 ;
        RECT 142.320 177.770 142.920 181.770 ;
        RECT 145.720 177.770 146.320 181.770 ;
        RECT 149.120 177.770 149.720 181.770 ;
        RECT 152.520 177.770 153.120 181.770 ;
      LAYER met4 ;
        RECT 112.120 202.175 147.960 203.775 ;
        RECT 112.120 198.875 147.960 200.475 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

