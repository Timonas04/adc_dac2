magic
tech sky130A
magscale 1 2
timestamp 1730846558
<< viali >>
rect 10241 39593 10275 39627
rect 11069 39389 11103 39423
rect 13185 39389 13219 39423
rect 10425 39321 10459 39355
rect 10057 39253 10091 39287
rect 10225 39253 10259 39287
rect 11253 39253 11287 39287
rect 13001 39253 13035 39287
rect 7573 39049 7607 39083
rect 7205 38981 7239 39015
rect 7405 38981 7439 39015
rect 7910 38981 7944 39015
rect 10140 38981 10174 39015
rect 6929 38913 6963 38947
rect 7113 38913 7147 38947
rect 13102 38913 13136 38947
rect 7665 38845 7699 38879
rect 9873 38845 9907 38879
rect 13369 38845 13403 38879
rect 7113 38709 7147 38743
rect 7389 38709 7423 38743
rect 9045 38709 9079 38743
rect 11253 38709 11287 38743
rect 11989 38709 12023 38743
rect 7849 38505 7883 38539
rect 8585 38505 8619 38539
rect 10793 38505 10827 38539
rect 12081 38505 12115 38539
rect 12265 38505 12299 38539
rect 8125 38437 8159 38471
rect 6101 38369 6135 38403
rect 11161 38369 11195 38403
rect 13921 38369 13955 38403
rect 8125 38301 8159 38335
rect 8309 38301 8343 38335
rect 8953 38301 8987 38335
rect 10609 38301 10643 38335
rect 10793 38301 10827 38335
rect 11069 38301 11103 38335
rect 11253 38301 11287 38335
rect 11621 38301 11655 38335
rect 11805 38301 11839 38335
rect 6368 38233 6402 38267
rect 8033 38233 8067 38267
rect 8401 38233 8435 38267
rect 9198 38233 9232 38267
rect 11897 38233 11931 38267
rect 13654 38233 13688 38267
rect 7481 38165 7515 38199
rect 7665 38165 7699 38199
rect 7833 38165 7867 38199
rect 8601 38165 8635 38199
rect 8769 38165 8803 38199
rect 10333 38165 10367 38199
rect 11713 38165 11747 38199
rect 12097 38165 12131 38199
rect 12541 38165 12575 38199
rect 6653 37961 6687 37995
rect 6821 37961 6855 37995
rect 7205 37961 7239 37995
rect 8131 37961 8165 37995
rect 8217 37961 8251 37995
rect 12081 37961 12115 37995
rect 12725 37961 12759 37995
rect 13093 37961 13127 37995
rect 7021 37893 7055 37927
rect 7757 37893 7791 37927
rect 11253 37893 11287 37927
rect 12909 37893 12943 37927
rect 13553 37893 13587 37927
rect 7113 37825 7147 37859
rect 7297 37825 7331 37859
rect 7573 37825 7607 37859
rect 7665 37825 7699 37859
rect 8033 37825 8067 37859
rect 8309 37825 8343 37859
rect 8776 37825 8810 37859
rect 11529 37825 11563 37859
rect 11713 37825 11747 37859
rect 11805 37825 11839 37859
rect 11897 37825 11931 37859
rect 12173 37825 12207 37859
rect 12357 37825 12391 37859
rect 12449 37825 12483 37859
rect 12817 37825 12851 37859
rect 13185 37825 13219 37859
rect 13369 37825 13403 37859
rect 8401 37757 8435 37791
rect 8861 37757 8895 37791
rect 7389 37689 7423 37723
rect 12173 37689 12207 37723
rect 12541 37689 12575 37723
rect 6837 37621 6871 37655
rect 7941 37621 7975 37655
rect 10977 37621 11011 37655
rect 6929 37417 6963 37451
rect 11529 37417 11563 37451
rect 11713 37417 11747 37451
rect 12725 37417 12759 37451
rect 10149 37349 10183 37383
rect 10701 37281 10735 37315
rect 11345 37281 11379 37315
rect 9873 37213 9907 37247
rect 9965 37213 9999 37247
rect 10425 37213 10459 37247
rect 10517 37213 10551 37247
rect 10793 37213 10827 37247
rect 11069 37213 11103 37247
rect 11253 37213 11287 37247
rect 12633 37213 12667 37247
rect 12817 37213 12851 37247
rect 7113 37145 7147 37179
rect 10149 37145 10183 37179
rect 10885 37145 10919 37179
rect 11697 37145 11731 37179
rect 11897 37145 11931 37179
rect 6745 37077 6779 37111
rect 6913 37077 6947 37111
rect 10241 37077 10275 37111
rect 9873 36873 9907 36907
rect 2957 36805 2991 36839
rect 3157 36805 3191 36839
rect 6644 36805 6678 36839
rect 4241 36737 4275 36771
rect 6377 36737 6411 36771
rect 9781 36737 9815 36771
rect 10057 36737 10091 36771
rect 10609 36737 10643 36771
rect 10701 36737 10735 36771
rect 3985 36669 4019 36703
rect 10885 36669 10919 36703
rect 2789 36533 2823 36567
rect 2973 36533 3007 36567
rect 5365 36533 5399 36567
rect 7757 36533 7791 36567
rect 10057 36533 10091 36567
rect 10793 36533 10827 36567
rect 2053 36329 2087 36363
rect 3985 36329 4019 36363
rect 4169 36329 4203 36363
rect 6101 36329 6135 36363
rect 7021 36329 7055 36363
rect 12265 36329 12299 36363
rect 10609 36261 10643 36295
rect 12541 36261 12575 36295
rect 4721 36193 4755 36227
rect 6745 36193 6779 36227
rect 11437 36193 11471 36227
rect 13921 36193 13955 36227
rect 1961 36125 1995 36159
rect 2145 36125 2179 36159
rect 3350 36125 3384 36159
rect 3617 36125 3651 36159
rect 4629 36125 4663 36159
rect 4813 36125 4847 36159
rect 4905 36125 4939 36159
rect 5273 36125 5307 36159
rect 5549 36125 5583 36159
rect 5641 36125 5675 36159
rect 5825 36125 5859 36159
rect 5917 36125 5951 36159
rect 6101 36125 6135 36159
rect 6377 36125 6411 36159
rect 6653 36125 6687 36159
rect 9137 36125 9171 36159
rect 9413 36125 9447 36159
rect 10333 36125 10367 36159
rect 10517 36125 10551 36159
rect 10701 36125 10735 36159
rect 10793 36125 10827 36159
rect 11253 36125 11287 36159
rect 11529 36125 11563 36159
rect 11897 36125 11931 36159
rect 4153 36057 4187 36091
rect 4353 36057 4387 36091
rect 5089 36057 5123 36091
rect 6193 36057 6227 36091
rect 8033 36057 8067 36091
rect 9321 36057 9355 36091
rect 11621 36057 11655 36091
rect 13654 36057 13688 36091
rect 2237 35989 2271 36023
rect 4445 35989 4479 36023
rect 5457 35989 5491 36023
rect 7941 35989 7975 36023
rect 8953 35989 8987 36023
rect 10977 35989 11011 36023
rect 11069 35989 11103 36023
rect 12265 35989 12299 36023
rect 12449 35989 12483 36023
rect 2881 35785 2915 35819
rect 7113 35785 7147 35819
rect 8309 35785 8343 35819
rect 8585 35785 8619 35819
rect 8953 35785 8987 35819
rect 9965 35785 9999 35819
rect 11345 35785 11379 35819
rect 14013 35785 14047 35819
rect 3249 35717 3283 35751
rect 4721 35717 4755 35751
rect 4905 35717 4939 35751
rect 7297 35717 7331 35751
rect 8426 35717 8460 35751
rect 10333 35717 10367 35751
rect 11713 35717 11747 35751
rect 12173 35717 12207 35751
rect 12373 35717 12407 35751
rect 12878 35717 12912 35751
rect 3065 35649 3099 35683
rect 4813 35649 4847 35683
rect 5457 35649 5491 35683
rect 5549 35649 5583 35683
rect 5641 35649 5675 35683
rect 5733 35649 5767 35683
rect 6745 35649 6779 35683
rect 7205 35649 7239 35683
rect 7389 35649 7423 35683
rect 7481 35649 7515 35683
rect 7665 35649 7699 35683
rect 7849 35649 7883 35683
rect 8217 35649 8251 35683
rect 8677 35649 8711 35683
rect 9229 35649 9263 35683
rect 9413 35649 9447 35683
rect 9597 35649 9631 35683
rect 9873 35649 9907 35683
rect 10149 35649 10183 35683
rect 10241 35649 10275 35683
rect 10517 35649 10551 35683
rect 10609 35649 10643 35683
rect 10793 35649 10827 35683
rect 12081 35649 12115 35683
rect 5089 35581 5123 35615
rect 6653 35581 6687 35615
rect 7941 35581 7975 35615
rect 8769 35581 8803 35615
rect 8953 35581 8987 35615
rect 11069 35581 11103 35615
rect 12633 35581 12667 35615
rect 11529 35513 11563 35547
rect 4537 35445 4571 35479
rect 5273 35445 5307 35479
rect 9873 35445 9907 35479
rect 11161 35445 11195 35479
rect 11713 35445 11747 35479
rect 12357 35445 12391 35479
rect 12541 35445 12575 35479
rect 2237 35241 2271 35275
rect 4169 35241 4203 35275
rect 5825 35241 5859 35275
rect 6009 35241 6043 35275
rect 8033 35241 8067 35275
rect 8401 35241 8435 35275
rect 8953 35241 8987 35275
rect 9781 35241 9815 35275
rect 9965 35241 9999 35275
rect 10149 35241 10183 35275
rect 10977 35241 11011 35275
rect 3801 35173 3835 35207
rect 6193 35173 6227 35207
rect 8677 35173 8711 35207
rect 10609 35173 10643 35207
rect 8309 35105 8343 35139
rect 9413 35105 9447 35139
rect 12541 35105 12575 35139
rect 12817 35105 12851 35139
rect 3617 35037 3651 35071
rect 4445 35037 4479 35071
rect 7665 35037 7699 35071
rect 7849 35037 7883 35071
rect 8217 35037 8251 35071
rect 8493 35037 8527 35071
rect 9137 35037 9171 35071
rect 9229 35037 9263 35071
rect 9505 35037 9539 35071
rect 9689 35037 9723 35071
rect 9873 35037 9907 35071
rect 10701 35037 10735 35071
rect 11253 35037 11287 35071
rect 11345 35037 11379 35071
rect 11437 35037 11471 35071
rect 11621 35037 11655 35071
rect 12455 35037 12489 35071
rect 12633 35037 12667 35071
rect 12725 35037 12759 35071
rect 12909 35037 12943 35071
rect 3350 34969 3384 35003
rect 4690 34969 4724 35003
rect 6469 34969 6503 35003
rect 10333 34969 10367 35003
rect 10425 34969 10459 35003
rect 4169 34901 4203 34935
rect 4353 34901 4387 34935
rect 10133 34901 10167 34935
rect 10701 34901 10735 34935
rect 3065 34697 3099 34731
rect 2605 34629 2639 34663
rect 12909 34629 12943 34663
rect 13185 34629 13219 34663
rect 7389 34561 7423 34595
rect 7573 34561 7607 34595
rect 12265 34561 12299 34595
rect 12541 34561 12575 34595
rect 12725 34561 12759 34595
rect 12817 34561 12851 34595
rect 13001 34561 13035 34595
rect 13093 34561 13127 34595
rect 13277 34561 13311 34595
rect 12173 34493 12207 34527
rect 12633 34493 12667 34527
rect 2881 34425 2915 34459
rect 7389 34357 7423 34391
rect 4629 34153 4663 34187
rect 5089 34153 5123 34187
rect 7205 34153 7239 34187
rect 7665 34153 7699 34187
rect 8217 34153 8251 34187
rect 10241 34153 10275 34187
rect 12449 34153 12483 34187
rect 4905 34085 4939 34119
rect 9229 34085 9263 34119
rect 10149 34085 10183 34119
rect 11805 34085 11839 34119
rect 6101 34017 6135 34051
rect 12357 34017 12391 34051
rect 14105 34017 14139 34051
rect 6929 33949 6963 33983
rect 7941 33949 7975 33983
rect 8217 33949 8251 33983
rect 9045 33949 9079 33983
rect 9505 33949 9539 33983
rect 9965 33949 9999 33983
rect 10149 33949 10183 33983
rect 10425 33949 10459 33983
rect 10793 33949 10827 33983
rect 11160 33949 11194 33983
rect 11253 33949 11287 33983
rect 12081 33949 12115 33983
rect 12633 33949 12667 33983
rect 12817 33949 12851 33983
rect 13185 33949 13219 33983
rect 13461 33949 13495 33983
rect 14361 33949 14395 33983
rect 4445 33881 4479 33915
rect 5057 33881 5091 33915
rect 5273 33881 5307 33915
rect 7189 33881 7223 33915
rect 7389 33881 7423 33915
rect 7649 33881 7683 33915
rect 7849 33881 7883 33915
rect 9321 33881 9355 33915
rect 10517 33881 10551 33915
rect 10609 33881 10643 33915
rect 10885 33881 10919 33915
rect 11989 33881 12023 33915
rect 12909 33881 12943 33915
rect 13277 33881 13311 33915
rect 13553 33881 13587 33915
rect 13737 33881 13771 33915
rect 13921 33881 13955 33915
rect 4645 33813 4679 33847
rect 4813 33813 4847 33847
rect 7021 33813 7055 33847
rect 7481 33813 7515 33847
rect 8033 33813 8067 33847
rect 12173 33813 12207 33847
rect 13093 33813 13127 33847
rect 15485 33813 15519 33847
rect 4537 33609 4571 33643
rect 11529 33609 11563 33643
rect 11713 33609 11747 33643
rect 2881 33473 2915 33507
rect 3137 33473 3171 33507
rect 4353 33473 4387 33507
rect 4537 33473 4571 33507
rect 4896 33473 4930 33507
rect 6929 33473 6963 33507
rect 7757 33473 7791 33507
rect 8401 33473 8435 33507
rect 8668 33473 8702 33507
rect 9873 33473 9907 33507
rect 10241 33473 10275 33507
rect 10793 33473 10827 33507
rect 11710 33473 11744 33507
rect 12081 33473 12115 33507
rect 13746 33473 13780 33507
rect 14013 33473 14047 33507
rect 4629 33405 4663 33439
rect 10057 33405 10091 33439
rect 12173 33405 12207 33439
rect 7665 33337 7699 33371
rect 9965 33337 9999 33371
rect 12633 33337 12667 33371
rect 4261 33269 4295 33303
rect 6009 33269 6043 33303
rect 9781 33269 9815 33303
rect 10057 33269 10091 33303
rect 10609 33269 10643 33303
rect 2973 33065 3007 33099
rect 3157 33065 3191 33099
rect 3801 33065 3835 33099
rect 8033 33065 8067 33099
rect 8769 33065 8803 33099
rect 9321 33065 9355 33099
rect 12817 33065 12851 33099
rect 13001 33065 13035 33099
rect 3525 32997 3559 33031
rect 9781 32997 9815 33031
rect 9965 32929 9999 32963
rect 10793 32929 10827 32963
rect 11161 32929 11195 32963
rect 11621 32929 11655 32963
rect 3985 32861 4019 32895
rect 4261 32861 4295 32895
rect 4629 32861 4663 32895
rect 5549 32861 5583 32895
rect 5733 32861 5767 32895
rect 6009 32861 6043 32895
rect 6653 32861 6687 32895
rect 6920 32861 6954 32895
rect 8125 32861 8159 32895
rect 8309 32861 8343 32895
rect 8401 32861 8435 32895
rect 8493 32861 8527 32895
rect 8953 32861 8987 32895
rect 9137 32861 9171 32895
rect 9229 32861 9263 32895
rect 10057 32861 10091 32895
rect 11253 32861 11287 32895
rect 12633 32861 12667 32895
rect 5917 32793 5951 32827
rect 9505 32793 9539 32827
rect 12969 32793 13003 32827
rect 13185 32793 13219 32827
rect 3157 32725 3191 32759
rect 4169 32725 4203 32759
rect 9137 32725 9171 32759
rect 3893 32521 3927 32555
rect 11345 32521 11379 32555
rect 3249 32453 3283 32487
rect 5733 32453 5767 32487
rect 12173 32453 12207 32487
rect 13001 32453 13035 32487
rect 3433 32385 3467 32419
rect 3985 32385 4019 32419
rect 4077 32385 4111 32419
rect 5273 32385 5307 32419
rect 5549 32385 5583 32419
rect 5825 32385 5859 32419
rect 10149 32385 10183 32419
rect 10977 32385 11011 32419
rect 11131 32385 11165 32419
rect 11621 32385 11655 32419
rect 4537 32317 4571 32351
rect 4261 32249 4295 32283
rect 3617 32181 3651 32215
rect 3709 32181 3743 32215
rect 5365 32181 5399 32215
rect 11713 32181 11747 32215
rect 4169 31977 4203 32011
rect 4813 31977 4847 32011
rect 3801 31909 3835 31943
rect 5733 31909 5767 31943
rect 5365 31841 5399 31875
rect 5825 31841 5859 31875
rect 7021 31841 7055 31875
rect 8585 31841 8619 31875
rect 10333 31841 10367 31875
rect 11161 31841 11195 31875
rect 12081 31841 12115 31875
rect 12541 31841 12575 31875
rect 13118 31841 13152 31875
rect 4445 31773 4479 31807
rect 4997 31773 5031 31807
rect 5181 31773 5215 31807
rect 5273 31773 5307 31807
rect 5549 31773 5583 31807
rect 6009 31773 6043 31807
rect 6193 31773 6227 31807
rect 6285 31773 6319 31807
rect 6929 31773 6963 31807
rect 8401 31773 8435 31807
rect 8493 31773 8527 31807
rect 8677 31773 8711 31807
rect 9413 31773 9447 31807
rect 9689 31773 9723 31807
rect 10241 31773 10275 31807
rect 10425 31773 10459 31807
rect 10537 31773 10571 31807
rect 10701 31773 10735 31807
rect 10793 31773 10827 31807
rect 10909 31773 10943 31807
rect 11436 31773 11470 31807
rect 11529 31773 11563 31807
rect 12173 31773 12207 31807
rect 12633 31773 12667 31807
rect 12909 31773 12943 31807
rect 13001 31773 13035 31807
rect 4169 31705 4203 31739
rect 4629 31705 4663 31739
rect 8033 31705 8067 31739
rect 9597 31705 9631 31739
rect 4353 31637 4387 31671
rect 6561 31637 6595 31671
rect 7941 31637 7975 31671
rect 8217 31637 8251 31671
rect 9229 31637 9263 31671
rect 9873 31637 9907 31671
rect 11069 31637 11103 31671
rect 13277 31637 13311 31671
rect 3341 31433 3375 31467
rect 4997 31433 5031 31467
rect 6193 31433 6227 31467
rect 7849 31433 7883 31467
rect 9321 31433 9355 31467
rect 4454 31365 4488 31399
rect 13360 31365 13394 31399
rect 5181 31297 5215 31331
rect 6009 31297 6043 31331
rect 6193 31297 6227 31331
rect 6469 31297 6503 31331
rect 6736 31297 6770 31331
rect 7941 31297 7975 31331
rect 8208 31297 8242 31331
rect 9873 31297 9907 31331
rect 10057 31297 10091 31331
rect 10149 31297 10183 31331
rect 4721 31229 4755 31263
rect 5457 31229 5491 31263
rect 13093 31229 13127 31263
rect 5365 31093 5399 31127
rect 9689 31093 9723 31127
rect 14473 31093 14507 31127
rect 6561 30889 6595 30923
rect 8217 30889 8251 30923
rect 9321 30889 9355 30923
rect 10609 30889 10643 30923
rect 9873 30821 9907 30855
rect 10057 30821 10091 30855
rect 12081 30821 12115 30855
rect 5457 30753 5491 30787
rect 6720 30753 6754 30787
rect 7205 30753 7239 30787
rect 7573 30753 7607 30787
rect 10425 30753 10459 30787
rect 11713 30753 11747 30787
rect 12541 30753 12575 30787
rect 14105 30753 14139 30787
rect 3801 30685 3835 30719
rect 3985 30685 4019 30719
rect 5273 30685 5307 30719
rect 8058 30685 8092 30719
rect 9446 30685 9480 30719
rect 9965 30685 9999 30719
rect 10241 30685 10275 30719
rect 10701 30685 10735 30719
rect 10977 30685 11011 30719
rect 11069 30685 11103 30719
rect 11253 30685 11287 30719
rect 11345 30685 11379 30719
rect 11805 30685 11839 30719
rect 12449 30685 12483 30719
rect 12817 30685 12851 30719
rect 13001 30685 13035 30719
rect 13093 30685 13127 30719
rect 13461 30685 13495 30719
rect 6929 30617 6963 30651
rect 7849 30617 7883 30651
rect 12909 30617 12943 30651
rect 13578 30617 13612 30651
rect 14350 30617 14384 30651
rect 3801 30549 3835 30583
rect 5089 30549 5123 30583
rect 6837 30549 6871 30583
rect 7941 30549 7975 30583
rect 9505 30549 9539 30583
rect 10793 30549 10827 30583
rect 11437 30549 11471 30583
rect 13369 30549 13403 30583
rect 13737 30549 13771 30583
rect 15485 30549 15519 30583
rect 5273 30345 5307 30379
rect 10885 30345 10919 30379
rect 13369 30345 13403 30379
rect 2973 30277 3007 30311
rect 3189 30277 3223 30311
rect 3433 30277 3467 30311
rect 3617 30277 3651 30311
rect 3801 30277 3835 30311
rect 12541 30277 12575 30311
rect 12633 30277 12667 30311
rect 13521 30277 13555 30311
rect 13737 30277 13771 30311
rect 14105 30277 14139 30311
rect 3893 30209 3927 30243
rect 4149 30209 4183 30243
rect 8493 30209 8527 30243
rect 8677 30209 8711 30243
rect 8953 30209 8987 30243
rect 9045 30209 9079 30243
rect 9229 30209 9263 30243
rect 9413 30209 9447 30243
rect 9689 30209 9723 30243
rect 11069 30209 11103 30243
rect 11253 30209 11287 30243
rect 11897 30209 11931 30243
rect 12081 30209 12115 30243
rect 12725 30209 12759 30243
rect 13829 30209 13863 30243
rect 13921 30209 13955 30243
rect 9505 30141 9539 30175
rect 3341 30073 3375 30107
rect 9137 30073 9171 30107
rect 12909 30073 12943 30107
rect 14105 30073 14139 30107
rect 3157 30005 3191 30039
rect 8493 30005 8527 30039
rect 8769 30005 8803 30039
rect 9413 30005 9447 30039
rect 9873 30005 9907 30039
rect 11253 30005 11287 30039
rect 11713 30005 11747 30039
rect 12081 30005 12115 30039
rect 12357 30005 12391 30039
rect 13553 30005 13587 30039
rect 8493 29801 8527 29835
rect 11345 29801 11379 29835
rect 5917 29733 5951 29767
rect 6745 29665 6779 29699
rect 7021 29665 7055 29699
rect 7481 29665 7515 29699
rect 8493 29665 8527 29699
rect 9781 29665 9815 29699
rect 10425 29665 10459 29699
rect 13553 29665 13587 29699
rect 2237 29597 2271 29631
rect 3985 29597 4019 29631
rect 4261 29597 4295 29631
rect 4905 29597 4939 29631
rect 4998 29597 5032 29631
rect 5181 29597 5215 29631
rect 5411 29597 5445 29631
rect 6192 29597 6226 29631
rect 6285 29597 6319 29631
rect 6653 29597 6687 29631
rect 7573 29597 7607 29631
rect 8585 29597 8619 29631
rect 9045 29597 9079 29631
rect 9505 29597 9539 29631
rect 10149 29597 10183 29631
rect 10517 29597 10551 29631
rect 10665 29597 10699 29631
rect 10793 29597 10827 29631
rect 10982 29597 11016 29631
rect 11253 29597 11287 29631
rect 11437 29597 11471 29631
rect 13185 29597 13219 29631
rect 13369 29597 13403 29631
rect 13461 29597 13495 29631
rect 13645 29597 13679 29631
rect 2504 29529 2538 29563
rect 5273 29529 5307 29563
rect 8309 29529 8343 29563
rect 10885 29529 10919 29563
rect 3617 29461 3651 29495
rect 3801 29461 3835 29495
rect 4169 29461 4203 29495
rect 5549 29461 5583 29495
rect 7941 29461 7975 29495
rect 8769 29461 8803 29495
rect 11161 29461 11195 29495
rect 13277 29461 13311 29495
rect 2513 29257 2547 29291
rect 2697 29257 2731 29291
rect 3417 29257 3451 29291
rect 6377 29257 6411 29291
rect 8401 29257 8435 29291
rect 8769 29257 8803 29291
rect 10609 29257 10643 29291
rect 10701 29257 10735 29291
rect 13093 29257 13127 29291
rect 13369 29257 13403 29291
rect 14841 29257 14875 29291
rect 3617 29189 3651 29223
rect 11529 29189 11563 29223
rect 12265 29189 12299 29223
rect 13706 29189 13740 29223
rect 4813 29121 4847 29155
rect 4997 29121 5031 29155
rect 5089 29121 5123 29155
rect 5365 29121 5399 29155
rect 7490 29121 7524 29155
rect 8309 29121 8343 29155
rect 8585 29121 8619 29155
rect 10241 29121 10275 29155
rect 10425 29121 10459 29155
rect 10977 29121 11011 29155
rect 11069 29121 11103 29155
rect 11161 29121 11195 29155
rect 11345 29121 11379 29155
rect 11805 29121 11839 29155
rect 11897 29121 11931 29155
rect 11989 29121 12023 29155
rect 12173 29121 12207 29155
rect 12540 29121 12574 29155
rect 12633 29121 12667 29155
rect 13001 29121 13035 29155
rect 5200 29053 5234 29087
rect 7757 29053 7791 29087
rect 12725 29053 12759 29087
rect 13210 29053 13244 29087
rect 13461 29053 13495 29087
rect 3065 28985 3099 29019
rect 3249 28985 3283 29019
rect 4905 28985 4939 29019
rect 2697 28917 2731 28951
rect 3433 28917 3467 28951
rect 4537 28713 4571 28747
rect 6193 28713 6227 28747
rect 7205 28713 7239 28747
rect 10517 28713 10551 28747
rect 10701 28713 10735 28747
rect 11161 28713 11195 28747
rect 13645 28645 13679 28679
rect 14105 28645 14139 28679
rect 6929 28577 6963 28611
rect 7046 28577 7080 28611
rect 12725 28577 12759 28611
rect 4077 28509 4111 28543
rect 4261 28509 4295 28543
rect 4721 28509 4755 28543
rect 4997 28509 5031 28543
rect 5089 28509 5123 28543
rect 5733 28509 5767 28543
rect 6285 28509 6319 28543
rect 6561 28509 6595 28543
rect 10241 28509 10275 28543
rect 10333 28509 10367 28543
rect 10609 28509 10643 28543
rect 10977 28509 11011 28543
rect 11805 28509 11839 28543
rect 13185 28509 13219 28543
rect 14289 28509 14323 28543
rect 5825 28441 5859 28475
rect 6009 28441 6043 28475
rect 6837 28441 6871 28475
rect 11897 28441 11931 28475
rect 13093 28441 13127 28475
rect 13645 28441 13679 28475
rect 4169 28373 4203 28407
rect 4905 28373 4939 28407
rect 6377 28373 6411 28407
rect 12909 28373 12943 28407
rect 3065 28169 3099 28203
rect 8769 28169 8803 28203
rect 10425 28169 10459 28203
rect 11529 28169 11563 28203
rect 13829 28169 13863 28203
rect 4721 28101 4755 28135
rect 8585 28101 8619 28135
rect 12716 28101 12750 28135
rect 3249 28033 3283 28067
rect 3525 28033 3559 28067
rect 3709 28033 3743 28067
rect 3985 28033 4019 28067
rect 4353 28033 4387 28067
rect 4445 28033 4479 28067
rect 6101 28033 6135 28067
rect 6193 28033 6227 28067
rect 6377 28033 6411 28067
rect 7113 28033 7147 28067
rect 7389 28033 7423 28067
rect 7573 28033 7607 28067
rect 8125 28033 8159 28067
rect 8309 28033 8343 28067
rect 9882 28033 9916 28067
rect 10609 28033 10643 28067
rect 10701 28033 10735 28067
rect 10977 28033 11011 28067
rect 11713 28033 11747 28067
rect 11897 28033 11931 28067
rect 3433 27965 3467 27999
rect 5457 27965 5491 27999
rect 5733 27965 5767 27999
rect 8217 27965 8251 27999
rect 10149 27965 10183 27999
rect 10885 27965 10919 27999
rect 11989 27965 12023 27999
rect 12449 27965 12483 27999
rect 3893 27829 3927 27863
rect 4077 27829 4111 27863
rect 4629 27829 4663 27863
rect 5917 27829 5951 27863
rect 6929 27829 6963 27863
rect 7573 27829 7607 27863
rect 8493 27829 8527 27863
rect 3617 27625 3651 27659
rect 8217 27625 8251 27659
rect 8585 27625 8619 27659
rect 8769 27557 8803 27591
rect 9597 27557 9631 27591
rect 9689 27557 9723 27591
rect 2237 27489 2271 27523
rect 6837 27489 6871 27523
rect 10149 27489 10183 27523
rect 11345 27489 11379 27523
rect 5641 27421 5675 27455
rect 6285 27421 6319 27455
rect 8953 27421 8987 27455
rect 9229 27421 9263 27455
rect 9965 27421 9999 27455
rect 11897 27421 11931 27455
rect 2504 27353 2538 27387
rect 3985 27353 4019 27387
rect 5396 27353 5430 27387
rect 5733 27353 5767 27387
rect 7104 27353 7138 27387
rect 8401 27353 8435 27387
rect 8617 27353 8651 27387
rect 9438 27353 9472 27387
rect 9689 27353 9723 27387
rect 10977 27353 11011 27387
rect 11529 27353 11563 27387
rect 4077 27285 4111 27319
rect 4261 27285 4295 27319
rect 9321 27285 9355 27319
rect 9873 27285 9907 27319
rect 11621 27285 11655 27319
rect 11713 27285 11747 27319
rect 2697 27081 2731 27115
rect 2881 27081 2915 27115
rect 3985 27081 4019 27115
rect 4277 27081 4311 27115
rect 4445 27081 4479 27115
rect 7573 27081 7607 27115
rect 7849 27081 7883 27115
rect 7941 27081 7975 27115
rect 8309 27081 8343 27115
rect 8677 27081 8711 27115
rect 9045 27081 9079 27115
rect 12817 27081 12851 27115
rect 13093 27081 13127 27115
rect 3617 27013 3651 27047
rect 4077 27013 4111 27047
rect 4782 27013 4816 27047
rect 6561 27013 6595 27047
rect 14298 27013 14332 27047
rect 1685 26945 1719 26979
rect 3249 26945 3283 26979
rect 3801 26945 3835 26979
rect 4537 26945 4571 26979
rect 7732 26945 7766 26979
rect 8493 26945 8527 26979
rect 8585 26945 8619 26979
rect 8861 26945 8895 26979
rect 8953 26945 8987 26979
rect 9137 26945 9171 26979
rect 10149 26945 10183 26979
rect 11897 26945 11931 26979
rect 12081 26945 12115 26979
rect 14565 26945 14599 26979
rect 7297 26877 7331 26911
rect 8217 26877 8251 26911
rect 12449 26877 12483 26911
rect 12725 26877 12759 26911
rect 12934 26877 12968 26911
rect 13185 26809 13219 26843
rect 1501 26741 1535 26775
rect 2881 26741 2915 26775
rect 4261 26741 4295 26775
rect 5917 26741 5951 26775
rect 12081 26741 12115 26775
rect 11621 26537 11655 26571
rect 11805 26537 11839 26571
rect 12081 26537 12115 26571
rect 13185 26537 13219 26571
rect 5273 26469 5307 26503
rect 8953 26401 8987 26435
rect 10333 26401 10367 26435
rect 10425 26401 10459 26435
rect 12725 26401 12759 26435
rect 4721 26333 4755 26367
rect 5549 26333 5583 26367
rect 6101 26333 6135 26367
rect 9137 26333 9171 26367
rect 10057 26333 10091 26367
rect 10793 26333 10827 26367
rect 10977 26333 11011 26367
rect 11161 26333 11195 26367
rect 11345 26333 11379 26367
rect 12265 26333 12299 26367
rect 12357 26333 12391 26367
rect 12817 26333 12851 26367
rect 5273 26265 5307 26299
rect 5457 26265 5491 26299
rect 6368 26265 6402 26299
rect 10542 26265 10576 26299
rect 10885 26265 10919 26299
rect 11253 26265 11287 26299
rect 11789 26265 11823 26299
rect 11989 26265 12023 26299
rect 12081 26265 12115 26299
rect 7481 26197 7515 26231
rect 10701 26197 10735 26231
rect 3893 25993 3927 26027
rect 4077 25993 4111 26027
rect 6561 25993 6595 26027
rect 9229 25993 9263 26027
rect 11345 25993 11379 26027
rect 13093 25993 13127 26027
rect 6377 25925 6411 25959
rect 9137 25925 9171 25959
rect 10232 25925 10266 25959
rect 6653 25857 6687 25891
rect 7757 25857 7791 25891
rect 7941 25857 7975 25891
rect 8401 25857 8435 25891
rect 9346 25857 9380 25891
rect 9965 25857 9999 25891
rect 11713 25857 11747 25891
rect 11980 25857 12014 25891
rect 4445 25789 4479 25823
rect 4629 25789 4663 25823
rect 5641 25789 5675 25823
rect 7665 25789 7699 25823
rect 8493 25789 8527 25823
rect 8769 25789 8803 25823
rect 8861 25789 8895 25823
rect 6377 25721 6411 25755
rect 4077 25653 4111 25687
rect 5273 25653 5307 25687
rect 6193 25653 6227 25687
rect 7021 25653 7055 25687
rect 7849 25653 7883 25687
rect 9505 25653 9539 25687
rect 10609 25449 10643 25483
rect 12173 25449 12207 25483
rect 7849 25381 7883 25415
rect 7665 25313 7699 25347
rect 11529 25313 11563 25347
rect 12014 25313 12048 25347
rect 4925 25245 4959 25279
rect 5181 25245 5215 25279
rect 5733 25245 5767 25279
rect 6000 25245 6034 25279
rect 7297 25245 7331 25279
rect 7573 25245 7607 25279
rect 8493 25245 8527 25279
rect 8953 25245 8987 25279
rect 9137 25245 9171 25279
rect 9229 25245 9263 25279
rect 11805 25245 11839 25279
rect 5457 25177 5491 25211
rect 5641 25177 5675 25211
rect 7205 25177 7239 25211
rect 7941 25177 7975 25211
rect 9496 25177 9530 25211
rect 3801 25109 3835 25143
rect 5273 25109 5307 25143
rect 7113 25109 7147 25143
rect 8953 25109 8987 25143
rect 11897 25109 11931 25143
rect 4169 24905 4203 24939
rect 5641 24905 5675 24939
rect 7941 24905 7975 24939
rect 5293 24769 5327 24803
rect 6009 24769 6043 24803
rect 7665 24769 7699 24803
rect 8289 24769 8323 24803
rect 5549 24701 5583 24735
rect 5917 24701 5951 24735
rect 6561 24701 6595 24735
rect 7297 24701 7331 24735
rect 7389 24701 7423 24735
rect 7757 24701 7791 24735
rect 8033 24701 8067 24735
rect 9413 24633 9447 24667
rect 7205 24565 7239 24599
rect 5457 24361 5491 24395
rect 6469 24361 6503 24395
rect 6561 24361 6595 24395
rect 8125 24361 8159 24395
rect 8217 24361 8251 24395
rect 5733 24293 5767 24327
rect 9229 24293 9263 24327
rect 4077 24225 4111 24259
rect 5825 24225 5859 24259
rect 8309 24225 8343 24259
rect 11621 24225 11655 24259
rect 11713 24225 11747 24259
rect 5641 24157 5675 24191
rect 5917 24157 5951 24191
rect 6101 24157 6135 24191
rect 6285 24157 6319 24191
rect 6377 24157 6411 24191
rect 6653 24157 6687 24191
rect 6745 24157 6779 24191
rect 8217 24157 8251 24191
rect 10425 24157 10459 24191
rect 11989 24157 12023 24191
rect 12081 24157 12115 24191
rect 12173 24157 12207 24191
rect 12357 24157 12391 24191
rect 7012 24089 7046 24123
rect 9045 24089 9079 24123
rect 4721 24021 4755 24055
rect 8585 24021 8619 24055
rect 9873 24021 9907 24055
rect 10977 24021 11011 24055
rect 4445 23817 4479 23851
rect 8033 23817 8067 23851
rect 11069 23817 11103 23851
rect 7665 23749 7699 23783
rect 3065 23681 3099 23715
rect 3321 23681 3355 23715
rect 7849 23681 7883 23715
rect 8125 23681 8159 23715
rect 8217 23681 8251 23715
rect 8401 23681 8435 23715
rect 9505 23681 9539 23715
rect 9772 23681 9806 23715
rect 10977 23681 11011 23715
rect 11161 23681 11195 23715
rect 13021 23681 13055 23715
rect 13277 23681 13311 23715
rect 8401 23545 8435 23579
rect 10885 23545 10919 23579
rect 7481 23477 7515 23511
rect 11897 23477 11931 23511
rect 3157 23273 3191 23307
rect 11897 23273 11931 23307
rect 11989 23273 12023 23307
rect 13277 23273 13311 23307
rect 3065 23137 3099 23171
rect 3801 23137 3835 23171
rect 12541 23137 12575 23171
rect 3341 23069 3375 23103
rect 3525 23069 3559 23103
rect 3617 23069 3651 23103
rect 5825 23069 5859 23103
rect 6653 23069 6687 23103
rect 8953 23069 8987 23103
rect 10517 23069 10551 23103
rect 10784 23069 10818 23103
rect 12725 23069 12759 23103
rect 13093 23069 13127 23103
rect 2820 23001 2854 23035
rect 4046 23001 4080 23035
rect 9220 23001 9254 23035
rect 12909 23001 12943 23035
rect 13001 23001 13035 23035
rect 1685 22933 1719 22967
rect 5181 22933 5215 22967
rect 5273 22933 5307 22967
rect 6101 22933 6135 22967
rect 10333 22933 10367 22967
rect 3617 22729 3651 22763
rect 6469 22729 6503 22763
rect 9873 22729 9907 22763
rect 11713 22729 11747 22763
rect 12265 22729 12299 22763
rect 3249 22661 3283 22695
rect 3785 22661 3819 22695
rect 3985 22661 4019 22695
rect 1501 22593 1535 22627
rect 3433 22593 3467 22627
rect 3525 22593 3559 22627
rect 4077 22593 4111 22627
rect 4813 22593 4847 22627
rect 4997 22593 5031 22627
rect 5917 22593 5951 22627
rect 6009 22593 6043 22627
rect 6469 22593 6503 22627
rect 6653 22593 6687 22627
rect 7481 22593 7515 22627
rect 7665 22593 7699 22627
rect 8493 22593 8527 22627
rect 8760 22593 8794 22627
rect 11621 22593 11655 22627
rect 11805 22593 11839 22627
rect 12173 22593 12207 22627
rect 12357 22593 12391 22627
rect 16221 22593 16255 22627
rect 4721 22525 4755 22559
rect 4905 22525 4939 22559
rect 5825 22525 5859 22559
rect 6101 22525 6135 22559
rect 6745 22525 6779 22559
rect 8401 22525 8435 22559
rect 12909 22525 12943 22559
rect 1685 22457 1719 22491
rect 3249 22457 3283 22491
rect 7757 22457 7791 22491
rect 13185 22457 13219 22491
rect 16405 22457 16439 22491
rect 3801 22389 3835 22423
rect 5641 22389 5675 22423
rect 7389 22389 7423 22423
rect 7573 22389 7607 22423
rect 13369 22389 13403 22423
rect 9873 22185 9907 22219
rect 16129 22185 16163 22219
rect 8769 22117 8803 22151
rect 12449 22117 12483 22151
rect 7389 22049 7423 22083
rect 10149 22049 10183 22083
rect 1409 21981 1443 22015
rect 1685 21981 1719 22015
rect 2881 21981 2915 22015
rect 5365 21981 5399 22015
rect 7021 21981 7055 22015
rect 7205 21981 7239 22015
rect 7294 21981 7328 22015
rect 9505 21981 9539 22015
rect 11621 21981 11655 22015
rect 11805 21981 11839 22015
rect 12357 21981 12391 22015
rect 13829 21981 13863 22015
rect 15945 21981 15979 22015
rect 16221 21981 16255 22015
rect 5632 21913 5666 21947
rect 6837 21913 6871 21947
rect 7656 21913 7690 21947
rect 9873 21913 9907 21947
rect 10416 21913 10450 21947
rect 11713 21913 11747 21947
rect 13562 21913 13596 21947
rect 2329 21845 2363 21879
rect 6745 21845 6779 21879
rect 10057 21845 10091 21879
rect 11529 21845 11563 21879
rect 12265 21845 12299 21879
rect 16405 21845 16439 21879
rect 2697 21641 2731 21675
rect 6101 21641 6135 21675
rect 7665 21641 7699 21675
rect 11345 21641 11379 21675
rect 11897 21641 11931 21675
rect 12173 21641 12207 21675
rect 12449 21641 12483 21675
rect 4988 21573 5022 21607
rect 7113 21573 7147 21607
rect 7849 21573 7883 21607
rect 13185 21573 13219 21607
rect 1685 21505 1719 21539
rect 2053 21505 2087 21539
rect 2789 21505 2823 21539
rect 3056 21505 3090 21539
rect 4261 21505 4295 21539
rect 4445 21505 4479 21539
rect 4721 21505 4755 21539
rect 6377 21505 6411 21539
rect 6561 21505 6595 21539
rect 6929 21505 6963 21539
rect 7389 21505 7423 21539
rect 7757 21505 7791 21539
rect 9689 21505 9723 21539
rect 9873 21505 9907 21539
rect 9965 21505 9999 21539
rect 11161 21505 11195 21539
rect 13553 21505 13587 21539
rect 14381 21505 14415 21539
rect 14648 21505 14682 21539
rect 1961 21437 1995 21471
rect 7665 21437 7699 21471
rect 10885 21437 10919 21471
rect 11529 21437 11563 21471
rect 11805 21437 11839 21471
rect 12014 21437 12048 21471
rect 13001 21437 13035 21471
rect 13369 21437 13403 21471
rect 16405 21437 16439 21471
rect 1777 21369 1811 21403
rect 6745 21369 6779 21403
rect 10333 21369 10367 21403
rect 10977 21369 11011 21403
rect 13461 21369 13495 21403
rect 15761 21369 15795 21403
rect 1869 21301 1903 21335
rect 4169 21301 4203 21335
rect 4261 21301 4295 21335
rect 6561 21301 6595 21335
rect 7297 21301 7331 21335
rect 7481 21301 7515 21335
rect 13369 21301 13403 21335
rect 15853 21301 15887 21335
rect 2789 21097 2823 21131
rect 3065 21097 3099 21131
rect 3249 21097 3283 21131
rect 3985 21097 4019 21131
rect 4629 21097 4663 21131
rect 4813 21097 4847 21131
rect 5825 21097 5859 21131
rect 6285 21097 6319 21131
rect 8585 21097 8619 21131
rect 10241 21097 10275 21131
rect 11805 21097 11839 21131
rect 12449 21097 12483 21131
rect 12909 21097 12943 21131
rect 13461 21097 13495 21131
rect 14841 21097 14875 21131
rect 16129 21097 16163 21131
rect 2973 21029 3007 21063
rect 6469 21029 6503 21063
rect 12817 21029 12851 21063
rect 13277 21029 13311 21063
rect 3157 20961 3191 20995
rect 13001 20961 13035 20995
rect 15393 20961 15427 20995
rect 1409 20893 1443 20927
rect 2881 20893 2915 20927
rect 3433 20893 3467 20927
rect 3617 20893 3651 20927
rect 4169 20893 4203 20927
rect 4537 20893 4571 20927
rect 4813 20893 4847 20927
rect 4997 20893 5031 20927
rect 5549 20893 5583 20927
rect 5733 20893 5767 20927
rect 6101 20893 6135 20927
rect 6377 20893 6411 20927
rect 7021 20893 7055 20927
rect 7297 20893 7331 20927
rect 7389 20893 7423 20927
rect 7573 20893 7607 20927
rect 8953 20893 8987 20927
rect 11713 20893 11747 20927
rect 12909 20893 12943 20927
rect 13369 20893 13403 20927
rect 13553 20893 13587 20927
rect 14105 20893 14139 20927
rect 14198 20893 14232 20927
rect 15209 20893 15243 20927
rect 15945 20893 15979 20927
rect 1654 20825 1688 20859
rect 4379 20825 4413 20859
rect 8401 20825 8435 20859
rect 5733 20757 5767 20791
rect 8601 20757 8635 20791
rect 8769 20757 8803 20791
rect 12265 20757 12299 20791
rect 12449 20757 12483 20791
rect 14473 20757 14507 20791
rect 15301 20757 15335 20791
rect 1501 20553 1535 20587
rect 3433 20553 3467 20587
rect 6193 20553 6227 20587
rect 6469 20553 6503 20587
rect 7021 20553 7055 20587
rect 8585 20553 8619 20587
rect 9889 20553 9923 20587
rect 14197 20553 14231 20587
rect 1777 20485 1811 20519
rect 1869 20485 1903 20519
rect 2007 20485 2041 20519
rect 9689 20485 9723 20519
rect 1685 20417 1719 20451
rect 2145 20417 2179 20451
rect 2513 20417 2547 20451
rect 2789 20417 2823 20451
rect 2973 20417 3007 20451
rect 3065 20417 3099 20451
rect 3709 20417 3743 20451
rect 4813 20417 4847 20451
rect 5080 20417 5114 20451
rect 6377 20417 6411 20451
rect 6653 20417 6687 20451
rect 6929 20417 6963 20451
rect 7113 20417 7147 20451
rect 7472 20417 7506 20451
rect 11529 20417 11563 20451
rect 13093 20417 13127 20451
rect 13277 20417 13311 20451
rect 13553 20417 13587 20451
rect 13737 20417 13771 20451
rect 13829 20417 13863 20451
rect 13921 20417 13955 20451
rect 14565 20417 14599 20451
rect 2881 20349 2915 20383
rect 3433 20349 3467 20383
rect 4629 20349 4663 20383
rect 6837 20349 6871 20383
rect 7205 20349 7239 20383
rect 9413 20349 9447 20383
rect 10149 20349 10183 20383
rect 11805 20349 11839 20383
rect 16221 20349 16255 20383
rect 2329 20281 2363 20315
rect 3249 20281 3283 20315
rect 10057 20281 10091 20315
rect 3617 20213 3651 20247
rect 4077 20213 4111 20247
rect 8861 20213 8895 20247
rect 9873 20213 9907 20247
rect 10793 20213 10827 20247
rect 11621 20213 11655 20247
rect 11713 20213 11747 20247
rect 13369 20213 13403 20247
rect 14381 20213 14415 20247
rect 15669 20213 15703 20247
rect 1593 20009 1627 20043
rect 5181 20009 5215 20043
rect 6193 20009 6227 20043
rect 6469 20009 6503 20043
rect 7757 20009 7791 20043
rect 8677 20009 8711 20043
rect 9137 20009 9171 20043
rect 15945 20009 15979 20043
rect 7481 19941 7515 19975
rect 11621 19941 11655 19975
rect 3157 19873 3191 19907
rect 3801 19873 3835 19907
rect 7389 19873 7423 19907
rect 11069 19873 11103 19907
rect 11253 19873 11287 19907
rect 13093 19873 13127 19907
rect 13369 19873 13403 19907
rect 1501 19805 1535 19839
rect 1961 19805 1995 19839
rect 2145 19805 2179 19839
rect 2329 19805 2363 19839
rect 3249 19805 3283 19839
rect 6101 19805 6135 19839
rect 6285 19805 6319 19839
rect 6653 19805 6687 19839
rect 6745 19805 6779 19839
rect 6929 19805 6963 19839
rect 7021 19805 7055 19839
rect 7113 19805 7147 19839
rect 7297 19805 7331 19839
rect 7573 19805 7607 19839
rect 8769 19805 8803 19839
rect 10517 19805 10551 19839
rect 11437 19805 11471 19839
rect 11805 19805 11839 19839
rect 11989 19805 12023 19839
rect 13001 19805 13035 19839
rect 13185 19805 13219 19839
rect 13277 19805 13311 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 14565 19805 14599 19839
rect 4046 19737 4080 19771
rect 10272 19737 10306 19771
rect 10977 19737 11011 19771
rect 14832 19737 14866 19771
rect 2145 19669 2179 19703
rect 2881 19669 2915 19703
rect 3617 19669 3651 19703
rect 10609 19669 10643 19703
rect 11897 19669 11931 19703
rect 13829 19669 13863 19703
rect 3157 19465 3191 19499
rect 3249 19465 3283 19499
rect 7021 19465 7055 19499
rect 7389 19465 7423 19499
rect 9229 19465 9263 19499
rect 11345 19465 11379 19499
rect 11529 19465 11563 19499
rect 11989 19465 12023 19499
rect 13369 19465 13403 19499
rect 13921 19465 13955 19499
rect 14933 19465 14967 19499
rect 15301 19465 15335 19499
rect 1676 19397 1710 19431
rect 3709 19397 3743 19431
rect 9873 19397 9907 19431
rect 10232 19397 10266 19431
rect 14565 19397 14599 19431
rect 1409 19329 1443 19363
rect 3617 19329 3651 19363
rect 3801 19329 3835 19363
rect 7481 19329 7515 19363
rect 7849 19329 7883 19363
rect 8116 19329 8150 19363
rect 9689 19329 9723 19363
rect 11897 19329 11931 19363
rect 12909 19329 12943 19363
rect 13185 19329 13219 19363
rect 13553 19329 13587 19363
rect 13737 19329 13771 19363
rect 14289 19329 14323 19363
rect 14381 19329 14415 19363
rect 3040 19261 3074 19295
rect 3525 19261 3559 19295
rect 7573 19261 7607 19295
rect 9965 19261 9999 19295
rect 12081 19261 12115 19295
rect 13093 19261 13127 19295
rect 14197 19261 14231 19295
rect 15393 19261 15427 19295
rect 15485 19261 15519 19295
rect 13001 19193 13035 19227
rect 13553 19193 13587 19227
rect 14749 19193 14783 19227
rect 2789 19125 2823 19159
rect 2881 19125 2915 19159
rect 9597 19125 9631 19159
rect 14289 19125 14323 19159
rect 2237 18921 2271 18955
rect 2329 18921 2363 18955
rect 6745 18921 6779 18955
rect 8033 18921 8067 18955
rect 12081 18921 12115 18955
rect 13369 18921 13403 18955
rect 13645 18921 13679 18955
rect 15025 18921 15059 18955
rect 6653 18853 6687 18887
rect 2421 18785 2455 18819
rect 2513 18785 2547 18819
rect 5273 18785 5307 18819
rect 7297 18785 7331 18819
rect 8677 18785 8711 18819
rect 9597 18785 9631 18819
rect 14473 18785 14507 18819
rect 14565 18785 14599 18819
rect 2145 18717 2179 18751
rect 3065 18717 3099 18751
rect 8493 18717 8527 18751
rect 9321 18717 9355 18751
rect 10793 18717 10827 18751
rect 11437 18717 11471 18751
rect 12357 18717 12391 18751
rect 12541 18717 12575 18751
rect 13277 18717 13311 18751
rect 13369 18717 13403 18751
rect 5540 18649 5574 18683
rect 8401 18649 8435 18683
rect 9413 18649 9447 18683
rect 12265 18649 12299 18683
rect 8953 18581 8987 18615
rect 11897 18581 11931 18615
rect 12065 18581 12099 18615
rect 12449 18581 12483 18615
rect 14657 18581 14691 18615
rect 2973 18377 3007 18411
rect 5089 18377 5123 18411
rect 5457 18377 5491 18411
rect 5825 18377 5859 18411
rect 6469 18377 6503 18411
rect 7497 18377 7531 18411
rect 9505 18377 9539 18411
rect 11529 18377 11563 18411
rect 13645 18377 13679 18411
rect 14933 18377 14967 18411
rect 5917 18309 5951 18343
rect 7297 18309 7331 18343
rect 10640 18309 10674 18343
rect 11805 18309 11839 18343
rect 11897 18309 11931 18343
rect 12265 18309 12299 18343
rect 2053 18241 2087 18275
rect 2605 18241 2639 18275
rect 2789 18241 2823 18275
rect 3709 18241 3743 18275
rect 3976 18241 4010 18275
rect 6837 18241 6871 18275
rect 6929 18241 6963 18275
rect 11713 18241 11747 18275
rect 12081 18241 12115 18275
rect 12449 18241 12483 18275
rect 12541 18241 12575 18275
rect 12725 18241 12759 18275
rect 12817 18241 12851 18275
rect 13277 18241 13311 18275
rect 13737 18241 13771 18275
rect 13921 18241 13955 18275
rect 14105 18241 14139 18275
rect 14381 18241 14415 18275
rect 14565 18241 14599 18275
rect 14657 18241 14691 18275
rect 14749 18241 14783 18275
rect 2145 18173 2179 18207
rect 2237 18173 2271 18207
rect 6101 18173 6135 18207
rect 7113 18173 7147 18207
rect 10885 18173 10919 18207
rect 13369 18173 13403 18207
rect 1685 18037 1719 18071
rect 2789 18037 2823 18071
rect 7481 18037 7515 18071
rect 7665 18037 7699 18071
rect 13461 18037 13495 18071
rect 2789 17833 2823 17867
rect 3341 17833 3375 17867
rect 3525 17833 3559 17867
rect 3893 17833 3927 17867
rect 8217 17833 8251 17867
rect 12909 17833 12943 17867
rect 13093 17833 13127 17867
rect 1409 17697 1443 17731
rect 4445 17697 4479 17731
rect 6653 17697 6687 17731
rect 14473 17697 14507 17731
rect 4353 17629 4387 17663
rect 8033 17629 8067 17663
rect 8217 17629 8251 17663
rect 12081 17629 12115 17663
rect 12265 17629 12299 17663
rect 14197 17629 14231 17663
rect 14289 17629 14323 17663
rect 14749 17629 14783 17663
rect 16405 17629 16439 17663
rect 12955 17595 12989 17629
rect 1676 17561 1710 17595
rect 3157 17561 3191 17595
rect 4261 17561 4295 17595
rect 7757 17561 7791 17595
rect 11897 17561 11931 17595
rect 12725 17561 12759 17595
rect 3357 17493 3391 17527
rect 7205 17493 7239 17527
rect 8401 17493 8435 17527
rect 14657 17493 14691 17527
rect 15853 17493 15887 17527
rect 1869 17289 1903 17323
rect 6193 17289 6227 17323
rect 6377 17289 6411 17323
rect 6745 17289 6779 17323
rect 7573 17289 7607 17323
rect 8309 17289 8343 17323
rect 8953 17289 8987 17323
rect 11253 17289 11287 17323
rect 12909 17289 12943 17323
rect 13277 17289 13311 17323
rect 16129 17289 16163 17323
rect 3801 17221 3835 17255
rect 4001 17221 4035 17255
rect 5080 17221 5114 17255
rect 8493 17221 8527 17255
rect 11897 17221 11931 17255
rect 14197 17221 14231 17255
rect 2237 17153 2271 17187
rect 2329 17153 2363 17187
rect 2596 17153 2630 17187
rect 7849 17153 7883 17187
rect 7941 17153 7975 17187
rect 8033 17153 8067 17187
rect 8217 17153 8251 17187
rect 8861 17153 8895 17187
rect 10140 17153 10174 17187
rect 11529 17153 11563 17187
rect 11713 17153 11747 17187
rect 11805 17153 11839 17187
rect 12015 17153 12049 17187
rect 12173 17153 12207 17187
rect 12449 17153 12483 17187
rect 13001 17153 13035 17187
rect 13093 17153 13127 17187
rect 14013 17153 14047 17187
rect 14289 17153 14323 17187
rect 14381 17153 14415 17187
rect 14749 17153 14783 17187
rect 15016 17153 15050 17187
rect 16221 17153 16255 17187
rect 2145 17085 2179 17119
rect 4813 17085 4847 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 9413 17085 9447 17119
rect 9873 17085 9907 17119
rect 13277 17085 13311 17119
rect 9137 17017 9171 17051
rect 12817 17017 12851 17051
rect 16405 17017 16439 17051
rect 2053 16949 2087 16983
rect 3709 16949 3743 16983
rect 3985 16949 4019 16983
rect 4169 16949 4203 16983
rect 8493 16949 8527 16983
rect 14565 16949 14599 16983
rect 2881 16745 2915 16779
rect 3525 16745 3559 16779
rect 7573 16745 7607 16779
rect 11989 16745 12023 16779
rect 13093 16745 13127 16779
rect 15117 16745 15151 16779
rect 16129 16745 16163 16779
rect 7205 16677 7239 16711
rect 8125 16677 8159 16711
rect 11253 16677 11287 16711
rect 2789 16609 2823 16643
rect 3985 16609 4019 16643
rect 9597 16609 9631 16643
rect 9873 16609 9907 16643
rect 11345 16609 11379 16643
rect 13277 16609 13311 16643
rect 13921 16609 13955 16643
rect 14473 16609 14507 16643
rect 14841 16609 14875 16643
rect 15669 16609 15703 16643
rect 3065 16541 3099 16575
rect 3157 16541 3191 16575
rect 3433 16541 3467 16575
rect 7113 16541 7147 16575
rect 10140 16541 10174 16575
rect 11529 16541 11563 16575
rect 11621 16541 11655 16575
rect 11805 16541 11839 16575
rect 11897 16541 11931 16575
rect 12173 16541 12207 16575
rect 12357 16541 12391 16575
rect 12449 16541 12483 16575
rect 12633 16541 12667 16575
rect 13001 16541 13035 16575
rect 13553 16541 13587 16575
rect 14105 16541 14139 16575
rect 14289 16541 14323 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 15485 16541 15519 16575
rect 15945 16541 15979 16575
rect 2421 16473 2455 16507
rect 2605 16473 2639 16507
rect 4230 16473 4264 16507
rect 7573 16473 7607 16507
rect 8493 16473 8527 16507
rect 13737 16473 13771 16507
rect 15577 16473 15611 16507
rect 5365 16405 5399 16439
rect 6469 16405 6503 16439
rect 7757 16405 7791 16439
rect 8033 16405 8067 16439
rect 8953 16405 8987 16439
rect 9321 16405 9355 16439
rect 9413 16405 9447 16439
rect 12541 16405 12575 16439
rect 13277 16405 13311 16439
rect 4077 16201 4111 16235
rect 7757 16201 7791 16235
rect 7849 16201 7883 16235
rect 9873 16201 9907 16235
rect 9965 16201 9999 16235
rect 12081 16201 12115 16235
rect 13619 16201 13653 16235
rect 4537 16133 4571 16167
rect 8309 16133 8343 16167
rect 8760 16133 8794 16167
rect 12817 16133 12851 16167
rect 13829 16133 13863 16167
rect 4445 16065 4479 16099
rect 6377 16065 6411 16099
rect 6644 16065 6678 16099
rect 8033 16065 8067 16099
rect 10517 16065 10551 16099
rect 11713 16065 11747 16099
rect 15577 16065 15611 16099
rect 16405 16065 16439 16099
rect 4629 15997 4663 16031
rect 8125 15997 8159 16031
rect 8493 15997 8527 16031
rect 12265 15929 12299 15963
rect 12449 15929 12483 15963
rect 8309 15861 8343 15895
rect 12081 15861 12115 15895
rect 12357 15861 12391 15895
rect 13461 15861 13495 15895
rect 13645 15861 13679 15895
rect 15761 15861 15795 15895
rect 15853 15861 15887 15895
rect 3157 15657 3191 15691
rect 6929 15657 6963 15691
rect 8953 15657 8987 15691
rect 9137 15657 9171 15691
rect 9413 15657 9447 15691
rect 12265 15657 12299 15691
rect 13921 15657 13955 15691
rect 16129 15657 16163 15691
rect 16405 15657 16439 15691
rect 3617 15589 3651 15623
rect 2237 15521 2271 15555
rect 2421 15521 2455 15555
rect 4629 15521 4663 15555
rect 6285 15521 6319 15555
rect 6469 15521 6503 15555
rect 7941 15521 7975 15555
rect 8125 15521 8159 15555
rect 9965 15521 9999 15555
rect 14749 15521 14783 15555
rect 2053 15453 2087 15487
rect 2329 15453 2363 15487
rect 2513 15453 2547 15487
rect 2605 15453 2639 15487
rect 2789 15453 2823 15487
rect 3065 15453 3099 15487
rect 3341 15453 3375 15487
rect 4445 15453 4479 15487
rect 9873 15453 9907 15487
rect 11345 15453 11379 15487
rect 11989 15453 12023 15487
rect 13185 15453 13219 15487
rect 13369 15453 13403 15487
rect 13461 15453 13495 15487
rect 13553 15453 13587 15487
rect 13737 15453 13771 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 14381 15453 14415 15487
rect 14473 15453 14507 15487
rect 16221 15453 16255 15487
rect 2697 15385 2731 15419
rect 9321 15385 9355 15419
rect 12081 15385 12115 15419
rect 12281 15385 12315 15419
rect 15016 15385 15050 15419
rect 1869 15317 1903 15351
rect 4077 15317 4111 15351
rect 4537 15317 4571 15351
rect 6561 15317 6595 15351
rect 7389 15317 7423 15351
rect 8769 15317 8803 15351
rect 9121 15317 9155 15351
rect 9781 15317 9815 15351
rect 12449 15317 12483 15351
rect 14657 15317 14691 15351
rect 2973 15113 3007 15147
rect 5549 15113 5583 15147
rect 7757 15113 7791 15147
rect 7941 15113 7975 15147
rect 9965 15113 9999 15147
rect 13093 15113 13127 15147
rect 14013 15113 14047 15147
rect 15117 15113 15151 15147
rect 15485 15113 15519 15147
rect 11100 15045 11134 15079
rect 11529 15045 11563 15079
rect 13461 15045 13495 15079
rect 13645 15045 13679 15079
rect 15577 15045 15611 15079
rect 1593 14977 1627 15011
rect 1860 14977 1894 15011
rect 3433 14977 3467 15011
rect 3709 14977 3743 15011
rect 4169 14977 4203 15011
rect 4425 14977 4459 15011
rect 6377 14977 6411 15011
rect 6644 14977 6678 15011
rect 9054 14977 9088 15011
rect 11345 14977 11379 15011
rect 11713 14977 11747 15011
rect 11805 14977 11839 15011
rect 11989 14977 12023 15011
rect 12357 14977 12391 15011
rect 12633 14977 12667 15011
rect 13001 14977 13035 15011
rect 13277 14977 13311 15011
rect 13553 14977 13587 15011
rect 13829 14977 13863 15011
rect 15945 14977 15979 15011
rect 9321 14909 9355 14943
rect 12173 14909 12207 14943
rect 12449 14909 12483 14943
rect 12541 14909 12575 14943
rect 15669 14909 15703 14943
rect 3985 14841 4019 14875
rect 11897 14841 11931 14875
rect 3525 14773 3559 14807
rect 16129 14773 16163 14807
rect 1777 14569 1811 14603
rect 2697 14569 2731 14603
rect 3157 14569 3191 14603
rect 6929 14569 6963 14603
rect 8953 14569 8987 14603
rect 9873 14569 9907 14603
rect 13093 14569 13127 14603
rect 16129 14569 16163 14603
rect 2329 14501 2363 14535
rect 7389 14433 7423 14467
rect 7481 14433 7515 14467
rect 8217 14433 8251 14467
rect 8309 14433 8343 14467
rect 9413 14433 9447 14467
rect 9597 14433 9631 14467
rect 11345 14433 11379 14467
rect 11989 14433 12023 14467
rect 12541 14433 12575 14467
rect 12725 14433 12759 14467
rect 14749 14433 14783 14467
rect 1961 14365 1995 14399
rect 2145 14365 2179 14399
rect 3065 14365 3099 14399
rect 3433 14365 3467 14399
rect 4261 14365 4295 14399
rect 6745 14365 6779 14399
rect 11253 14365 11287 14399
rect 12265 14365 12299 14399
rect 12357 14365 12391 14399
rect 12633 14365 12667 14399
rect 12909 14365 12943 14399
rect 13185 14365 13219 14399
rect 13369 14365 13403 14399
rect 13553 14365 13587 14399
rect 16221 14365 16255 14399
rect 2697 14297 2731 14331
rect 4506 14297 4540 14331
rect 11008 14297 11042 14331
rect 12081 14297 12115 14331
rect 15016 14297 15050 14331
rect 2881 14229 2915 14263
rect 3617 14229 3651 14263
rect 5641 14229 5675 14263
rect 7297 14229 7331 14263
rect 7757 14229 7791 14263
rect 8125 14229 8159 14263
rect 9321 14229 9355 14263
rect 13277 14229 13311 14263
rect 13737 14229 13771 14263
rect 16405 14229 16439 14263
rect 1961 14025 1995 14059
rect 3709 14025 3743 14059
rect 4077 14025 4111 14059
rect 12173 14025 12207 14059
rect 12541 14025 12575 14059
rect 13737 14025 13771 14059
rect 15025 14025 15059 14059
rect 4905 13957 4939 13991
rect 6561 13957 6595 13991
rect 7297 13957 7331 13991
rect 13369 13957 13403 13991
rect 15485 13957 15519 13991
rect 1869 13889 1903 13923
rect 2697 13889 2731 13923
rect 4169 13889 4203 13923
rect 8125 13889 8159 13923
rect 8392 13889 8426 13923
rect 9965 13889 9999 13923
rect 10057 13889 10091 13923
rect 10425 13889 10459 13923
rect 11069 13889 11103 13923
rect 11621 13889 11655 13923
rect 12173 13889 12207 13923
rect 12357 13889 12391 13923
rect 12449 13889 12483 13923
rect 12633 13889 12667 13923
rect 12731 13889 12765 13923
rect 12903 13889 12937 13923
rect 13185 13889 13219 13923
rect 13461 13889 13495 13923
rect 13553 13889 13587 13923
rect 13829 13889 13863 13923
rect 14013 13889 14047 13923
rect 14105 13889 14139 13923
rect 14197 13889 14231 13923
rect 15393 13889 15427 13923
rect 15853 13889 15887 13923
rect 16405 13889 16439 13923
rect 2053 13821 2087 13855
rect 2789 13821 2823 13855
rect 2881 13821 2915 13855
rect 3433 13821 3467 13855
rect 3617 13821 3651 13855
rect 10149 13821 10183 13855
rect 15577 13821 15611 13855
rect 9505 13753 9539 13787
rect 9597 13753 9631 13787
rect 14473 13753 14507 13787
rect 1501 13685 1535 13719
rect 2329 13685 2363 13719
rect 12909 13685 12943 13719
rect 2789 13481 2823 13515
rect 13185 13481 13219 13515
rect 13553 13481 13587 13515
rect 13737 13481 13771 13515
rect 7941 13413 7975 13447
rect 3801 13345 3835 13379
rect 6377 13345 6411 13379
rect 8677 13345 8711 13379
rect 9505 13345 9539 13379
rect 11345 13345 11379 13379
rect 12357 13345 12391 13379
rect 13461 13345 13495 13379
rect 1409 13277 1443 13311
rect 6561 13277 6595 13311
rect 10609 13277 10643 13311
rect 11621 13277 11655 13311
rect 12541 13277 12575 13311
rect 12633 13277 12667 13311
rect 12909 13277 12943 13311
rect 13001 13277 13035 13311
rect 13093 13277 13127 13311
rect 13277 13277 13311 13311
rect 13369 13277 13403 13311
rect 14289 13277 14323 13311
rect 14657 13277 14691 13311
rect 15761 13277 15795 13311
rect 16405 13277 16439 13311
rect 1654 13209 1688 13243
rect 4068 13209 4102 13243
rect 6828 13209 6862 13243
rect 14473 13209 14507 13243
rect 14565 13209 14599 13243
rect 5181 13141 5215 13175
rect 5733 13141 5767 13175
rect 6101 13141 6135 13175
rect 6193 13141 6227 13175
rect 8033 13141 8067 13175
rect 8401 13141 8435 13175
rect 8493 13141 8527 13175
rect 8953 13141 8987 13175
rect 12265 13141 12299 13175
rect 14841 13141 14875 13175
rect 15577 13141 15611 13175
rect 15853 13141 15887 13175
rect 1501 12937 1535 12971
rect 3341 12937 3375 12971
rect 3893 12937 3927 12971
rect 4261 12937 4295 12971
rect 6469 12937 6503 12971
rect 9045 12937 9079 12971
rect 9505 12937 9539 12971
rect 9873 12937 9907 12971
rect 11529 12937 11563 12971
rect 11897 12937 11931 12971
rect 13369 12937 13403 12971
rect 14105 12937 14139 12971
rect 16221 12937 16255 12971
rect 11008 12869 11042 12903
rect 14381 12869 14415 12903
rect 15108 12869 15142 12903
rect 1685 12801 1719 12835
rect 1961 12801 1995 12835
rect 2228 12801 2262 12835
rect 7113 12801 7147 12835
rect 7205 12801 7239 12835
rect 7297 12801 7331 12835
rect 7481 12801 7515 12835
rect 7573 12801 7607 12835
rect 9413 12801 9447 12835
rect 11989 12801 12023 12835
rect 13001 12801 13035 12835
rect 13185 12801 13219 12835
rect 13461 12801 13495 12835
rect 13645 12801 13679 12835
rect 13737 12801 13771 12835
rect 13829 12801 13863 12835
rect 14197 12801 14231 12835
rect 14473 12801 14507 12835
rect 14565 12801 14599 12835
rect 14841 12801 14875 12835
rect 16497 12801 16531 12835
rect 3617 12733 3651 12767
rect 3801 12733 3835 12767
rect 8125 12733 8159 12767
rect 8677 12733 8711 12767
rect 9597 12733 9631 12767
rect 11253 12733 11287 12767
rect 12081 12733 12115 12767
rect 7757 12665 7791 12699
rect 16313 12665 16347 12699
rect 13001 12597 13035 12631
rect 14749 12597 14783 12631
rect 6745 12393 6779 12427
rect 10333 12393 10367 12427
rect 13921 12393 13955 12427
rect 15209 12393 15243 12427
rect 16405 12325 16439 12359
rect 8033 12257 8067 12291
rect 8953 12257 8987 12291
rect 10977 12257 11011 12291
rect 11897 12257 11931 12291
rect 13277 12257 13311 12291
rect 15669 12257 15703 12291
rect 15761 12257 15795 12291
rect 1685 12189 1719 12223
rect 2053 12189 2087 12223
rect 2697 12189 2731 12223
rect 4077 12189 4111 12223
rect 4169 12189 4203 12223
rect 4261 12189 4295 12223
rect 4445 12189 4479 12223
rect 4721 12189 4755 12223
rect 5365 12189 5399 12223
rect 7757 12189 7791 12223
rect 8677 12189 8711 12223
rect 11161 12189 11195 12223
rect 12081 12189 12115 12223
rect 12173 12189 12207 12223
rect 13553 12189 13587 12223
rect 13737 12189 13771 12223
rect 14565 12189 14599 12223
rect 16221 12189 16255 12223
rect 4537 12121 4571 12155
rect 5632 12121 5666 12155
rect 9220 12121 9254 12155
rect 12449 12121 12483 12155
rect 15577 12121 15611 12155
rect 1501 12053 1535 12087
rect 1869 12053 1903 12087
rect 2513 12053 2547 12087
rect 3801 12053 3835 12087
rect 4905 12053 4939 12087
rect 7389 12053 7423 12087
rect 7849 12053 7883 12087
rect 8585 12053 8619 12087
rect 10425 12053 10459 12087
rect 11805 12053 11839 12087
rect 11897 12053 11931 12087
rect 15117 12053 15151 12087
rect 6193 11849 6227 11883
rect 8309 11849 8343 11883
rect 9045 11849 9079 11883
rect 9505 11849 9539 11883
rect 9965 11849 9999 11883
rect 11529 11849 11563 11883
rect 14749 11849 14783 11883
rect 15485 11849 15519 11883
rect 15945 11849 15979 11883
rect 1685 11781 1719 11815
rect 1869 11781 1903 11815
rect 7196 11781 7230 11815
rect 9137 11781 9171 11815
rect 11100 11781 11134 11815
rect 11897 11781 11931 11815
rect 3341 11713 3375 11747
rect 3608 11713 3642 11747
rect 4813 11713 4847 11747
rect 5080 11713 5114 11747
rect 6929 11713 6963 11747
rect 11345 11713 11379 11747
rect 11713 11713 11747 11747
rect 11805 11713 11839 11747
rect 12081 11713 12115 11747
rect 12173 11713 12207 11747
rect 12357 11713 12391 11747
rect 12633 11713 12667 11747
rect 14657 11713 14691 11747
rect 14841 11713 14875 11747
rect 16129 11713 16163 11747
rect 16221 11713 16255 11747
rect 2973 11645 3007 11679
rect 3249 11645 3283 11679
rect 8953 11645 8987 11679
rect 15577 11645 15611 11679
rect 15669 11645 15703 11679
rect 16405 11577 16439 11611
rect 2053 11509 2087 11543
rect 4721 11509 4755 11543
rect 12265 11509 12299 11543
rect 15117 11509 15151 11543
rect 1501 11305 1535 11339
rect 4169 11305 4203 11339
rect 4997 11305 5031 11339
rect 6929 11305 6963 11339
rect 8585 11305 8619 11339
rect 9689 11305 9723 11339
rect 13921 11305 13955 11339
rect 14657 11305 14691 11339
rect 16221 11305 16255 11339
rect 16313 11305 16347 11339
rect 3157 11237 3191 11271
rect 7573 11169 7607 11203
rect 7941 11169 7975 11203
rect 8125 11169 8159 11203
rect 10149 11169 10183 11203
rect 10333 11169 10367 11203
rect 12357 11169 12391 11203
rect 13461 11169 13495 11203
rect 13553 11169 13587 11203
rect 14841 11169 14875 11203
rect 1685 11101 1719 11135
rect 1777 11101 1811 11135
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 4353 11101 4387 11135
rect 4537 11101 4571 11135
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 5457 11101 5491 11135
rect 8217 11101 8251 11135
rect 11805 11101 11839 11135
rect 11897 11101 11931 11135
rect 12173 11101 12207 11135
rect 12265 11101 12299 11135
rect 12449 11101 12483 11135
rect 12725 11101 12759 11135
rect 12817 11101 12851 11135
rect 12909 11101 12943 11135
rect 13001 11101 13035 11135
rect 13185 11101 13219 11135
rect 13369 11101 13403 11135
rect 13737 11101 13771 11135
rect 14105 11101 14139 11135
rect 14289 11101 14323 11135
rect 14473 11101 14507 11135
rect 15108 11101 15142 11135
rect 16497 11101 16531 11135
rect 2044 11033 2078 11067
rect 5724 11033 5758 11067
rect 7389 11033 7423 11067
rect 11989 11033 12023 11067
rect 14381 11033 14415 11067
rect 6837 10965 6871 10999
rect 7297 10965 7331 10999
rect 10057 10965 10091 10999
rect 11621 10965 11655 10999
rect 12541 10965 12575 10999
rect 1685 10761 1719 10795
rect 3709 10761 3743 10795
rect 6377 10761 6411 10795
rect 7941 10761 7975 10795
rect 12173 10761 12207 10795
rect 14013 10761 14047 10795
rect 4445 10693 4479 10727
rect 4782 10693 4816 10727
rect 12357 10693 12391 10727
rect 12541 10693 12575 10727
rect 12633 10693 12667 10727
rect 1961 10625 1995 10659
rect 2053 10625 2087 10659
rect 2145 10625 2179 10659
rect 2329 10625 2363 10659
rect 2697 10625 2731 10659
rect 2786 10625 2820 10659
rect 2902 10631 2936 10665
rect 3065 10625 3099 10659
rect 3157 10625 3191 10659
rect 3249 10625 3283 10659
rect 3433 10625 3467 10659
rect 3525 10625 3559 10659
rect 3801 10625 3835 10659
rect 3985 10625 4019 10659
rect 4077 10625 4111 10659
rect 4169 10625 4203 10659
rect 4537 10625 4571 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 7757 10625 7791 10659
rect 8125 10625 8159 10659
rect 8217 10625 8251 10659
rect 8401 10625 8435 10659
rect 8493 10625 8527 10659
rect 9321 10625 9355 10659
rect 9781 10625 9815 10659
rect 11529 10625 11563 10659
rect 12265 10625 12299 10659
rect 12909 10625 12943 10659
rect 13185 10625 13219 10659
rect 13553 10625 13587 10659
rect 13645 10625 13679 10659
rect 13921 10625 13955 10659
rect 14565 10625 14599 10659
rect 14832 10625 14866 10659
rect 16221 10625 16255 10659
rect 6837 10557 6871 10591
rect 7021 10557 7055 10591
rect 9413 10557 9447 10591
rect 9597 10557 9631 10591
rect 10333 10557 10367 10591
rect 11161 10557 11195 10591
rect 12633 10557 12667 10591
rect 13277 10557 13311 10591
rect 14381 10557 14415 10591
rect 12265 10489 12299 10523
rect 13829 10489 13863 10523
rect 2421 10421 2455 10455
rect 5917 10421 5951 10455
rect 8953 10421 8987 10455
rect 10609 10421 10643 10455
rect 12817 10421 12851 10455
rect 14197 10421 14231 10455
rect 15945 10421 15979 10455
rect 16405 10421 16439 10455
rect 1777 10217 1811 10251
rect 5365 10217 5399 10251
rect 8217 10217 8251 10251
rect 10517 10217 10551 10251
rect 12081 10217 12115 10251
rect 14933 10217 14967 10251
rect 10609 10149 10643 10183
rect 13645 10149 13679 10183
rect 1869 10081 1903 10115
rect 13461 10081 13495 10115
rect 14749 10081 14783 10115
rect 15393 10081 15427 10115
rect 15485 10081 15519 10115
rect 16313 10081 16347 10115
rect 4813 10013 4847 10047
rect 4905 10013 4939 10047
rect 5089 10013 5123 10047
rect 5181 10013 5215 10047
rect 8401 10013 8435 10047
rect 8493 10013 8527 10047
rect 8677 10013 8711 10047
rect 8769 10013 8803 10047
rect 9137 10013 9171 10047
rect 11722 10013 11756 10047
rect 11989 10013 12023 10047
rect 13553 10013 13587 10047
rect 13737 10013 13771 10047
rect 1409 9945 1443 9979
rect 1593 9945 1627 9979
rect 2136 9945 2170 9979
rect 3801 9945 3835 9979
rect 9404 9945 9438 9979
rect 13194 9945 13228 9979
rect 3249 9877 3283 9911
rect 14105 9877 14139 9911
rect 15301 9877 15335 9911
rect 15761 9877 15795 9911
rect 10149 9673 10183 9707
rect 10517 9673 10551 9707
rect 3341 9605 3375 9639
rect 4721 9605 4755 9639
rect 8944 9605 8978 9639
rect 14197 9605 14231 9639
rect 1685 9537 1719 9571
rect 2053 9537 2087 9571
rect 3525 9537 3559 9571
rect 4813 9537 4847 9571
rect 4997 9537 5031 9571
rect 6101 9537 6135 9571
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 6929 9537 6963 9571
rect 7021 9537 7055 9571
rect 7472 9537 7506 9571
rect 8677 9537 8711 9571
rect 14105 9537 14139 9571
rect 16497 9537 16531 9571
rect 3985 9469 4019 9503
rect 5181 9469 5215 9503
rect 7205 9469 7239 9503
rect 10609 9469 10643 9503
rect 10701 9469 10735 9503
rect 1869 9401 1903 9435
rect 8585 9401 8619 9435
rect 10057 9401 10091 9435
rect 16313 9401 16347 9435
rect 1501 9333 1535 9367
rect 3709 9333 3743 9367
rect 6469 9333 6503 9367
rect 6009 9129 6043 9163
rect 7573 9129 7607 9163
rect 9873 9129 9907 9163
rect 10885 9129 10919 9163
rect 1501 9061 1535 9095
rect 13001 9061 13035 9095
rect 4629 8993 4663 9027
rect 8033 8993 8067 9027
rect 8217 8993 8251 9027
rect 9505 8993 9539 9027
rect 1685 8925 1719 8959
rect 1961 8925 1995 8959
rect 2145 8925 2179 8959
rect 2237 8925 2271 8959
rect 2329 8925 2363 8959
rect 2973 8925 3007 8959
rect 3893 8925 3927 8959
rect 4077 8925 4111 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 6101 8925 6135 8959
rect 10149 8925 10183 8959
rect 11069 8925 11103 8959
rect 11161 8925 11195 8959
rect 11437 8925 11471 8959
rect 11529 8925 11563 8959
rect 11805 8925 11839 8959
rect 12449 8925 12483 8959
rect 12817 8925 12851 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 14381 8925 14415 8959
rect 14473 8925 14507 8959
rect 4537 8857 4571 8891
rect 4874 8857 4908 8891
rect 6368 8857 6402 8891
rect 7941 8857 7975 8891
rect 8953 8857 8987 8891
rect 9689 8857 9723 8891
rect 10333 8857 10367 8891
rect 10517 8857 10551 8891
rect 11253 8857 11287 8891
rect 12633 8857 12667 8891
rect 12725 8857 12759 8891
rect 13277 8857 13311 8891
rect 13461 8857 13495 8891
rect 2605 8789 2639 8823
rect 2789 8789 2823 8823
rect 7481 8789 7515 8823
rect 9873 8789 9907 8823
rect 13093 8789 13127 8823
rect 14749 8789 14783 8823
rect 2053 8585 2087 8619
rect 3525 8585 3559 8619
rect 14657 8585 14691 8619
rect 1685 8517 1719 8551
rect 1869 8517 1903 8551
rect 2412 8517 2446 8551
rect 3809 8517 3843 8551
rect 3985 8517 4019 8551
rect 6377 8517 6411 8551
rect 7389 8517 7423 8551
rect 9321 8517 9355 8551
rect 13093 8517 13127 8551
rect 3617 8449 3651 8483
rect 4077 8449 4111 8483
rect 4261 8449 4295 8483
rect 4353 8449 4387 8483
rect 4445 8449 4479 8483
rect 4813 8449 4847 8483
rect 5069 8449 5103 8483
rect 7941 8449 7975 8483
rect 8217 8449 8251 8483
rect 8585 8449 8619 8483
rect 8769 8449 8803 8483
rect 9045 8449 9079 8483
rect 9781 8449 9815 8483
rect 10701 8449 10735 8483
rect 10885 8449 10919 8483
rect 12173 8449 12207 8483
rect 12265 8449 12299 8483
rect 13533 8449 13567 8483
rect 16221 8449 16255 8483
rect 2145 8381 2179 8415
rect 4721 8381 4755 8415
rect 7113 8381 7147 8415
rect 9137 8381 9171 8415
rect 10517 8381 10551 8415
rect 13277 8381 13311 8415
rect 6193 8313 6227 8347
rect 16405 8313 16439 8347
rect 2789 8041 2823 8075
rect 4537 8041 4571 8075
rect 6377 8041 6411 8075
rect 8769 8041 8803 8075
rect 13185 8041 13219 8075
rect 13645 8041 13679 8075
rect 4353 7973 4387 8007
rect 1409 7905 1443 7939
rect 4997 7905 5031 7939
rect 6837 7905 6871 7939
rect 7021 7905 7055 7939
rect 3157 7837 3191 7871
rect 3801 7837 3835 7871
rect 3893 7837 3927 7871
rect 4077 7837 4111 7871
rect 4169 7837 4203 7871
rect 4813 7837 4847 7871
rect 4905 7837 4939 7871
rect 6745 7837 6779 7871
rect 7389 7837 7423 7871
rect 8953 7837 8987 7871
rect 9229 7837 9263 7871
rect 10885 7837 10919 7871
rect 12541 7837 12575 7871
rect 12725 7837 12759 7871
rect 12817 7837 12851 7871
rect 12909 7837 12943 7871
rect 13461 7837 13495 7871
rect 14105 7837 14139 7871
rect 1676 7769 1710 7803
rect 4629 7769 4663 7803
rect 7656 7769 7690 7803
rect 9496 7769 9530 7803
rect 11152 7769 11186 7803
rect 13277 7769 13311 7803
rect 14372 7769 14406 7803
rect 2973 7701 3007 7735
rect 9045 7701 9079 7735
rect 10609 7701 10643 7735
rect 12265 7701 12299 7735
rect 15485 7701 15519 7735
rect 1593 7497 1627 7531
rect 3341 7497 3375 7531
rect 8033 7497 8067 7531
rect 8401 7497 8435 7531
rect 9137 7497 9171 7531
rect 9597 7497 9631 7531
rect 11529 7497 11563 7531
rect 15209 7497 15243 7531
rect 2329 7429 2363 7463
rect 2513 7429 2547 7463
rect 3065 7429 3099 7463
rect 4353 7429 4387 7463
rect 9321 7429 9355 7463
rect 10701 7429 10735 7463
rect 1869 7361 1903 7395
rect 1961 7361 1995 7395
rect 2053 7361 2087 7395
rect 2237 7361 2271 7395
rect 2697 7361 2731 7395
rect 2789 7361 2823 7395
rect 2973 7361 3007 7395
rect 3181 7361 3215 7395
rect 4261 7361 4295 7395
rect 4445 7361 4479 7395
rect 4997 7361 5031 7395
rect 5181 7361 5215 7395
rect 6929 7361 6963 7395
rect 7021 7361 7055 7395
rect 7205 7361 7239 7395
rect 7297 7361 7331 7395
rect 9689 7361 9723 7395
rect 10977 7361 11011 7395
rect 11805 7361 11839 7395
rect 11897 7361 11931 7395
rect 11989 7361 12023 7395
rect 12173 7361 12207 7395
rect 12357 7361 12391 7395
rect 12541 7361 12575 7395
rect 12817 7361 12851 7395
rect 13001 7361 13035 7395
rect 13277 7361 13311 7395
rect 13461 7361 13495 7395
rect 14473 7361 14507 7395
rect 14657 7361 14691 7395
rect 14749 7361 14783 7395
rect 14841 7361 14875 7395
rect 15393 7361 15427 7395
rect 8493 7293 8527 7327
rect 8677 7293 8711 7327
rect 9965 7293 9999 7327
rect 10793 7293 10827 7327
rect 12725 7293 12759 7327
rect 6745 7225 6779 7259
rect 15117 7225 15151 7259
rect 4813 7157 4847 7191
rect 8953 7157 8987 7191
rect 9137 7157 9171 7191
rect 11161 7157 11195 7191
rect 12909 7157 12943 7191
rect 13645 7157 13679 7191
rect 5457 6953 5491 6987
rect 9505 6953 9539 6987
rect 13921 6953 13955 6987
rect 2053 6817 2087 6851
rect 10057 6817 10091 6851
rect 10885 6817 10919 6851
rect 4445 6749 4479 6783
rect 4629 6749 4663 6783
rect 4721 6749 4755 6783
rect 4813 6749 4847 6783
rect 5273 6749 5307 6783
rect 5549 6749 5583 6783
rect 7389 6749 7423 6783
rect 7757 6749 7791 6783
rect 7849 6749 7883 6783
rect 7941 6749 7975 6783
rect 8125 6749 8159 6783
rect 14289 6749 14323 6783
rect 14473 6749 14507 6783
rect 14565 6749 14599 6783
rect 14657 6749 14691 6783
rect 15025 6749 15059 6783
rect 2320 6681 2354 6715
rect 3985 6681 4019 6715
rect 4169 6681 4203 6715
rect 7144 6681 7178 6715
rect 7481 6681 7515 6715
rect 9873 6681 9907 6715
rect 10333 6681 10367 6715
rect 11161 6681 11195 6715
rect 13553 6681 13587 6715
rect 13737 6681 13771 6715
rect 14933 6681 14967 6715
rect 15270 6681 15304 6715
rect 3433 6613 3467 6647
rect 3801 6613 3835 6647
rect 5089 6613 5123 6647
rect 6009 6613 6043 6647
rect 9965 6613 9999 6647
rect 11253 6613 11287 6647
rect 16405 6613 16439 6647
rect 2697 6409 2731 6443
rect 4537 6409 4571 6443
rect 6929 6409 6963 6443
rect 7389 6409 7423 6443
rect 9045 6409 9079 6443
rect 14197 6409 14231 6443
rect 16497 6409 16531 6443
rect 6653 6341 6687 6375
rect 7205 6341 7239 6375
rect 14565 6341 14599 6375
rect 15384 6341 15418 6375
rect 2973 6273 3007 6307
rect 3065 6273 3099 6307
rect 3157 6273 3191 6307
rect 3341 6273 3375 6307
rect 3433 6273 3467 6307
rect 4169 6273 4203 6307
rect 4353 6273 4387 6307
rect 4629 6273 4663 6307
rect 4885 6273 4919 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 7021 6273 7055 6307
rect 8953 6273 8987 6307
rect 9229 6273 9263 6307
rect 9413 6273 9447 6307
rect 10221 6273 10255 6307
rect 12633 6273 12667 6307
rect 12909 6273 12943 6307
rect 13093 6273 13127 6307
rect 13829 6273 13863 6307
rect 14013 6273 14047 6307
rect 14473 6273 14507 6307
rect 14657 6273 14691 6307
rect 14841 6273 14875 6307
rect 9965 6205 9999 6239
rect 12817 6205 12851 6239
rect 13277 6205 13311 6239
rect 15117 6205 15151 6239
rect 12449 6137 12483 6171
rect 14289 6137 14323 6171
rect 3617 6069 3651 6103
rect 6009 6069 6043 6103
rect 11345 6069 11379 6103
rect 8769 5865 8803 5899
rect 9873 5865 9907 5899
rect 13737 5797 13771 5831
rect 9965 5729 9999 5763
rect 10425 5729 10459 5763
rect 1685 5661 1719 5695
rect 2237 5661 2271 5695
rect 3065 5661 3099 5695
rect 3157 5661 3191 5695
rect 3249 5661 3283 5695
rect 3433 5661 3467 5695
rect 8217 5661 8251 5695
rect 8585 5661 8619 5695
rect 9229 5661 9263 5695
rect 9413 5661 9447 5695
rect 9505 5661 9539 5695
rect 9597 5661 9631 5695
rect 10333 5661 10367 5695
rect 12081 5661 12115 5695
rect 12357 5661 12391 5695
rect 16221 5661 16255 5695
rect 2053 5593 2087 5627
rect 7297 5593 7331 5627
rect 7481 5593 7515 5627
rect 8401 5593 8435 5627
rect 8493 5593 8527 5627
rect 10149 5593 10183 5627
rect 10670 5593 10704 5627
rect 12265 5593 12299 5627
rect 12624 5593 12658 5627
rect 14197 5593 14231 5627
rect 14381 5593 14415 5627
rect 1501 5525 1535 5559
rect 1869 5525 1903 5559
rect 2789 5525 2823 5559
rect 7665 5525 7699 5559
rect 11805 5525 11839 5559
rect 11897 5525 11931 5559
rect 14565 5525 14599 5559
rect 16405 5525 16439 5559
rect 3709 5321 3743 5355
rect 11713 5321 11747 5355
rect 13001 5321 13035 5355
rect 14933 5321 14967 5355
rect 2504 5253 2538 5287
rect 6193 5253 6227 5287
rect 10977 5253 11011 5287
rect 11989 5253 12023 5287
rect 15301 5253 15335 5287
rect 1777 5185 1811 5219
rect 1869 5185 1903 5219
rect 1961 5185 1995 5219
rect 2145 5185 2179 5219
rect 3893 5185 3927 5219
rect 4077 5185 4111 5219
rect 4537 5185 4571 5219
rect 4629 5185 4663 5219
rect 4721 5185 4755 5219
rect 4905 5185 4939 5219
rect 5089 5185 5123 5219
rect 5273 5185 5307 5219
rect 5365 5185 5399 5219
rect 5457 5185 5491 5219
rect 5825 5185 5859 5219
rect 6009 5185 6043 5219
rect 7196 5185 7230 5219
rect 8677 5185 8711 5219
rect 8944 5185 8978 5219
rect 10517 5185 10551 5219
rect 10609 5185 10643 5219
rect 10701 5185 10735 5219
rect 10885 5185 10919 5219
rect 11161 5185 11195 5219
rect 11345 5185 11379 5219
rect 11897 5185 11931 5219
rect 12081 5185 12115 5219
rect 12265 5185 12299 5219
rect 12357 5185 12391 5219
rect 12541 5185 12575 5219
rect 12633 5185 12667 5219
rect 12725 5185 12759 5219
rect 13553 5185 13587 5219
rect 13820 5185 13854 5219
rect 15209 5185 15243 5219
rect 15393 5185 15427 5219
rect 15577 5185 15611 5219
rect 2237 5117 2271 5151
rect 6929 5117 6963 5151
rect 10241 5049 10275 5083
rect 1501 4981 1535 5015
rect 3617 4981 3651 5015
rect 4261 4981 4295 5015
rect 5733 4981 5767 5015
rect 8309 4981 8343 5015
rect 10057 4981 10091 5015
rect 15025 4981 15059 5015
rect 2789 4777 2823 4811
rect 3433 4777 3467 4811
rect 6929 4777 6963 4811
rect 7205 4777 7239 4811
rect 14105 4777 14139 4811
rect 8953 4709 8987 4743
rect 15117 4641 15151 4675
rect 1409 4573 1443 4607
rect 2881 4573 2915 4607
rect 3157 4573 3191 4607
rect 3249 4573 3283 4607
rect 4077 4573 4111 4607
rect 4344 4573 4378 4607
rect 5549 4573 5583 4607
rect 5816 4573 5850 4607
rect 7481 4573 7515 4607
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 7849 4573 7883 4607
rect 9229 4573 9263 4607
rect 9321 4573 9355 4607
rect 9413 4573 9447 4607
rect 9597 4573 9631 4607
rect 10333 4573 10367 4607
rect 13553 4573 13587 4607
rect 14381 4573 14415 4607
rect 14473 4573 14507 4607
rect 14565 4573 14599 4607
rect 14749 4573 14783 4607
rect 1654 4505 1688 4539
rect 3065 4505 3099 4539
rect 8401 4505 8435 4539
rect 8585 4505 8619 4539
rect 8769 4505 8803 4539
rect 13737 4505 13771 4539
rect 15362 4505 15396 4539
rect 5457 4437 5491 4471
rect 10149 4437 10183 4471
rect 13921 4437 13955 4471
rect 16497 4437 16531 4471
rect 4537 4233 4571 4267
rect 3157 4165 3191 4199
rect 4169 4165 4203 4199
rect 4353 4165 4387 4199
rect 6929 4165 6963 4199
rect 7849 4165 7883 4199
rect 11161 4165 11195 4199
rect 13277 4165 13311 4199
rect 1685 4097 1719 4131
rect 2329 4097 2363 4131
rect 2697 4097 2731 4131
rect 2973 4097 3007 4131
rect 3249 4097 3283 4131
rect 3341 4097 3375 4131
rect 3617 4097 3651 4131
rect 6745 4097 6779 4131
rect 7021 4097 7055 4131
rect 7113 4097 7147 4131
rect 7665 4097 7699 4131
rect 7941 4097 7975 4131
rect 8033 4097 8067 4131
rect 10517 4097 10551 4131
rect 10609 4097 10643 4131
rect 10701 4097 10735 4131
rect 10885 4097 10919 4131
rect 11345 4097 11379 4131
rect 11713 4097 11747 4131
rect 11805 4097 11839 4131
rect 11897 4097 11931 4131
rect 12081 4097 12115 4131
rect 12449 4097 12483 4131
rect 12541 4097 12575 4131
rect 12633 4097 12667 4131
rect 12817 4097 12851 4131
rect 13093 4097 13127 4131
rect 14013 4097 14047 4131
rect 14105 4097 14139 4131
rect 14197 4097 14231 4131
rect 14381 4097 14415 4131
rect 14473 4097 14507 4131
rect 14657 4097 14691 4131
rect 14749 4097 14783 4131
rect 14841 4097 14875 4131
rect 15485 4097 15519 4131
rect 15853 4097 15887 4131
rect 16497 4097 16531 4131
rect 10977 4029 11011 4063
rect 12909 4029 12943 4063
rect 15117 4029 15151 4063
rect 3801 3961 3835 3995
rect 7297 3961 7331 3995
rect 8217 3961 8251 3995
rect 11529 3961 11563 3995
rect 13829 3961 13863 3995
rect 15669 3961 15703 3995
rect 16037 3961 16071 3995
rect 1501 3893 1535 3927
rect 2145 3893 2179 3927
rect 2513 3893 2547 3927
rect 3525 3893 3559 3927
rect 10241 3893 10275 3927
rect 12173 3893 12207 3927
rect 16313 3893 16347 3927
rect 6745 3689 6779 3723
rect 13001 3689 13035 3723
rect 16221 3621 16255 3655
rect 1777 3485 1811 3519
rect 1869 3485 1903 3519
rect 1961 3485 1995 3519
rect 2145 3485 2179 3519
rect 2697 3485 2731 3519
rect 3065 3485 3099 3519
rect 3157 3485 3191 3519
rect 3249 3485 3283 3519
rect 3433 3485 3467 3519
rect 3893 3485 3927 3519
rect 4077 3485 4111 3519
rect 4169 3485 4203 3519
rect 4261 3485 4295 3519
rect 4629 3485 4663 3519
rect 4813 3485 4847 3519
rect 4905 3485 4939 3519
rect 4997 3485 5031 3519
rect 5365 3485 5399 3519
rect 7297 3485 7331 3519
rect 7389 3485 7423 3519
rect 7481 3485 7515 3519
rect 7665 3485 7699 3519
rect 8401 3485 8435 3519
rect 8493 3485 8527 3519
rect 8585 3485 8619 3519
rect 8769 3485 8803 3519
rect 9689 3485 9723 3519
rect 9781 3485 9815 3519
rect 9873 3485 9907 3519
rect 10057 3485 10091 3519
rect 10149 3485 10183 3519
rect 10405 3485 10439 3519
rect 11621 3485 11655 3519
rect 13369 3485 13403 3519
rect 13461 3485 13495 3519
rect 13553 3485 13587 3519
rect 13737 3485 13771 3519
rect 14197 3485 14231 3519
rect 14381 3485 14415 3519
rect 14473 3485 14507 3519
rect 14565 3485 14599 3519
rect 14933 3485 14967 3519
rect 15117 3482 15151 3516
rect 15209 3485 15243 3519
rect 15301 3485 15335 3519
rect 15669 3485 15703 3519
rect 16037 3485 16071 3519
rect 5273 3417 5307 3451
rect 5610 3417 5644 3451
rect 11888 3417 11922 3451
rect 1501 3349 1535 3383
rect 2513 3349 2547 3383
rect 2789 3349 2823 3383
rect 4537 3349 4571 3383
rect 7021 3349 7055 3383
rect 8125 3349 8159 3383
rect 9413 3349 9447 3383
rect 11529 3349 11563 3383
rect 13093 3349 13127 3383
rect 14841 3349 14875 3383
rect 15577 3349 15611 3383
rect 15853 3349 15887 3383
rect 1961 3145 1995 3179
rect 4169 3145 4203 3179
rect 5733 3145 5767 3179
rect 9413 3145 9447 3179
rect 10977 3145 11011 3179
rect 14289 3145 14323 3179
rect 16037 3145 16071 3179
rect 1593 3077 1627 3111
rect 1777 3077 1811 3111
rect 4528 3077 4562 3111
rect 5917 3077 5951 3111
rect 7582 3077 7616 3111
rect 11345 3077 11379 3111
rect 11805 3077 11839 3111
rect 11897 3077 11931 3111
rect 2329 3009 2363 3043
rect 2596 3009 2630 3043
rect 3801 3009 3835 3043
rect 3985 3009 4019 3043
rect 4261 3009 4295 3043
rect 6101 3009 6135 3043
rect 7849 3009 7883 3043
rect 8033 3009 8067 3043
rect 8289 3009 8323 3043
rect 9505 3009 9539 3043
rect 9761 3009 9795 3043
rect 11161 3009 11195 3043
rect 11713 3009 11747 3043
rect 12081 3009 12115 3043
rect 12716 3009 12750 3043
rect 13921 3009 13955 3043
rect 14105 3009 14139 3043
rect 14924 3009 14958 3043
rect 16129 3009 16163 3043
rect 12449 2941 12483 2975
rect 14657 2941 14691 2975
rect 10885 2873 10919 2907
rect 13829 2873 13863 2907
rect 3709 2805 3743 2839
rect 5641 2805 5675 2839
rect 6469 2805 6503 2839
rect 11529 2805 11563 2839
rect 16313 2805 16347 2839
rect 2789 2601 2823 2635
rect 3065 2601 3099 2635
rect 7573 2601 7607 2635
rect 8769 2601 8803 2635
rect 14473 2601 14507 2635
rect 14933 2601 14967 2635
rect 5273 2533 5307 2567
rect 7113 2533 7147 2567
rect 15117 2465 15151 2499
rect 1409 2397 1443 2431
rect 3249 2397 3283 2431
rect 4261 2397 4295 2431
rect 4721 2397 4755 2431
rect 5089 2397 5123 2431
rect 5457 2397 5491 2431
rect 5825 2397 5859 2431
rect 6193 2397 6227 2431
rect 6561 2397 6595 2431
rect 6745 2397 6779 2431
rect 6837 2397 6871 2431
rect 6929 2397 6963 2431
rect 7389 2397 7423 2431
rect 7941 2397 7975 2431
rect 8033 2397 8067 2431
rect 8585 2397 8619 2431
rect 9413 2397 9447 2431
rect 10057 2397 10091 2431
rect 10425 2397 10459 2431
rect 11345 2397 11379 2431
rect 11989 2397 12023 2431
rect 12633 2397 12667 2431
rect 13001 2397 13035 2431
rect 13921 2397 13955 2431
rect 14289 2397 14323 2431
rect 15384 2397 15418 2431
rect 1654 2329 1688 2363
rect 3433 2329 3467 2363
rect 7205 2329 7239 2363
rect 8401 2329 8435 2363
rect 14105 2329 14139 2363
rect 14565 2329 14599 2363
rect 14749 2329 14783 2363
rect 4077 2261 4111 2295
rect 4537 2261 4571 2295
rect 4905 2261 4939 2295
rect 5641 2261 5675 2295
rect 6009 2261 6043 2295
rect 7757 2261 7791 2295
rect 8217 2261 8251 2295
rect 9229 2261 9263 2295
rect 9873 2261 9907 2295
rect 10609 2261 10643 2295
rect 11161 2261 11195 2295
rect 11805 2261 11839 2295
rect 12449 2261 12483 2295
rect 13185 2261 13219 2295
rect 13737 2261 13771 2295
rect 16497 2261 16531 2295
<< metal1 >>
rect 1104 39738 16836 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 16836 39738
rect 1104 39664 16836 39686
rect 8662 39584 8668 39636
rect 8720 39624 8726 39636
rect 10229 39627 10287 39633
rect 10229 39624 10241 39627
rect 8720 39596 10241 39624
rect 8720 39584 8726 39596
rect 10229 39593 10241 39596
rect 10275 39593 10287 39627
rect 10229 39587 10287 39593
rect 10962 39380 10968 39432
rect 11020 39420 11026 39432
rect 11057 39423 11115 39429
rect 11057 39420 11069 39423
rect 11020 39392 11069 39420
rect 11020 39380 11026 39392
rect 11057 39389 11069 39392
rect 11103 39389 11115 39423
rect 11057 39383 11115 39389
rect 12894 39380 12900 39432
rect 12952 39420 12958 39432
rect 13173 39423 13231 39429
rect 13173 39420 13185 39423
rect 12952 39392 13185 39420
rect 12952 39380 12958 39392
rect 13173 39389 13185 39392
rect 13219 39389 13231 39423
rect 13173 39383 13231 39389
rect 8202 39312 8208 39364
rect 8260 39352 8266 39364
rect 10413 39355 10471 39361
rect 10413 39352 10425 39355
rect 8260 39324 10425 39352
rect 8260 39312 8266 39324
rect 10413 39321 10425 39324
rect 10459 39321 10471 39355
rect 10413 39315 10471 39321
rect 10042 39244 10048 39296
rect 10100 39244 10106 39296
rect 10213 39287 10271 39293
rect 10213 39253 10225 39287
rect 10259 39284 10271 39287
rect 10778 39284 10784 39296
rect 10259 39256 10784 39284
rect 10259 39253 10271 39256
rect 10213 39247 10271 39253
rect 10778 39244 10784 39256
rect 10836 39244 10842 39296
rect 11241 39287 11299 39293
rect 11241 39253 11253 39287
rect 11287 39284 11299 39287
rect 11330 39284 11336 39296
rect 11287 39256 11336 39284
rect 11287 39253 11299 39256
rect 11241 39247 11299 39253
rect 11330 39244 11336 39256
rect 11388 39244 11394 39296
rect 12618 39244 12624 39296
rect 12676 39284 12682 39296
rect 12989 39287 13047 39293
rect 12989 39284 13001 39287
rect 12676 39256 13001 39284
rect 12676 39244 12682 39256
rect 12989 39253 13001 39256
rect 13035 39253 13047 39287
rect 12989 39247 13047 39253
rect 1104 39194 16836 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 16836 39194
rect 1104 39120 16836 39142
rect 7561 39083 7619 39089
rect 7561 39049 7573 39083
rect 7607 39049 7619 39083
rect 7561 39043 7619 39049
rect 7006 38972 7012 39024
rect 7064 39012 7070 39024
rect 7193 39015 7251 39021
rect 7193 39012 7205 39015
rect 7064 38984 7205 39012
rect 7064 38972 7070 38984
rect 7193 38981 7205 38984
rect 7239 38981 7251 39015
rect 7193 38975 7251 38981
rect 6914 38904 6920 38956
rect 6972 38904 6978 38956
rect 7098 38904 7104 38956
rect 7156 38904 7162 38956
rect 7208 38944 7236 38975
rect 7374 38972 7380 39024
rect 7432 39021 7438 39024
rect 7432 39015 7451 39021
rect 7439 38981 7451 39015
rect 7576 39012 7604 39043
rect 10042 39040 10048 39092
rect 10100 39080 10106 39092
rect 10100 39052 10180 39080
rect 10100 39040 10106 39052
rect 10152 39021 10180 39052
rect 7898 39015 7956 39021
rect 7898 39012 7910 39015
rect 7576 38984 7910 39012
rect 7432 38975 7451 38981
rect 7898 38981 7910 38984
rect 7944 38981 7956 39015
rect 7898 38975 7956 38981
rect 10128 39015 10186 39021
rect 10128 38981 10140 39015
rect 10174 38981 10186 39015
rect 10128 38975 10186 38981
rect 7432 38972 7438 38975
rect 8202 38944 8208 38956
rect 7208 38916 8208 38944
rect 8202 38904 8208 38916
rect 8260 38904 8266 38956
rect 12710 38904 12716 38956
rect 12768 38944 12774 38956
rect 13090 38947 13148 38953
rect 13090 38944 13102 38947
rect 12768 38916 13102 38944
rect 12768 38904 12774 38916
rect 13090 38913 13102 38916
rect 13136 38913 13148 38947
rect 13090 38907 13148 38913
rect 6086 38836 6092 38888
rect 6144 38876 6150 38888
rect 7653 38879 7711 38885
rect 7653 38876 7665 38879
rect 6144 38848 7665 38876
rect 6144 38836 6150 38848
rect 7653 38845 7665 38848
rect 7699 38845 7711 38879
rect 7653 38839 7711 38845
rect 9766 38836 9772 38888
rect 9824 38876 9830 38888
rect 9861 38879 9919 38885
rect 9861 38876 9873 38879
rect 9824 38848 9873 38876
rect 9824 38836 9830 38848
rect 9861 38845 9873 38848
rect 9907 38845 9919 38879
rect 9861 38839 9919 38845
rect 13357 38879 13415 38885
rect 13357 38845 13369 38879
rect 13403 38876 13415 38879
rect 13906 38876 13912 38888
rect 13403 38848 13912 38876
rect 13403 38845 13415 38848
rect 13357 38839 13415 38845
rect 13906 38836 13912 38848
rect 13964 38836 13970 38888
rect 7098 38700 7104 38752
rect 7156 38700 7162 38752
rect 7377 38743 7435 38749
rect 7377 38709 7389 38743
rect 7423 38740 7435 38743
rect 7926 38740 7932 38752
rect 7423 38712 7932 38740
rect 7423 38709 7435 38712
rect 7377 38703 7435 38709
rect 7926 38700 7932 38712
rect 7984 38700 7990 38752
rect 8294 38700 8300 38752
rect 8352 38740 8358 38752
rect 9033 38743 9091 38749
rect 9033 38740 9045 38743
rect 8352 38712 9045 38740
rect 8352 38700 8358 38712
rect 9033 38709 9045 38712
rect 9079 38709 9091 38743
rect 9033 38703 9091 38709
rect 11054 38700 11060 38752
rect 11112 38740 11118 38752
rect 11241 38743 11299 38749
rect 11241 38740 11253 38743
rect 11112 38712 11253 38740
rect 11112 38700 11118 38712
rect 11241 38709 11253 38712
rect 11287 38709 11299 38743
rect 11241 38703 11299 38709
rect 11977 38743 12035 38749
rect 11977 38709 11989 38743
rect 12023 38740 12035 38743
rect 12066 38740 12072 38752
rect 12023 38712 12072 38740
rect 12023 38709 12035 38712
rect 11977 38703 12035 38709
rect 12066 38700 12072 38712
rect 12124 38700 12130 38752
rect 1104 38650 16836 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 16836 38650
rect 1104 38576 16836 38598
rect 7742 38496 7748 38548
rect 7800 38536 7806 38548
rect 7837 38539 7895 38545
rect 7837 38536 7849 38539
rect 7800 38508 7849 38536
rect 7800 38496 7806 38508
rect 7837 38505 7849 38508
rect 7883 38505 7895 38539
rect 7837 38499 7895 38505
rect 7926 38496 7932 38548
rect 7984 38536 7990 38548
rect 8573 38539 8631 38545
rect 8573 38536 8585 38539
rect 7984 38508 8585 38536
rect 7984 38496 7990 38508
rect 8573 38505 8585 38508
rect 8619 38536 8631 38539
rect 8662 38536 8668 38548
rect 8619 38508 8668 38536
rect 8619 38505 8631 38508
rect 8573 38499 8631 38505
rect 8662 38496 8668 38508
rect 8720 38496 8726 38548
rect 10778 38496 10784 38548
rect 10836 38496 10842 38548
rect 12069 38539 12127 38545
rect 12069 38505 12081 38539
rect 12115 38536 12127 38539
rect 12158 38536 12164 38548
rect 12115 38508 12164 38536
rect 12115 38505 12127 38508
rect 12069 38499 12127 38505
rect 12158 38496 12164 38508
rect 12216 38496 12222 38548
rect 12253 38539 12311 38545
rect 12253 38505 12265 38539
rect 12299 38536 12311 38539
rect 12710 38536 12716 38548
rect 12299 38508 12716 38536
rect 12299 38505 12311 38508
rect 12253 38499 12311 38505
rect 12710 38496 12716 38508
rect 12768 38496 12774 38548
rect 7374 38428 7380 38480
rect 7432 38468 7438 38480
rect 8113 38471 8171 38477
rect 8113 38468 8125 38471
rect 7432 38440 8125 38468
rect 7432 38428 7438 38440
rect 8113 38437 8125 38440
rect 8159 38437 8171 38471
rect 8113 38431 8171 38437
rect 6086 38360 6092 38412
rect 6144 38360 6150 38412
rect 11149 38403 11207 38409
rect 11149 38400 11161 38403
rect 7668 38372 8340 38400
rect 6356 38267 6414 38273
rect 6356 38233 6368 38267
rect 6402 38264 6414 38267
rect 6638 38264 6644 38276
rect 6402 38236 6644 38264
rect 6402 38233 6414 38236
rect 6356 38227 6414 38233
rect 6638 38224 6644 38236
rect 6696 38224 6702 38276
rect 7668 38208 7696 38372
rect 8110 38292 8116 38344
rect 8168 38292 8174 38344
rect 8312 38341 8340 38372
rect 10796 38372 11161 38400
rect 8297 38335 8355 38341
rect 8297 38301 8309 38335
rect 8343 38301 8355 38335
rect 8297 38295 8355 38301
rect 8478 38292 8484 38344
rect 8536 38332 8542 38344
rect 8941 38335 8999 38341
rect 8941 38332 8953 38335
rect 8536 38304 8953 38332
rect 8536 38292 8542 38304
rect 8941 38301 8953 38304
rect 8987 38332 8999 38335
rect 9766 38332 9772 38344
rect 8987 38304 9772 38332
rect 8987 38301 8999 38304
rect 8941 38295 8999 38301
rect 9766 38292 9772 38304
rect 9824 38292 9830 38344
rect 10594 38292 10600 38344
rect 10652 38292 10658 38344
rect 10796 38341 10824 38372
rect 11149 38369 11161 38372
rect 11195 38369 11207 38403
rect 11149 38363 11207 38369
rect 13906 38360 13912 38412
rect 13964 38360 13970 38412
rect 10781 38335 10839 38341
rect 10781 38301 10793 38335
rect 10827 38301 10839 38335
rect 10781 38295 10839 38301
rect 11054 38292 11060 38344
rect 11112 38292 11118 38344
rect 11241 38335 11299 38341
rect 11241 38301 11253 38335
rect 11287 38332 11299 38335
rect 11514 38332 11520 38344
rect 11287 38304 11520 38332
rect 11287 38301 11299 38304
rect 11241 38295 11299 38301
rect 11514 38292 11520 38304
rect 11572 38332 11578 38344
rect 11609 38335 11667 38341
rect 11609 38332 11621 38335
rect 11572 38304 11621 38332
rect 11572 38292 11578 38304
rect 11609 38301 11621 38304
rect 11655 38301 11667 38335
rect 11609 38295 11667 38301
rect 11793 38335 11851 38341
rect 11793 38301 11805 38335
rect 11839 38332 11851 38335
rect 12158 38332 12164 38344
rect 11839 38304 12164 38332
rect 11839 38301 11851 38304
rect 11793 38295 11851 38301
rect 12158 38292 12164 38304
rect 12216 38292 12222 38344
rect 8021 38267 8079 38273
rect 8021 38233 8033 38267
rect 8067 38233 8079 38267
rect 8021 38227 8079 38233
rect 7469 38199 7527 38205
rect 7469 38165 7481 38199
rect 7515 38196 7527 38199
rect 7558 38196 7564 38208
rect 7515 38168 7564 38196
rect 7515 38165 7527 38168
rect 7469 38159 7527 38165
rect 7558 38156 7564 38168
rect 7616 38156 7622 38208
rect 7650 38156 7656 38208
rect 7708 38156 7714 38208
rect 7834 38205 7840 38208
rect 7821 38199 7840 38205
rect 7821 38165 7833 38199
rect 7821 38159 7840 38165
rect 7834 38156 7840 38159
rect 7892 38156 7898 38208
rect 8036 38196 8064 38227
rect 8202 38224 8208 38276
rect 8260 38264 8266 38276
rect 8389 38267 8447 38273
rect 8389 38264 8401 38267
rect 8260 38236 8401 38264
rect 8260 38224 8266 38236
rect 8389 38233 8401 38236
rect 8435 38233 8447 38267
rect 9186 38267 9244 38273
rect 9186 38264 9198 38267
rect 8389 38227 8447 38233
rect 8772 38236 9198 38264
rect 8294 38196 8300 38208
rect 8036 38168 8300 38196
rect 8294 38156 8300 38168
rect 8352 38156 8358 38208
rect 8570 38156 8576 38208
rect 8628 38205 8634 38208
rect 8772 38205 8800 38236
rect 9186 38233 9198 38236
rect 9232 38233 9244 38267
rect 9186 38227 9244 38233
rect 11882 38224 11888 38276
rect 11940 38224 11946 38276
rect 13078 38224 13084 38276
rect 13136 38264 13142 38276
rect 13642 38267 13700 38273
rect 13642 38264 13654 38267
rect 13136 38236 13654 38264
rect 13136 38224 13142 38236
rect 13642 38233 13654 38236
rect 13688 38233 13700 38267
rect 13642 38227 13700 38233
rect 8628 38199 8647 38205
rect 8635 38165 8647 38199
rect 8628 38159 8647 38165
rect 8757 38199 8815 38205
rect 8757 38165 8769 38199
rect 8803 38165 8815 38199
rect 8757 38159 8815 38165
rect 8628 38156 8634 38159
rect 10318 38156 10324 38208
rect 10376 38156 10382 38208
rect 11701 38199 11759 38205
rect 11701 38165 11713 38199
rect 11747 38196 11759 38199
rect 12085 38199 12143 38205
rect 12085 38196 12097 38199
rect 11747 38168 12097 38196
rect 11747 38165 11759 38168
rect 11701 38159 11759 38165
rect 12085 38165 12097 38168
rect 12131 38165 12143 38199
rect 12085 38159 12143 38165
rect 12342 38156 12348 38208
rect 12400 38196 12406 38208
rect 12529 38199 12587 38205
rect 12529 38196 12541 38199
rect 12400 38168 12541 38196
rect 12400 38156 12406 38168
rect 12529 38165 12541 38168
rect 12575 38165 12587 38199
rect 12529 38159 12587 38165
rect 1104 38106 16836 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 16836 38106
rect 1104 38032 16836 38054
rect 6638 37952 6644 38004
rect 6696 37952 6702 38004
rect 6809 37995 6867 38001
rect 6809 37961 6821 37995
rect 6855 37992 6867 37995
rect 7098 37992 7104 38004
rect 6855 37964 7104 37992
rect 6855 37961 6867 37964
rect 6809 37955 6867 37961
rect 7098 37952 7104 37964
rect 7156 37952 7162 38004
rect 7190 37952 7196 38004
rect 7248 37952 7254 38004
rect 7650 37952 7656 38004
rect 7708 37952 7714 38004
rect 8110 37992 8116 38004
rect 8168 38001 8174 38004
rect 8077 37964 8116 37992
rect 8110 37952 8116 37964
rect 8168 37955 8177 38001
rect 8205 37995 8263 38001
rect 8205 37961 8217 37995
rect 8251 37992 8263 37995
rect 8754 37992 8760 38004
rect 8251 37964 8760 37992
rect 8251 37961 8263 37964
rect 8205 37955 8263 37961
rect 8168 37952 8174 37955
rect 8754 37952 8760 37964
rect 8812 37992 8818 38004
rect 9950 37992 9956 38004
rect 8812 37964 9956 37992
rect 8812 37952 8818 37964
rect 9950 37952 9956 37964
rect 10008 37992 10014 38004
rect 10318 37992 10324 38004
rect 10008 37964 10324 37992
rect 10008 37952 10014 37964
rect 10318 37952 10324 37964
rect 10376 37952 10382 38004
rect 10594 37952 10600 38004
rect 10652 37992 10658 38004
rect 12069 37995 12127 38001
rect 12069 37992 12081 37995
rect 10652 37964 12081 37992
rect 10652 37952 10658 37964
rect 12069 37961 12081 37964
rect 12115 37961 12127 37995
rect 12069 37955 12127 37961
rect 12250 37952 12256 38004
rect 12308 37992 12314 38004
rect 12713 37995 12771 38001
rect 12713 37992 12725 37995
rect 12308 37964 12725 37992
rect 12308 37952 12314 37964
rect 12713 37961 12725 37964
rect 12759 37961 12771 37995
rect 12713 37955 12771 37961
rect 13078 37952 13084 38004
rect 13136 37952 13142 38004
rect 7006 37884 7012 37936
rect 7064 37884 7070 37936
rect 7668 37924 7696 37952
rect 7116 37896 7696 37924
rect 7745 37927 7803 37933
rect 7116 37865 7144 37896
rect 7745 37893 7757 37927
rect 7791 37924 7803 37927
rect 7834 37924 7840 37936
rect 7791 37896 7840 37924
rect 7791 37893 7803 37896
rect 7745 37887 7803 37893
rect 7834 37884 7840 37896
rect 7892 37924 7898 37936
rect 7892 37896 8340 37924
rect 7892 37884 7898 37896
rect 7101 37859 7159 37865
rect 7101 37825 7113 37859
rect 7147 37825 7159 37859
rect 7101 37819 7159 37825
rect 7285 37859 7343 37865
rect 7285 37825 7297 37859
rect 7331 37856 7343 37859
rect 7558 37856 7564 37868
rect 7331 37828 7564 37856
rect 7331 37825 7343 37828
rect 7285 37819 7343 37825
rect 7558 37816 7564 37828
rect 7616 37816 7622 37868
rect 7650 37816 7656 37868
rect 7708 37816 7714 37868
rect 8312 37865 8340 37896
rect 8021 37859 8079 37865
rect 8021 37825 8033 37859
rect 8067 37856 8079 37859
rect 8297 37859 8355 37865
rect 8067 37828 8156 37856
rect 8067 37825 8079 37828
rect 8021 37819 8079 37825
rect 7377 37723 7435 37729
rect 7377 37689 7389 37723
rect 7423 37720 7435 37723
rect 8128 37720 8156 37828
rect 8297 37825 8309 37859
rect 8343 37856 8355 37859
rect 8343 37828 8699 37856
rect 8343 37825 8355 37828
rect 8297 37819 8355 37825
rect 8389 37791 8447 37797
rect 8389 37757 8401 37791
rect 8435 37788 8447 37791
rect 8570 37788 8576 37800
rect 8435 37760 8576 37788
rect 8435 37757 8447 37760
rect 8389 37751 8447 37757
rect 8570 37748 8576 37760
rect 8628 37748 8634 37800
rect 8671 37788 8699 37828
rect 8754 37816 8760 37868
rect 8812 37865 8818 37868
rect 8812 37856 8822 37865
rect 8812 37828 8857 37856
rect 8812 37819 8822 37828
rect 8812 37816 8818 37819
rect 8849 37791 8907 37797
rect 8849 37788 8861 37791
rect 8671 37760 8861 37788
rect 8849 37757 8861 37760
rect 8895 37788 8907 37791
rect 10612 37788 10640 37952
rect 11241 37927 11299 37933
rect 11241 37893 11253 37927
rect 11287 37924 11299 37927
rect 12618 37924 12624 37936
rect 11287 37896 12624 37924
rect 11287 37893 11299 37896
rect 11241 37887 11299 37893
rect 12618 37884 12624 37896
rect 12676 37884 12682 37936
rect 12897 37927 12955 37933
rect 12897 37893 12909 37927
rect 12943 37924 12955 37927
rect 13541 37927 13599 37933
rect 13541 37924 13553 37927
rect 12943 37896 13553 37924
rect 12943 37893 12955 37896
rect 12897 37887 12955 37893
rect 13541 37893 13553 37896
rect 13587 37893 13599 37927
rect 13541 37887 13599 37893
rect 11054 37816 11060 37868
rect 11112 37856 11118 37868
rect 11517 37859 11575 37865
rect 11517 37856 11529 37859
rect 11112 37828 11529 37856
rect 11112 37816 11118 37828
rect 11517 37825 11529 37828
rect 11563 37825 11575 37859
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 11517 37819 11575 37825
rect 11624 37828 11713 37856
rect 8895 37760 10640 37788
rect 8895 37757 8907 37760
rect 8849 37751 8907 37757
rect 11238 37748 11244 37800
rect 11296 37788 11302 37800
rect 11624 37788 11652 37828
rect 11701 37825 11713 37828
rect 11747 37825 11759 37859
rect 11701 37819 11759 37825
rect 11793 37859 11851 37865
rect 11793 37825 11805 37859
rect 11839 37825 11851 37859
rect 11793 37819 11851 37825
rect 11885 37859 11943 37865
rect 11885 37825 11897 37859
rect 11931 37825 11943 37859
rect 11885 37819 11943 37825
rect 11808 37788 11836 37819
rect 11296 37760 11652 37788
rect 11716 37760 11836 37788
rect 11900 37788 11928 37819
rect 12066 37816 12072 37868
rect 12124 37856 12130 37868
rect 12161 37859 12219 37865
rect 12161 37856 12173 37859
rect 12124 37828 12173 37856
rect 12124 37816 12130 37828
rect 12161 37825 12173 37828
rect 12207 37825 12219 37859
rect 12161 37819 12219 37825
rect 12342 37816 12348 37868
rect 12400 37816 12406 37868
rect 12437 37859 12495 37865
rect 12437 37825 12449 37859
rect 12483 37856 12495 37859
rect 12483 37828 12572 37856
rect 12483 37825 12495 37828
rect 12437 37819 12495 37825
rect 12544 37788 12572 37828
rect 12802 37816 12808 37868
rect 12860 37816 12866 37868
rect 13173 37859 13231 37865
rect 13173 37825 13185 37859
rect 13219 37825 13231 37859
rect 13173 37819 13231 37825
rect 12618 37788 12624 37800
rect 11900 37760 12624 37788
rect 11296 37748 11302 37760
rect 11716 37732 11744 37760
rect 12618 37748 12624 37760
rect 12676 37788 12682 37800
rect 13188 37788 13216 37819
rect 13354 37816 13360 37868
rect 13412 37816 13418 37868
rect 12676 37760 13216 37788
rect 12676 37748 12682 37760
rect 8294 37720 8300 37732
rect 7423 37692 8300 37720
rect 7423 37689 7435 37692
rect 7377 37683 7435 37689
rect 8294 37680 8300 37692
rect 8352 37680 8358 37732
rect 11698 37680 11704 37732
rect 11756 37680 11762 37732
rect 12158 37680 12164 37732
rect 12216 37680 12222 37732
rect 12529 37723 12587 37729
rect 12529 37720 12541 37723
rect 12406 37692 12541 37720
rect 6822 37612 6828 37664
rect 6880 37612 6886 37664
rect 6914 37612 6920 37664
rect 6972 37652 6978 37664
rect 7929 37655 7987 37661
rect 7929 37652 7941 37655
rect 6972 37624 7941 37652
rect 6972 37612 6978 37624
rect 7929 37621 7941 37624
rect 7975 37621 7987 37655
rect 7929 37615 7987 37621
rect 10870 37612 10876 37664
rect 10928 37652 10934 37664
rect 10965 37655 11023 37661
rect 10965 37652 10977 37655
rect 10928 37624 10977 37652
rect 10928 37612 10934 37624
rect 10965 37621 10977 37624
rect 11011 37621 11023 37655
rect 10965 37615 11023 37621
rect 11146 37612 11152 37664
rect 11204 37652 11210 37664
rect 11882 37652 11888 37664
rect 11204 37624 11888 37652
rect 11204 37612 11210 37624
rect 11882 37612 11888 37624
rect 11940 37652 11946 37664
rect 12406 37652 12434 37692
rect 12529 37689 12541 37692
rect 12575 37689 12587 37723
rect 12529 37683 12587 37689
rect 11940 37624 12434 37652
rect 11940 37612 11946 37624
rect 1104 37562 16836 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 16836 37562
rect 1104 37488 16836 37510
rect 6822 37408 6828 37460
rect 6880 37448 6886 37460
rect 6917 37451 6975 37457
rect 6917 37448 6929 37451
rect 6880 37420 6929 37448
rect 6880 37408 6886 37420
rect 6917 37417 6929 37420
rect 6963 37448 6975 37451
rect 8662 37448 8668 37460
rect 6963 37420 8668 37448
rect 6963 37417 6975 37420
rect 6917 37411 6975 37417
rect 8662 37408 8668 37420
rect 8720 37408 8726 37460
rect 11514 37408 11520 37460
rect 11572 37408 11578 37460
rect 11698 37408 11704 37460
rect 11756 37408 11762 37460
rect 12713 37451 12771 37457
rect 12713 37417 12725 37451
rect 12759 37448 12771 37451
rect 12802 37448 12808 37460
rect 12759 37420 12808 37448
rect 12759 37417 12771 37420
rect 12713 37411 12771 37417
rect 12802 37408 12808 37420
rect 12860 37408 12866 37460
rect 10137 37383 10195 37389
rect 10137 37349 10149 37383
rect 10183 37380 10195 37383
rect 10594 37380 10600 37392
rect 10183 37352 10600 37380
rect 10183 37349 10195 37352
rect 10137 37343 10195 37349
rect 10594 37340 10600 37352
rect 10652 37340 10658 37392
rect 10870 37340 10876 37392
rect 10928 37380 10934 37392
rect 10928 37352 11376 37380
rect 10928 37340 10934 37352
rect 11348 37321 11376 37352
rect 10689 37315 10747 37321
rect 9968 37284 10548 37312
rect 9968 37256 9996 37284
rect 7006 37204 7012 37256
rect 7064 37204 7070 37256
rect 9858 37204 9864 37256
rect 9916 37204 9922 37256
rect 9950 37204 9956 37256
rect 10008 37204 10014 37256
rect 10520 37253 10548 37284
rect 10689 37281 10701 37315
rect 10735 37312 10747 37315
rect 11333 37315 11391 37321
rect 10735 37284 11100 37312
rect 10735 37281 10747 37284
rect 10689 37275 10747 37281
rect 11072 37256 11100 37284
rect 11333 37281 11345 37315
rect 11379 37281 11391 37315
rect 11333 37275 11391 37281
rect 11698 37272 11704 37324
rect 11756 37312 11762 37324
rect 12342 37312 12348 37324
rect 11756 37284 12348 37312
rect 11756 37272 11762 37284
rect 12342 37272 12348 37284
rect 12400 37312 12406 37324
rect 12400 37284 12848 37312
rect 12400 37272 12406 37284
rect 10413 37247 10471 37253
rect 10413 37244 10425 37247
rect 10060 37216 10425 37244
rect 7024 37176 7052 37204
rect 7101 37179 7159 37185
rect 7101 37176 7113 37179
rect 7024 37148 7113 37176
rect 7101 37145 7113 37148
rect 7147 37145 7159 37179
rect 9876 37176 9904 37204
rect 10060 37176 10088 37216
rect 10413 37213 10425 37216
rect 10459 37213 10471 37247
rect 10413 37207 10471 37213
rect 10505 37247 10563 37253
rect 10505 37213 10517 37247
rect 10551 37213 10563 37247
rect 10505 37207 10563 37213
rect 10778 37204 10784 37256
rect 10836 37204 10842 37256
rect 11054 37204 11060 37256
rect 11112 37204 11118 37256
rect 11238 37204 11244 37256
rect 11296 37204 11302 37256
rect 12618 37244 12624 37256
rect 11808 37216 12624 37244
rect 9876 37148 10088 37176
rect 10137 37179 10195 37185
rect 7101 37139 7159 37145
rect 10137 37145 10149 37179
rect 10183 37176 10195 37179
rect 10873 37179 10931 37185
rect 10873 37176 10885 37179
rect 10183 37148 10885 37176
rect 10183 37145 10195 37148
rect 10137 37139 10195 37145
rect 10873 37145 10885 37148
rect 10919 37145 10931 37179
rect 10873 37139 10931 37145
rect 11685 37179 11743 37185
rect 11685 37145 11697 37179
rect 11731 37176 11743 37179
rect 11808 37176 11836 37216
rect 12618 37204 12624 37216
rect 12676 37204 12682 37256
rect 12820 37253 12848 37284
rect 12805 37247 12863 37253
rect 12805 37213 12817 37247
rect 12851 37244 12863 37247
rect 13354 37244 13360 37256
rect 12851 37216 13360 37244
rect 12851 37213 12863 37216
rect 12805 37207 12863 37213
rect 13354 37204 13360 37216
rect 13412 37204 13418 37256
rect 11731 37148 11836 37176
rect 11885 37179 11943 37185
rect 11731 37145 11743 37148
rect 11685 37139 11743 37145
rect 11885 37145 11897 37179
rect 11931 37176 11943 37179
rect 12066 37176 12072 37188
rect 11931 37148 12072 37176
rect 11931 37145 11943 37148
rect 11885 37139 11943 37145
rect 6730 37068 6736 37120
rect 6788 37068 6794 37120
rect 6901 37111 6959 37117
rect 6901 37077 6913 37111
rect 6947 37108 6959 37111
rect 7006 37108 7012 37120
rect 6947 37080 7012 37108
rect 6947 37077 6959 37080
rect 6901 37071 6959 37077
rect 7006 37068 7012 37080
rect 7064 37068 7070 37120
rect 10042 37068 10048 37120
rect 10100 37108 10106 37120
rect 10229 37111 10287 37117
rect 10229 37108 10241 37111
rect 10100 37080 10241 37108
rect 10100 37068 10106 37080
rect 10229 37077 10241 37080
rect 10275 37077 10287 37111
rect 10229 37071 10287 37077
rect 11238 37068 11244 37120
rect 11296 37108 11302 37120
rect 11900 37108 11928 37139
rect 12066 37136 12072 37148
rect 12124 37136 12130 37188
rect 12636 37176 12664 37204
rect 12986 37176 12992 37188
rect 12636 37148 12992 37176
rect 12986 37136 12992 37148
rect 13044 37136 13050 37188
rect 11296 37080 11928 37108
rect 11296 37068 11302 37080
rect 1104 37018 16836 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 16836 37018
rect 1104 36944 16836 36966
rect 9861 36907 9919 36913
rect 9861 36873 9873 36907
rect 9907 36904 9919 36907
rect 9950 36904 9956 36916
rect 9907 36876 9956 36904
rect 9907 36873 9919 36876
rect 9861 36867 9919 36873
rect 9950 36864 9956 36876
rect 10008 36864 10014 36916
rect 2958 36845 2964 36848
rect 2945 36839 2964 36845
rect 2945 36805 2957 36839
rect 2945 36799 2964 36805
rect 2958 36796 2964 36799
rect 3016 36796 3022 36848
rect 3145 36839 3203 36845
rect 3145 36805 3157 36839
rect 3191 36805 3203 36839
rect 3145 36799 3203 36805
rect 6632 36839 6690 36845
rect 6632 36805 6644 36839
rect 6678 36836 6690 36839
rect 6730 36836 6736 36848
rect 6678 36808 6736 36836
rect 6678 36805 6690 36808
rect 6632 36799 6690 36805
rect 2038 36660 2044 36712
rect 2096 36700 2102 36712
rect 3160 36700 3188 36799
rect 6730 36796 6736 36808
rect 6788 36796 6794 36848
rect 9030 36796 9036 36848
rect 9088 36836 9094 36848
rect 11146 36836 11152 36848
rect 9088 36808 11152 36836
rect 9088 36796 9094 36808
rect 11146 36796 11152 36808
rect 11204 36796 11210 36848
rect 4062 36728 4068 36780
rect 4120 36768 4126 36780
rect 4229 36771 4287 36777
rect 4229 36768 4241 36771
rect 4120 36740 4241 36768
rect 4120 36728 4126 36740
rect 4229 36737 4241 36740
rect 4275 36737 4287 36771
rect 4229 36731 4287 36737
rect 6086 36728 6092 36780
rect 6144 36768 6150 36780
rect 6365 36771 6423 36777
rect 6365 36768 6377 36771
rect 6144 36740 6377 36768
rect 6144 36728 6150 36740
rect 6365 36737 6377 36740
rect 6411 36737 6423 36771
rect 6365 36731 6423 36737
rect 9769 36771 9827 36777
rect 9769 36737 9781 36771
rect 9815 36737 9827 36771
rect 9769 36731 9827 36737
rect 2096 36672 3188 36700
rect 2096 36660 2102 36672
rect 3602 36660 3608 36712
rect 3660 36700 3666 36712
rect 3973 36703 4031 36709
rect 3973 36700 3985 36703
rect 3660 36672 3985 36700
rect 3660 36660 3666 36672
rect 3973 36669 3985 36672
rect 4019 36669 4031 36703
rect 9784 36700 9812 36731
rect 10042 36728 10048 36780
rect 10100 36728 10106 36780
rect 10410 36728 10416 36780
rect 10468 36768 10474 36780
rect 10597 36771 10655 36777
rect 10597 36768 10609 36771
rect 10468 36740 10609 36768
rect 10468 36728 10474 36740
rect 10597 36737 10609 36740
rect 10643 36737 10655 36771
rect 10597 36731 10655 36737
rect 10689 36771 10747 36777
rect 10689 36737 10701 36771
rect 10735 36768 10747 36771
rect 11238 36768 11244 36780
rect 10735 36740 11244 36768
rect 10735 36737 10747 36740
rect 10689 36731 10747 36737
rect 11238 36728 11244 36740
rect 11296 36728 11302 36780
rect 9858 36700 9864 36712
rect 9784 36672 9864 36700
rect 3973 36663 4031 36669
rect 9858 36660 9864 36672
rect 9916 36700 9922 36712
rect 10226 36700 10232 36712
rect 9916 36672 10232 36700
rect 9916 36660 9922 36672
rect 10226 36660 10232 36672
rect 10284 36660 10290 36712
rect 10873 36703 10931 36709
rect 10873 36669 10885 36703
rect 10919 36700 10931 36703
rect 11698 36700 11704 36712
rect 10919 36672 11704 36700
rect 10919 36669 10931 36672
rect 10873 36663 10931 36669
rect 11698 36660 11704 36672
rect 11756 36660 11762 36712
rect 7926 36592 7932 36644
rect 7984 36632 7990 36644
rect 8202 36632 8208 36644
rect 7984 36604 8208 36632
rect 7984 36592 7990 36604
rect 8202 36592 8208 36604
rect 8260 36632 8266 36644
rect 12158 36632 12164 36644
rect 8260 36604 12164 36632
rect 8260 36592 8266 36604
rect 12158 36592 12164 36604
rect 12216 36592 12222 36644
rect 2774 36524 2780 36576
rect 2832 36524 2838 36576
rect 2961 36567 3019 36573
rect 2961 36533 2973 36567
rect 3007 36564 3019 36567
rect 3970 36564 3976 36576
rect 3007 36536 3976 36564
rect 3007 36533 3019 36536
rect 2961 36527 3019 36533
rect 3970 36524 3976 36536
rect 4028 36524 4034 36576
rect 5350 36524 5356 36576
rect 5408 36524 5414 36576
rect 7282 36524 7288 36576
rect 7340 36564 7346 36576
rect 7745 36567 7803 36573
rect 7745 36564 7757 36567
rect 7340 36536 7757 36564
rect 7340 36524 7346 36536
rect 7745 36533 7757 36536
rect 7791 36533 7803 36567
rect 7745 36527 7803 36533
rect 10045 36567 10103 36573
rect 10045 36533 10057 36567
rect 10091 36564 10103 36567
rect 10502 36564 10508 36576
rect 10091 36536 10508 36564
rect 10091 36533 10103 36536
rect 10045 36527 10103 36533
rect 10502 36524 10508 36536
rect 10560 36524 10566 36576
rect 10778 36524 10784 36576
rect 10836 36524 10842 36576
rect 1104 36474 16836 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 16836 36474
rect 1104 36400 16836 36422
rect 2038 36320 2044 36372
rect 2096 36320 2102 36372
rect 3973 36363 4031 36369
rect 3973 36329 3985 36363
rect 4019 36360 4031 36363
rect 4062 36360 4068 36372
rect 4019 36332 4068 36360
rect 4019 36329 4031 36332
rect 3973 36323 4031 36329
rect 4062 36320 4068 36332
rect 4120 36320 4126 36372
rect 4154 36320 4160 36372
rect 4212 36320 4218 36372
rect 6089 36363 6147 36369
rect 6089 36360 6101 36363
rect 4264 36332 6101 36360
rect 1949 36159 2007 36165
rect 1949 36125 1961 36159
rect 1995 36125 2007 36159
rect 1949 36119 2007 36125
rect 1964 36088 1992 36119
rect 2130 36116 2136 36168
rect 2188 36116 2194 36168
rect 2774 36116 2780 36168
rect 2832 36156 2838 36168
rect 3338 36159 3396 36165
rect 3338 36156 3350 36159
rect 2832 36128 3350 36156
rect 2832 36116 2838 36128
rect 3338 36125 3350 36128
rect 3384 36125 3396 36159
rect 3338 36119 3396 36125
rect 3602 36116 3608 36168
rect 3660 36116 3666 36168
rect 4141 36091 4199 36097
rect 1964 36060 2268 36088
rect 2240 36029 2268 36060
rect 4141 36057 4153 36091
rect 4187 36088 4199 36091
rect 4264 36088 4292 36332
rect 6089 36329 6101 36332
rect 6135 36329 6147 36363
rect 6089 36323 6147 36329
rect 7006 36320 7012 36372
rect 7064 36320 7070 36372
rect 10042 36320 10048 36372
rect 10100 36360 10106 36372
rect 11422 36360 11428 36372
rect 10100 36332 11428 36360
rect 10100 36320 10106 36332
rect 4632 36264 5764 36292
rect 4522 36116 4528 36168
rect 4580 36156 4586 36168
rect 4632 36165 4660 36264
rect 4706 36184 4712 36236
rect 4764 36224 4770 36236
rect 4764 36196 5304 36224
rect 4764 36184 4770 36196
rect 4617 36159 4675 36165
rect 4617 36156 4629 36159
rect 4580 36128 4629 36156
rect 4580 36116 4586 36128
rect 4617 36125 4629 36128
rect 4663 36125 4675 36159
rect 4617 36119 4675 36125
rect 4798 36116 4804 36168
rect 4856 36116 4862 36168
rect 4890 36116 4896 36168
rect 4948 36116 4954 36168
rect 5276 36165 5304 36196
rect 5261 36159 5319 36165
rect 5261 36125 5273 36159
rect 5307 36156 5319 36159
rect 5350 36156 5356 36168
rect 5307 36128 5356 36156
rect 5307 36125 5319 36128
rect 5261 36119 5319 36125
rect 5350 36116 5356 36128
rect 5408 36116 5414 36168
rect 5460 36158 5488 36264
rect 5736 36224 5764 36264
rect 6733 36227 6791 36233
rect 5736 36196 6408 36224
rect 5537 36159 5595 36165
rect 5537 36158 5549 36159
rect 5460 36130 5549 36158
rect 5537 36125 5549 36130
rect 5583 36125 5595 36159
rect 5537 36119 5595 36125
rect 5626 36116 5632 36168
rect 5684 36116 5690 36168
rect 5736 36156 5764 36196
rect 5813 36159 5871 36165
rect 5813 36156 5825 36159
rect 5736 36128 5825 36156
rect 5813 36125 5825 36128
rect 5859 36125 5871 36159
rect 5813 36119 5871 36125
rect 5902 36116 5908 36168
rect 5960 36116 5966 36168
rect 6380 36165 6408 36196
rect 6733 36193 6745 36227
rect 6779 36224 6791 36227
rect 6914 36224 6920 36236
rect 6779 36196 6920 36224
rect 6779 36193 6791 36196
rect 6733 36187 6791 36193
rect 6914 36184 6920 36196
rect 6972 36184 6978 36236
rect 6089 36159 6147 36165
rect 6089 36125 6101 36159
rect 6135 36156 6147 36159
rect 6365 36159 6423 36165
rect 6135 36128 6316 36156
rect 6135 36125 6147 36128
rect 6089 36119 6147 36125
rect 4187 36060 4292 36088
rect 4341 36091 4399 36097
rect 4187 36057 4199 36060
rect 4141 36051 4199 36057
rect 4341 36057 4353 36091
rect 4387 36088 4399 36091
rect 5077 36091 5135 36097
rect 5077 36088 5089 36091
rect 4387 36060 5089 36088
rect 4387 36057 4399 36060
rect 4341 36051 4399 36057
rect 5077 36057 5089 36060
rect 5123 36088 5135 36091
rect 5166 36088 5172 36100
rect 5123 36060 5172 36088
rect 5123 36057 5135 36060
rect 5077 36051 5135 36057
rect 5166 36048 5172 36060
rect 5224 36048 5230 36100
rect 5368 36088 5396 36116
rect 6181 36091 6239 36097
rect 6181 36088 6193 36091
rect 5368 36060 6193 36088
rect 6181 36057 6193 36060
rect 6227 36057 6239 36091
rect 6181 36051 6239 36057
rect 2225 36023 2283 36029
rect 2225 35989 2237 36023
rect 2271 36020 2283 36023
rect 3234 36020 3240 36032
rect 2271 35992 3240 36020
rect 2271 35989 2283 35992
rect 2225 35983 2283 35989
rect 3234 35980 3240 35992
rect 3292 35980 3298 36032
rect 4433 36023 4491 36029
rect 4433 35989 4445 36023
rect 4479 36020 4491 36023
rect 4614 36020 4620 36032
rect 4479 35992 4620 36020
rect 4479 35989 4491 35992
rect 4433 35983 4491 35989
rect 4614 35980 4620 35992
rect 4672 35980 4678 36032
rect 4982 35980 4988 36032
rect 5040 36020 5046 36032
rect 5350 36020 5356 36032
rect 5040 35992 5356 36020
rect 5040 35980 5046 35992
rect 5350 35980 5356 35992
rect 5408 36020 5414 36032
rect 5445 36023 5503 36029
rect 5445 36020 5457 36023
rect 5408 35992 5457 36020
rect 5408 35980 5414 35992
rect 5445 35989 5457 35992
rect 5491 36020 5503 36023
rect 6288 36020 6316 36128
rect 6365 36125 6377 36159
rect 6411 36125 6423 36159
rect 6365 36119 6423 36125
rect 6641 36159 6699 36165
rect 6641 36125 6653 36159
rect 6687 36156 6699 36159
rect 7190 36156 7196 36168
rect 6687 36128 7196 36156
rect 6687 36125 6699 36128
rect 6641 36119 6699 36125
rect 7190 36116 7196 36128
rect 7248 36116 7254 36168
rect 9122 36116 9128 36168
rect 9180 36116 9186 36168
rect 9401 36159 9459 36165
rect 9401 36125 9413 36159
rect 9447 36156 9459 36159
rect 9950 36156 9956 36168
rect 9447 36128 9956 36156
rect 9447 36125 9459 36128
rect 9401 36119 9459 36125
rect 9950 36116 9956 36128
rect 10008 36116 10014 36168
rect 10336 36165 10364 36332
rect 11422 36320 11428 36332
rect 11480 36320 11486 36372
rect 12158 36320 12164 36372
rect 12216 36360 12222 36372
rect 12253 36363 12311 36369
rect 12253 36360 12265 36363
rect 12216 36332 12265 36360
rect 12216 36320 12222 36332
rect 12253 36329 12265 36332
rect 12299 36329 12311 36363
rect 12253 36323 12311 36329
rect 10597 36295 10655 36301
rect 10597 36261 10609 36295
rect 10643 36292 10655 36295
rect 10778 36292 10784 36304
rect 10643 36264 10784 36292
rect 10643 36261 10655 36264
rect 10597 36255 10655 36261
rect 10778 36252 10784 36264
rect 10836 36252 10842 36304
rect 12066 36252 12072 36304
rect 12124 36292 12130 36304
rect 12529 36295 12587 36301
rect 12529 36292 12541 36295
rect 12124 36264 12541 36292
rect 12124 36252 12130 36264
rect 12529 36261 12541 36264
rect 12575 36261 12587 36295
rect 12529 36255 12587 36261
rect 10980 36196 11376 36224
rect 10321 36159 10379 36165
rect 10321 36125 10333 36159
rect 10367 36125 10379 36159
rect 10321 36119 10379 36125
rect 10505 36159 10563 36165
rect 10505 36125 10517 36159
rect 10551 36156 10563 36159
rect 10594 36156 10600 36168
rect 10551 36128 10600 36156
rect 10551 36125 10563 36128
rect 10505 36119 10563 36125
rect 10594 36116 10600 36128
rect 10652 36116 10658 36168
rect 10689 36159 10747 36165
rect 10689 36125 10701 36159
rect 10735 36125 10747 36159
rect 10689 36119 10747 36125
rect 10781 36159 10839 36165
rect 10781 36125 10793 36159
rect 10827 36158 10839 36159
rect 10980 36158 11008 36196
rect 10827 36130 11008 36158
rect 10827 36125 10839 36130
rect 10781 36119 10839 36125
rect 7098 36048 7104 36100
rect 7156 36088 7162 36100
rect 8021 36091 8079 36097
rect 8021 36088 8033 36091
rect 7156 36060 8033 36088
rect 7156 36048 7162 36060
rect 8021 36057 8033 36060
rect 8067 36057 8079 36091
rect 8021 36051 8079 36057
rect 8570 36048 8576 36100
rect 8628 36088 8634 36100
rect 9309 36091 9367 36097
rect 9309 36088 9321 36091
rect 8628 36060 9321 36088
rect 8628 36048 8634 36060
rect 9309 36057 9321 36060
rect 9355 36057 9367 36091
rect 10704 36088 10732 36119
rect 11146 36116 11152 36168
rect 11204 36156 11210 36168
rect 11241 36159 11299 36165
rect 11241 36156 11253 36159
rect 11204 36128 11253 36156
rect 11204 36116 11210 36128
rect 11241 36125 11253 36128
rect 11287 36125 11299 36159
rect 11348 36156 11376 36196
rect 11422 36184 11428 36236
rect 11480 36184 11486 36236
rect 13906 36184 13912 36236
rect 13964 36184 13970 36236
rect 11348 36128 11468 36156
rect 11241 36119 11299 36125
rect 11330 36088 11336 36100
rect 10704 36060 11336 36088
rect 9309 36051 9367 36057
rect 11330 36048 11336 36060
rect 11388 36048 11394 36100
rect 11440 36088 11468 36128
rect 11514 36116 11520 36168
rect 11572 36116 11578 36168
rect 11885 36159 11943 36165
rect 11885 36125 11897 36159
rect 11931 36156 11943 36159
rect 13078 36156 13084 36168
rect 11931 36128 13084 36156
rect 11931 36125 11943 36128
rect 11885 36119 11943 36125
rect 13078 36116 13084 36128
rect 13136 36116 13142 36168
rect 11609 36091 11667 36097
rect 11609 36088 11621 36091
rect 11440 36060 11621 36088
rect 11609 36057 11621 36060
rect 11655 36057 11667 36091
rect 11609 36051 11667 36057
rect 12802 36048 12808 36100
rect 12860 36088 12866 36100
rect 13642 36091 13700 36097
rect 13642 36088 13654 36091
rect 12860 36060 13654 36088
rect 12860 36048 12866 36060
rect 13642 36057 13654 36060
rect 13688 36057 13700 36091
rect 13642 36051 13700 36057
rect 5491 35992 6316 36020
rect 5491 35989 5503 35992
rect 5445 35983 5503 35989
rect 7466 35980 7472 36032
rect 7524 36020 7530 36032
rect 7929 36023 7987 36029
rect 7929 36020 7941 36023
rect 7524 35992 7941 36020
rect 7524 35980 7530 35992
rect 7929 35989 7941 35992
rect 7975 36020 7987 36023
rect 8202 36020 8208 36032
rect 7975 35992 8208 36020
rect 7975 35989 7987 35992
rect 7929 35983 7987 35989
rect 8202 35980 8208 35992
rect 8260 35980 8266 36032
rect 8941 36023 8999 36029
rect 8941 35989 8953 36023
rect 8987 36020 8999 36023
rect 9030 36020 9036 36032
rect 8987 35992 9036 36020
rect 8987 35989 8999 35992
rect 8941 35983 8999 35989
rect 9030 35980 9036 35992
rect 9088 35980 9094 36032
rect 10594 35980 10600 36032
rect 10652 36020 10658 36032
rect 10965 36023 11023 36029
rect 10965 36020 10977 36023
rect 10652 35992 10977 36020
rect 10652 35980 10658 35992
rect 10965 35989 10977 35992
rect 11011 35989 11023 36023
rect 10965 35983 11023 35989
rect 11054 35980 11060 36032
rect 11112 35980 11118 36032
rect 12250 35980 12256 36032
rect 12308 35980 12314 36032
rect 12434 35980 12440 36032
rect 12492 35980 12498 36032
rect 1104 35930 16836 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 16836 35930
rect 1104 35856 16836 35878
rect 2869 35819 2927 35825
rect 2869 35785 2881 35819
rect 2915 35816 2927 35819
rect 2958 35816 2964 35828
rect 2915 35788 2964 35816
rect 2915 35785 2927 35788
rect 2869 35779 2927 35785
rect 2958 35776 2964 35788
rect 3016 35776 3022 35828
rect 4798 35776 4804 35828
rect 4856 35816 4862 35828
rect 4856 35788 4936 35816
rect 4856 35776 4862 35788
rect 3234 35708 3240 35760
rect 3292 35748 3298 35760
rect 4522 35748 4528 35760
rect 3292 35720 4528 35748
rect 3292 35708 3298 35720
rect 4522 35708 4528 35720
rect 4580 35748 4586 35760
rect 4908 35757 4936 35788
rect 5258 35776 5264 35828
rect 5316 35816 5322 35828
rect 5534 35816 5540 35828
rect 5316 35788 5540 35816
rect 5316 35776 5322 35788
rect 5534 35776 5540 35788
rect 5592 35776 5598 35828
rect 7101 35819 7159 35825
rect 7101 35785 7113 35819
rect 7147 35816 7159 35819
rect 8297 35819 8355 35825
rect 8297 35816 8309 35819
rect 7147 35788 8309 35816
rect 7147 35785 7159 35788
rect 7101 35779 7159 35785
rect 8297 35785 8309 35788
rect 8343 35785 8355 35819
rect 8297 35779 8355 35785
rect 8570 35776 8576 35828
rect 8628 35776 8634 35828
rect 8941 35819 8999 35825
rect 8941 35785 8953 35819
rect 8987 35816 8999 35819
rect 9122 35816 9128 35828
rect 8987 35788 9128 35816
rect 8987 35785 8999 35788
rect 8941 35779 8999 35785
rect 9122 35776 9128 35788
rect 9180 35776 9186 35828
rect 9950 35776 9956 35828
rect 10008 35776 10014 35828
rect 10226 35776 10232 35828
rect 10284 35816 10290 35828
rect 11333 35819 11391 35825
rect 10284 35788 11192 35816
rect 10284 35776 10290 35788
rect 4709 35751 4767 35757
rect 4709 35748 4721 35751
rect 4580 35720 4721 35748
rect 4580 35708 4586 35720
rect 4709 35717 4721 35720
rect 4755 35717 4767 35751
rect 4709 35711 4767 35717
rect 4893 35751 4951 35757
rect 4893 35717 4905 35751
rect 4939 35748 4951 35751
rect 7285 35751 7343 35757
rect 4939 35720 5764 35748
rect 4939 35717 4951 35720
rect 4893 35711 4951 35717
rect 5736 35692 5764 35720
rect 7285 35717 7297 35751
rect 7331 35748 7343 35751
rect 8414 35751 8472 35757
rect 8414 35748 8426 35751
rect 7331 35720 8426 35748
rect 7331 35717 7343 35720
rect 7285 35711 7343 35717
rect 8414 35717 8426 35720
rect 8460 35717 8472 35751
rect 8588 35748 8616 35776
rect 8588 35720 9628 35748
rect 8414 35711 8472 35717
rect 2130 35640 2136 35692
rect 2188 35680 2194 35692
rect 3053 35683 3111 35689
rect 3053 35680 3065 35683
rect 2188 35652 3065 35680
rect 2188 35640 2194 35652
rect 3053 35649 3065 35652
rect 3099 35649 3111 35683
rect 3053 35643 3111 35649
rect 3068 35612 3096 35643
rect 4798 35640 4804 35692
rect 4856 35640 4862 35692
rect 5445 35683 5503 35689
rect 5445 35649 5457 35683
rect 5491 35649 5503 35683
rect 5445 35643 5503 35649
rect 5077 35615 5135 35621
rect 5077 35612 5089 35615
rect 3068 35584 5089 35612
rect 5077 35581 5089 35584
rect 5123 35612 5135 35615
rect 5350 35612 5356 35624
rect 5123 35584 5356 35612
rect 5123 35581 5135 35584
rect 5077 35575 5135 35581
rect 5350 35572 5356 35584
rect 5408 35572 5414 35624
rect 5460 35612 5488 35643
rect 5534 35640 5540 35692
rect 5592 35640 5598 35692
rect 5626 35640 5632 35692
rect 5684 35640 5690 35692
rect 5718 35640 5724 35692
rect 5776 35640 5782 35692
rect 6730 35640 6736 35692
rect 6788 35640 6794 35692
rect 7190 35640 7196 35692
rect 7248 35640 7254 35692
rect 7377 35683 7435 35689
rect 7377 35649 7389 35683
rect 7423 35680 7435 35683
rect 7466 35680 7472 35692
rect 7423 35652 7472 35680
rect 7423 35649 7435 35652
rect 7377 35643 7435 35649
rect 7466 35640 7472 35652
rect 7524 35640 7530 35692
rect 7653 35683 7711 35689
rect 7653 35649 7665 35683
rect 7699 35649 7711 35683
rect 7653 35643 7711 35649
rect 7837 35683 7895 35689
rect 7837 35649 7849 35683
rect 7883 35680 7895 35683
rect 8205 35683 8263 35689
rect 8205 35680 8217 35683
rect 7883 35652 8217 35680
rect 7883 35649 7895 35652
rect 7837 35643 7895 35649
rect 8205 35649 8217 35652
rect 8251 35649 8263 35683
rect 8205 35643 8263 35649
rect 8665 35683 8723 35689
rect 8665 35649 8677 35683
rect 8711 35680 8723 35683
rect 9217 35683 9275 35689
rect 8711 35652 8892 35680
rect 8711 35649 8723 35652
rect 8665 35643 8723 35649
rect 5994 35612 6000 35624
rect 5460 35584 6000 35612
rect 5994 35572 6000 35584
rect 6052 35612 6058 35624
rect 6641 35615 6699 35621
rect 6641 35612 6653 35615
rect 6052 35584 6653 35612
rect 6052 35572 6058 35584
rect 6641 35581 6653 35584
rect 6687 35581 6699 35615
rect 7208 35612 7236 35640
rect 7668 35612 7696 35643
rect 7208 35584 7696 35612
rect 6641 35575 6699 35581
rect 4154 35436 4160 35488
rect 4212 35476 4218 35488
rect 4525 35479 4583 35485
rect 4525 35476 4537 35479
rect 4212 35448 4537 35476
rect 4212 35436 4218 35448
rect 4525 35445 4537 35448
rect 4571 35476 4583 35479
rect 4706 35476 4712 35488
rect 4571 35448 4712 35476
rect 4571 35445 4583 35448
rect 4525 35439 4583 35445
rect 4706 35436 4712 35448
rect 4764 35436 4770 35488
rect 5261 35479 5319 35485
rect 5261 35445 5273 35479
rect 5307 35476 5319 35479
rect 5350 35476 5356 35488
rect 5307 35448 5356 35476
rect 5307 35445 5319 35448
rect 5261 35439 5319 35445
rect 5350 35436 5356 35448
rect 5408 35436 5414 35488
rect 7668 35476 7696 35584
rect 7929 35615 7987 35621
rect 7929 35581 7941 35615
rect 7975 35612 7987 35615
rect 8018 35612 8024 35624
rect 7975 35584 8024 35612
rect 7975 35581 7987 35584
rect 7929 35575 7987 35581
rect 8018 35572 8024 35584
rect 8076 35572 8082 35624
rect 8220 35612 8248 35643
rect 8757 35615 8815 35621
rect 8757 35612 8769 35615
rect 8220 35584 8769 35612
rect 8757 35581 8769 35584
rect 8803 35581 8815 35615
rect 8757 35575 8815 35581
rect 7834 35504 7840 35556
rect 7892 35544 7898 35556
rect 8864 35544 8892 35652
rect 9217 35649 9229 35683
rect 9263 35649 9275 35683
rect 9217 35643 9275 35649
rect 9401 35683 9459 35689
rect 9401 35649 9413 35683
rect 9447 35680 9459 35683
rect 9490 35680 9496 35692
rect 9447 35652 9496 35680
rect 9447 35649 9459 35652
rect 9401 35643 9459 35649
rect 8938 35572 8944 35624
rect 8996 35572 9002 35624
rect 9232 35612 9260 35643
rect 9490 35640 9496 35652
rect 9548 35640 9554 35692
rect 9600 35689 9628 35720
rect 10318 35708 10324 35760
rect 10376 35748 10382 35760
rect 11054 35748 11060 35760
rect 10376 35720 11060 35748
rect 10376 35708 10382 35720
rect 11054 35708 11060 35720
rect 11112 35708 11118 35760
rect 11164 35748 11192 35788
rect 11333 35785 11345 35819
rect 11379 35816 11391 35819
rect 11514 35816 11520 35828
rect 11379 35788 11520 35816
rect 11379 35785 11391 35788
rect 11333 35779 11391 35785
rect 11514 35776 11520 35788
rect 11572 35776 11578 35828
rect 13078 35776 13084 35828
rect 13136 35816 13142 35828
rect 14001 35819 14059 35825
rect 14001 35816 14013 35819
rect 13136 35788 14013 35816
rect 13136 35776 13142 35788
rect 14001 35785 14013 35788
rect 14047 35785 14059 35819
rect 14001 35779 14059 35785
rect 11422 35748 11428 35760
rect 11164 35720 11428 35748
rect 11422 35708 11428 35720
rect 11480 35748 11486 35760
rect 11701 35751 11759 35757
rect 11701 35748 11713 35751
rect 11480 35720 11713 35748
rect 11480 35708 11486 35720
rect 11701 35717 11713 35720
rect 11747 35717 11759 35751
rect 11701 35711 11759 35717
rect 12158 35708 12164 35760
rect 12216 35708 12222 35760
rect 12342 35708 12348 35760
rect 12400 35757 12406 35760
rect 12400 35751 12419 35757
rect 12407 35717 12419 35751
rect 12400 35711 12419 35717
rect 12400 35708 12406 35711
rect 12526 35708 12532 35760
rect 12584 35748 12590 35760
rect 12866 35751 12924 35757
rect 12866 35748 12878 35751
rect 12584 35720 12878 35748
rect 12584 35708 12590 35720
rect 12866 35717 12878 35720
rect 12912 35717 12924 35751
rect 12866 35711 12924 35717
rect 9585 35683 9643 35689
rect 9585 35649 9597 35683
rect 9631 35649 9643 35683
rect 9585 35643 9643 35649
rect 9861 35683 9919 35689
rect 9861 35649 9873 35683
rect 9907 35680 9919 35683
rect 9950 35680 9956 35692
rect 9907 35652 9956 35680
rect 9907 35649 9919 35652
rect 9861 35643 9919 35649
rect 9950 35640 9956 35652
rect 10008 35640 10014 35692
rect 10137 35683 10195 35689
rect 10137 35649 10149 35683
rect 10183 35649 10195 35683
rect 10137 35643 10195 35649
rect 9674 35612 9680 35624
rect 9232 35584 9680 35612
rect 7892 35516 8892 35544
rect 7892 35504 7898 35516
rect 8110 35476 8116 35488
rect 7668 35448 8116 35476
rect 8110 35436 8116 35448
rect 8168 35436 8174 35488
rect 8202 35436 8208 35488
rect 8260 35476 8266 35488
rect 9232 35476 9260 35584
rect 9674 35572 9680 35584
rect 9732 35572 9738 35624
rect 9766 35572 9772 35624
rect 9824 35612 9830 35624
rect 10152 35612 10180 35643
rect 10226 35640 10232 35692
rect 10284 35640 10290 35692
rect 10502 35640 10508 35692
rect 10560 35640 10566 35692
rect 10594 35640 10600 35692
rect 10652 35640 10658 35692
rect 10781 35683 10839 35689
rect 10781 35649 10793 35683
rect 10827 35680 10839 35683
rect 12066 35680 12072 35692
rect 10827 35652 11008 35680
rect 10827 35649 10839 35652
rect 10781 35643 10839 35649
rect 10980 35624 11008 35652
rect 11164 35652 12072 35680
rect 9824 35584 10180 35612
rect 9824 35572 9830 35584
rect 10962 35572 10968 35624
rect 11020 35572 11026 35624
rect 11057 35615 11115 35621
rect 11057 35581 11069 35615
rect 11103 35581 11115 35615
rect 11057 35575 11115 35581
rect 10870 35504 10876 35556
rect 10928 35544 10934 35556
rect 11072 35544 11100 35575
rect 10928 35516 11100 35544
rect 10928 35504 10934 35516
rect 8260 35448 9260 35476
rect 8260 35436 8266 35448
rect 9858 35436 9864 35488
rect 9916 35436 9922 35488
rect 11164 35485 11192 35652
rect 12066 35640 12072 35652
rect 12124 35640 12130 35692
rect 12434 35612 12440 35624
rect 11716 35584 12440 35612
rect 11330 35504 11336 35556
rect 11388 35544 11394 35556
rect 11517 35547 11575 35553
rect 11517 35544 11529 35547
rect 11388 35516 11529 35544
rect 11388 35504 11394 35516
rect 11517 35513 11529 35516
rect 11563 35513 11575 35547
rect 11517 35507 11575 35513
rect 11716 35485 11744 35584
rect 12434 35572 12440 35584
rect 12492 35572 12498 35624
rect 12618 35572 12624 35624
rect 12676 35572 12682 35624
rect 11149 35479 11207 35485
rect 11149 35445 11161 35479
rect 11195 35445 11207 35479
rect 11149 35439 11207 35445
rect 11701 35479 11759 35485
rect 11701 35445 11713 35479
rect 11747 35445 11759 35479
rect 11701 35439 11759 35445
rect 12250 35436 12256 35488
rect 12308 35476 12314 35488
rect 12345 35479 12403 35485
rect 12345 35476 12357 35479
rect 12308 35448 12357 35476
rect 12308 35436 12314 35448
rect 12345 35445 12357 35448
rect 12391 35445 12403 35479
rect 12345 35439 12403 35445
rect 12529 35479 12587 35485
rect 12529 35445 12541 35479
rect 12575 35476 12587 35479
rect 12802 35476 12808 35488
rect 12575 35448 12808 35476
rect 12575 35445 12587 35448
rect 12529 35439 12587 35445
rect 12802 35436 12808 35448
rect 12860 35436 12866 35488
rect 1104 35386 16836 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 16836 35386
rect 1104 35312 16836 35334
rect 2130 35232 2136 35284
rect 2188 35272 2194 35284
rect 2225 35275 2283 35281
rect 2225 35272 2237 35275
rect 2188 35244 2237 35272
rect 2188 35232 2194 35244
rect 2225 35241 2237 35244
rect 2271 35241 2283 35275
rect 2225 35235 2283 35241
rect 4157 35275 4215 35281
rect 4157 35241 4169 35275
rect 4203 35272 4215 35275
rect 4614 35272 4620 35284
rect 4203 35244 4620 35272
rect 4203 35241 4215 35244
rect 4157 35235 4215 35241
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 5718 35232 5724 35284
rect 5776 35272 5782 35284
rect 5813 35275 5871 35281
rect 5813 35272 5825 35275
rect 5776 35244 5825 35272
rect 5776 35232 5782 35244
rect 5813 35241 5825 35244
rect 5859 35241 5871 35275
rect 5813 35235 5871 35241
rect 5994 35232 6000 35284
rect 6052 35232 6058 35284
rect 8018 35232 8024 35284
rect 8076 35232 8082 35284
rect 8386 35232 8392 35284
rect 8444 35232 8450 35284
rect 8588 35244 8800 35272
rect 3789 35207 3847 35213
rect 3789 35173 3801 35207
rect 3835 35204 3847 35207
rect 4062 35204 4068 35216
rect 3835 35176 4068 35204
rect 3835 35173 3847 35176
rect 3789 35167 3847 35173
rect 4062 35164 4068 35176
rect 4120 35164 4126 35216
rect 5902 35164 5908 35216
rect 5960 35204 5966 35216
rect 6181 35207 6239 35213
rect 6181 35204 6193 35207
rect 5960 35176 6193 35204
rect 5960 35164 5966 35176
rect 6181 35173 6193 35176
rect 6227 35204 6239 35207
rect 6822 35204 6828 35216
rect 6227 35176 6828 35204
rect 6227 35173 6239 35176
rect 6181 35167 6239 35173
rect 6822 35164 6828 35176
rect 6880 35164 6886 35216
rect 3602 35028 3608 35080
rect 3660 35028 3666 35080
rect 4433 35071 4491 35077
rect 4433 35037 4445 35071
rect 4479 35068 4491 35071
rect 6086 35068 6092 35080
rect 4479 35040 6092 35068
rect 4479 35037 4491 35040
rect 4433 35031 4491 35037
rect 6086 35028 6092 35040
rect 6144 35028 6150 35080
rect 7558 35028 7564 35080
rect 7616 35068 7622 35080
rect 7653 35071 7711 35077
rect 7653 35068 7665 35071
rect 7616 35040 7665 35068
rect 7616 35028 7622 35040
rect 7653 35037 7665 35040
rect 7699 35037 7711 35071
rect 7653 35031 7711 35037
rect 7834 35028 7840 35080
rect 7892 35028 7898 35080
rect 8036 35068 8064 35232
rect 8110 35096 8116 35148
rect 8168 35136 8174 35148
rect 8297 35139 8355 35145
rect 8297 35136 8309 35139
rect 8168 35108 8309 35136
rect 8168 35096 8174 35108
rect 8297 35105 8309 35108
rect 8343 35105 8355 35139
rect 8297 35099 8355 35105
rect 8205 35071 8263 35077
rect 8205 35068 8217 35071
rect 8036 35040 8217 35068
rect 8205 35037 8217 35040
rect 8251 35037 8263 35071
rect 8205 35031 8263 35037
rect 8481 35071 8539 35077
rect 8481 35037 8493 35071
rect 8527 35068 8539 35071
rect 8588 35068 8616 35244
rect 8665 35207 8723 35213
rect 8665 35173 8677 35207
rect 8711 35173 8723 35207
rect 8772 35204 8800 35244
rect 8938 35232 8944 35284
rect 8996 35232 9002 35284
rect 9766 35232 9772 35284
rect 9824 35232 9830 35284
rect 9950 35232 9956 35284
rect 10008 35232 10014 35284
rect 10137 35275 10195 35281
rect 10137 35241 10149 35275
rect 10183 35272 10195 35275
rect 10226 35272 10232 35284
rect 10183 35244 10232 35272
rect 10183 35241 10195 35244
rect 10137 35235 10195 35241
rect 10226 35232 10232 35244
rect 10284 35272 10290 35284
rect 10965 35275 11023 35281
rect 10965 35272 10977 35275
rect 10284 35244 10977 35272
rect 10284 35232 10290 35244
rect 10965 35241 10977 35244
rect 11011 35241 11023 35275
rect 10965 35235 11023 35241
rect 12342 35232 12348 35284
rect 12400 35272 12406 35284
rect 12400 35244 12848 35272
rect 12400 35232 12406 35244
rect 9306 35204 9312 35216
rect 8772 35176 9312 35204
rect 8665 35167 8723 35173
rect 8527 35040 8616 35068
rect 8680 35068 8708 35167
rect 9306 35164 9312 35176
rect 9364 35204 9370 35216
rect 10410 35204 10416 35216
rect 9364 35176 10416 35204
rect 9364 35164 9370 35176
rect 10410 35164 10416 35176
rect 10468 35164 10474 35216
rect 10597 35207 10655 35213
rect 10597 35173 10609 35207
rect 10643 35204 10655 35207
rect 10778 35204 10784 35216
rect 10643 35176 10784 35204
rect 10643 35173 10655 35176
rect 10597 35167 10655 35173
rect 10778 35164 10784 35176
rect 10836 35164 10842 35216
rect 9401 35139 9459 35145
rect 9401 35105 9413 35139
rect 9447 35136 9459 35139
rect 9447 35108 9674 35136
rect 9447 35105 9459 35108
rect 9401 35099 9459 35105
rect 9646 35080 9674 35108
rect 9950 35096 9956 35148
rect 10008 35136 10014 35148
rect 12250 35136 12256 35148
rect 10008 35108 12256 35136
rect 10008 35096 10014 35108
rect 12250 35096 12256 35108
rect 12308 35096 12314 35148
rect 12820 35145 12848 35244
rect 12529 35139 12587 35145
rect 12529 35105 12541 35139
rect 12575 35136 12587 35139
rect 12805 35139 12863 35145
rect 12575 35108 12756 35136
rect 12575 35105 12587 35108
rect 12529 35099 12587 35105
rect 9125 35071 9183 35077
rect 9125 35068 9137 35071
rect 8680 35040 9137 35068
rect 8527 35037 8539 35040
rect 8481 35031 8539 35037
rect 9125 35037 9137 35040
rect 9171 35037 9183 35071
rect 9125 35031 9183 35037
rect 9217 35071 9275 35077
rect 9217 35037 9229 35071
rect 9263 35037 9275 35071
rect 9217 35031 9275 35037
rect 3050 34960 3056 35012
rect 3108 35000 3114 35012
rect 3338 35003 3396 35009
rect 3338 35000 3350 35003
rect 3108 34972 3350 35000
rect 3108 34960 3114 34972
rect 3338 34969 3350 34972
rect 3384 34969 3396 35003
rect 4678 35003 4736 35009
rect 4678 35000 4690 35003
rect 3338 34963 3396 34969
rect 4356 34972 4690 35000
rect 4154 34892 4160 34944
rect 4212 34892 4218 34944
rect 4356 34941 4384 34972
rect 4678 34969 4690 34972
rect 4724 34969 4736 35003
rect 4678 34963 4736 34969
rect 5534 34960 5540 35012
rect 5592 35000 5598 35012
rect 6457 35003 6515 35009
rect 6457 35000 6469 35003
rect 5592 34972 6469 35000
rect 5592 34960 5598 34972
rect 6457 34969 6469 34972
rect 6503 34969 6515 35003
rect 6457 34963 6515 34969
rect 6730 34960 6736 35012
rect 6788 35000 6794 35012
rect 8294 35000 8300 35012
rect 6788 34972 8300 35000
rect 6788 34960 6794 34972
rect 8294 34960 8300 34972
rect 8352 35000 8358 35012
rect 9232 35000 9260 35031
rect 9490 35028 9496 35080
rect 9548 35028 9554 35080
rect 9646 35040 9680 35080
rect 9674 35028 9680 35040
rect 9732 35028 9738 35080
rect 9861 35071 9919 35077
rect 9861 35037 9873 35071
rect 9907 35068 9919 35071
rect 9907 35040 10456 35068
rect 9907 35037 9919 35040
rect 9861 35031 9919 35037
rect 8352 34972 9260 35000
rect 9692 35000 9720 35028
rect 10428 35012 10456 35040
rect 10502 35028 10508 35080
rect 10560 35068 10566 35080
rect 10689 35071 10747 35077
rect 10689 35068 10701 35071
rect 10560 35040 10701 35068
rect 10560 35028 10566 35040
rect 10689 35037 10701 35040
rect 10735 35037 10747 35071
rect 10689 35031 10747 35037
rect 11241 35071 11299 35077
rect 11241 35037 11253 35071
rect 11287 35037 11299 35071
rect 11241 35031 11299 35037
rect 10226 35000 10232 35012
rect 9692 34972 10232 35000
rect 8352 34960 8358 34972
rect 10226 34960 10232 34972
rect 10284 34960 10290 35012
rect 10318 34960 10324 35012
rect 10376 34960 10382 35012
rect 10410 34960 10416 35012
rect 10468 34960 10474 35012
rect 4341 34935 4399 34941
rect 4341 34901 4353 34935
rect 4387 34901 4399 34935
rect 4341 34895 4399 34901
rect 10121 34935 10179 34941
rect 10121 34901 10133 34935
rect 10167 34932 10179 34935
rect 10689 34935 10747 34941
rect 10689 34932 10701 34935
rect 10167 34904 10701 34932
rect 10167 34901 10179 34904
rect 10121 34895 10179 34901
rect 10689 34901 10701 34904
rect 10735 34901 10747 34935
rect 11256 34932 11284 35031
rect 11330 35028 11336 35080
rect 11388 35028 11394 35080
rect 11425 35071 11483 35077
rect 11425 35037 11437 35071
rect 11471 35068 11483 35071
rect 11514 35068 11520 35080
rect 11471 35040 11520 35068
rect 11471 35037 11483 35040
rect 11425 35031 11483 35037
rect 11514 35028 11520 35040
rect 11572 35028 11578 35080
rect 11606 35028 11612 35080
rect 11664 35028 11670 35080
rect 12728 35077 12756 35108
rect 12805 35105 12817 35139
rect 12851 35105 12863 35139
rect 12805 35099 12863 35105
rect 12443 35071 12501 35077
rect 12443 35037 12455 35071
rect 12489 35037 12501 35071
rect 12443 35031 12501 35037
rect 12621 35071 12679 35077
rect 12621 35037 12633 35071
rect 12667 35037 12679 35071
rect 12621 35031 12679 35037
rect 12713 35071 12771 35077
rect 12713 35037 12725 35071
rect 12759 35037 12771 35071
rect 12713 35031 12771 35037
rect 12897 35071 12955 35077
rect 12897 35037 12909 35071
rect 12943 35068 12955 35071
rect 12986 35068 12992 35080
rect 12943 35040 12992 35068
rect 12943 35037 12955 35040
rect 12897 35031 12955 35037
rect 12066 34960 12072 35012
rect 12124 35000 12130 35012
rect 12452 35000 12480 35031
rect 12124 34972 12480 35000
rect 12124 34960 12130 34972
rect 12434 34932 12440 34944
rect 11256 34904 12440 34932
rect 10689 34895 10747 34901
rect 12434 34892 12440 34904
rect 12492 34892 12498 34944
rect 12636 34932 12664 35031
rect 12986 35028 12992 35040
rect 13044 35028 13050 35080
rect 12710 34932 12716 34944
rect 12636 34904 12716 34932
rect 12710 34892 12716 34904
rect 12768 34892 12774 34944
rect 1104 34842 16836 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 16836 34842
rect 1104 34768 16836 34790
rect 3050 34688 3056 34740
rect 3108 34688 3114 34740
rect 8386 34688 8392 34740
rect 8444 34728 8450 34740
rect 11146 34728 11152 34740
rect 8444 34700 11152 34728
rect 8444 34688 8450 34700
rect 11146 34688 11152 34700
rect 11204 34688 11210 34740
rect 2130 34620 2136 34672
rect 2188 34660 2194 34672
rect 2593 34663 2651 34669
rect 2593 34660 2605 34663
rect 2188 34632 2605 34660
rect 2188 34620 2194 34632
rect 2593 34629 2605 34632
rect 2639 34629 2651 34663
rect 2593 34623 2651 34629
rect 10686 34620 10692 34672
rect 10744 34660 10750 34672
rect 11330 34660 11336 34672
rect 10744 34632 11336 34660
rect 10744 34620 10750 34632
rect 11330 34620 11336 34632
rect 11388 34620 11394 34672
rect 12897 34663 12955 34669
rect 12897 34660 12909 34663
rect 12728 34632 12909 34660
rect 12728 34604 12756 34632
rect 12897 34629 12909 34632
rect 12943 34629 12955 34663
rect 13170 34660 13176 34672
rect 12897 34623 12955 34629
rect 13004 34632 13176 34660
rect 7377 34595 7435 34601
rect 7377 34561 7389 34595
rect 7423 34592 7435 34595
rect 7466 34592 7472 34604
rect 7423 34564 7472 34592
rect 7423 34561 7435 34564
rect 7377 34555 7435 34561
rect 7466 34552 7472 34564
rect 7524 34552 7530 34604
rect 7561 34595 7619 34601
rect 7561 34561 7573 34595
rect 7607 34592 7619 34595
rect 8202 34592 8208 34604
rect 7607 34564 8208 34592
rect 7607 34561 7619 34564
rect 7561 34555 7619 34561
rect 8202 34552 8208 34564
rect 8260 34552 8266 34604
rect 12250 34552 12256 34604
rect 12308 34552 12314 34604
rect 12526 34552 12532 34604
rect 12584 34552 12590 34604
rect 12710 34552 12716 34604
rect 12768 34552 12774 34604
rect 12802 34552 12808 34604
rect 12860 34552 12866 34604
rect 13004 34601 13032 34632
rect 13170 34620 13176 34632
rect 13228 34620 13234 34672
rect 12989 34595 13047 34601
rect 12989 34561 13001 34595
rect 13035 34561 13047 34595
rect 12989 34555 13047 34561
rect 13078 34552 13084 34604
rect 13136 34552 13142 34604
rect 13265 34595 13323 34601
rect 13265 34561 13277 34595
rect 13311 34592 13323 34595
rect 13354 34592 13360 34604
rect 13311 34564 13360 34592
rect 13311 34561 13323 34564
rect 13265 34555 13323 34561
rect 13354 34552 13360 34564
rect 13412 34552 13418 34604
rect 12161 34527 12219 34533
rect 12161 34493 12173 34527
rect 12207 34524 12219 34527
rect 12434 34524 12440 34536
rect 12207 34496 12440 34524
rect 12207 34493 12219 34496
rect 12161 34487 12219 34493
rect 2866 34416 2872 34468
rect 2924 34456 2930 34468
rect 4154 34456 4160 34468
rect 2924 34428 4160 34456
rect 2924 34416 2930 34428
rect 4154 34416 4160 34428
rect 4212 34416 4218 34468
rect 7282 34416 7288 34468
rect 7340 34456 7346 34468
rect 8662 34456 8668 34468
rect 7340 34428 8668 34456
rect 7340 34416 7346 34428
rect 8662 34416 8668 34428
rect 8720 34456 8726 34468
rect 9214 34456 9220 34468
rect 8720 34428 9220 34456
rect 8720 34416 8726 34428
rect 9214 34416 9220 34428
rect 9272 34416 9278 34468
rect 12360 34456 12388 34496
rect 12434 34484 12440 34496
rect 12492 34484 12498 34536
rect 12621 34527 12679 34533
rect 12621 34493 12633 34527
rect 12667 34524 12679 34527
rect 12894 34524 12900 34536
rect 12667 34496 12900 34524
rect 12667 34493 12679 34496
rect 12621 34487 12679 34493
rect 12894 34484 12900 34496
rect 12952 34484 12958 34536
rect 12802 34456 12808 34468
rect 12360 34428 12808 34456
rect 12802 34416 12808 34428
rect 12860 34416 12866 34468
rect 7190 34348 7196 34400
rect 7248 34388 7254 34400
rect 7377 34391 7435 34397
rect 7377 34388 7389 34391
rect 7248 34360 7389 34388
rect 7248 34348 7254 34360
rect 7377 34357 7389 34360
rect 7423 34357 7435 34391
rect 7377 34351 7435 34357
rect 9030 34348 9036 34400
rect 9088 34388 9094 34400
rect 12342 34388 12348 34400
rect 9088 34360 12348 34388
rect 9088 34348 9094 34360
rect 12342 34348 12348 34360
rect 12400 34348 12406 34400
rect 12710 34348 12716 34400
rect 12768 34388 12774 34400
rect 12986 34388 12992 34400
rect 12768 34360 12992 34388
rect 12768 34348 12774 34360
rect 12986 34348 12992 34360
rect 13044 34348 13050 34400
rect 1104 34298 16836 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 16836 34298
rect 1104 34224 16836 34246
rect 4522 34144 4528 34196
rect 4580 34184 4586 34196
rect 4617 34187 4675 34193
rect 4617 34184 4629 34187
rect 4580 34156 4629 34184
rect 4580 34144 4586 34156
rect 4617 34153 4629 34156
rect 4663 34153 4675 34187
rect 4617 34147 4675 34153
rect 5077 34187 5135 34193
rect 5077 34153 5089 34187
rect 5123 34184 5135 34187
rect 5902 34184 5908 34196
rect 5123 34156 5908 34184
rect 5123 34153 5135 34156
rect 5077 34147 5135 34153
rect 4154 34076 4160 34128
rect 4212 34116 4218 34128
rect 4893 34119 4951 34125
rect 4893 34116 4905 34119
rect 4212 34088 4905 34116
rect 4212 34076 4218 34088
rect 4893 34085 4905 34088
rect 4939 34085 4951 34119
rect 4893 34079 4951 34085
rect 4430 34008 4436 34060
rect 4488 34048 4494 34060
rect 5092 34048 5120 34147
rect 5902 34144 5908 34156
rect 5960 34144 5966 34196
rect 7193 34187 7251 34193
rect 7193 34153 7205 34187
rect 7239 34184 7251 34187
rect 7282 34184 7288 34196
rect 7239 34156 7288 34184
rect 7239 34153 7251 34156
rect 7193 34147 7251 34153
rect 7282 34144 7288 34156
rect 7340 34144 7346 34196
rect 7653 34187 7711 34193
rect 7653 34153 7665 34187
rect 7699 34184 7711 34187
rect 7834 34184 7840 34196
rect 7699 34156 7840 34184
rect 7699 34153 7711 34156
rect 7653 34147 7711 34153
rect 7834 34144 7840 34156
rect 7892 34144 7898 34196
rect 8202 34144 8208 34196
rect 8260 34144 8266 34196
rect 10229 34187 10287 34193
rect 10229 34153 10241 34187
rect 10275 34184 10287 34187
rect 10410 34184 10416 34196
rect 10275 34156 10416 34184
rect 10275 34153 10287 34156
rect 10229 34147 10287 34153
rect 10410 34144 10416 34156
rect 10468 34144 10474 34196
rect 12437 34187 12495 34193
rect 12437 34153 12449 34187
rect 12483 34184 12495 34187
rect 12526 34184 12532 34196
rect 12483 34156 12532 34184
rect 12483 34153 12495 34156
rect 12437 34147 12495 34153
rect 12526 34144 12532 34156
rect 12584 34144 12590 34196
rect 13078 34144 13084 34196
rect 13136 34184 13142 34196
rect 13722 34184 13728 34196
rect 13136 34156 13728 34184
rect 13136 34144 13142 34156
rect 13722 34144 13728 34156
rect 13780 34144 13786 34196
rect 7374 34076 7380 34128
rect 7432 34116 7438 34128
rect 7926 34116 7932 34128
rect 7432 34088 7932 34116
rect 7432 34076 7438 34088
rect 7926 34076 7932 34088
rect 7984 34116 7990 34128
rect 9217 34119 9275 34125
rect 9217 34116 9229 34119
rect 7984 34088 9229 34116
rect 7984 34076 7990 34088
rect 9217 34085 9229 34088
rect 9263 34085 9275 34119
rect 9217 34079 9275 34085
rect 10137 34119 10195 34125
rect 10137 34085 10149 34119
rect 10183 34085 10195 34119
rect 10137 34079 10195 34085
rect 11793 34119 11851 34125
rect 11793 34085 11805 34119
rect 11839 34116 11851 34119
rect 12710 34116 12716 34128
rect 11839 34088 12716 34116
rect 11839 34085 11851 34088
rect 11793 34079 11851 34085
rect 4488 34020 5120 34048
rect 4488 34008 4494 34020
rect 6086 34008 6092 34060
rect 6144 34008 6150 34060
rect 10042 34048 10048 34060
rect 6932 34020 10048 34048
rect 4338 33940 4344 33992
rect 4396 33980 4402 33992
rect 4706 33980 4712 33992
rect 4396 33952 4712 33980
rect 4396 33940 4402 33952
rect 4706 33940 4712 33952
rect 4764 33940 4770 33992
rect 6932 33989 6960 34020
rect 10042 34008 10048 34020
rect 10100 34008 10106 34060
rect 10152 34048 10180 34079
rect 12710 34076 12716 34088
rect 12768 34076 12774 34128
rect 12986 34076 12992 34128
rect 13044 34116 13050 34128
rect 13354 34116 13360 34128
rect 13044 34088 13360 34116
rect 13044 34076 13050 34088
rect 13354 34076 13360 34088
rect 13412 34076 13418 34128
rect 12345 34051 12403 34057
rect 12345 34048 12357 34051
rect 10152 34020 10824 34048
rect 6917 33983 6975 33989
rect 6917 33949 6929 33983
rect 6963 33949 6975 33983
rect 6917 33943 6975 33949
rect 7006 33940 7012 33992
rect 7064 33980 7070 33992
rect 7929 33983 7987 33989
rect 7929 33980 7941 33983
rect 7064 33952 7941 33980
rect 7064 33940 7070 33952
rect 3970 33872 3976 33924
rect 4028 33912 4034 33924
rect 4433 33915 4491 33921
rect 4433 33912 4445 33915
rect 4028 33884 4445 33912
rect 4028 33872 4034 33884
rect 4433 33881 4445 33884
rect 4479 33881 4491 33915
rect 4724 33912 4752 33940
rect 5045 33915 5103 33921
rect 5045 33912 5057 33915
rect 4724 33884 5057 33912
rect 4433 33875 4491 33881
rect 5045 33881 5057 33884
rect 5091 33881 5103 33915
rect 5045 33875 5103 33881
rect 5261 33915 5319 33921
rect 5261 33881 5273 33915
rect 5307 33912 5319 33915
rect 5442 33912 5448 33924
rect 5307 33884 5448 33912
rect 5307 33881 5319 33884
rect 5261 33875 5319 33881
rect 5442 33872 5448 33884
rect 5500 33872 5506 33924
rect 7190 33921 7196 33924
rect 7177 33915 7196 33921
rect 7177 33881 7189 33915
rect 7177 33875 7196 33881
rect 7190 33872 7196 33875
rect 7248 33872 7254 33924
rect 7374 33872 7380 33924
rect 7432 33872 7438 33924
rect 7668 33921 7696 33952
rect 7929 33949 7941 33952
rect 7975 33949 7987 33983
rect 7929 33943 7987 33949
rect 8018 33940 8024 33992
rect 8076 33980 8082 33992
rect 8205 33983 8263 33989
rect 8205 33980 8217 33983
rect 8076 33952 8217 33980
rect 8076 33940 8082 33952
rect 8205 33949 8217 33952
rect 8251 33949 8263 33983
rect 8205 33943 8263 33949
rect 9030 33940 9036 33992
rect 9088 33940 9094 33992
rect 9493 33983 9551 33989
rect 9493 33949 9505 33983
rect 9539 33980 9551 33983
rect 9858 33980 9864 33992
rect 9539 33952 9864 33980
rect 9539 33949 9551 33952
rect 9493 33943 9551 33949
rect 9858 33940 9864 33952
rect 9916 33940 9922 33992
rect 9950 33940 9956 33992
rect 10008 33940 10014 33992
rect 10137 33983 10195 33989
rect 10137 33949 10149 33983
rect 10183 33949 10195 33983
rect 10137 33943 10195 33949
rect 7637 33915 7696 33921
rect 7637 33881 7649 33915
rect 7683 33884 7696 33915
rect 7837 33915 7895 33921
rect 7683 33881 7695 33884
rect 7637 33875 7695 33881
rect 7837 33881 7849 33915
rect 7883 33881 7895 33915
rect 7837 33875 7895 33881
rect 4614 33804 4620 33856
rect 4672 33853 4678 33856
rect 4672 33847 4691 33853
rect 4679 33813 4691 33847
rect 4672 33807 4691 33813
rect 4672 33804 4678 33807
rect 4798 33804 4804 33856
rect 4856 33804 4862 33856
rect 6914 33804 6920 33856
rect 6972 33844 6978 33856
rect 7009 33847 7067 33853
rect 7009 33844 7021 33847
rect 6972 33816 7021 33844
rect 6972 33804 6978 33816
rect 7009 33813 7021 33816
rect 7055 33813 7067 33847
rect 7009 33807 7067 33813
rect 7466 33804 7472 33856
rect 7524 33804 7530 33856
rect 7852 33844 7880 33875
rect 9214 33872 9220 33924
rect 9272 33912 9278 33924
rect 9309 33915 9367 33921
rect 9309 33912 9321 33915
rect 9272 33884 9321 33912
rect 9272 33872 9278 33884
rect 9309 33881 9321 33884
rect 9355 33881 9367 33915
rect 10152 33912 10180 33943
rect 10410 33940 10416 33992
rect 10468 33940 10474 33992
rect 10796 33989 10824 34020
rect 11256 34020 12357 34048
rect 11256 33992 11284 34020
rect 12345 34017 12357 34020
rect 12391 34048 12403 34051
rect 12434 34048 12440 34060
rect 12391 34020 12440 34048
rect 12391 34017 12403 34020
rect 12345 34011 12403 34017
rect 12434 34008 12440 34020
rect 12492 34008 12498 34060
rect 12636 34020 13216 34048
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33949 10839 33983
rect 11146 33980 11152 33992
rect 11107 33952 11152 33980
rect 10781 33943 10839 33949
rect 11146 33940 11152 33952
rect 11204 33940 11210 33992
rect 11238 33940 11244 33992
rect 11296 33940 11302 33992
rect 12069 33983 12127 33989
rect 12069 33949 12081 33983
rect 12115 33980 12127 33983
rect 12250 33980 12256 33992
rect 12115 33952 12256 33980
rect 12115 33949 12127 33952
rect 12069 33943 12127 33949
rect 12250 33940 12256 33952
rect 12308 33940 12314 33992
rect 12636 33989 12664 34020
rect 13188 33992 13216 34020
rect 13906 34008 13912 34060
rect 13964 34048 13970 34060
rect 14093 34051 14151 34057
rect 14093 34048 14105 34051
rect 13964 34020 14105 34048
rect 13964 34008 13970 34020
rect 14093 34017 14105 34020
rect 14139 34017 14151 34051
rect 14093 34011 14151 34017
rect 12621 33983 12679 33989
rect 12621 33949 12633 33983
rect 12667 33949 12679 33983
rect 12621 33943 12679 33949
rect 12802 33940 12808 33992
rect 12860 33940 12866 33992
rect 13170 33940 13176 33992
rect 13228 33940 13234 33992
rect 13449 33983 13507 33989
rect 13449 33949 13461 33983
rect 13495 33980 13507 33983
rect 14349 33983 14407 33989
rect 14349 33980 14361 33983
rect 13495 33952 14361 33980
rect 13495 33949 13507 33952
rect 13449 33943 13507 33949
rect 14349 33949 14361 33952
rect 14395 33949 14407 33983
rect 14349 33943 14407 33949
rect 10505 33915 10563 33921
rect 10505 33912 10517 33915
rect 10152 33884 10517 33912
rect 9309 33875 9367 33881
rect 10505 33881 10517 33884
rect 10551 33881 10563 33915
rect 10505 33875 10563 33881
rect 10597 33915 10655 33921
rect 10597 33881 10609 33915
rect 10643 33912 10655 33915
rect 10873 33915 10931 33921
rect 10873 33912 10885 33915
rect 10643 33884 10885 33912
rect 10643 33881 10655 33884
rect 10597 33875 10655 33881
rect 10873 33881 10885 33884
rect 10919 33881 10931 33915
rect 10873 33875 10931 33881
rect 11977 33915 12035 33921
rect 11977 33881 11989 33915
rect 12023 33912 12035 33915
rect 12023 33884 12296 33912
rect 12023 33881 12035 33884
rect 11977 33875 12035 33881
rect 8021 33847 8079 33853
rect 8021 33844 8033 33847
rect 7852 33816 8033 33844
rect 8021 33813 8033 33816
rect 8067 33844 8079 33847
rect 8110 33844 8116 33856
rect 8067 33816 8116 33844
rect 8067 33813 8079 33816
rect 8021 33807 8079 33813
rect 8110 33804 8116 33816
rect 8168 33804 8174 33856
rect 10520 33844 10548 33875
rect 11992 33844 12020 33875
rect 10520 33816 12020 33844
rect 12066 33804 12072 33856
rect 12124 33844 12130 33856
rect 12161 33847 12219 33853
rect 12161 33844 12173 33847
rect 12124 33816 12173 33844
rect 12124 33804 12130 33816
rect 12161 33813 12173 33816
rect 12207 33813 12219 33847
rect 12268 33844 12296 33884
rect 12342 33872 12348 33924
rect 12400 33912 12406 33924
rect 12897 33915 12955 33921
rect 12897 33912 12909 33915
rect 12400 33884 12909 33912
rect 12400 33872 12406 33884
rect 12897 33881 12909 33884
rect 12943 33912 12955 33915
rect 13265 33915 13323 33921
rect 12943 33884 13216 33912
rect 12943 33881 12955 33884
rect 12897 33875 12955 33881
rect 13188 33856 13216 33884
rect 13265 33881 13277 33915
rect 13311 33912 13323 33915
rect 13541 33915 13599 33921
rect 13541 33912 13553 33915
rect 13311 33884 13553 33912
rect 13311 33881 13323 33884
rect 13265 33875 13323 33881
rect 13541 33881 13553 33884
rect 13587 33881 13599 33915
rect 13541 33875 13599 33881
rect 13722 33872 13728 33924
rect 13780 33872 13786 33924
rect 13909 33915 13967 33921
rect 13909 33881 13921 33915
rect 13955 33881 13967 33915
rect 13909 33875 13967 33881
rect 12986 33844 12992 33856
rect 12268 33816 12992 33844
rect 12161 33807 12219 33813
rect 12986 33804 12992 33816
rect 13044 33804 13050 33856
rect 13078 33804 13084 33856
rect 13136 33804 13142 33856
rect 13170 33804 13176 33856
rect 13228 33804 13234 33856
rect 13354 33804 13360 33856
rect 13412 33844 13418 33856
rect 13924 33844 13952 33875
rect 15473 33847 15531 33853
rect 15473 33844 15485 33847
rect 13412 33816 15485 33844
rect 13412 33804 13418 33816
rect 15473 33813 15485 33816
rect 15519 33813 15531 33847
rect 15473 33807 15531 33813
rect 1104 33754 16836 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 16836 33754
rect 1104 33680 16836 33702
rect 4522 33600 4528 33652
rect 4580 33600 4586 33652
rect 9950 33640 9956 33652
rect 6932 33612 9956 33640
rect 3602 33572 3608 33584
rect 2884 33544 3608 33572
rect 2884 33513 2912 33544
rect 3602 33532 3608 33544
rect 3660 33572 3666 33584
rect 4614 33572 4620 33584
rect 3660 33544 4620 33572
rect 3660 33532 3666 33544
rect 4614 33532 4620 33544
rect 4672 33532 4678 33584
rect 6086 33572 6092 33584
rect 4816 33544 6092 33572
rect 2869 33507 2927 33513
rect 2869 33473 2881 33507
rect 2915 33473 2927 33507
rect 2869 33467 2927 33473
rect 2958 33464 2964 33516
rect 3016 33504 3022 33516
rect 3125 33507 3183 33513
rect 3125 33504 3137 33507
rect 3016 33476 3137 33504
rect 3016 33464 3022 33476
rect 3125 33473 3137 33476
rect 3171 33473 3183 33507
rect 3125 33467 3183 33473
rect 4338 33464 4344 33516
rect 4396 33464 4402 33516
rect 4430 33464 4436 33516
rect 4488 33504 4494 33516
rect 4525 33507 4583 33513
rect 4525 33504 4537 33507
rect 4488 33476 4537 33504
rect 4488 33464 4494 33476
rect 4525 33473 4537 33476
rect 4571 33473 4583 33507
rect 4816 33504 4844 33544
rect 6086 33532 6092 33544
rect 6144 33532 6150 33584
rect 4890 33513 4896 33516
rect 4525 33467 4583 33473
rect 4632 33476 4844 33504
rect 4632 33445 4660 33476
rect 4884 33467 4896 33513
rect 4948 33504 4954 33516
rect 4948 33476 4984 33504
rect 4890 33464 4896 33467
rect 4948 33464 4954 33476
rect 6822 33464 6828 33516
rect 6880 33504 6886 33516
rect 6932 33513 6960 33612
rect 9950 33600 9956 33612
rect 10008 33640 10014 33652
rect 10778 33640 10784 33652
rect 10008 33612 10784 33640
rect 10008 33600 10014 33612
rect 10778 33600 10784 33612
rect 10836 33600 10842 33652
rect 11517 33643 11575 33649
rect 11517 33609 11529 33643
rect 11563 33640 11575 33643
rect 11606 33640 11612 33652
rect 11563 33612 11612 33640
rect 11563 33609 11575 33612
rect 11517 33603 11575 33609
rect 11606 33600 11612 33612
rect 11664 33600 11670 33652
rect 11698 33600 11704 33652
rect 11756 33600 11762 33652
rect 10134 33572 10140 33584
rect 8496 33544 10140 33572
rect 8496 33516 8524 33544
rect 10134 33532 10140 33544
rect 10192 33572 10198 33584
rect 12618 33572 12624 33584
rect 10192 33544 12624 33572
rect 10192 33532 10198 33544
rect 12618 33532 12624 33544
rect 12676 33532 12682 33584
rect 6917 33507 6975 33513
rect 6917 33504 6929 33507
rect 6880 33476 6929 33504
rect 6880 33464 6886 33476
rect 6917 33473 6929 33476
rect 6963 33473 6975 33507
rect 6917 33467 6975 33473
rect 7745 33507 7803 33513
rect 7745 33473 7757 33507
rect 7791 33504 7803 33507
rect 8294 33504 8300 33516
rect 7791 33476 8300 33504
rect 7791 33473 7803 33476
rect 7745 33467 7803 33473
rect 8294 33464 8300 33476
rect 8352 33464 8358 33516
rect 8389 33507 8447 33513
rect 8389 33473 8401 33507
rect 8435 33504 8447 33507
rect 8478 33504 8484 33516
rect 8435 33476 8484 33504
rect 8435 33473 8447 33476
rect 8389 33467 8447 33473
rect 8478 33464 8484 33476
rect 8536 33464 8542 33516
rect 8662 33513 8668 33516
rect 8656 33467 8668 33513
rect 8662 33464 8668 33467
rect 8720 33464 8726 33516
rect 9861 33507 9919 33513
rect 9861 33504 9873 33507
rect 9784 33476 9873 33504
rect 4617 33439 4675 33445
rect 4617 33405 4629 33439
rect 4663 33405 4675 33439
rect 4617 33399 4675 33405
rect 7650 33328 7656 33380
rect 7708 33328 7714 33380
rect 3878 33260 3884 33312
rect 3936 33300 3942 33312
rect 4249 33303 4307 33309
rect 4249 33300 4261 33303
rect 3936 33272 4261 33300
rect 3936 33260 3942 33272
rect 4249 33269 4261 33272
rect 4295 33269 4307 33303
rect 4249 33263 4307 33269
rect 4338 33260 4344 33312
rect 4396 33300 4402 33312
rect 4798 33300 4804 33312
rect 4396 33272 4804 33300
rect 4396 33260 4402 33272
rect 4798 33260 4804 33272
rect 4856 33260 4862 33312
rect 5902 33260 5908 33312
rect 5960 33300 5966 33312
rect 5997 33303 6055 33309
rect 5997 33300 6009 33303
rect 5960 33272 6009 33300
rect 5960 33260 5966 33272
rect 5997 33269 6009 33272
rect 6043 33269 6055 33303
rect 5997 33263 6055 33269
rect 8754 33260 8760 33312
rect 8812 33300 8818 33312
rect 9490 33300 9496 33312
rect 8812 33272 9496 33300
rect 8812 33260 8818 33272
rect 9490 33260 9496 33272
rect 9548 33300 9554 33312
rect 9784 33309 9812 33476
rect 9861 33473 9873 33476
rect 9907 33473 9919 33507
rect 9861 33467 9919 33473
rect 9950 33464 9956 33516
rect 10008 33504 10014 33516
rect 10229 33507 10287 33513
rect 10229 33504 10241 33507
rect 10008 33476 10241 33504
rect 10008 33464 10014 33476
rect 10229 33473 10241 33476
rect 10275 33473 10287 33507
rect 10229 33467 10287 33473
rect 10778 33464 10784 33516
rect 10836 33464 10842 33516
rect 11698 33507 11756 33513
rect 11698 33473 11710 33507
rect 11744 33504 11756 33507
rect 11974 33504 11980 33516
rect 11744 33476 11980 33504
rect 11744 33473 11756 33476
rect 11698 33467 11756 33473
rect 11974 33464 11980 33476
rect 12032 33464 12038 33516
rect 12069 33507 12127 33513
rect 12069 33473 12081 33507
rect 12115 33504 12127 33507
rect 12250 33504 12256 33516
rect 12115 33476 12256 33504
rect 12115 33473 12127 33476
rect 12069 33467 12127 33473
rect 12250 33464 12256 33476
rect 12308 33504 12314 33516
rect 12308 33476 12434 33504
rect 12308 33464 12314 33476
rect 10045 33439 10103 33445
rect 10045 33405 10057 33439
rect 10091 33436 10103 33439
rect 11238 33436 11244 33448
rect 10091 33408 11244 33436
rect 10091 33405 10103 33408
rect 10045 33399 10103 33405
rect 11238 33396 11244 33408
rect 11296 33396 11302 33448
rect 12158 33396 12164 33448
rect 12216 33396 12222 33448
rect 9953 33371 10011 33377
rect 9953 33337 9965 33371
rect 9999 33368 10011 33371
rect 10410 33368 10416 33380
rect 9999 33340 10416 33368
rect 9999 33337 10011 33340
rect 9953 33331 10011 33337
rect 10410 33328 10416 33340
rect 10468 33328 10474 33380
rect 12406 33368 12434 33476
rect 12802 33464 12808 33516
rect 12860 33504 12866 33516
rect 13734 33507 13792 33513
rect 13734 33504 13746 33507
rect 12860 33476 13746 33504
rect 12860 33464 12866 33476
rect 13734 33473 13746 33476
rect 13780 33473 13792 33507
rect 13734 33467 13792 33473
rect 13906 33464 13912 33516
rect 13964 33504 13970 33516
rect 14001 33507 14059 33513
rect 14001 33504 14013 33507
rect 13964 33476 14013 33504
rect 13964 33464 13970 33476
rect 14001 33473 14013 33476
rect 14047 33473 14059 33507
rect 14001 33467 14059 33473
rect 12621 33371 12679 33377
rect 12621 33368 12633 33371
rect 12406 33340 12633 33368
rect 12621 33337 12633 33340
rect 12667 33337 12679 33371
rect 12621 33331 12679 33337
rect 9769 33303 9827 33309
rect 9769 33300 9781 33303
rect 9548 33272 9781 33300
rect 9548 33260 9554 33272
rect 9769 33269 9781 33272
rect 9815 33269 9827 33303
rect 9769 33263 9827 33269
rect 10045 33303 10103 33309
rect 10045 33269 10057 33303
rect 10091 33300 10103 33303
rect 10502 33300 10508 33312
rect 10091 33272 10508 33300
rect 10091 33269 10103 33272
rect 10045 33263 10103 33269
rect 10502 33260 10508 33272
rect 10560 33260 10566 33312
rect 10594 33260 10600 33312
rect 10652 33260 10658 33312
rect 10778 33260 10784 33312
rect 10836 33300 10842 33312
rect 12710 33300 12716 33312
rect 10836 33272 12716 33300
rect 10836 33260 10842 33272
rect 12710 33260 12716 33272
rect 12768 33260 12774 33312
rect 1104 33210 16836 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 16836 33210
rect 1104 33136 16836 33158
rect 2958 33056 2964 33108
rect 3016 33056 3022 33108
rect 3145 33099 3203 33105
rect 3145 33065 3157 33099
rect 3191 33096 3203 33099
rect 3789 33099 3847 33105
rect 3789 33096 3801 33099
rect 3191 33068 3801 33096
rect 3191 33065 3203 33068
rect 3145 33059 3203 33065
rect 3789 33065 3801 33068
rect 3835 33065 3847 33099
rect 6822 33096 6828 33108
rect 3789 33059 3847 33065
rect 5736 33068 6828 33096
rect 3513 33031 3571 33037
rect 3513 32997 3525 33031
rect 3559 33028 3571 33031
rect 4062 33028 4068 33040
rect 3559 33000 4068 33028
rect 3559 32997 3571 33000
rect 3513 32991 3571 32997
rect 4062 32988 4068 33000
rect 4120 32988 4126 33040
rect 4798 32960 4804 32972
rect 4264 32932 4804 32960
rect 4264 32904 4292 32932
rect 4798 32920 4804 32932
rect 4856 32920 4862 32972
rect 3878 32852 3884 32904
rect 3936 32892 3942 32904
rect 3973 32895 4031 32901
rect 3973 32892 3985 32895
rect 3936 32864 3985 32892
rect 3936 32852 3942 32864
rect 3973 32861 3985 32864
rect 4019 32861 4031 32895
rect 3973 32855 4031 32861
rect 3988 32824 4016 32855
rect 4246 32852 4252 32904
rect 4304 32852 4310 32904
rect 4614 32852 4620 32904
rect 4672 32852 4678 32904
rect 5534 32852 5540 32904
rect 5592 32852 5598 32904
rect 5736 32901 5764 33068
rect 6822 33056 6828 33068
rect 6880 33056 6886 33108
rect 8018 33056 8024 33108
rect 8076 33056 8082 33108
rect 8662 33056 8668 33108
rect 8720 33096 8726 33108
rect 8757 33099 8815 33105
rect 8757 33096 8769 33099
rect 8720 33068 8769 33096
rect 8720 33056 8726 33068
rect 8757 33065 8769 33068
rect 8803 33065 8815 33099
rect 8757 33059 8815 33065
rect 9306 33056 9312 33108
rect 9364 33096 9370 33108
rect 9858 33096 9864 33108
rect 9364 33068 9864 33096
rect 9364 33056 9370 33068
rect 9858 33056 9864 33068
rect 9916 33056 9922 33108
rect 12802 33056 12808 33108
rect 12860 33056 12866 33108
rect 12989 33099 13047 33105
rect 12989 33065 13001 33099
rect 13035 33096 13047 33099
rect 13078 33096 13084 33108
rect 13035 33068 13084 33096
rect 13035 33065 13047 33068
rect 12989 33059 13047 33065
rect 8294 32988 8300 33040
rect 8352 33028 8358 33040
rect 9398 33028 9404 33040
rect 8352 33000 9404 33028
rect 8352 32988 8358 33000
rect 9398 32988 9404 33000
rect 9456 33028 9462 33040
rect 9769 33031 9827 33037
rect 9769 33028 9781 33031
rect 9456 33000 9781 33028
rect 9456 32988 9462 33000
rect 9769 32997 9781 33000
rect 9815 33028 9827 33031
rect 9815 33000 11192 33028
rect 9815 32997 9827 33000
rect 9769 32991 9827 32997
rect 11164 32972 11192 33000
rect 8128 32932 9168 32960
rect 5721 32895 5779 32901
rect 5721 32861 5733 32895
rect 5767 32861 5779 32895
rect 5721 32855 5779 32861
rect 5997 32895 6055 32901
rect 5997 32861 6009 32895
rect 6043 32892 6055 32895
rect 6086 32892 6092 32904
rect 6043 32864 6092 32892
rect 6043 32861 6055 32864
rect 5997 32855 6055 32861
rect 6086 32852 6092 32864
rect 6144 32892 6150 32904
rect 6454 32892 6460 32904
rect 6144 32864 6460 32892
rect 6144 32852 6150 32864
rect 6454 32852 6460 32864
rect 6512 32892 6518 32904
rect 6914 32901 6920 32904
rect 6641 32895 6699 32901
rect 6641 32892 6653 32895
rect 6512 32864 6653 32892
rect 6512 32852 6518 32864
rect 6641 32861 6653 32864
rect 6687 32861 6699 32895
rect 6908 32892 6920 32901
rect 6875 32864 6920 32892
rect 6641 32855 6699 32861
rect 6908 32855 6920 32864
rect 6914 32852 6920 32855
rect 6972 32852 6978 32904
rect 7374 32852 7380 32904
rect 7432 32892 7438 32904
rect 8128 32901 8156 32932
rect 8113 32895 8171 32901
rect 8113 32892 8125 32895
rect 7432 32864 8125 32892
rect 7432 32852 7438 32864
rect 8113 32861 8125 32864
rect 8159 32861 8171 32895
rect 8113 32855 8171 32861
rect 8294 32852 8300 32904
rect 8352 32852 8358 32904
rect 8389 32895 8447 32901
rect 8389 32861 8401 32895
rect 8435 32861 8447 32895
rect 8389 32855 8447 32861
rect 8481 32895 8539 32901
rect 8481 32861 8493 32895
rect 8527 32892 8539 32895
rect 8754 32892 8760 32904
rect 8527 32864 8760 32892
rect 8527 32861 8539 32864
rect 8481 32855 8539 32861
rect 4338 32824 4344 32836
rect 3988 32796 4344 32824
rect 4338 32784 4344 32796
rect 4396 32784 4402 32836
rect 5905 32827 5963 32833
rect 5905 32793 5917 32827
rect 5951 32824 5963 32827
rect 7006 32824 7012 32836
rect 5951 32796 7012 32824
rect 5951 32793 5963 32796
rect 5905 32787 5963 32793
rect 7006 32784 7012 32796
rect 7064 32784 7070 32836
rect 7466 32784 7472 32836
rect 7524 32824 7530 32836
rect 8404 32824 8432 32855
rect 8754 32852 8760 32864
rect 8812 32852 8818 32904
rect 8941 32895 8999 32901
rect 8941 32861 8953 32895
rect 8987 32892 8999 32895
rect 9030 32892 9036 32904
rect 8987 32864 9036 32892
rect 8987 32861 8999 32864
rect 8941 32855 8999 32861
rect 7524 32796 8432 32824
rect 7524 32784 7530 32796
rect 8570 32784 8576 32836
rect 8628 32824 8634 32836
rect 8956 32824 8984 32855
rect 9030 32852 9036 32864
rect 9088 32852 9094 32904
rect 9140 32901 9168 32932
rect 9950 32920 9956 32972
rect 10008 32920 10014 32972
rect 10134 32920 10140 32972
rect 10192 32960 10198 32972
rect 10781 32963 10839 32969
rect 10781 32960 10793 32963
rect 10192 32932 10793 32960
rect 10192 32920 10198 32932
rect 10781 32929 10793 32932
rect 10827 32960 10839 32963
rect 10870 32960 10876 32972
rect 10827 32932 10876 32960
rect 10827 32929 10839 32932
rect 10781 32923 10839 32929
rect 10870 32920 10876 32932
rect 10928 32920 10934 32972
rect 11146 32920 11152 32972
rect 11204 32920 11210 32972
rect 11609 32963 11667 32969
rect 11609 32929 11621 32963
rect 11655 32960 11667 32963
rect 12158 32960 12164 32972
rect 11655 32932 12164 32960
rect 11655 32929 11667 32932
rect 11609 32923 11667 32929
rect 12158 32920 12164 32932
rect 12216 32920 12222 32972
rect 13004 32960 13032 33059
rect 13078 33056 13084 33068
rect 13136 33056 13142 33108
rect 12406 32932 13032 32960
rect 9125 32895 9183 32901
rect 9125 32861 9137 32895
rect 9171 32861 9183 32895
rect 9125 32855 9183 32861
rect 9217 32895 9275 32901
rect 9217 32861 9229 32895
rect 9263 32861 9275 32895
rect 9217 32855 9275 32861
rect 9232 32824 9260 32855
rect 10042 32852 10048 32904
rect 10100 32852 10106 32904
rect 10594 32892 10600 32904
rect 10244 32864 10600 32892
rect 10244 32836 10272 32864
rect 10594 32852 10600 32864
rect 10652 32892 10658 32904
rect 11241 32895 11299 32901
rect 11241 32892 11253 32895
rect 10652 32864 11253 32892
rect 10652 32852 10658 32864
rect 11241 32861 11253 32864
rect 11287 32861 11299 32895
rect 11241 32855 11299 32861
rect 9493 32827 9551 32833
rect 9493 32824 9505 32827
rect 8628 32796 8984 32824
rect 9048 32796 9505 32824
rect 8628 32784 8634 32796
rect 3145 32759 3203 32765
rect 3145 32725 3157 32759
rect 3191 32756 3203 32759
rect 3510 32756 3516 32768
rect 3191 32728 3516 32756
rect 3191 32725 3203 32728
rect 3145 32719 3203 32725
rect 3510 32716 3516 32728
rect 3568 32756 3574 32768
rect 3970 32756 3976 32768
rect 3568 32728 3976 32756
rect 3568 32716 3574 32728
rect 3970 32716 3976 32728
rect 4028 32716 4034 32768
rect 4062 32716 4068 32768
rect 4120 32756 4126 32768
rect 4157 32759 4215 32765
rect 4157 32756 4169 32759
rect 4120 32728 4169 32756
rect 4120 32716 4126 32728
rect 4157 32725 4169 32728
rect 4203 32756 4215 32759
rect 5810 32756 5816 32768
rect 4203 32728 5816 32756
rect 4203 32725 4215 32728
rect 4157 32719 4215 32725
rect 5810 32716 5816 32728
rect 5868 32716 5874 32768
rect 6270 32716 6276 32768
rect 6328 32756 6334 32768
rect 9048 32756 9076 32796
rect 9493 32793 9505 32796
rect 9539 32824 9551 32827
rect 10226 32824 10232 32836
rect 9539 32796 10232 32824
rect 9539 32793 9551 32796
rect 9493 32787 9551 32793
rect 10226 32784 10232 32796
rect 10284 32784 10290 32836
rect 6328 32728 9076 32756
rect 6328 32716 6334 32728
rect 9122 32716 9128 32768
rect 9180 32716 9186 32768
rect 9214 32716 9220 32768
rect 9272 32756 9278 32768
rect 12406 32756 12434 32932
rect 12621 32895 12679 32901
rect 12621 32861 12633 32895
rect 12667 32892 12679 32895
rect 13906 32892 13912 32904
rect 12667 32864 13912 32892
rect 12667 32861 12679 32864
rect 12621 32855 12679 32861
rect 13906 32852 13912 32864
rect 13964 32852 13970 32904
rect 12894 32784 12900 32836
rect 12952 32833 12958 32836
rect 12952 32827 13015 32833
rect 12952 32793 12969 32827
rect 13003 32793 13015 32827
rect 12952 32787 13015 32793
rect 12952 32784 12958 32787
rect 13170 32784 13176 32836
rect 13228 32784 13234 32836
rect 9272 32728 12434 32756
rect 9272 32716 9278 32728
rect 1104 32666 16836 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 16836 32666
rect 1104 32592 16836 32614
rect 3881 32555 3939 32561
rect 3881 32521 3893 32555
rect 3927 32552 3939 32555
rect 4246 32552 4252 32564
rect 3927 32524 4252 32552
rect 3927 32521 3939 32524
rect 3881 32515 3939 32521
rect 4246 32512 4252 32524
rect 4304 32512 4310 32564
rect 5166 32512 5172 32564
rect 5224 32552 5230 32564
rect 7650 32552 7656 32564
rect 5224 32524 7656 32552
rect 5224 32512 5230 32524
rect 7650 32512 7656 32524
rect 7708 32552 7714 32564
rect 10502 32552 10508 32564
rect 7708 32524 10508 32552
rect 7708 32512 7714 32524
rect 10502 32512 10508 32524
rect 10560 32512 10566 32564
rect 11333 32555 11391 32561
rect 11333 32521 11345 32555
rect 11379 32552 11391 32555
rect 11698 32552 11704 32564
rect 11379 32524 11704 32552
rect 11379 32521 11391 32524
rect 11333 32515 11391 32521
rect 11698 32512 11704 32524
rect 11756 32512 11762 32564
rect 3237 32487 3295 32493
rect 3237 32453 3249 32487
rect 3283 32484 3295 32487
rect 4154 32484 4160 32496
rect 3283 32456 4160 32484
rect 3283 32453 3295 32456
rect 3237 32447 3295 32453
rect 4154 32444 4160 32456
rect 4212 32444 4218 32496
rect 5721 32487 5779 32493
rect 5721 32453 5733 32487
rect 5767 32484 5779 32487
rect 6270 32484 6276 32496
rect 5767 32456 6276 32484
rect 5767 32453 5779 32456
rect 5721 32447 5779 32453
rect 6270 32444 6276 32456
rect 6328 32444 6334 32496
rect 10042 32444 10048 32496
rect 10100 32484 10106 32496
rect 11882 32484 11888 32496
rect 10100 32456 11888 32484
rect 10100 32444 10106 32456
rect 11882 32444 11888 32456
rect 11940 32484 11946 32496
rect 12161 32487 12219 32493
rect 12161 32484 12173 32487
rect 11940 32456 12173 32484
rect 11940 32444 11946 32456
rect 12161 32453 12173 32456
rect 12207 32453 12219 32487
rect 12161 32447 12219 32453
rect 12989 32487 13047 32493
rect 12989 32453 13001 32487
rect 13035 32484 13047 32487
rect 13906 32484 13912 32496
rect 13035 32456 13912 32484
rect 13035 32453 13047 32456
rect 12989 32447 13047 32453
rect 13906 32444 13912 32456
rect 13964 32444 13970 32496
rect 3421 32419 3479 32425
rect 3421 32385 3433 32419
rect 3467 32385 3479 32419
rect 3421 32379 3479 32385
rect 3436 32348 3464 32379
rect 3970 32376 3976 32428
rect 4028 32376 4034 32428
rect 4065 32419 4123 32425
rect 4065 32385 4077 32419
rect 4111 32416 4123 32419
rect 4338 32416 4344 32428
rect 4111 32388 4344 32416
rect 4111 32385 4123 32388
rect 4065 32379 4123 32385
rect 4338 32376 4344 32388
rect 4396 32416 4402 32428
rect 4396 32388 4844 32416
rect 4396 32376 4402 32388
rect 4525 32351 4583 32357
rect 3436 32320 4292 32348
rect 4264 32289 4292 32320
rect 4525 32317 4537 32351
rect 4571 32348 4583 32351
rect 4614 32348 4620 32360
rect 4571 32320 4620 32348
rect 4571 32317 4583 32320
rect 4525 32311 4583 32317
rect 4614 32308 4620 32320
rect 4672 32308 4678 32360
rect 4816 32348 4844 32388
rect 5258 32376 5264 32428
rect 5316 32376 5322 32428
rect 5537 32419 5595 32425
rect 5537 32385 5549 32419
rect 5583 32385 5595 32419
rect 5537 32379 5595 32385
rect 5813 32419 5871 32425
rect 5813 32385 5825 32419
rect 5859 32416 5871 32419
rect 5902 32416 5908 32428
rect 5859 32388 5908 32416
rect 5859 32385 5871 32388
rect 5813 32379 5871 32385
rect 5442 32348 5448 32360
rect 4816 32320 5448 32348
rect 5442 32308 5448 32320
rect 5500 32348 5506 32360
rect 5552 32348 5580 32379
rect 5902 32376 5908 32388
rect 5960 32376 5966 32428
rect 10134 32376 10140 32428
rect 10192 32376 10198 32428
rect 10226 32376 10232 32428
rect 10284 32416 10290 32428
rect 11146 32425 11152 32428
rect 10965 32419 11023 32425
rect 10965 32416 10977 32419
rect 10284 32388 10977 32416
rect 10284 32376 10290 32388
rect 10965 32385 10977 32388
rect 11011 32385 11023 32419
rect 10965 32379 11023 32385
rect 11119 32419 11152 32425
rect 11119 32385 11131 32419
rect 11119 32379 11152 32385
rect 11146 32376 11152 32379
rect 11204 32376 11210 32428
rect 11238 32376 11244 32428
rect 11296 32416 11302 32428
rect 11609 32419 11667 32425
rect 11609 32416 11621 32419
rect 11296 32388 11621 32416
rect 11296 32376 11302 32388
rect 11609 32385 11621 32388
rect 11655 32385 11667 32419
rect 11609 32379 11667 32385
rect 5994 32348 6000 32360
rect 5500 32320 6000 32348
rect 5500 32308 5506 32320
rect 5994 32308 6000 32320
rect 6052 32308 6058 32360
rect 4249 32283 4307 32289
rect 4249 32249 4261 32283
rect 4295 32280 4307 32283
rect 4798 32280 4804 32292
rect 4295 32252 4804 32280
rect 4295 32249 4307 32252
rect 4249 32243 4307 32249
rect 4798 32240 4804 32252
rect 4856 32240 4862 32292
rect 3602 32172 3608 32224
rect 3660 32172 3666 32224
rect 3694 32172 3700 32224
rect 3752 32172 3758 32224
rect 4982 32172 4988 32224
rect 5040 32212 5046 32224
rect 5353 32215 5411 32221
rect 5353 32212 5365 32215
rect 5040 32184 5365 32212
rect 5040 32172 5046 32184
rect 5353 32181 5365 32184
rect 5399 32181 5411 32215
rect 11164 32212 11192 32376
rect 11422 32212 11428 32224
rect 11164 32184 11428 32212
rect 5353 32175 5411 32181
rect 11422 32172 11428 32184
rect 11480 32212 11486 32224
rect 11701 32215 11759 32221
rect 11701 32212 11713 32215
rect 11480 32184 11713 32212
rect 11480 32172 11486 32184
rect 11701 32181 11713 32184
rect 11747 32181 11759 32215
rect 11701 32175 11759 32181
rect 1104 32122 16836 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 16836 32122
rect 1104 32048 16836 32070
rect 3602 31968 3608 32020
rect 3660 32008 3666 32020
rect 4157 32011 4215 32017
rect 4157 32008 4169 32011
rect 3660 31980 4169 32008
rect 3660 31968 3666 31980
rect 4157 31977 4169 31980
rect 4203 31977 4215 32011
rect 4157 31971 4215 31977
rect 4706 31968 4712 32020
rect 4764 32008 4770 32020
rect 4801 32011 4859 32017
rect 4801 32008 4813 32011
rect 4764 31980 4813 32008
rect 4764 31968 4770 31980
rect 4801 31977 4813 31980
rect 4847 31977 4859 32011
rect 5902 32008 5908 32020
rect 4801 31971 4859 31977
rect 4908 31980 5908 32008
rect 3694 31900 3700 31952
rect 3752 31940 3758 31952
rect 3789 31943 3847 31949
rect 3789 31940 3801 31943
rect 3752 31912 3801 31940
rect 3752 31900 3758 31912
rect 3789 31909 3801 31912
rect 3835 31909 3847 31943
rect 3789 31903 3847 31909
rect 4908 31872 4936 31980
rect 5902 31968 5908 31980
rect 5960 31968 5966 32020
rect 7006 31968 7012 32020
rect 7064 32008 7070 32020
rect 7064 31980 9720 32008
rect 7064 31968 7070 31980
rect 5166 31900 5172 31952
rect 5224 31940 5230 31952
rect 5224 31912 5304 31940
rect 5224 31900 5230 31912
rect 4356 31844 4936 31872
rect 2958 31764 2964 31816
rect 3016 31804 3022 31816
rect 3016 31776 3924 31804
rect 3016 31764 3022 31776
rect 3896 31736 3924 31776
rect 4157 31739 4215 31745
rect 4157 31736 4169 31739
rect 3896 31708 4169 31736
rect 4157 31705 4169 31708
rect 4203 31705 4215 31739
rect 4356 31736 4384 31844
rect 4433 31807 4491 31813
rect 4433 31773 4445 31807
rect 4479 31804 4491 31807
rect 4890 31804 4896 31816
rect 4479 31776 4896 31804
rect 4479 31773 4491 31776
rect 4433 31767 4491 31773
rect 4890 31764 4896 31776
rect 4948 31764 4954 31816
rect 4982 31764 4988 31816
rect 5040 31764 5046 31816
rect 5276 31813 5304 31912
rect 5442 31900 5448 31952
rect 5500 31940 5506 31952
rect 5721 31943 5779 31949
rect 5721 31940 5733 31943
rect 5500 31912 5733 31940
rect 5500 31900 5506 31912
rect 5721 31909 5733 31912
rect 5767 31909 5779 31943
rect 5721 31903 5779 31909
rect 6178 31900 6184 31952
rect 6236 31940 6242 31952
rect 6236 31912 8616 31940
rect 6236 31900 6242 31912
rect 5350 31832 5356 31884
rect 5408 31832 5414 31884
rect 5813 31875 5871 31881
rect 5813 31872 5825 31875
rect 5552 31844 5825 31872
rect 5552 31813 5580 31844
rect 5813 31841 5825 31844
rect 5859 31841 5871 31875
rect 5813 31835 5871 31841
rect 5902 31832 5908 31884
rect 5960 31872 5966 31884
rect 5960 31844 6224 31872
rect 5960 31832 5966 31844
rect 5169 31807 5227 31813
rect 5169 31804 5181 31807
rect 5147 31776 5181 31804
rect 5169 31773 5181 31776
rect 5215 31773 5227 31807
rect 5169 31767 5227 31773
rect 5261 31807 5319 31813
rect 5261 31773 5273 31807
rect 5307 31804 5319 31807
rect 5537 31807 5595 31813
rect 5307 31776 5341 31804
rect 5307 31773 5319 31776
rect 5261 31767 5319 31773
rect 5537 31773 5549 31807
rect 5583 31773 5595 31807
rect 5537 31767 5595 31773
rect 4617 31739 4675 31745
rect 4617 31736 4629 31739
rect 4356 31708 4629 31736
rect 4157 31699 4215 31705
rect 4617 31705 4629 31708
rect 4663 31705 4675 31739
rect 4617 31699 4675 31705
rect 4798 31696 4804 31748
rect 4856 31736 4862 31748
rect 5184 31736 5212 31767
rect 4856 31708 5212 31736
rect 5276 31736 5304 31767
rect 5994 31764 6000 31816
rect 6052 31764 6058 31816
rect 6196 31813 6224 31844
rect 7006 31832 7012 31884
rect 7064 31832 7070 31884
rect 8588 31881 8616 31912
rect 8573 31875 8631 31881
rect 8573 31841 8585 31875
rect 8619 31841 8631 31875
rect 8573 31835 8631 31841
rect 6181 31807 6239 31813
rect 6181 31773 6193 31807
rect 6227 31773 6239 31807
rect 6181 31767 6239 31773
rect 6270 31764 6276 31816
rect 6328 31764 6334 31816
rect 6914 31764 6920 31816
rect 6972 31764 6978 31816
rect 8389 31807 8447 31813
rect 8389 31804 8401 31807
rect 7024 31776 8401 31804
rect 5350 31736 5356 31748
rect 5276 31708 5356 31736
rect 4856 31696 4862 31708
rect 5350 31696 5356 31708
rect 5408 31696 5414 31748
rect 6822 31696 6828 31748
rect 6880 31736 6886 31748
rect 7024 31736 7052 31776
rect 8389 31773 8401 31776
rect 8435 31773 8447 31807
rect 8389 31767 8447 31773
rect 8478 31764 8484 31816
rect 8536 31764 8542 31816
rect 8665 31807 8723 31813
rect 8665 31773 8677 31807
rect 8711 31804 8723 31807
rect 9306 31804 9312 31816
rect 8711 31776 9312 31804
rect 8711 31773 8723 31776
rect 8665 31767 8723 31773
rect 9306 31764 9312 31776
rect 9364 31804 9370 31816
rect 9692 31813 9720 31980
rect 10612 31912 12204 31940
rect 10321 31875 10379 31881
rect 10321 31841 10333 31875
rect 10367 31872 10379 31875
rect 10367 31844 10548 31872
rect 10367 31841 10379 31844
rect 10321 31835 10379 31841
rect 9401 31807 9459 31813
rect 9401 31804 9413 31807
rect 9364 31776 9413 31804
rect 9364 31764 9370 31776
rect 9401 31773 9413 31776
rect 9447 31773 9459 31807
rect 9401 31767 9459 31773
rect 9677 31807 9735 31813
rect 9677 31773 9689 31807
rect 9723 31773 9735 31807
rect 9677 31767 9735 31773
rect 10226 31764 10232 31816
rect 10284 31764 10290 31816
rect 10520 31813 10548 31844
rect 10413 31807 10471 31813
rect 10413 31804 10425 31807
rect 10391 31776 10425 31804
rect 10413 31773 10425 31776
rect 10459 31773 10471 31807
rect 10520 31807 10583 31813
rect 10520 31776 10537 31807
rect 10413 31767 10471 31773
rect 10525 31773 10537 31776
rect 10571 31773 10583 31807
rect 10525 31767 10583 31773
rect 6880 31708 7052 31736
rect 8021 31739 8079 31745
rect 6880 31696 6886 31708
rect 8021 31705 8033 31739
rect 8067 31736 8079 31739
rect 9585 31739 9643 31745
rect 8067 31708 9444 31736
rect 8067 31705 8079 31708
rect 8021 31699 8079 31705
rect 9416 31680 9444 31708
rect 9585 31705 9597 31739
rect 9631 31705 9643 31739
rect 10428 31736 10456 31767
rect 10612 31736 10640 31912
rect 11149 31875 11207 31881
rect 11149 31872 11161 31875
rect 10704 31844 11161 31872
rect 10704 31813 10732 31844
rect 11149 31841 11161 31844
rect 11195 31841 11207 31875
rect 11149 31835 11207 31841
rect 12069 31875 12127 31881
rect 12069 31841 12081 31875
rect 12115 31841 12127 31875
rect 12069 31835 12127 31841
rect 10689 31807 10747 31813
rect 10689 31773 10701 31807
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 10781 31807 10839 31813
rect 10781 31773 10793 31807
rect 10827 31773 10839 31807
rect 10897 31807 10955 31813
rect 10897 31804 10909 31807
rect 10781 31767 10839 31773
rect 10888 31773 10909 31804
rect 10943 31773 10955 31807
rect 11422 31804 11428 31816
rect 11383 31776 11428 31804
rect 10888 31767 10955 31773
rect 10796 31736 10824 31767
rect 10428 31708 10824 31736
rect 9585 31699 9643 31705
rect 4338 31628 4344 31680
rect 4396 31628 4402 31680
rect 6546 31628 6552 31680
rect 6604 31628 6610 31680
rect 7926 31628 7932 31680
rect 7984 31628 7990 31680
rect 8110 31628 8116 31680
rect 8168 31668 8174 31680
rect 8205 31671 8263 31677
rect 8205 31668 8217 31671
rect 8168 31640 8217 31668
rect 8168 31628 8174 31640
rect 8205 31637 8217 31640
rect 8251 31637 8263 31671
rect 8205 31631 8263 31637
rect 9122 31628 9128 31680
rect 9180 31668 9186 31680
rect 9217 31671 9275 31677
rect 9217 31668 9229 31671
rect 9180 31640 9229 31668
rect 9180 31628 9186 31640
rect 9217 31637 9229 31640
rect 9263 31637 9275 31671
rect 9217 31631 9275 31637
rect 9398 31628 9404 31680
rect 9456 31628 9462 31680
rect 9490 31628 9496 31680
rect 9548 31668 9554 31680
rect 9600 31668 9628 31699
rect 9861 31671 9919 31677
rect 9861 31668 9873 31671
rect 9548 31640 9873 31668
rect 9548 31628 9554 31640
rect 9861 31637 9873 31640
rect 9907 31668 9919 31671
rect 10888 31668 10916 31767
rect 11422 31764 11428 31776
rect 11480 31764 11486 31816
rect 11514 31764 11520 31816
rect 11572 31804 11578 31816
rect 12084 31804 12112 31835
rect 12176 31813 12204 31912
rect 12529 31875 12587 31881
rect 12529 31841 12541 31875
rect 12575 31872 12587 31875
rect 13106 31875 13164 31881
rect 13106 31872 13118 31875
rect 12575 31844 13118 31872
rect 12575 31841 12587 31844
rect 12529 31835 12587 31841
rect 13106 31841 13118 31844
rect 13152 31841 13164 31875
rect 13106 31835 13164 31841
rect 11572 31776 12112 31804
rect 12161 31807 12219 31813
rect 11572 31764 11578 31776
rect 12161 31773 12173 31807
rect 12207 31804 12219 31807
rect 12434 31804 12440 31816
rect 12207 31776 12440 31804
rect 12207 31773 12219 31776
rect 12161 31767 12219 31773
rect 12434 31764 12440 31776
rect 12492 31764 12498 31816
rect 12618 31764 12624 31816
rect 12676 31764 12682 31816
rect 12894 31764 12900 31816
rect 12952 31764 12958 31816
rect 12986 31764 12992 31816
rect 13044 31764 13050 31816
rect 9907 31640 10916 31668
rect 9907 31637 9919 31640
rect 9861 31631 9919 31637
rect 11054 31628 11060 31680
rect 11112 31628 11118 31680
rect 13265 31671 13323 31677
rect 13265 31637 13277 31671
rect 13311 31668 13323 31671
rect 13354 31668 13360 31680
rect 13311 31640 13360 31668
rect 13311 31637 13323 31640
rect 13265 31631 13323 31637
rect 13354 31628 13360 31640
rect 13412 31628 13418 31680
rect 1104 31578 16836 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 16836 31578
rect 1104 31504 16836 31526
rect 3329 31467 3387 31473
rect 3329 31433 3341 31467
rect 3375 31433 3387 31467
rect 3329 31427 3387 31433
rect 3344 31328 3372 31427
rect 4706 31424 4712 31476
rect 4764 31424 4770 31476
rect 4798 31424 4804 31476
rect 4856 31464 4862 31476
rect 4985 31467 5043 31473
rect 4985 31464 4997 31467
rect 4856 31436 4997 31464
rect 4856 31424 4862 31436
rect 4985 31433 4997 31436
rect 5031 31433 5043 31467
rect 4985 31427 5043 31433
rect 6181 31467 6239 31473
rect 6181 31433 6193 31467
rect 6227 31464 6239 31467
rect 7006 31464 7012 31476
rect 6227 31436 7012 31464
rect 6227 31433 6239 31436
rect 6181 31427 6239 31433
rect 7006 31424 7012 31436
rect 7064 31424 7070 31476
rect 7837 31467 7895 31473
rect 7837 31464 7849 31467
rect 7795 31436 7849 31464
rect 7837 31433 7849 31436
rect 7883 31464 7895 31467
rect 8478 31464 8484 31476
rect 7883 31436 8484 31464
rect 7883 31433 7895 31436
rect 7837 31427 7895 31433
rect 4338 31356 4344 31408
rect 4396 31396 4402 31408
rect 4442 31399 4500 31405
rect 4442 31396 4454 31399
rect 4396 31368 4454 31396
rect 4396 31356 4402 31368
rect 4442 31365 4454 31368
rect 4488 31365 4500 31399
rect 4442 31359 4500 31365
rect 4724 31328 4752 31424
rect 6822 31396 6828 31408
rect 6012 31368 6828 31396
rect 5166 31328 5172 31340
rect 3344 31300 5172 31328
rect 5166 31288 5172 31300
rect 5224 31288 5230 31340
rect 6012 31337 6040 31368
rect 6822 31356 6828 31368
rect 6880 31356 6886 31408
rect 6914 31356 6920 31408
rect 6972 31396 6978 31408
rect 7852 31396 7880 31427
rect 8478 31424 8484 31436
rect 8536 31424 8542 31476
rect 9306 31424 9312 31476
rect 9364 31424 9370 31476
rect 10870 31396 10876 31408
rect 6972 31368 7880 31396
rect 7944 31368 10876 31396
rect 6972 31356 6978 31368
rect 5997 31331 6055 31337
rect 5997 31297 6009 31331
rect 6043 31297 6055 31331
rect 5997 31291 6055 31297
rect 6178 31288 6184 31340
rect 6236 31328 6242 31340
rect 6362 31328 6368 31340
rect 6236 31300 6368 31328
rect 6236 31288 6242 31300
rect 6362 31288 6368 31300
rect 6420 31288 6426 31340
rect 6454 31288 6460 31340
rect 6512 31288 6518 31340
rect 6730 31337 6736 31340
rect 6724 31291 6736 31337
rect 6730 31288 6736 31291
rect 6788 31288 6794 31340
rect 7944 31337 7972 31368
rect 10870 31356 10876 31368
rect 10928 31356 10934 31408
rect 13170 31396 13176 31408
rect 12406 31368 13176 31396
rect 8202 31337 8208 31340
rect 7929 31331 7987 31337
rect 7929 31297 7941 31331
rect 7975 31297 7987 31331
rect 7929 31291 7987 31297
rect 8196 31291 8208 31337
rect 8202 31288 8208 31291
rect 8260 31288 8266 31340
rect 9122 31288 9128 31340
rect 9180 31328 9186 31340
rect 9861 31331 9919 31337
rect 9861 31328 9873 31331
rect 9180 31300 9873 31328
rect 9180 31288 9186 31300
rect 9861 31297 9873 31300
rect 9907 31297 9919 31331
rect 9861 31291 9919 31297
rect 9950 31288 9956 31340
rect 10008 31328 10014 31340
rect 10045 31331 10103 31337
rect 10045 31328 10057 31331
rect 10008 31300 10057 31328
rect 10008 31288 10014 31300
rect 10045 31297 10057 31300
rect 10091 31297 10103 31331
rect 10045 31291 10103 31297
rect 10137 31331 10195 31337
rect 10137 31297 10149 31331
rect 10183 31328 10195 31331
rect 11514 31328 11520 31340
rect 10183 31300 11520 31328
rect 10183 31297 10195 31300
rect 10137 31291 10195 31297
rect 11514 31288 11520 31300
rect 11572 31328 11578 31340
rect 12406 31328 12434 31368
rect 13170 31356 13176 31368
rect 13228 31356 13234 31408
rect 13354 31405 13360 31408
rect 13348 31359 13360 31405
rect 13354 31356 13360 31359
rect 13412 31356 13418 31408
rect 13538 31356 13544 31408
rect 13596 31356 13602 31408
rect 13556 31328 13584 31356
rect 11572 31300 12434 31328
rect 13004 31300 13584 31328
rect 11572 31288 11578 31300
rect 13004 31272 13032 31300
rect 4706 31220 4712 31272
rect 4764 31220 4770 31272
rect 5445 31263 5503 31269
rect 5445 31229 5457 31263
rect 5491 31260 5503 31263
rect 5626 31260 5632 31272
rect 5491 31232 5632 31260
rect 5491 31229 5503 31232
rect 5445 31223 5503 31229
rect 5626 31220 5632 31232
rect 5684 31220 5690 31272
rect 9398 31220 9404 31272
rect 9456 31260 9462 31272
rect 12986 31260 12992 31272
rect 9456 31232 12992 31260
rect 9456 31220 9462 31232
rect 12986 31220 12992 31232
rect 13044 31220 13050 31272
rect 13081 31263 13139 31269
rect 13081 31229 13093 31263
rect 13127 31260 13139 31263
rect 13127 31229 13149 31260
rect 13081 31223 13149 31229
rect 8938 31152 8944 31204
rect 8996 31192 9002 31204
rect 12618 31192 12624 31204
rect 8996 31164 12624 31192
rect 8996 31152 9002 31164
rect 12618 31152 12624 31164
rect 12676 31192 12682 31204
rect 12802 31192 12808 31204
rect 12676 31164 12808 31192
rect 12676 31152 12682 31164
rect 12802 31152 12808 31164
rect 12860 31152 12866 31204
rect 5353 31127 5411 31133
rect 5353 31093 5365 31127
rect 5399 31124 5411 31127
rect 5534 31124 5540 31136
rect 5399 31096 5540 31124
rect 5399 31093 5411 31096
rect 5353 31087 5411 31093
rect 5534 31084 5540 31096
rect 5592 31084 5598 31136
rect 9677 31127 9735 31133
rect 9677 31093 9689 31127
rect 9723 31124 9735 31127
rect 10686 31124 10692 31136
rect 9723 31096 10692 31124
rect 9723 31093 9735 31096
rect 9677 31087 9735 31093
rect 10686 31084 10692 31096
rect 10744 31084 10750 31136
rect 10778 31084 10784 31136
rect 10836 31124 10842 31136
rect 12986 31124 12992 31136
rect 10836 31096 12992 31124
rect 10836 31084 10842 31096
rect 12986 31084 12992 31096
rect 13044 31084 13050 31136
rect 13121 31124 13149 31223
rect 14090 31124 14096 31136
rect 13121 31096 14096 31124
rect 14090 31084 14096 31096
rect 14148 31084 14154 31136
rect 14458 31084 14464 31136
rect 14516 31084 14522 31136
rect 1104 31034 16836 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 16836 31034
rect 1104 30960 16836 30982
rect 6549 30923 6607 30929
rect 6549 30889 6561 30923
rect 6595 30920 6607 30923
rect 6730 30920 6736 30932
rect 6595 30892 6736 30920
rect 6595 30889 6607 30892
rect 6549 30883 6607 30889
rect 6730 30880 6736 30892
rect 6788 30880 6794 30932
rect 8202 30880 8208 30932
rect 8260 30880 8266 30932
rect 9309 30923 9367 30929
rect 9309 30889 9321 30923
rect 9355 30920 9367 30923
rect 9398 30920 9404 30932
rect 9355 30892 9404 30920
rect 9355 30889 9367 30892
rect 9309 30883 9367 30889
rect 9398 30880 9404 30892
rect 9456 30880 9462 30932
rect 10597 30923 10655 30929
rect 10597 30889 10609 30923
rect 10643 30920 10655 30923
rect 11054 30920 11060 30932
rect 10643 30892 11060 30920
rect 10643 30889 10655 30892
rect 10597 30883 10655 30889
rect 11054 30880 11060 30892
rect 11112 30880 11118 30932
rect 12802 30880 12808 30932
rect 12860 30920 12866 30932
rect 13262 30920 13268 30932
rect 12860 30892 13268 30920
rect 12860 30880 12866 30892
rect 13262 30880 13268 30892
rect 13320 30880 13326 30932
rect 8938 30852 8944 30864
rect 7576 30824 8944 30852
rect 3694 30744 3700 30796
rect 3752 30784 3758 30796
rect 3752 30756 4016 30784
rect 3752 30744 3758 30756
rect 3789 30719 3847 30725
rect 3789 30685 3801 30719
rect 3835 30716 3847 30719
rect 3878 30716 3884 30728
rect 3835 30688 3884 30716
rect 3835 30685 3847 30688
rect 3789 30679 3847 30685
rect 3878 30676 3884 30688
rect 3936 30676 3942 30728
rect 3988 30725 4016 30756
rect 5166 30744 5172 30796
rect 5224 30784 5230 30796
rect 5445 30787 5503 30793
rect 5445 30784 5457 30787
rect 5224 30756 5457 30784
rect 5224 30744 5230 30756
rect 5445 30753 5457 30756
rect 5491 30753 5503 30787
rect 5445 30747 5503 30753
rect 6546 30744 6552 30796
rect 6604 30784 6610 30796
rect 7576 30793 7604 30824
rect 8938 30812 8944 30824
rect 8996 30812 9002 30864
rect 9861 30855 9919 30861
rect 9861 30821 9873 30855
rect 9907 30852 9919 30855
rect 10045 30855 10103 30861
rect 10045 30852 10057 30855
rect 9907 30824 10057 30852
rect 9907 30821 9919 30824
rect 9861 30815 9919 30821
rect 10045 30821 10057 30824
rect 10091 30821 10103 30855
rect 10778 30852 10784 30864
rect 10045 30815 10103 30821
rect 10152 30824 10784 30852
rect 6708 30787 6766 30793
rect 6708 30784 6720 30787
rect 6604 30756 6720 30784
rect 6604 30744 6610 30756
rect 6708 30753 6720 30756
rect 6754 30753 6766 30787
rect 6708 30747 6766 30753
rect 7193 30787 7251 30793
rect 7193 30753 7205 30787
rect 7239 30784 7251 30787
rect 7561 30787 7619 30793
rect 7561 30784 7573 30787
rect 7239 30756 7573 30784
rect 7239 30753 7251 30756
rect 7193 30747 7251 30753
rect 7561 30753 7573 30756
rect 7607 30753 7619 30787
rect 10152 30784 10180 30824
rect 10778 30812 10784 30824
rect 10836 30812 10842 30864
rect 12069 30855 12127 30861
rect 12069 30852 12081 30855
rect 11348 30824 12081 30852
rect 7561 30747 7619 30753
rect 8680 30756 10180 30784
rect 10413 30787 10471 30793
rect 3973 30719 4031 30725
rect 3973 30685 3985 30719
rect 4019 30685 4031 30719
rect 3973 30679 4031 30685
rect 5261 30719 5319 30725
rect 5261 30685 5273 30719
rect 5307 30716 5319 30719
rect 5350 30716 5356 30728
rect 5307 30688 5356 30716
rect 5307 30685 5319 30688
rect 5261 30679 5319 30685
rect 5350 30676 5356 30688
rect 5408 30676 5414 30728
rect 8018 30676 8024 30728
rect 8076 30725 8082 30728
rect 8076 30719 8104 30725
rect 8092 30685 8104 30719
rect 8076 30679 8104 30685
rect 8076 30676 8082 30679
rect 6917 30651 6975 30657
rect 6917 30617 6929 30651
rect 6963 30648 6975 30651
rect 7837 30651 7895 30657
rect 7837 30648 7849 30651
rect 6963 30620 7849 30648
rect 6963 30617 6975 30620
rect 6917 30611 6975 30617
rect 7837 30617 7849 30620
rect 7883 30648 7895 30651
rect 8386 30648 8392 30660
rect 7883 30620 8392 30648
rect 7883 30617 7895 30620
rect 7837 30611 7895 30617
rect 8386 30608 8392 30620
rect 8444 30608 8450 30660
rect 3142 30540 3148 30592
rect 3200 30580 3206 30592
rect 3789 30583 3847 30589
rect 3789 30580 3801 30583
rect 3200 30552 3801 30580
rect 3200 30540 3206 30552
rect 3789 30549 3801 30552
rect 3835 30549 3847 30583
rect 3789 30543 3847 30549
rect 4798 30540 4804 30592
rect 4856 30580 4862 30592
rect 5077 30583 5135 30589
rect 5077 30580 5089 30583
rect 4856 30552 5089 30580
rect 4856 30540 4862 30552
rect 5077 30549 5089 30552
rect 5123 30549 5135 30583
rect 5077 30543 5135 30549
rect 6825 30583 6883 30589
rect 6825 30549 6837 30583
rect 6871 30580 6883 30583
rect 7006 30580 7012 30592
rect 6871 30552 7012 30580
rect 6871 30549 6883 30552
rect 6825 30543 6883 30549
rect 7006 30540 7012 30552
rect 7064 30580 7070 30592
rect 7926 30580 7932 30592
rect 7064 30552 7932 30580
rect 7064 30540 7070 30552
rect 7926 30540 7932 30552
rect 7984 30580 7990 30592
rect 8680 30580 8708 30756
rect 10413 30753 10425 30787
rect 10459 30784 10471 30787
rect 11146 30784 11152 30796
rect 10459 30756 11152 30784
rect 10459 30753 10471 30756
rect 10413 30747 10471 30753
rect 11146 30744 11152 30756
rect 11204 30744 11210 30796
rect 11348 30728 11376 30824
rect 12069 30821 12081 30824
rect 12115 30821 12127 30855
rect 12069 30815 12127 30821
rect 12986 30812 12992 30864
rect 13044 30852 13050 30864
rect 13446 30852 13452 30864
rect 13044 30824 13452 30852
rect 13044 30812 13050 30824
rect 13446 30812 13452 30824
rect 13504 30812 13510 30864
rect 11698 30744 11704 30796
rect 11756 30744 11762 30796
rect 12158 30744 12164 30796
rect 12216 30784 12222 30796
rect 12529 30787 12587 30793
rect 12529 30784 12541 30787
rect 12216 30756 12541 30784
rect 12216 30744 12222 30756
rect 12529 30753 12541 30756
rect 12575 30753 12587 30787
rect 13998 30784 14004 30796
rect 12529 30747 12587 30753
rect 13004 30756 14004 30784
rect 9306 30676 9312 30728
rect 9364 30716 9370 30728
rect 9434 30719 9492 30725
rect 9434 30716 9446 30719
rect 9364 30688 9446 30716
rect 9364 30676 9370 30688
rect 9434 30685 9446 30688
rect 9480 30685 9492 30719
rect 9434 30679 9492 30685
rect 9950 30676 9956 30728
rect 10008 30676 10014 30728
rect 10226 30676 10232 30728
rect 10284 30676 10290 30728
rect 10686 30676 10692 30728
rect 10744 30676 10750 30728
rect 10962 30676 10968 30728
rect 11020 30676 11026 30728
rect 11057 30719 11115 30725
rect 11057 30685 11069 30719
rect 11103 30685 11115 30719
rect 11241 30719 11299 30725
rect 11241 30716 11253 30719
rect 11057 30679 11115 30685
rect 11164 30688 11253 30716
rect 11072 30648 11100 30679
rect 9646 30620 11100 30648
rect 7984 30552 8708 30580
rect 7984 30540 7990 30552
rect 9306 30540 9312 30592
rect 9364 30580 9370 30592
rect 9490 30580 9496 30592
rect 9364 30552 9496 30580
rect 9364 30540 9370 30552
rect 9490 30540 9496 30552
rect 9548 30580 9554 30592
rect 9646 30580 9674 30620
rect 9548 30552 9674 30580
rect 9548 30540 9554 30552
rect 10778 30540 10784 30592
rect 10836 30540 10842 30592
rect 11164 30580 11192 30688
rect 11241 30685 11253 30688
rect 11287 30685 11299 30719
rect 11241 30679 11299 30685
rect 11330 30676 11336 30728
rect 11388 30676 11394 30728
rect 11790 30676 11796 30728
rect 11848 30676 11854 30728
rect 12434 30676 12440 30728
rect 12492 30676 12498 30728
rect 12802 30676 12808 30728
rect 12860 30676 12866 30728
rect 13004 30725 13032 30756
rect 13998 30744 14004 30756
rect 14056 30744 14062 30796
rect 14090 30744 14096 30796
rect 14148 30744 14154 30796
rect 12989 30719 13047 30725
rect 12989 30685 13001 30719
rect 13035 30685 13047 30719
rect 12989 30679 13047 30685
rect 13081 30719 13139 30725
rect 13081 30685 13093 30719
rect 13127 30716 13139 30719
rect 13262 30716 13268 30728
rect 13127 30688 13268 30716
rect 13127 30685 13139 30688
rect 13081 30679 13139 30685
rect 13262 30676 13268 30688
rect 13320 30676 13326 30728
rect 13446 30676 13452 30728
rect 13504 30676 13510 30728
rect 12897 30651 12955 30657
rect 12897 30617 12909 30651
rect 12943 30648 12955 30651
rect 13566 30651 13624 30657
rect 13566 30648 13578 30651
rect 12943 30620 13578 30648
rect 12943 30617 12955 30620
rect 12897 30611 12955 30617
rect 13566 30617 13578 30620
rect 13612 30617 13624 30651
rect 14338 30651 14396 30657
rect 14338 30648 14350 30651
rect 13566 30611 13624 30617
rect 13740 30620 14350 30648
rect 11238 30580 11244 30592
rect 11164 30552 11244 30580
rect 11238 30540 11244 30552
rect 11296 30580 11302 30592
rect 11425 30583 11483 30589
rect 11425 30580 11437 30583
rect 11296 30552 11437 30580
rect 11296 30540 11302 30552
rect 11425 30549 11437 30552
rect 11471 30549 11483 30583
rect 11425 30543 11483 30549
rect 13078 30540 13084 30592
rect 13136 30580 13142 30592
rect 13740 30589 13768 30620
rect 14338 30617 14350 30620
rect 14384 30617 14396 30651
rect 14338 30611 14396 30617
rect 13357 30583 13415 30589
rect 13357 30580 13369 30583
rect 13136 30552 13369 30580
rect 13136 30540 13142 30552
rect 13357 30549 13369 30552
rect 13403 30549 13415 30583
rect 13357 30543 13415 30549
rect 13725 30583 13783 30589
rect 13725 30549 13737 30583
rect 13771 30549 13783 30583
rect 13725 30543 13783 30549
rect 14090 30540 14096 30592
rect 14148 30580 14154 30592
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 14148 30552 15485 30580
rect 14148 30540 14154 30552
rect 15473 30549 15485 30552
rect 15519 30549 15531 30583
rect 15473 30543 15531 30549
rect 1104 30490 16836 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 16836 30490
rect 1104 30416 16836 30438
rect 3878 30376 3884 30388
rect 3620 30348 3884 30376
rect 2958 30268 2964 30320
rect 3016 30268 3022 30320
rect 3620 30317 3648 30348
rect 3878 30336 3884 30348
rect 3936 30336 3942 30388
rect 5261 30379 5319 30385
rect 5261 30345 5273 30379
rect 5307 30376 5319 30379
rect 5350 30376 5356 30388
rect 5307 30348 5356 30376
rect 5307 30345 5319 30348
rect 5261 30339 5319 30345
rect 5350 30336 5356 30348
rect 5408 30376 5414 30388
rect 5534 30376 5540 30388
rect 5408 30348 5540 30376
rect 5408 30336 5414 30348
rect 5534 30336 5540 30348
rect 5592 30336 5598 30388
rect 8478 30336 8484 30388
rect 8536 30376 8542 30388
rect 8536 30348 9076 30376
rect 8536 30336 8542 30348
rect 3177 30311 3235 30317
rect 3177 30277 3189 30311
rect 3223 30308 3235 30311
rect 3421 30311 3479 30317
rect 3421 30308 3433 30311
rect 3223 30280 3433 30308
rect 3223 30277 3235 30280
rect 3177 30271 3235 30277
rect 3421 30277 3433 30280
rect 3467 30277 3479 30311
rect 3421 30271 3479 30277
rect 3605 30311 3663 30317
rect 3605 30277 3617 30311
rect 3651 30277 3663 30311
rect 3605 30271 3663 30277
rect 3694 30268 3700 30320
rect 3752 30308 3758 30320
rect 3789 30311 3847 30317
rect 3789 30308 3801 30311
rect 3752 30280 3801 30308
rect 3752 30268 3758 30280
rect 3789 30277 3801 30280
rect 3835 30277 3847 30311
rect 4706 30308 4712 30320
rect 3789 30271 3847 30277
rect 3896 30280 4712 30308
rect 3896 30249 3924 30280
rect 4706 30268 4712 30280
rect 4764 30268 4770 30320
rect 6362 30268 6368 30320
rect 6420 30308 6426 30320
rect 6420 30280 8708 30308
rect 6420 30268 6426 30280
rect 3881 30243 3939 30249
rect 3881 30209 3893 30243
rect 3927 30209 3939 30243
rect 4137 30243 4195 30249
rect 4137 30240 4149 30243
rect 3881 30203 3939 30209
rect 3988 30212 4149 30240
rect 3988 30172 4016 30212
rect 4137 30209 4149 30212
rect 4183 30209 4195 30243
rect 4137 30203 4195 30209
rect 8294 30200 8300 30252
rect 8352 30240 8358 30252
rect 8680 30249 8708 30280
rect 9048 30249 9076 30348
rect 9950 30336 9956 30388
rect 10008 30376 10014 30388
rect 10873 30379 10931 30385
rect 10873 30376 10885 30379
rect 10008 30348 10885 30376
rect 10008 30336 10014 30348
rect 10873 30345 10885 30348
rect 10919 30345 10931 30379
rect 10873 30339 10931 30345
rect 12544 30348 12756 30376
rect 12544 30317 12572 30348
rect 12529 30311 12587 30317
rect 12529 30277 12541 30311
rect 12575 30277 12587 30311
rect 12529 30271 12587 30277
rect 12618 30268 12624 30320
rect 12676 30268 12682 30320
rect 12728 30308 12756 30348
rect 12802 30336 12808 30388
rect 12860 30376 12866 30388
rect 13354 30376 13360 30388
rect 12860 30348 13360 30376
rect 12860 30336 12866 30348
rect 13354 30336 13360 30348
rect 13412 30336 13418 30388
rect 13170 30308 13176 30320
rect 12728 30280 13176 30308
rect 13170 30268 13176 30280
rect 13228 30308 13234 30320
rect 13509 30311 13567 30317
rect 13509 30308 13521 30311
rect 13228 30280 13521 30308
rect 13228 30268 13234 30280
rect 13509 30277 13521 30280
rect 13555 30277 13567 30311
rect 13509 30271 13567 30277
rect 13725 30311 13783 30317
rect 13725 30277 13737 30311
rect 13771 30308 13783 30311
rect 14090 30308 14096 30320
rect 13771 30280 14096 30308
rect 13771 30277 13783 30280
rect 13725 30271 13783 30277
rect 8481 30243 8539 30249
rect 8481 30240 8493 30243
rect 8352 30212 8493 30240
rect 8352 30200 8358 30212
rect 8481 30209 8493 30212
rect 8527 30209 8539 30243
rect 8481 30203 8539 30209
rect 8665 30243 8723 30249
rect 8665 30209 8677 30243
rect 8711 30240 8723 30243
rect 8941 30243 8999 30249
rect 8941 30240 8953 30243
rect 8711 30212 8953 30240
rect 8711 30209 8723 30212
rect 8665 30203 8723 30209
rect 8941 30209 8953 30212
rect 8987 30209 8999 30243
rect 8941 30203 8999 30209
rect 9033 30243 9091 30249
rect 9033 30209 9045 30243
rect 9079 30209 9091 30243
rect 9033 30203 9091 30209
rect 3344 30144 4016 30172
rect 8496 30172 8524 30203
rect 9048 30172 9076 30203
rect 9122 30200 9128 30252
rect 9180 30240 9186 30252
rect 9217 30243 9275 30249
rect 9217 30240 9229 30243
rect 9180 30212 9229 30240
rect 9180 30200 9186 30212
rect 9217 30209 9229 30212
rect 9263 30209 9275 30243
rect 9217 30203 9275 30209
rect 9398 30200 9404 30252
rect 9456 30200 9462 30252
rect 9677 30243 9735 30249
rect 9677 30209 9689 30243
rect 9723 30240 9735 30243
rect 9858 30240 9864 30252
rect 9723 30212 9864 30240
rect 9723 30209 9735 30212
rect 9677 30203 9735 30209
rect 9858 30200 9864 30212
rect 9916 30200 9922 30252
rect 11054 30200 11060 30252
rect 11112 30200 11118 30252
rect 11241 30243 11299 30249
rect 11241 30209 11253 30243
rect 11287 30240 11299 30243
rect 11330 30240 11336 30252
rect 11287 30212 11336 30240
rect 11287 30209 11299 30212
rect 11241 30203 11299 30209
rect 11330 30200 11336 30212
rect 11388 30200 11394 30252
rect 11790 30200 11796 30252
rect 11848 30240 11854 30252
rect 11885 30243 11943 30249
rect 11885 30240 11897 30243
rect 11848 30212 11897 30240
rect 11848 30200 11854 30212
rect 11885 30209 11897 30212
rect 11931 30209 11943 30243
rect 11885 30203 11943 30209
rect 12069 30243 12127 30249
rect 12069 30209 12081 30243
rect 12115 30240 12127 30243
rect 12158 30240 12164 30252
rect 12115 30212 12164 30240
rect 12115 30209 12127 30212
rect 12069 30203 12127 30209
rect 9493 30175 9551 30181
rect 9493 30172 9505 30175
rect 8496 30144 8984 30172
rect 9048 30144 9505 30172
rect 3344 30113 3372 30144
rect 3329 30107 3387 30113
rect 3329 30073 3341 30107
rect 3375 30073 3387 30107
rect 3329 30067 3387 30073
rect 5626 30064 5632 30116
rect 5684 30104 5690 30116
rect 6270 30104 6276 30116
rect 5684 30076 6276 30104
rect 5684 30064 5690 30076
rect 6270 30064 6276 30076
rect 6328 30104 6334 30116
rect 8956 30104 8984 30144
rect 9493 30141 9505 30144
rect 9539 30141 9551 30175
rect 11900 30172 11928 30203
rect 12158 30200 12164 30212
rect 12216 30200 12222 30252
rect 12434 30200 12440 30252
rect 12492 30240 12498 30252
rect 12713 30243 12771 30249
rect 12713 30240 12725 30243
rect 12492 30212 12725 30240
rect 12492 30200 12498 30212
rect 12713 30209 12725 30212
rect 12759 30240 12771 30243
rect 13740 30240 13768 30271
rect 14090 30268 14096 30280
rect 14148 30268 14154 30320
rect 12759 30212 13768 30240
rect 13817 30243 13875 30249
rect 12759 30209 12771 30212
rect 12713 30203 12771 30209
rect 13817 30209 13829 30243
rect 13863 30209 13875 30243
rect 13817 30203 13875 30209
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30240 13967 30243
rect 14458 30240 14464 30252
rect 13955 30212 14464 30240
rect 13955 30209 13967 30212
rect 13909 30203 13967 30209
rect 11900 30144 12940 30172
rect 9493 30135 9551 30141
rect 9125 30107 9183 30113
rect 9125 30104 9137 30107
rect 6328 30076 8892 30104
rect 8956 30076 9137 30104
rect 6328 30064 6334 30076
rect 3142 29996 3148 30048
rect 3200 29996 3206 30048
rect 8478 29996 8484 30048
rect 8536 29996 8542 30048
rect 8754 29996 8760 30048
rect 8812 29996 8818 30048
rect 8864 30036 8892 30076
rect 9125 30073 9137 30076
rect 9171 30104 9183 30107
rect 9306 30104 9312 30116
rect 9171 30076 9312 30104
rect 9171 30073 9183 30076
rect 9125 30067 9183 30073
rect 9306 30064 9312 30076
rect 9364 30064 9370 30116
rect 9582 30104 9588 30116
rect 9416 30076 9588 30104
rect 9416 30045 9444 30076
rect 9582 30064 9588 30076
rect 9640 30064 9646 30116
rect 12434 30104 12440 30116
rect 12084 30076 12440 30104
rect 9401 30039 9459 30045
rect 9401 30036 9413 30039
rect 8864 30008 9413 30036
rect 9401 30005 9413 30008
rect 9447 30005 9459 30039
rect 9401 29999 9459 30005
rect 9490 29996 9496 30048
rect 9548 30036 9554 30048
rect 9861 30039 9919 30045
rect 9861 30036 9873 30039
rect 9548 30008 9873 30036
rect 9548 29996 9554 30008
rect 9861 30005 9873 30008
rect 9907 30005 9919 30039
rect 9861 29999 9919 30005
rect 11238 29996 11244 30048
rect 11296 29996 11302 30048
rect 11422 29996 11428 30048
rect 11480 30036 11486 30048
rect 12084 30045 12112 30076
rect 12434 30064 12440 30076
rect 12492 30064 12498 30116
rect 12912 30113 12940 30144
rect 13170 30132 13176 30184
rect 13228 30172 13234 30184
rect 13722 30172 13728 30184
rect 13228 30144 13728 30172
rect 13228 30132 13234 30144
rect 13722 30132 13728 30144
rect 13780 30172 13786 30184
rect 13832 30172 13860 30203
rect 13780 30144 13860 30172
rect 13780 30132 13786 30144
rect 12897 30107 12955 30113
rect 12897 30073 12909 30107
rect 12943 30104 12955 30107
rect 13630 30104 13636 30116
rect 12943 30076 13636 30104
rect 12943 30073 12955 30076
rect 12897 30067 12955 30073
rect 13630 30064 13636 30076
rect 13688 30064 13694 30116
rect 11701 30039 11759 30045
rect 11701 30036 11713 30039
rect 11480 30008 11713 30036
rect 11480 29996 11486 30008
rect 11701 30005 11713 30008
rect 11747 30005 11759 30039
rect 11701 29999 11759 30005
rect 12069 30039 12127 30045
rect 12069 30005 12081 30039
rect 12115 30005 12127 30039
rect 12069 29999 12127 30005
rect 12342 29996 12348 30048
rect 12400 29996 12406 30048
rect 12618 29996 12624 30048
rect 12676 30036 12682 30048
rect 13541 30039 13599 30045
rect 13541 30036 13553 30039
rect 12676 30008 13553 30036
rect 12676 29996 12682 30008
rect 13541 30005 13553 30008
rect 13587 30036 13599 30039
rect 13924 30036 13952 30203
rect 14458 30200 14464 30212
rect 14516 30200 14522 30252
rect 13998 30064 14004 30116
rect 14056 30104 14062 30116
rect 14093 30107 14151 30113
rect 14093 30104 14105 30107
rect 14056 30076 14105 30104
rect 14056 30064 14062 30076
rect 14093 30073 14105 30076
rect 14139 30073 14151 30107
rect 14093 30067 14151 30073
rect 13587 30008 13952 30036
rect 13587 30005 13599 30008
rect 13541 29999 13599 30005
rect 1104 29946 16836 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 16836 29946
rect 1104 29872 16836 29894
rect 8478 29792 8484 29844
rect 8536 29792 8542 29844
rect 10410 29792 10416 29844
rect 10468 29832 10474 29844
rect 10468 29804 11192 29832
rect 10468 29792 10474 29804
rect 5905 29767 5963 29773
rect 5905 29733 5917 29767
rect 5951 29764 5963 29767
rect 9398 29764 9404 29776
rect 5951 29736 7512 29764
rect 5951 29733 5963 29736
rect 5905 29727 5963 29733
rect 3694 29656 3700 29708
rect 3752 29696 3758 29708
rect 3752 29668 4292 29696
rect 3752 29656 3758 29668
rect 2222 29588 2228 29640
rect 2280 29588 2286 29640
rect 4264 29637 4292 29668
rect 4706 29656 4712 29708
rect 4764 29696 4770 29708
rect 5810 29696 5816 29708
rect 4764 29668 5029 29696
rect 4764 29656 4770 29668
rect 5001 29637 5029 29668
rect 5184 29668 5816 29696
rect 5184 29637 5212 29668
rect 5810 29656 5816 29668
rect 5868 29656 5874 29708
rect 3973 29631 4031 29637
rect 3973 29597 3985 29631
rect 4019 29597 4031 29631
rect 3973 29591 4031 29597
rect 4249 29631 4307 29637
rect 4249 29597 4261 29631
rect 4295 29597 4307 29631
rect 4249 29591 4307 29597
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29597 4951 29631
rect 4893 29591 4951 29597
rect 4986 29631 5044 29637
rect 4986 29597 4998 29631
rect 5032 29597 5044 29631
rect 4986 29591 5044 29597
rect 5169 29631 5227 29637
rect 5169 29597 5181 29631
rect 5215 29597 5227 29631
rect 5169 29591 5227 29597
rect 5399 29631 5457 29637
rect 5399 29597 5411 29631
rect 5445 29628 5457 29631
rect 5920 29628 5948 29727
rect 6733 29699 6791 29705
rect 6733 29665 6745 29699
rect 6779 29665 6791 29699
rect 6733 29659 6791 29665
rect 5445 29600 5948 29628
rect 5445 29597 5457 29600
rect 5399 29591 5457 29597
rect 2498 29569 2504 29572
rect 2492 29523 2504 29569
rect 2498 29520 2504 29523
rect 2556 29520 2562 29572
rect 3988 29560 4016 29591
rect 4908 29560 4936 29591
rect 6178 29588 6184 29640
rect 6236 29588 6242 29640
rect 6270 29588 6276 29640
rect 6328 29588 6334 29640
rect 6362 29588 6368 29640
rect 6420 29628 6426 29640
rect 6641 29631 6699 29637
rect 6641 29628 6653 29631
rect 6420 29600 6653 29628
rect 6420 29588 6426 29600
rect 6641 29597 6653 29600
rect 6687 29597 6699 29631
rect 6748 29628 6776 29659
rect 7006 29656 7012 29708
rect 7064 29656 7070 29708
rect 7484 29705 7512 29736
rect 8496 29736 9404 29764
rect 8496 29705 8524 29736
rect 9398 29724 9404 29736
rect 9456 29724 9462 29776
rect 11164 29764 11192 29804
rect 11238 29792 11244 29844
rect 11296 29832 11302 29844
rect 11333 29835 11391 29841
rect 11333 29832 11345 29835
rect 11296 29804 11345 29832
rect 11296 29792 11302 29804
rect 11333 29801 11345 29804
rect 11379 29801 11391 29835
rect 11333 29795 11391 29801
rect 12894 29764 12900 29776
rect 10336 29736 11100 29764
rect 11164 29736 12900 29764
rect 7469 29699 7527 29705
rect 7469 29665 7481 29699
rect 7515 29665 7527 29699
rect 7469 29659 7527 29665
rect 8481 29699 8539 29705
rect 8481 29665 8493 29699
rect 8527 29665 8539 29699
rect 8481 29659 8539 29665
rect 8754 29656 8760 29708
rect 8812 29696 8818 29708
rect 9769 29699 9827 29705
rect 9769 29696 9781 29699
rect 8812 29668 9781 29696
rect 8812 29656 8818 29668
rect 9769 29665 9781 29668
rect 9815 29665 9827 29699
rect 9769 29659 9827 29665
rect 6822 29628 6828 29640
rect 6748 29600 6828 29628
rect 6641 29591 6699 29597
rect 6822 29588 6828 29600
rect 6880 29628 6886 29640
rect 7374 29628 7380 29640
rect 6880 29600 7380 29628
rect 6880 29588 6886 29600
rect 7374 29588 7380 29600
rect 7432 29588 7438 29640
rect 7561 29631 7619 29637
rect 7561 29597 7573 29631
rect 7607 29628 7619 29631
rect 7607 29600 8524 29628
rect 7607 29597 7619 29600
rect 7561 29591 7619 29597
rect 3620 29532 4936 29560
rect 5261 29563 5319 29569
rect 3620 29504 3648 29532
rect 5261 29529 5273 29563
rect 5307 29560 5319 29563
rect 8297 29563 8355 29569
rect 5307 29532 5396 29560
rect 5307 29529 5319 29532
rect 5261 29523 5319 29529
rect 5368 29504 5396 29532
rect 8297 29529 8309 29563
rect 8343 29529 8355 29563
rect 8496 29560 8524 29600
rect 8570 29588 8576 29640
rect 8628 29588 8634 29640
rect 9033 29631 9091 29637
rect 9033 29628 9045 29631
rect 8680 29600 9045 29628
rect 8680 29572 8708 29600
rect 9033 29597 9045 29600
rect 9079 29597 9091 29631
rect 9033 29591 9091 29597
rect 9490 29588 9496 29640
rect 9548 29588 9554 29640
rect 10137 29631 10195 29637
rect 10137 29597 10149 29631
rect 10183 29628 10195 29631
rect 10336 29628 10364 29736
rect 10410 29656 10416 29708
rect 10468 29656 10474 29708
rect 10686 29637 10692 29640
rect 10183 29600 10364 29628
rect 10505 29631 10563 29637
rect 10183 29597 10195 29600
rect 10137 29591 10195 29597
rect 10505 29597 10517 29631
rect 10551 29597 10563 29631
rect 10505 29591 10563 29597
rect 10653 29631 10692 29637
rect 10653 29597 10665 29631
rect 10653 29591 10692 29597
rect 8662 29560 8668 29572
rect 8496 29532 8668 29560
rect 8297 29523 8355 29529
rect 3602 29452 3608 29504
rect 3660 29452 3666 29504
rect 3786 29452 3792 29504
rect 3844 29452 3850 29504
rect 3878 29452 3884 29504
rect 3936 29492 3942 29504
rect 4157 29495 4215 29501
rect 4157 29492 4169 29495
rect 3936 29464 4169 29492
rect 3936 29452 3942 29464
rect 4157 29461 4169 29464
rect 4203 29492 4215 29495
rect 5350 29492 5356 29504
rect 4203 29464 5356 29492
rect 4203 29461 4215 29464
rect 4157 29455 4215 29461
rect 5350 29452 5356 29464
rect 5408 29452 5414 29504
rect 5534 29452 5540 29504
rect 5592 29452 5598 29504
rect 7929 29495 7987 29501
rect 7929 29461 7941 29495
rect 7975 29492 7987 29495
rect 8312 29492 8340 29523
rect 8662 29520 8668 29532
rect 8720 29520 8726 29572
rect 10226 29560 10232 29572
rect 8772 29532 10232 29560
rect 8772 29501 8800 29532
rect 10226 29520 10232 29532
rect 10284 29560 10290 29572
rect 10520 29560 10548 29591
rect 10686 29588 10692 29591
rect 10744 29588 10750 29640
rect 10778 29588 10784 29640
rect 10836 29588 10842 29640
rect 10970 29631 11028 29637
rect 10970 29597 10982 29631
rect 11016 29597 11028 29631
rect 11072 29628 11100 29736
rect 12894 29724 12900 29736
rect 12952 29764 12958 29776
rect 13170 29764 13176 29776
rect 12952 29736 13176 29764
rect 12952 29724 12958 29736
rect 13170 29724 13176 29736
rect 13228 29724 13234 29776
rect 13541 29699 13599 29705
rect 13541 29696 13553 29699
rect 13372 29668 13553 29696
rect 11241 29631 11299 29637
rect 11072 29600 11192 29628
rect 10970 29591 11028 29597
rect 10284 29532 10548 29560
rect 10284 29520 10290 29532
rect 10870 29520 10876 29572
rect 10928 29520 10934 29572
rect 7975 29464 8340 29492
rect 8757 29495 8815 29501
rect 7975 29461 7987 29464
rect 7929 29455 7987 29461
rect 8757 29461 8769 29495
rect 8803 29461 8815 29495
rect 8757 29455 8815 29461
rect 10594 29452 10600 29504
rect 10652 29492 10658 29504
rect 10980 29492 11008 29591
rect 11164 29501 11192 29600
rect 11241 29597 11253 29631
rect 11287 29597 11299 29631
rect 11241 29591 11299 29597
rect 11425 29631 11483 29637
rect 11425 29597 11437 29631
rect 11471 29628 11483 29631
rect 11974 29628 11980 29640
rect 11471 29600 11980 29628
rect 11471 29597 11483 29600
rect 11425 29591 11483 29597
rect 11256 29560 11284 29591
rect 11974 29588 11980 29600
rect 12032 29588 12038 29640
rect 12342 29588 12348 29640
rect 12400 29628 12406 29640
rect 13372 29637 13400 29668
rect 13541 29665 13553 29668
rect 13587 29665 13599 29699
rect 13541 29659 13599 29665
rect 13173 29631 13231 29637
rect 13173 29628 13185 29631
rect 12400 29600 13185 29628
rect 12400 29588 12406 29600
rect 13173 29597 13185 29600
rect 13219 29597 13231 29631
rect 13173 29591 13231 29597
rect 13357 29631 13415 29637
rect 13357 29597 13369 29631
rect 13403 29597 13415 29631
rect 13357 29591 13415 29597
rect 13446 29588 13452 29640
rect 13504 29588 13510 29640
rect 13630 29588 13636 29640
rect 13688 29628 13694 29640
rect 14826 29628 14832 29640
rect 13688 29600 14832 29628
rect 13688 29588 13694 29600
rect 14826 29588 14832 29600
rect 14884 29588 14890 29640
rect 11606 29560 11612 29572
rect 11256 29532 11612 29560
rect 11606 29520 11612 29532
rect 11664 29560 11670 29572
rect 12158 29560 12164 29572
rect 11664 29532 12164 29560
rect 11664 29520 11670 29532
rect 12158 29520 12164 29532
rect 12216 29520 12222 29572
rect 10652 29464 11008 29492
rect 11149 29495 11207 29501
rect 10652 29452 10658 29464
rect 11149 29461 11161 29495
rect 11195 29461 11207 29495
rect 11149 29455 11207 29461
rect 12894 29452 12900 29504
rect 12952 29492 12958 29504
rect 13265 29495 13323 29501
rect 13265 29492 13277 29495
rect 12952 29464 13277 29492
rect 12952 29452 12958 29464
rect 13265 29461 13277 29464
rect 13311 29461 13323 29495
rect 13265 29455 13323 29461
rect 1104 29402 16836 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 16836 29402
rect 1104 29328 16836 29350
rect 2498 29248 2504 29300
rect 2556 29248 2562 29300
rect 2685 29291 2743 29297
rect 2685 29257 2697 29291
rect 2731 29288 2743 29291
rect 2958 29288 2964 29300
rect 2731 29260 2964 29288
rect 2731 29257 2743 29260
rect 2685 29251 2743 29257
rect 2958 29248 2964 29260
rect 3016 29248 3022 29300
rect 3405 29291 3463 29297
rect 3405 29257 3417 29291
rect 3451 29288 3463 29291
rect 3694 29288 3700 29300
rect 3451 29260 3700 29288
rect 3451 29257 3463 29260
rect 3405 29251 3463 29257
rect 3694 29248 3700 29260
rect 3752 29248 3758 29300
rect 4706 29248 4712 29300
rect 4764 29288 4770 29300
rect 4764 29260 6316 29288
rect 4764 29248 4770 29260
rect 3602 29180 3608 29232
rect 3660 29180 3666 29232
rect 5534 29220 5540 29232
rect 5092 29192 5540 29220
rect 4798 29112 4804 29164
rect 4856 29112 4862 29164
rect 4890 29112 4896 29164
rect 4948 29152 4954 29164
rect 5092 29161 5120 29192
rect 5534 29180 5540 29192
rect 5592 29180 5598 29232
rect 6288 29220 6316 29260
rect 6362 29248 6368 29300
rect 6420 29288 6426 29300
rect 8389 29291 8447 29297
rect 8389 29288 8401 29291
rect 6420 29260 8401 29288
rect 6420 29248 6426 29260
rect 8389 29257 8401 29260
rect 8435 29257 8447 29291
rect 8389 29251 8447 29257
rect 8757 29291 8815 29297
rect 8757 29257 8769 29291
rect 8803 29288 8815 29291
rect 9398 29288 9404 29300
rect 8803 29260 9404 29288
rect 8803 29257 8815 29260
rect 8757 29251 8815 29257
rect 9398 29248 9404 29260
rect 9456 29248 9462 29300
rect 10594 29248 10600 29300
rect 10652 29248 10658 29300
rect 10686 29248 10692 29300
rect 10744 29248 10750 29300
rect 12986 29248 12992 29300
rect 13044 29288 13050 29300
rect 13081 29291 13139 29297
rect 13081 29288 13093 29291
rect 13044 29260 13093 29288
rect 13044 29248 13050 29260
rect 13081 29257 13093 29260
rect 13127 29257 13139 29291
rect 13081 29251 13139 29257
rect 13357 29291 13415 29297
rect 13357 29257 13369 29291
rect 13403 29257 13415 29291
rect 13357 29251 13415 29257
rect 11422 29220 11428 29232
rect 6288 29192 8248 29220
rect 4985 29155 5043 29161
rect 4985 29152 4997 29155
rect 4948 29124 4997 29152
rect 4948 29112 4954 29124
rect 4985 29121 4997 29124
rect 5031 29121 5043 29155
rect 4985 29115 5043 29121
rect 5077 29155 5135 29161
rect 5077 29121 5089 29155
rect 5123 29121 5135 29155
rect 5077 29115 5135 29121
rect 5350 29112 5356 29164
rect 5408 29112 5414 29164
rect 7190 29112 7196 29164
rect 7248 29152 7254 29164
rect 7478 29155 7536 29161
rect 7478 29152 7490 29155
rect 7248 29124 7490 29152
rect 7248 29112 7254 29124
rect 7478 29121 7490 29124
rect 7524 29121 7536 29155
rect 8220 29152 8248 29192
rect 11164 29192 11428 29220
rect 8294 29152 8300 29164
rect 8220 29124 8300 29152
rect 7478 29115 7536 29121
rect 8294 29112 8300 29124
rect 8352 29112 8358 29164
rect 8478 29112 8484 29164
rect 8536 29152 8542 29164
rect 8573 29155 8631 29161
rect 8573 29152 8585 29155
rect 8536 29124 8585 29152
rect 8536 29112 8542 29124
rect 8573 29121 8585 29124
rect 8619 29121 8631 29155
rect 8573 29115 8631 29121
rect 10226 29112 10232 29164
rect 10284 29112 10290 29164
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29152 10471 29155
rect 10594 29152 10600 29164
rect 10459 29124 10600 29152
rect 10459 29121 10471 29124
rect 10413 29115 10471 29121
rect 10594 29112 10600 29124
rect 10652 29152 10658 29164
rect 11164 29161 11192 29192
rect 11422 29180 11428 29192
rect 11480 29180 11486 29232
rect 11517 29223 11575 29229
rect 11517 29189 11529 29223
rect 11563 29189 11575 29223
rect 11517 29183 11575 29189
rect 10965 29155 11023 29161
rect 10965 29152 10977 29155
rect 10652 29124 10977 29152
rect 10652 29112 10658 29124
rect 10965 29121 10977 29124
rect 11011 29121 11023 29155
rect 10965 29115 11023 29121
rect 11057 29155 11115 29161
rect 11057 29121 11069 29155
rect 11103 29121 11115 29155
rect 11057 29115 11115 29121
rect 11149 29155 11207 29161
rect 11149 29121 11161 29155
rect 11195 29121 11207 29155
rect 11149 29115 11207 29121
rect 11333 29155 11391 29161
rect 11333 29121 11345 29155
rect 11379 29152 11391 29155
rect 11532 29152 11560 29183
rect 11698 29180 11704 29232
rect 11756 29220 11762 29232
rect 12253 29223 12311 29229
rect 12253 29220 12265 29223
rect 11756 29192 11928 29220
rect 11756 29180 11762 29192
rect 11379 29124 11560 29152
rect 11379 29121 11391 29124
rect 11333 29115 11391 29121
rect 5188 29087 5246 29093
rect 5188 29053 5200 29087
rect 5234 29084 5246 29087
rect 5442 29084 5448 29096
rect 5234 29056 5448 29084
rect 5234 29053 5246 29056
rect 5188 29047 5246 29053
rect 5442 29044 5448 29056
rect 5500 29044 5506 29096
rect 7742 29044 7748 29096
rect 7800 29044 7806 29096
rect 10244 29084 10272 29112
rect 11072 29084 11100 29115
rect 11790 29112 11796 29164
rect 11848 29112 11854 29164
rect 11900 29161 11928 29192
rect 11992 29192 12265 29220
rect 11992 29164 12020 29192
rect 12253 29189 12265 29192
rect 12299 29189 12311 29223
rect 12710 29220 12716 29232
rect 12253 29183 12311 29189
rect 12544 29192 12716 29220
rect 11885 29155 11943 29161
rect 11885 29121 11897 29155
rect 11931 29121 11943 29155
rect 11885 29115 11943 29121
rect 11974 29112 11980 29164
rect 12032 29112 12038 29164
rect 12158 29112 12164 29164
rect 12216 29112 12222 29164
rect 12544 29161 12572 29192
rect 12710 29180 12716 29192
rect 12768 29180 12774 29232
rect 13372 29220 13400 29251
rect 14826 29248 14832 29300
rect 14884 29248 14890 29300
rect 13694 29223 13752 29229
rect 13694 29220 13706 29223
rect 13372 29192 13706 29220
rect 13694 29189 13706 29192
rect 13740 29189 13752 29223
rect 13694 29183 13752 29189
rect 12528 29155 12586 29161
rect 12528 29121 12540 29155
rect 12574 29121 12586 29155
rect 12528 29115 12586 29121
rect 12621 29155 12679 29161
rect 12621 29121 12633 29155
rect 12667 29121 12679 29155
rect 12621 29115 12679 29121
rect 10244 29056 11100 29084
rect 12066 29044 12072 29096
rect 12124 29084 12130 29096
rect 12636 29084 12664 29115
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 12989 29155 13047 29161
rect 12989 29152 13001 29155
rect 12860 29124 13001 29152
rect 12860 29112 12866 29124
rect 12989 29121 13001 29124
rect 13035 29152 13047 29155
rect 13078 29152 13084 29164
rect 13035 29124 13084 29152
rect 13035 29121 13047 29124
rect 12989 29115 13047 29121
rect 13078 29112 13084 29124
rect 13136 29112 13142 29164
rect 12124 29056 12664 29084
rect 12124 29044 12130 29056
rect 12710 29044 12716 29096
rect 12768 29044 12774 29096
rect 12894 29044 12900 29096
rect 12952 29084 12958 29096
rect 13198 29087 13256 29093
rect 13198 29084 13210 29087
rect 12952 29056 13210 29084
rect 12952 29044 12958 29056
rect 13198 29053 13210 29056
rect 13244 29053 13256 29087
rect 13198 29047 13256 29053
rect 13446 29044 13452 29096
rect 13504 29044 13510 29096
rect 3053 29019 3111 29025
rect 3053 28985 3065 29019
rect 3099 29016 3111 29019
rect 3234 29016 3240 29028
rect 3099 28988 3240 29016
rect 3099 28985 3111 28988
rect 3053 28979 3111 28985
rect 3234 28976 3240 28988
rect 3292 28976 3298 29028
rect 3786 29016 3792 29028
rect 3344 28988 3792 29016
rect 2685 28951 2743 28957
rect 2685 28917 2697 28951
rect 2731 28948 2743 28951
rect 3344 28948 3372 28988
rect 3786 28976 3792 28988
rect 3844 28976 3850 29028
rect 4893 29019 4951 29025
rect 4893 28985 4905 29019
rect 4939 29016 4951 29019
rect 6730 29016 6736 29028
rect 4939 28988 6736 29016
rect 4939 28985 4951 28988
rect 4893 28979 4951 28985
rect 6730 28976 6736 28988
rect 6788 28976 6794 29028
rect 2731 28920 3372 28948
rect 3421 28951 3479 28957
rect 2731 28917 2743 28920
rect 2685 28911 2743 28917
rect 3421 28917 3433 28951
rect 3467 28948 3479 28951
rect 3878 28948 3884 28960
rect 3467 28920 3884 28948
rect 3467 28917 3479 28920
rect 3421 28911 3479 28917
rect 3878 28908 3884 28920
rect 3936 28908 3942 28960
rect 1104 28858 16836 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 16836 28858
rect 1104 28784 16836 28806
rect 4525 28747 4583 28753
rect 4525 28713 4537 28747
rect 4571 28744 4583 28747
rect 4798 28744 4804 28756
rect 4571 28716 4804 28744
rect 4571 28713 4583 28716
rect 4525 28707 4583 28713
rect 4798 28704 4804 28716
rect 4856 28704 4862 28756
rect 5810 28704 5816 28756
rect 5868 28744 5874 28756
rect 6181 28747 6239 28753
rect 6181 28744 6193 28747
rect 5868 28716 6193 28744
rect 5868 28704 5874 28716
rect 6181 28713 6193 28716
rect 6227 28713 6239 28747
rect 6181 28707 6239 28713
rect 7190 28704 7196 28756
rect 7248 28704 7254 28756
rect 10226 28704 10232 28756
rect 10284 28744 10290 28756
rect 10505 28747 10563 28753
rect 10505 28744 10517 28747
rect 10284 28716 10517 28744
rect 10284 28704 10290 28716
rect 10505 28713 10517 28716
rect 10551 28744 10563 28747
rect 10689 28747 10747 28753
rect 10689 28744 10701 28747
rect 10551 28716 10701 28744
rect 10551 28713 10563 28716
rect 10505 28707 10563 28713
rect 10689 28713 10701 28716
rect 10735 28713 10747 28747
rect 10689 28707 10747 28713
rect 11054 28704 11060 28756
rect 11112 28744 11118 28756
rect 11149 28747 11207 28753
rect 11149 28744 11161 28747
rect 11112 28716 11161 28744
rect 11112 28704 11118 28716
rect 11149 28713 11161 28716
rect 11195 28713 11207 28747
rect 11149 28707 11207 28713
rect 4246 28636 4252 28688
rect 4304 28676 4310 28688
rect 5350 28676 5356 28688
rect 4304 28648 5356 28676
rect 4304 28636 4310 28648
rect 5350 28636 5356 28648
rect 5408 28636 5414 28688
rect 7834 28676 7840 28688
rect 6932 28648 7840 28676
rect 6932 28620 6960 28648
rect 7834 28636 7840 28648
rect 7892 28636 7898 28688
rect 13354 28636 13360 28688
rect 13412 28676 13418 28688
rect 13633 28679 13691 28685
rect 13633 28676 13645 28679
rect 13412 28648 13645 28676
rect 13412 28636 13418 28648
rect 13633 28645 13645 28648
rect 13679 28676 13691 28679
rect 14093 28679 14151 28685
rect 14093 28676 14105 28679
rect 13679 28648 14105 28676
rect 13679 28645 13691 28648
rect 13633 28639 13691 28645
rect 14093 28645 14105 28648
rect 14139 28645 14151 28679
rect 14093 28639 14151 28645
rect 3970 28568 3976 28620
rect 4028 28608 4034 28620
rect 4028 28580 5212 28608
rect 4028 28568 4034 28580
rect 4062 28500 4068 28552
rect 4120 28500 4126 28552
rect 4246 28500 4252 28552
rect 4304 28500 4310 28552
rect 4338 28500 4344 28552
rect 4396 28540 4402 28552
rect 4706 28540 4712 28552
rect 4396 28512 4712 28540
rect 4396 28500 4402 28512
rect 4706 28500 4712 28512
rect 4764 28500 4770 28552
rect 5000 28549 5028 28580
rect 4985 28543 5043 28549
rect 4985 28509 4997 28543
rect 5031 28509 5043 28543
rect 4985 28503 5043 28509
rect 5077 28543 5135 28549
rect 5077 28509 5089 28543
rect 5123 28509 5135 28543
rect 5077 28503 5135 28509
rect 5092 28472 5120 28503
rect 4908 28444 5120 28472
rect 5184 28472 5212 28580
rect 6914 28568 6920 28620
rect 6972 28568 6978 28620
rect 7006 28568 7012 28620
rect 7064 28617 7070 28620
rect 7064 28611 7092 28617
rect 7080 28577 7092 28611
rect 7064 28571 7092 28577
rect 12713 28611 12771 28617
rect 12713 28577 12725 28611
rect 12759 28608 12771 28611
rect 13446 28608 13452 28620
rect 12759 28580 13452 28608
rect 12759 28577 12771 28580
rect 12713 28571 12771 28577
rect 7064 28568 7070 28571
rect 5721 28543 5779 28549
rect 5721 28509 5733 28543
rect 5767 28540 5779 28543
rect 6273 28543 6331 28549
rect 6273 28540 6285 28543
rect 5767 28512 6285 28540
rect 5767 28509 5779 28512
rect 5721 28503 5779 28509
rect 6273 28509 6285 28512
rect 6319 28509 6331 28543
rect 6273 28503 6331 28509
rect 6549 28543 6607 28549
rect 6549 28509 6561 28543
rect 6595 28540 6607 28543
rect 8202 28540 8208 28552
rect 6595 28512 8208 28540
rect 6595 28509 6607 28512
rect 6549 28503 6607 28509
rect 8202 28500 8208 28512
rect 8260 28500 8266 28552
rect 10229 28543 10287 28549
rect 10229 28509 10241 28543
rect 10275 28509 10287 28543
rect 10229 28503 10287 28509
rect 10321 28543 10379 28549
rect 10321 28509 10333 28543
rect 10367 28540 10379 28543
rect 10502 28540 10508 28552
rect 10367 28512 10508 28540
rect 10367 28509 10379 28512
rect 10321 28503 10379 28509
rect 5813 28475 5871 28481
rect 5813 28472 5825 28475
rect 5184 28444 5825 28472
rect 3694 28364 3700 28416
rect 3752 28404 3758 28416
rect 4157 28407 4215 28413
rect 4157 28404 4169 28407
rect 3752 28376 4169 28404
rect 3752 28364 3758 28376
rect 4157 28373 4169 28376
rect 4203 28373 4215 28407
rect 4157 28367 4215 28373
rect 4798 28364 4804 28416
rect 4856 28404 4862 28416
rect 4908 28413 4936 28444
rect 5813 28441 5825 28444
rect 5859 28441 5871 28475
rect 5813 28435 5871 28441
rect 5997 28475 6055 28481
rect 5997 28441 6009 28475
rect 6043 28441 6055 28475
rect 5997 28435 6055 28441
rect 6825 28475 6883 28481
rect 6825 28441 6837 28475
rect 6871 28472 6883 28475
rect 7926 28472 7932 28484
rect 6871 28444 7932 28472
rect 6871 28441 6883 28444
rect 6825 28435 6883 28441
rect 4893 28407 4951 28413
rect 4893 28404 4905 28407
rect 4856 28376 4905 28404
rect 4856 28364 4862 28376
rect 4893 28373 4905 28376
rect 4939 28404 4951 28407
rect 6012 28404 6040 28435
rect 7926 28432 7932 28444
rect 7984 28472 7990 28484
rect 8386 28472 8392 28484
rect 7984 28444 8392 28472
rect 7984 28432 7990 28444
rect 8386 28432 8392 28444
rect 8444 28432 8450 28484
rect 10244 28472 10272 28503
rect 10502 28500 10508 28512
rect 10560 28500 10566 28552
rect 10594 28500 10600 28552
rect 10652 28500 10658 28552
rect 10965 28543 11023 28549
rect 10965 28509 10977 28543
rect 11011 28540 11023 28543
rect 11514 28540 11520 28552
rect 11011 28512 11520 28540
rect 11011 28509 11023 28512
rect 10965 28503 11023 28509
rect 11514 28500 11520 28512
rect 11572 28500 11578 28552
rect 11793 28543 11851 28549
rect 11793 28509 11805 28543
rect 11839 28540 11851 28543
rect 12728 28540 12756 28571
rect 13446 28568 13452 28580
rect 13504 28568 13510 28620
rect 11839 28512 12434 28540
rect 11839 28509 11851 28512
rect 11793 28503 11851 28509
rect 12406 28484 12434 28512
rect 10686 28472 10692 28484
rect 10244 28444 10692 28472
rect 10686 28432 10692 28444
rect 10744 28432 10750 28484
rect 11422 28432 11428 28484
rect 11480 28472 11486 28484
rect 11882 28472 11888 28484
rect 11480 28444 11888 28472
rect 11480 28432 11486 28444
rect 11882 28432 11888 28444
rect 11940 28432 11946 28484
rect 12342 28432 12348 28484
rect 12400 28472 12434 28484
rect 12544 28512 12756 28540
rect 12544 28472 12572 28512
rect 13170 28500 13176 28552
rect 13228 28500 13234 28552
rect 13814 28500 13820 28552
rect 13872 28540 13878 28552
rect 14277 28543 14335 28549
rect 14277 28540 14289 28543
rect 13872 28512 14289 28540
rect 13872 28500 13878 28512
rect 14277 28509 14289 28512
rect 14323 28509 14335 28543
rect 14277 28503 14335 28509
rect 12400 28444 12572 28472
rect 12400 28432 12406 28444
rect 12618 28432 12624 28484
rect 12676 28472 12682 28484
rect 13081 28475 13139 28481
rect 13081 28472 13093 28475
rect 12676 28444 13093 28472
rect 12676 28432 12682 28444
rect 13081 28441 13093 28444
rect 13127 28472 13139 28475
rect 13538 28472 13544 28484
rect 13127 28444 13544 28472
rect 13127 28441 13139 28444
rect 13081 28435 13139 28441
rect 13538 28432 13544 28444
rect 13596 28432 13602 28484
rect 13633 28475 13691 28481
rect 13633 28441 13645 28475
rect 13679 28472 13691 28475
rect 13722 28472 13728 28484
rect 13679 28444 13728 28472
rect 13679 28441 13691 28444
rect 13633 28435 13691 28441
rect 13722 28432 13728 28444
rect 13780 28432 13786 28484
rect 4939 28376 6040 28404
rect 4939 28373 4951 28376
rect 4893 28367 4951 28373
rect 6270 28364 6276 28416
rect 6328 28404 6334 28416
rect 6365 28407 6423 28413
rect 6365 28404 6377 28407
rect 6328 28376 6377 28404
rect 6328 28364 6334 28376
rect 6365 28373 6377 28376
rect 6411 28373 6423 28407
rect 6365 28367 6423 28373
rect 12894 28364 12900 28416
rect 12952 28364 12958 28416
rect 1104 28314 16836 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 16836 28314
rect 1104 28240 16836 28262
rect 3053 28203 3111 28209
rect 3053 28169 3065 28203
rect 3099 28200 3111 28203
rect 3602 28200 3608 28212
rect 3099 28172 3608 28200
rect 3099 28169 3111 28172
rect 3053 28163 3111 28169
rect 3602 28160 3608 28172
rect 3660 28200 3666 28212
rect 4062 28200 4068 28212
rect 3660 28172 4068 28200
rect 3660 28160 3666 28172
rect 4062 28160 4068 28172
rect 4120 28160 4126 28212
rect 8662 28160 8668 28212
rect 8720 28200 8726 28212
rect 8757 28203 8815 28209
rect 8757 28200 8769 28203
rect 8720 28172 8769 28200
rect 8720 28160 8726 28172
rect 8757 28169 8769 28172
rect 8803 28169 8815 28203
rect 8757 28163 8815 28169
rect 10413 28203 10471 28209
rect 10413 28169 10425 28203
rect 10459 28200 10471 28203
rect 10594 28200 10600 28212
rect 10459 28172 10600 28200
rect 10459 28169 10471 28172
rect 10413 28163 10471 28169
rect 10594 28160 10600 28172
rect 10652 28160 10658 28212
rect 11514 28160 11520 28212
rect 11572 28160 11578 28212
rect 13722 28160 13728 28212
rect 13780 28200 13786 28212
rect 13817 28203 13875 28209
rect 13817 28200 13829 28203
rect 13780 28172 13829 28200
rect 13780 28160 13786 28172
rect 13817 28169 13829 28172
rect 13863 28169 13875 28203
rect 13817 28163 13875 28169
rect 4246 28132 4252 28144
rect 3988 28104 4252 28132
rect 3234 28024 3240 28076
rect 3292 28064 3298 28076
rect 3513 28067 3571 28073
rect 3513 28064 3525 28067
rect 3292 28036 3525 28064
rect 3292 28024 3298 28036
rect 3513 28033 3525 28036
rect 3559 28033 3571 28067
rect 3513 28027 3571 28033
rect 3697 28067 3755 28073
rect 3697 28033 3709 28067
rect 3743 28064 3755 28067
rect 3878 28064 3884 28076
rect 3743 28036 3884 28064
rect 3743 28033 3755 28036
rect 3697 28027 3755 28033
rect 3421 27999 3479 28005
rect 3421 27965 3433 27999
rect 3467 27996 3479 27999
rect 3712 27996 3740 28027
rect 3878 28024 3884 28036
rect 3936 28024 3942 28076
rect 3988 28073 4016 28104
rect 4246 28092 4252 28104
rect 4304 28092 4310 28144
rect 4709 28135 4767 28141
rect 4709 28101 4721 28135
rect 4755 28132 4767 28135
rect 5258 28132 5264 28144
rect 4755 28104 5264 28132
rect 4755 28101 4767 28104
rect 4709 28095 4767 28101
rect 5258 28092 5264 28104
rect 5316 28092 5322 28144
rect 6270 28132 6276 28144
rect 6104 28104 6276 28132
rect 3973 28067 4031 28073
rect 3973 28033 3985 28067
rect 4019 28033 4031 28067
rect 3973 28027 4031 28033
rect 3467 27968 3740 27996
rect 3467 27965 3479 27968
rect 3421 27959 3479 27965
rect 3786 27956 3792 28008
rect 3844 27996 3850 28008
rect 3988 27996 4016 28027
rect 4338 28024 4344 28076
rect 4396 28024 4402 28076
rect 6104 28073 6132 28104
rect 6270 28092 6276 28104
rect 6328 28092 6334 28144
rect 7742 28132 7748 28144
rect 6380 28104 7748 28132
rect 6380 28076 6408 28104
rect 7742 28092 7748 28104
rect 7800 28092 7806 28144
rect 8478 28132 8484 28144
rect 8128 28104 8484 28132
rect 4433 28067 4491 28073
rect 4433 28033 4445 28067
rect 4479 28064 4491 28067
rect 6089 28067 6147 28073
rect 6089 28064 6101 28067
rect 4479 28036 6101 28064
rect 4479 28033 4491 28036
rect 4433 28027 4491 28033
rect 6089 28033 6101 28036
rect 6135 28033 6147 28067
rect 6089 28027 6147 28033
rect 6181 28067 6239 28073
rect 6181 28033 6193 28067
rect 6227 28033 6239 28067
rect 6181 28027 6239 28033
rect 3844 27968 4016 27996
rect 3844 27956 3850 27968
rect 4614 27956 4620 28008
rect 4672 27996 4678 28008
rect 5445 27999 5503 28005
rect 5445 27996 5457 27999
rect 4672 27968 5457 27996
rect 4672 27956 4678 27968
rect 5445 27965 5457 27968
rect 5491 27965 5503 27999
rect 5445 27959 5503 27965
rect 5718 27956 5724 28008
rect 5776 27956 5782 28008
rect 3694 27888 3700 27940
rect 3752 27928 3758 27940
rect 6196 27928 6224 28027
rect 6362 28024 6368 28076
rect 6420 28024 6426 28076
rect 6730 28024 6736 28076
rect 6788 28064 6794 28076
rect 7101 28067 7159 28073
rect 7101 28064 7113 28067
rect 6788 28036 7113 28064
rect 6788 28024 6794 28036
rect 7101 28033 7113 28036
rect 7147 28033 7159 28067
rect 7101 28027 7159 28033
rect 7374 28024 7380 28076
rect 7432 28064 7438 28076
rect 8128 28073 8156 28104
rect 8478 28092 8484 28104
rect 8536 28092 8542 28144
rect 8573 28135 8631 28141
rect 8573 28101 8585 28135
rect 8619 28132 8631 28135
rect 8619 28104 10272 28132
rect 8619 28101 8631 28104
rect 8573 28095 8631 28101
rect 7561 28067 7619 28073
rect 7432 28036 7512 28064
rect 7432 28024 7438 28036
rect 3752 27900 6224 27928
rect 7484 27928 7512 28036
rect 7561 28033 7573 28067
rect 7607 28033 7619 28067
rect 7561 28027 7619 28033
rect 8113 28067 8171 28073
rect 8113 28033 8125 28067
rect 8159 28033 8171 28067
rect 8113 28027 8171 28033
rect 7576 27996 7604 28027
rect 8294 28024 8300 28076
rect 8352 28024 8358 28076
rect 9858 28024 9864 28076
rect 9916 28073 9922 28076
rect 9916 28027 9928 28073
rect 10244 28064 10272 28104
rect 10318 28092 10324 28144
rect 10376 28132 10382 28144
rect 12704 28135 12762 28141
rect 10376 28104 11836 28132
rect 10376 28092 10382 28104
rect 10410 28064 10416 28076
rect 10244 28036 10416 28064
rect 9916 28024 9922 28027
rect 10410 28024 10416 28036
rect 10468 28024 10474 28076
rect 10502 28024 10508 28076
rect 10560 28064 10566 28076
rect 10597 28067 10655 28073
rect 10597 28064 10609 28067
rect 10560 28036 10609 28064
rect 10560 28024 10566 28036
rect 10597 28033 10609 28036
rect 10643 28033 10655 28067
rect 10597 28027 10655 28033
rect 10686 28024 10692 28076
rect 10744 28024 10750 28076
rect 10980 28073 11008 28104
rect 10965 28067 11023 28073
rect 10965 28033 10977 28067
rect 11011 28033 11023 28067
rect 10965 28027 11023 28033
rect 11698 28024 11704 28076
rect 11756 28024 11762 28076
rect 8205 27999 8263 28005
rect 8205 27996 8217 27999
rect 7576 27968 8217 27996
rect 8205 27965 8217 27968
rect 8251 27965 8263 27999
rect 8205 27959 8263 27965
rect 10134 27956 10140 28008
rect 10192 27956 10198 28008
rect 10873 27999 10931 28005
rect 10873 27965 10885 27999
rect 10919 27996 10931 27999
rect 11716 27996 11744 28024
rect 10919 27968 11744 27996
rect 11808 27996 11836 28104
rect 12704 28101 12716 28135
rect 12750 28132 12762 28135
rect 12894 28132 12900 28144
rect 12750 28104 12900 28132
rect 12750 28101 12762 28104
rect 12704 28095 12762 28101
rect 12894 28092 12900 28104
rect 12952 28092 12958 28144
rect 11885 28067 11943 28073
rect 11885 28033 11897 28067
rect 11931 28064 11943 28067
rect 12066 28064 12072 28076
rect 11931 28036 12072 28064
rect 11931 28033 11943 28036
rect 11885 28027 11943 28033
rect 12066 28024 12072 28036
rect 12124 28024 12130 28076
rect 11977 27999 12035 28005
rect 11977 27996 11989 27999
rect 11808 27968 11989 27996
rect 10919 27965 10931 27968
rect 10873 27959 10931 27965
rect 11977 27965 11989 27968
rect 12023 27965 12035 27999
rect 11977 27959 12035 27965
rect 12342 27956 12348 28008
rect 12400 27996 12406 28008
rect 12437 27999 12495 28005
rect 12437 27996 12449 27999
rect 12400 27968 12449 27996
rect 12400 27956 12406 27968
rect 12437 27965 12449 27968
rect 12483 27965 12495 27999
rect 12437 27959 12495 27965
rect 8386 27928 8392 27940
rect 7484 27900 8392 27928
rect 3752 27888 3758 27900
rect 8386 27888 8392 27900
rect 8444 27888 8450 27940
rect 3878 27820 3884 27872
rect 3936 27820 3942 27872
rect 3970 27820 3976 27872
rect 4028 27860 4034 27872
rect 4065 27863 4123 27869
rect 4065 27860 4077 27863
rect 4028 27832 4077 27860
rect 4028 27820 4034 27832
rect 4065 27829 4077 27832
rect 4111 27829 4123 27863
rect 4065 27823 4123 27829
rect 4617 27863 4675 27869
rect 4617 27829 4629 27863
rect 4663 27860 4675 27863
rect 4706 27860 4712 27872
rect 4663 27832 4712 27860
rect 4663 27829 4675 27832
rect 4617 27823 4675 27829
rect 4706 27820 4712 27832
rect 4764 27820 4770 27872
rect 5905 27863 5963 27869
rect 5905 27829 5917 27863
rect 5951 27860 5963 27863
rect 6270 27860 6276 27872
rect 5951 27832 6276 27860
rect 5951 27829 5963 27832
rect 5905 27823 5963 27829
rect 6270 27820 6276 27832
rect 6328 27820 6334 27872
rect 6914 27820 6920 27872
rect 6972 27820 6978 27872
rect 7558 27820 7564 27872
rect 7616 27820 7622 27872
rect 7926 27820 7932 27872
rect 7984 27860 7990 27872
rect 8481 27863 8539 27869
rect 8481 27860 8493 27863
rect 7984 27832 8493 27860
rect 7984 27820 7990 27832
rect 8481 27829 8493 27832
rect 8527 27860 8539 27863
rect 9122 27860 9128 27872
rect 8527 27832 9128 27860
rect 8527 27829 8539 27832
rect 8481 27823 8539 27829
rect 9122 27820 9128 27832
rect 9180 27820 9186 27872
rect 1104 27770 16836 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 16836 27770
rect 1104 27696 16836 27718
rect 3605 27659 3663 27665
rect 3605 27625 3617 27659
rect 3651 27656 3663 27659
rect 3970 27656 3976 27668
rect 3651 27628 3976 27656
rect 3651 27625 3663 27628
rect 3605 27619 3663 27625
rect 3970 27616 3976 27628
rect 4028 27616 4034 27668
rect 5718 27656 5724 27668
rect 4080 27628 5724 27656
rect 4080 27600 4108 27628
rect 5718 27616 5724 27628
rect 5776 27616 5782 27668
rect 8205 27659 8263 27665
rect 8205 27625 8217 27659
rect 8251 27656 8263 27659
rect 8478 27656 8484 27668
rect 8251 27628 8484 27656
rect 8251 27625 8263 27628
rect 8205 27619 8263 27625
rect 8478 27616 8484 27628
rect 8536 27616 8542 27668
rect 8573 27659 8631 27665
rect 8573 27625 8585 27659
rect 8619 27656 8631 27659
rect 9490 27656 9496 27668
rect 8619 27628 9496 27656
rect 8619 27625 8631 27628
rect 8573 27619 8631 27625
rect 9490 27616 9496 27628
rect 9548 27616 9554 27668
rect 9858 27656 9864 27668
rect 9600 27628 9864 27656
rect 4062 27548 4068 27600
rect 4120 27548 4126 27600
rect 8294 27548 8300 27600
rect 8352 27588 8358 27600
rect 8757 27591 8815 27597
rect 8757 27588 8769 27591
rect 8352 27560 8769 27588
rect 8352 27548 8358 27560
rect 8757 27557 8769 27560
rect 8803 27588 8815 27591
rect 8938 27588 8944 27600
rect 8803 27560 8944 27588
rect 8803 27557 8815 27560
rect 8757 27551 8815 27557
rect 8938 27548 8944 27560
rect 8996 27548 9002 27600
rect 9600 27597 9628 27628
rect 9858 27616 9864 27628
rect 9916 27616 9922 27668
rect 9585 27591 9643 27597
rect 9048 27560 9536 27588
rect 2222 27480 2228 27532
rect 2280 27480 2286 27532
rect 6362 27520 6368 27532
rect 5828 27492 6368 27520
rect 2240 27452 2268 27480
rect 5828 27464 5856 27492
rect 6362 27480 6368 27492
rect 6420 27520 6426 27532
rect 6825 27523 6883 27529
rect 6825 27520 6837 27523
rect 6420 27492 6837 27520
rect 6420 27480 6426 27492
rect 6825 27489 6837 27492
rect 6871 27489 6883 27523
rect 8662 27520 8668 27532
rect 6825 27483 6883 27489
rect 8404 27492 8668 27520
rect 3050 27452 3056 27464
rect 2240 27424 3056 27452
rect 3050 27412 3056 27424
rect 3108 27452 3114 27464
rect 4614 27452 4620 27464
rect 3108 27424 4620 27452
rect 3108 27412 3114 27424
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 5629 27455 5687 27461
rect 5629 27421 5641 27455
rect 5675 27452 5687 27455
rect 5810 27452 5816 27464
rect 5675 27424 5816 27452
rect 5675 27421 5687 27424
rect 5629 27415 5687 27421
rect 5810 27412 5816 27424
rect 5868 27412 5874 27464
rect 6270 27412 6276 27464
rect 6328 27412 6334 27464
rect 2492 27387 2550 27393
rect 2492 27353 2504 27387
rect 2538 27384 2550 27387
rect 2682 27384 2688 27396
rect 2538 27356 2688 27384
rect 2538 27353 2550 27356
rect 2492 27347 2550 27353
rect 2682 27344 2688 27356
rect 2740 27344 2746 27396
rect 3510 27344 3516 27396
rect 3568 27384 3574 27396
rect 3973 27387 4031 27393
rect 3973 27384 3985 27387
rect 3568 27356 3985 27384
rect 3568 27344 3574 27356
rect 3973 27353 3985 27356
rect 4019 27353 4031 27387
rect 3973 27347 4031 27353
rect 5384 27387 5442 27393
rect 5384 27353 5396 27387
rect 5430 27384 5442 27387
rect 5721 27387 5779 27393
rect 5721 27384 5733 27387
rect 5430 27356 5733 27384
rect 5430 27353 5442 27356
rect 5384 27347 5442 27353
rect 5721 27353 5733 27356
rect 5767 27353 5779 27387
rect 5721 27347 5779 27353
rect 7092 27387 7150 27393
rect 7092 27353 7104 27387
rect 7138 27384 7150 27387
rect 7466 27384 7472 27396
rect 7138 27356 7472 27384
rect 7138 27353 7150 27356
rect 7092 27347 7150 27353
rect 7466 27344 7472 27356
rect 7524 27344 7530 27396
rect 8404 27393 8432 27492
rect 8662 27480 8668 27492
rect 8720 27480 8726 27532
rect 9048 27520 9076 27560
rect 8864 27492 9076 27520
rect 9508 27520 9536 27560
rect 9585 27557 9597 27591
rect 9631 27557 9643 27591
rect 9585 27551 9643 27557
rect 9674 27548 9680 27600
rect 9732 27548 9738 27600
rect 9508 27492 9996 27520
rect 8389 27387 8447 27393
rect 8389 27353 8401 27387
rect 8435 27353 8447 27387
rect 8389 27347 8447 27353
rect 8570 27344 8576 27396
rect 8628 27393 8634 27396
rect 8628 27387 8663 27393
rect 8651 27384 8663 27387
rect 8864 27384 8892 27492
rect 8941 27455 8999 27461
rect 8941 27421 8953 27455
rect 8987 27421 8999 27455
rect 8941 27415 8999 27421
rect 8651 27356 8892 27384
rect 8651 27353 8663 27356
rect 8628 27347 8663 27353
rect 8628 27344 8634 27347
rect 2958 27276 2964 27328
rect 3016 27316 3022 27328
rect 4062 27316 4068 27328
rect 3016 27288 4068 27316
rect 3016 27276 3022 27288
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 4249 27319 4307 27325
rect 4249 27285 4261 27319
rect 4295 27316 4307 27319
rect 4798 27316 4804 27328
rect 4295 27288 4804 27316
rect 4295 27285 4307 27288
rect 4249 27279 4307 27285
rect 4798 27276 4804 27288
rect 4856 27276 4862 27328
rect 8202 27276 8208 27328
rect 8260 27316 8266 27328
rect 8956 27316 8984 27415
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9217 27455 9275 27461
rect 9217 27452 9229 27455
rect 9180 27424 9229 27452
rect 9180 27412 9186 27424
rect 9217 27421 9229 27424
rect 9263 27452 9275 27455
rect 9306 27452 9312 27464
rect 9263 27424 9312 27452
rect 9263 27421 9275 27424
rect 9217 27415 9275 27421
rect 9306 27412 9312 27424
rect 9364 27412 9370 27464
rect 9968 27461 9996 27492
rect 10134 27480 10140 27532
rect 10192 27480 10198 27532
rect 10778 27520 10784 27532
rect 10244 27492 10784 27520
rect 9953 27455 10011 27461
rect 9953 27421 9965 27455
rect 9999 27452 10011 27455
rect 10244 27452 10272 27492
rect 10778 27480 10784 27492
rect 10836 27520 10842 27532
rect 11333 27523 11391 27529
rect 11333 27520 11345 27523
rect 10836 27492 11345 27520
rect 10836 27480 10842 27492
rect 11333 27489 11345 27492
rect 11379 27489 11391 27523
rect 11333 27483 11391 27489
rect 9999 27424 10272 27452
rect 9999 27421 10011 27424
rect 9953 27415 10011 27421
rect 11146 27412 11152 27464
rect 11204 27452 11210 27464
rect 11698 27452 11704 27464
rect 11204 27424 11704 27452
rect 11204 27412 11210 27424
rect 11698 27412 11704 27424
rect 11756 27452 11762 27464
rect 11885 27455 11943 27461
rect 11885 27452 11897 27455
rect 11756 27424 11897 27452
rect 11756 27412 11762 27424
rect 11885 27421 11897 27424
rect 11931 27421 11943 27455
rect 11885 27415 11943 27421
rect 9030 27344 9036 27396
rect 9088 27384 9094 27396
rect 9426 27387 9484 27393
rect 9426 27384 9438 27387
rect 9088 27356 9438 27384
rect 9088 27344 9094 27356
rect 9426 27353 9438 27356
rect 9472 27353 9484 27387
rect 9426 27347 9484 27353
rect 9582 27344 9588 27396
rect 9640 27384 9646 27396
rect 9677 27387 9735 27393
rect 9677 27384 9689 27387
rect 9640 27356 9689 27384
rect 9640 27344 9646 27356
rect 9677 27353 9689 27356
rect 9723 27353 9735 27387
rect 9677 27347 9735 27353
rect 10226 27344 10232 27396
rect 10284 27384 10290 27396
rect 10965 27387 11023 27393
rect 10965 27384 10977 27387
rect 10284 27356 10977 27384
rect 10284 27344 10290 27356
rect 10965 27353 10977 27356
rect 11011 27384 11023 27387
rect 11422 27384 11428 27396
rect 11011 27356 11428 27384
rect 11011 27353 11023 27356
rect 10965 27347 11023 27353
rect 11422 27344 11428 27356
rect 11480 27344 11486 27396
rect 11517 27387 11575 27393
rect 11517 27353 11529 27387
rect 11563 27384 11575 27387
rect 11790 27384 11796 27396
rect 11563 27356 11796 27384
rect 11563 27353 11575 27356
rect 11517 27347 11575 27353
rect 11790 27344 11796 27356
rect 11848 27384 11854 27396
rect 12250 27384 12256 27396
rect 11848 27356 12256 27384
rect 11848 27344 11854 27356
rect 12250 27344 12256 27356
rect 12308 27344 12314 27396
rect 8260 27288 8984 27316
rect 8260 27276 8266 27288
rect 9306 27276 9312 27328
rect 9364 27276 9370 27328
rect 9766 27276 9772 27328
rect 9824 27316 9830 27328
rect 9861 27319 9919 27325
rect 9861 27316 9873 27319
rect 9824 27288 9873 27316
rect 9824 27276 9830 27288
rect 9861 27285 9873 27288
rect 9907 27316 9919 27319
rect 10594 27316 10600 27328
rect 9907 27288 10600 27316
rect 9907 27285 9919 27288
rect 9861 27279 9919 27285
rect 10594 27276 10600 27288
rect 10652 27276 10658 27328
rect 11606 27276 11612 27328
rect 11664 27276 11670 27328
rect 11701 27319 11759 27325
rect 11701 27285 11713 27319
rect 11747 27316 11759 27319
rect 12066 27316 12072 27328
rect 11747 27288 12072 27316
rect 11747 27285 11759 27288
rect 11701 27279 11759 27285
rect 12066 27276 12072 27288
rect 12124 27276 12130 27328
rect 1104 27226 16836 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 16836 27226
rect 1104 27152 16836 27174
rect 2682 27072 2688 27124
rect 2740 27072 2746 27124
rect 2869 27115 2927 27121
rect 2869 27081 2881 27115
rect 2915 27112 2927 27115
rect 2958 27112 2964 27124
rect 2915 27084 2964 27112
rect 2915 27081 2927 27084
rect 2869 27075 2927 27081
rect 2958 27072 2964 27084
rect 3016 27072 3022 27124
rect 3973 27115 4031 27121
rect 3973 27081 3985 27115
rect 4019 27112 4031 27115
rect 4265 27115 4323 27121
rect 4265 27112 4277 27115
rect 4019 27084 4277 27112
rect 4019 27081 4031 27084
rect 3973 27075 4031 27081
rect 4265 27081 4277 27084
rect 4311 27081 4323 27115
rect 4265 27075 4323 27081
rect 4433 27115 4491 27121
rect 4433 27081 4445 27115
rect 4479 27081 4491 27115
rect 4433 27075 4491 27081
rect 3602 27044 3608 27056
rect 3252 27016 3608 27044
rect 3252 26985 3280 27016
rect 3602 27004 3608 27016
rect 3660 27004 3666 27056
rect 4062 27004 4068 27056
rect 4120 27004 4126 27056
rect 4448 27044 4476 27075
rect 7466 27072 7472 27124
rect 7524 27112 7530 27124
rect 7561 27115 7619 27121
rect 7561 27112 7573 27115
rect 7524 27084 7573 27112
rect 7524 27072 7530 27084
rect 7561 27081 7573 27084
rect 7607 27081 7619 27115
rect 7561 27075 7619 27081
rect 7834 27072 7840 27124
rect 7892 27072 7898 27124
rect 7926 27072 7932 27124
rect 7984 27072 7990 27124
rect 8297 27115 8355 27121
rect 8297 27081 8309 27115
rect 8343 27112 8355 27115
rect 8386 27112 8392 27124
rect 8343 27084 8392 27112
rect 8343 27081 8355 27084
rect 8297 27075 8355 27081
rect 8386 27072 8392 27084
rect 8444 27072 8450 27124
rect 8478 27072 8484 27124
rect 8536 27112 8542 27124
rect 8665 27115 8723 27121
rect 8665 27112 8677 27115
rect 8536 27084 8677 27112
rect 8536 27072 8542 27084
rect 8665 27081 8677 27084
rect 8711 27081 8723 27115
rect 8665 27075 8723 27081
rect 9030 27072 9036 27124
rect 9088 27072 9094 27124
rect 10410 27072 10416 27124
rect 10468 27112 10474 27124
rect 12618 27112 12624 27124
rect 10468 27084 12624 27112
rect 10468 27072 10474 27084
rect 12618 27072 12624 27084
rect 12676 27112 12682 27124
rect 12805 27115 12863 27121
rect 12805 27112 12817 27115
rect 12676 27084 12817 27112
rect 12676 27072 12682 27084
rect 12805 27081 12817 27084
rect 12851 27081 12863 27115
rect 12805 27075 12863 27081
rect 13081 27115 13139 27121
rect 13081 27081 13093 27115
rect 13127 27081 13139 27115
rect 13081 27075 13139 27081
rect 4770 27047 4828 27053
rect 4770 27044 4782 27047
rect 4448 27016 4782 27044
rect 4770 27013 4782 27016
rect 4816 27013 4828 27047
rect 4770 27007 4828 27013
rect 5534 27004 5540 27056
rect 5592 27044 5598 27056
rect 6549 27047 6607 27053
rect 6549 27044 6561 27047
rect 5592 27016 6561 27044
rect 5592 27004 5598 27016
rect 6549 27013 6561 27016
rect 6595 27044 6607 27047
rect 10226 27044 10232 27056
rect 6595 27016 10232 27044
rect 6595 27013 6607 27016
rect 6549 27007 6607 27013
rect 10226 27004 10232 27016
rect 10284 27004 10290 27056
rect 10686 27004 10692 27056
rect 10744 27044 10750 27056
rect 12434 27044 12440 27056
rect 10744 27016 12440 27044
rect 10744 27004 10750 27016
rect 12434 27004 12440 27016
rect 12492 27044 12498 27056
rect 12710 27044 12716 27056
rect 12492 27016 12716 27044
rect 12492 27004 12498 27016
rect 12710 27004 12716 27016
rect 12768 27004 12774 27056
rect 13096 27044 13124 27075
rect 14286 27047 14344 27053
rect 14286 27044 14298 27047
rect 13096 27016 14298 27044
rect 14286 27013 14298 27016
rect 14332 27013 14344 27047
rect 14286 27007 14344 27013
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 3237 26979 3295 26985
rect 1719 26948 2774 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 2746 26908 2774 26948
rect 3237 26945 3249 26979
rect 3283 26945 3295 26979
rect 3237 26939 3295 26945
rect 3786 26936 3792 26988
rect 3844 26976 3850 26988
rect 4525 26979 4583 26985
rect 3844 26948 4476 26976
rect 3844 26936 3850 26948
rect 4062 26908 4068 26920
rect 2746 26880 4068 26908
rect 4062 26868 4068 26880
rect 4120 26868 4126 26920
rect 3694 26800 3700 26852
rect 3752 26840 3758 26852
rect 3752 26812 4292 26840
rect 3752 26800 3758 26812
rect 842 26732 848 26784
rect 900 26772 906 26784
rect 1489 26775 1547 26781
rect 1489 26772 1501 26775
rect 900 26744 1501 26772
rect 900 26732 906 26744
rect 1489 26741 1501 26744
rect 1535 26741 1547 26775
rect 1489 26735 1547 26741
rect 2869 26775 2927 26781
rect 2869 26741 2881 26775
rect 2915 26772 2927 26775
rect 3878 26772 3884 26784
rect 2915 26744 3884 26772
rect 2915 26741 2927 26744
rect 2869 26735 2927 26741
rect 3878 26732 3884 26744
rect 3936 26732 3942 26784
rect 4264 26781 4292 26812
rect 4249 26775 4307 26781
rect 4249 26741 4261 26775
rect 4295 26741 4307 26775
rect 4448 26772 4476 26948
rect 4525 26945 4537 26979
rect 4571 26976 4583 26979
rect 4614 26976 4620 26988
rect 4571 26948 4620 26976
rect 4571 26945 4583 26948
rect 4525 26939 4583 26945
rect 4614 26936 4620 26948
rect 4672 26936 4678 26988
rect 7558 26936 7564 26988
rect 7616 26976 7622 26988
rect 7720 26979 7778 26985
rect 7720 26976 7732 26979
rect 7616 26948 7732 26976
rect 7616 26936 7622 26948
rect 7720 26945 7732 26948
rect 7766 26945 7778 26979
rect 7720 26939 7778 26945
rect 8478 26936 8484 26988
rect 8536 26936 8542 26988
rect 8573 26979 8631 26985
rect 8573 26945 8585 26979
rect 8619 26945 8631 26979
rect 8573 26939 8631 26945
rect 5810 26868 5816 26920
rect 5868 26908 5874 26920
rect 7285 26911 7343 26917
rect 7285 26908 7297 26911
rect 5868 26880 7297 26908
rect 5868 26868 5874 26880
rect 7285 26877 7297 26880
rect 7331 26877 7343 26911
rect 7285 26871 7343 26877
rect 8202 26868 8208 26920
rect 8260 26868 8266 26920
rect 8588 26908 8616 26939
rect 8662 26936 8668 26988
rect 8720 26976 8726 26988
rect 8849 26979 8907 26985
rect 8849 26976 8861 26979
rect 8720 26948 8861 26976
rect 8720 26936 8726 26948
rect 8849 26945 8861 26948
rect 8895 26945 8907 26979
rect 8849 26939 8907 26945
rect 8864 26908 8892 26939
rect 8938 26936 8944 26988
rect 8996 26936 9002 26988
rect 9125 26979 9183 26985
rect 9125 26945 9137 26979
rect 9171 26976 9183 26979
rect 9674 26976 9680 26988
rect 9171 26948 9680 26976
rect 9171 26945 9183 26948
rect 9125 26939 9183 26945
rect 9674 26936 9680 26948
rect 9732 26936 9738 26988
rect 10134 26936 10140 26988
rect 10192 26936 10198 26988
rect 11606 26936 11612 26988
rect 11664 26976 11670 26988
rect 11885 26979 11943 26985
rect 11885 26976 11897 26979
rect 11664 26948 11897 26976
rect 11664 26936 11670 26948
rect 11885 26945 11897 26948
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 12066 26936 12072 26988
rect 12124 26936 12130 26988
rect 13814 26976 13820 26988
rect 12176 26948 13820 26976
rect 9582 26908 9588 26920
rect 8588 26880 8708 26908
rect 8864 26880 9588 26908
rect 5905 26775 5963 26781
rect 5905 26772 5917 26775
rect 4448 26744 5917 26772
rect 4249 26735 4307 26741
rect 5905 26741 5917 26744
rect 5951 26741 5963 26775
rect 5905 26735 5963 26741
rect 8386 26732 8392 26784
rect 8444 26772 8450 26784
rect 8680 26772 8708 26880
rect 9582 26868 9588 26880
rect 9640 26868 9646 26920
rect 12176 26908 12204 26948
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 13906 26936 13912 26988
rect 13964 26976 13970 26988
rect 14553 26979 14611 26985
rect 14553 26976 14565 26979
rect 13964 26948 14565 26976
rect 13964 26936 13970 26948
rect 14553 26945 14565 26948
rect 14599 26945 14611 26979
rect 14553 26939 14611 26945
rect 9692 26880 12204 26908
rect 9122 26800 9128 26852
rect 9180 26840 9186 26852
rect 9692 26840 9720 26880
rect 12434 26868 12440 26920
rect 12492 26868 12498 26920
rect 12710 26868 12716 26920
rect 12768 26868 12774 26920
rect 12922 26911 12980 26917
rect 12922 26877 12934 26911
rect 12968 26908 12980 26911
rect 13078 26908 13084 26920
rect 12968 26880 13084 26908
rect 12968 26877 12980 26880
rect 12922 26871 12980 26877
rect 13078 26868 13084 26880
rect 13136 26868 13142 26920
rect 9180 26812 9720 26840
rect 9180 26800 9186 26812
rect 11698 26800 11704 26852
rect 11756 26840 11762 26852
rect 13173 26843 13231 26849
rect 13173 26840 13185 26843
rect 11756 26812 13185 26840
rect 11756 26800 11762 26812
rect 13173 26809 13185 26812
rect 13219 26809 13231 26843
rect 13173 26803 13231 26809
rect 9766 26772 9772 26784
rect 8444 26744 9772 26772
rect 8444 26732 8450 26744
rect 9766 26732 9772 26744
rect 9824 26732 9830 26784
rect 12069 26775 12127 26781
rect 12069 26741 12081 26775
rect 12115 26772 12127 26775
rect 12158 26772 12164 26784
rect 12115 26744 12164 26772
rect 12115 26741 12127 26744
rect 12069 26735 12127 26741
rect 12158 26732 12164 26744
rect 12216 26732 12222 26784
rect 1104 26682 16836 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 16836 26682
rect 1104 26608 16836 26630
rect 7006 26528 7012 26580
rect 7064 26568 7070 26580
rect 7834 26568 7840 26580
rect 7064 26540 7840 26568
rect 7064 26528 7070 26540
rect 7834 26528 7840 26540
rect 7892 26568 7898 26580
rect 9306 26568 9312 26580
rect 7892 26540 9312 26568
rect 7892 26528 7898 26540
rect 9306 26528 9312 26540
rect 9364 26528 9370 26580
rect 11606 26528 11612 26580
rect 11664 26528 11670 26580
rect 11698 26528 11704 26580
rect 11756 26568 11762 26580
rect 11793 26571 11851 26577
rect 11793 26568 11805 26571
rect 11756 26540 11805 26568
rect 11756 26528 11762 26540
rect 11793 26537 11805 26540
rect 11839 26537 11851 26571
rect 11793 26531 11851 26537
rect 5258 26460 5264 26512
rect 5316 26460 5322 26512
rect 11422 26500 11428 26512
rect 10336 26472 11428 26500
rect 10336 26444 10364 26472
rect 11422 26460 11428 26472
rect 11480 26460 11486 26512
rect 8202 26392 8208 26444
rect 8260 26432 8266 26444
rect 8941 26435 8999 26441
rect 8941 26432 8953 26435
rect 8260 26404 8953 26432
rect 8260 26392 8266 26404
rect 8941 26401 8953 26404
rect 8987 26432 8999 26435
rect 8987 26404 10088 26432
rect 8987 26401 8999 26404
rect 8941 26395 8999 26401
rect 4614 26324 4620 26376
rect 4672 26364 4678 26376
rect 4709 26367 4767 26373
rect 4709 26364 4721 26367
rect 4672 26336 4721 26364
rect 4672 26324 4678 26336
rect 4709 26333 4721 26336
rect 4755 26333 4767 26367
rect 4709 26327 4767 26333
rect 4798 26324 4804 26376
rect 4856 26364 4862 26376
rect 5537 26367 5595 26373
rect 5537 26364 5549 26367
rect 4856 26336 5549 26364
rect 4856 26324 4862 26336
rect 5537 26333 5549 26336
rect 5583 26333 5595 26367
rect 5537 26327 5595 26333
rect 5810 26324 5816 26376
rect 5868 26364 5874 26376
rect 6089 26367 6147 26373
rect 6089 26364 6101 26367
rect 5868 26336 6101 26364
rect 5868 26324 5874 26336
rect 6089 26333 6101 26336
rect 6135 26333 6147 26367
rect 6914 26364 6920 26376
rect 6089 26327 6147 26333
rect 6196 26336 6920 26364
rect 5261 26299 5319 26305
rect 5261 26265 5273 26299
rect 5307 26296 5319 26299
rect 5350 26296 5356 26308
rect 5307 26268 5356 26296
rect 5307 26265 5319 26268
rect 5261 26259 5319 26265
rect 5350 26256 5356 26268
rect 5408 26256 5414 26308
rect 5445 26299 5503 26305
rect 5445 26265 5457 26299
rect 5491 26296 5503 26299
rect 6196 26296 6224 26336
rect 6914 26324 6920 26336
rect 6972 26324 6978 26376
rect 9122 26324 9128 26376
rect 9180 26324 9186 26376
rect 10060 26373 10088 26404
rect 10318 26392 10324 26444
rect 10376 26392 10382 26444
rect 10410 26392 10416 26444
rect 10468 26392 10474 26444
rect 10045 26367 10103 26373
rect 10045 26333 10057 26367
rect 10091 26364 10103 26367
rect 10686 26364 10692 26376
rect 10091 26336 10692 26364
rect 10091 26333 10103 26336
rect 10045 26327 10103 26333
rect 10686 26324 10692 26336
rect 10744 26324 10750 26376
rect 10778 26324 10784 26376
rect 10836 26324 10842 26376
rect 10965 26367 11023 26373
rect 10965 26333 10977 26367
rect 11011 26333 11023 26367
rect 10965 26327 11023 26333
rect 6362 26305 6368 26308
rect 5491 26268 6224 26296
rect 5491 26265 5503 26268
rect 5445 26259 5503 26265
rect 6356 26259 6368 26305
rect 4246 26188 4252 26240
rect 4304 26228 4310 26240
rect 5460 26228 5488 26259
rect 6362 26256 6368 26259
rect 6420 26256 6426 26308
rect 10530 26299 10588 26305
rect 10530 26265 10542 26299
rect 10576 26296 10588 26299
rect 10873 26299 10931 26305
rect 10873 26296 10885 26299
rect 10576 26268 10885 26296
rect 10576 26265 10588 26268
rect 10530 26259 10588 26265
rect 10873 26265 10885 26268
rect 10919 26265 10931 26299
rect 10980 26296 11008 26327
rect 11146 26324 11152 26376
rect 11204 26324 11210 26376
rect 11333 26367 11391 26373
rect 11333 26333 11345 26367
rect 11379 26364 11391 26367
rect 11624 26364 11652 26528
rect 11808 26432 11836 26531
rect 12066 26528 12072 26580
rect 12124 26528 12130 26580
rect 12250 26528 12256 26580
rect 12308 26568 12314 26580
rect 12308 26540 12434 26568
rect 12308 26528 12314 26540
rect 12406 26432 12434 26540
rect 13078 26528 13084 26580
rect 13136 26568 13142 26580
rect 13173 26571 13231 26577
rect 13173 26568 13185 26571
rect 13136 26540 13185 26568
rect 13136 26528 13142 26540
rect 13173 26537 13185 26540
rect 13219 26537 13231 26571
rect 13173 26531 13231 26537
rect 12713 26435 12771 26441
rect 12713 26432 12725 26435
rect 11808 26404 12204 26432
rect 11379 26336 11652 26364
rect 12176 26364 12204 26404
rect 12360 26404 12725 26432
rect 12360 26373 12388 26404
rect 12713 26401 12725 26404
rect 12759 26401 12771 26435
rect 12713 26395 12771 26401
rect 12253 26367 12311 26373
rect 12253 26364 12265 26367
rect 12176 26336 12265 26364
rect 11379 26333 11391 26336
rect 11333 26327 11391 26333
rect 12253 26333 12265 26336
rect 12299 26333 12311 26367
rect 12253 26327 12311 26333
rect 12345 26367 12403 26373
rect 12345 26333 12357 26367
rect 12391 26333 12403 26367
rect 12345 26327 12403 26333
rect 12805 26367 12863 26373
rect 12805 26333 12817 26367
rect 12851 26333 12863 26367
rect 12805 26327 12863 26333
rect 11790 26305 11796 26308
rect 11241 26299 11299 26305
rect 11241 26296 11253 26299
rect 10980 26268 11253 26296
rect 10873 26259 10931 26265
rect 11241 26265 11253 26268
rect 11287 26265 11299 26299
rect 11241 26259 11299 26265
rect 11777 26299 11796 26305
rect 11777 26265 11789 26299
rect 11777 26259 11796 26265
rect 11790 26256 11796 26259
rect 11848 26256 11854 26308
rect 11974 26256 11980 26308
rect 12032 26296 12038 26308
rect 12069 26299 12127 26305
rect 12069 26296 12081 26299
rect 12032 26268 12081 26296
rect 12032 26256 12038 26268
rect 12069 26265 12081 26268
rect 12115 26265 12127 26299
rect 12268 26296 12296 26327
rect 12820 26296 12848 26327
rect 12268 26268 12848 26296
rect 12069 26259 12127 26265
rect 4304 26200 5488 26228
rect 7469 26231 7527 26237
rect 4304 26188 4310 26200
rect 7469 26197 7481 26231
rect 7515 26228 7527 26231
rect 7926 26228 7932 26240
rect 7515 26200 7932 26228
rect 7515 26197 7527 26200
rect 7469 26191 7527 26197
rect 7926 26188 7932 26200
rect 7984 26188 7990 26240
rect 10686 26188 10692 26240
rect 10744 26188 10750 26240
rect 1104 26138 16836 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 16836 26138
rect 1104 26064 16836 26086
rect 3510 25984 3516 26036
rect 3568 26024 3574 26036
rect 3881 26027 3939 26033
rect 3881 26024 3893 26027
rect 3568 25996 3893 26024
rect 3568 25984 3574 25996
rect 3881 25993 3893 25996
rect 3927 25993 3939 26027
rect 3881 25987 3939 25993
rect 4065 26027 4123 26033
rect 4065 25993 4077 26027
rect 4111 26024 4123 26027
rect 4706 26024 4712 26036
rect 4111 25996 4712 26024
rect 4111 25993 4123 25996
rect 4065 25987 4123 25993
rect 4706 25984 4712 25996
rect 4764 25984 4770 26036
rect 6549 26027 6607 26033
rect 6549 25993 6561 26027
rect 6595 26024 6607 26027
rect 9217 26027 9275 26033
rect 6595 25996 8432 26024
rect 6595 25993 6607 25996
rect 6549 25987 6607 25993
rect 6365 25959 6423 25965
rect 6365 25925 6377 25959
rect 6411 25956 6423 25959
rect 8202 25956 8208 25968
rect 6411 25928 8208 25956
rect 6411 25925 6423 25928
rect 6365 25919 6423 25925
rect 8202 25916 8208 25928
rect 8260 25916 8266 25968
rect 8404 25956 8432 25996
rect 9217 25993 9229 26027
rect 9263 26024 9275 26027
rect 9306 26024 9312 26036
rect 9263 25996 9312 26024
rect 9263 25993 9275 25996
rect 9217 25987 9275 25993
rect 9306 25984 9312 25996
rect 9364 25984 9370 26036
rect 11146 25984 11152 26036
rect 11204 26024 11210 26036
rect 11333 26027 11391 26033
rect 11333 26024 11345 26027
rect 11204 25996 11345 26024
rect 11204 25984 11210 25996
rect 11333 25993 11345 25996
rect 11379 25993 11391 26027
rect 11333 25987 11391 25993
rect 11974 25984 11980 26036
rect 12032 26024 12038 26036
rect 13081 26027 13139 26033
rect 13081 26024 13093 26027
rect 12032 25996 13093 26024
rect 12032 25984 12038 25996
rect 13081 25993 13093 25996
rect 13127 25993 13139 26027
rect 13081 25987 13139 25993
rect 9030 25956 9036 25968
rect 8404 25928 9036 25956
rect 9030 25916 9036 25928
rect 9088 25956 9094 25968
rect 9125 25959 9183 25965
rect 9125 25956 9137 25959
rect 9088 25928 9137 25956
rect 9088 25916 9094 25928
rect 9125 25925 9137 25928
rect 9171 25925 9183 25959
rect 9125 25919 9183 25925
rect 10220 25959 10278 25965
rect 10220 25925 10232 25959
rect 10266 25956 10278 25959
rect 10686 25956 10692 25968
rect 10266 25928 10692 25956
rect 10266 25925 10278 25928
rect 10220 25919 10278 25925
rect 10686 25916 10692 25928
rect 10744 25916 10750 25968
rect 12342 25956 12348 25968
rect 11716 25928 12348 25956
rect 6641 25891 6699 25897
rect 6641 25857 6653 25891
rect 6687 25888 6699 25891
rect 7006 25888 7012 25900
rect 6687 25860 7012 25888
rect 6687 25857 6699 25860
rect 6641 25851 6699 25857
rect 7006 25848 7012 25860
rect 7064 25848 7070 25900
rect 7745 25891 7803 25897
rect 7745 25857 7757 25891
rect 7791 25888 7803 25891
rect 7834 25888 7840 25900
rect 7791 25860 7840 25888
rect 7791 25857 7803 25860
rect 7745 25851 7803 25857
rect 7834 25848 7840 25860
rect 7892 25848 7898 25900
rect 7926 25848 7932 25900
rect 7984 25848 7990 25900
rect 8386 25848 8392 25900
rect 8444 25848 8450 25900
rect 9334 25891 9392 25897
rect 9334 25888 9346 25891
rect 8772 25860 9346 25888
rect 4433 25823 4491 25829
rect 4433 25789 4445 25823
rect 4479 25820 4491 25823
rect 4614 25820 4620 25832
rect 4479 25792 4620 25820
rect 4479 25789 4491 25792
rect 4433 25783 4491 25789
rect 4614 25780 4620 25792
rect 4672 25780 4678 25832
rect 5626 25780 5632 25832
rect 5684 25780 5690 25832
rect 7653 25823 7711 25829
rect 7653 25789 7665 25823
rect 7699 25820 7711 25823
rect 7944 25820 7972 25848
rect 7699 25792 7972 25820
rect 7699 25789 7711 25792
rect 7653 25783 7711 25789
rect 8478 25780 8484 25832
rect 8536 25780 8542 25832
rect 8772 25829 8800 25860
rect 9334 25857 9346 25860
rect 9380 25857 9392 25891
rect 9334 25851 9392 25857
rect 9953 25891 10011 25897
rect 9953 25857 9965 25891
rect 9999 25888 10011 25891
rect 10042 25888 10048 25900
rect 9999 25860 10048 25888
rect 9999 25857 10011 25860
rect 9953 25851 10011 25857
rect 10042 25848 10048 25860
rect 10100 25848 10106 25900
rect 11716 25897 11744 25928
rect 12342 25916 12348 25928
rect 12400 25956 12406 25968
rect 13262 25956 13268 25968
rect 12400 25928 13268 25956
rect 12400 25916 12406 25928
rect 13262 25916 13268 25928
rect 13320 25956 13326 25968
rect 13722 25956 13728 25968
rect 13320 25928 13728 25956
rect 13320 25916 13326 25928
rect 13722 25916 13728 25928
rect 13780 25916 13786 25968
rect 11974 25897 11980 25900
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 11968 25851 11980 25897
rect 11974 25848 11980 25851
rect 12032 25848 12038 25900
rect 8757 25823 8815 25829
rect 8757 25789 8769 25823
rect 8803 25789 8815 25823
rect 8757 25783 8815 25789
rect 8849 25823 8907 25829
rect 8849 25789 8861 25823
rect 8895 25789 8907 25823
rect 8849 25783 8907 25789
rect 6362 25712 6368 25764
rect 6420 25712 6426 25764
rect 8202 25712 8208 25764
rect 8260 25752 8266 25764
rect 8864 25752 8892 25783
rect 8260 25724 8892 25752
rect 8260 25712 8266 25724
rect 4065 25687 4123 25693
rect 4065 25653 4077 25687
rect 4111 25684 4123 25687
rect 4246 25684 4252 25696
rect 4111 25656 4252 25684
rect 4111 25653 4123 25656
rect 4065 25647 4123 25653
rect 4246 25644 4252 25656
rect 4304 25644 4310 25696
rect 4706 25644 4712 25696
rect 4764 25684 4770 25696
rect 5261 25687 5319 25693
rect 5261 25684 5273 25687
rect 4764 25656 5273 25684
rect 4764 25644 4770 25656
rect 5261 25653 5273 25656
rect 5307 25684 5319 25687
rect 5350 25684 5356 25696
rect 5307 25656 5356 25684
rect 5307 25653 5319 25656
rect 5261 25647 5319 25653
rect 5350 25644 5356 25656
rect 5408 25644 5414 25696
rect 5994 25644 6000 25696
rect 6052 25684 6058 25696
rect 6181 25687 6239 25693
rect 6181 25684 6193 25687
rect 6052 25656 6193 25684
rect 6052 25644 6058 25656
rect 6181 25653 6193 25656
rect 6227 25653 6239 25687
rect 6181 25647 6239 25653
rect 7006 25644 7012 25696
rect 7064 25644 7070 25696
rect 7558 25644 7564 25696
rect 7616 25684 7622 25696
rect 7837 25687 7895 25693
rect 7837 25684 7849 25687
rect 7616 25656 7849 25684
rect 7616 25644 7622 25656
rect 7837 25653 7849 25656
rect 7883 25653 7895 25687
rect 7837 25647 7895 25653
rect 9490 25644 9496 25696
rect 9548 25644 9554 25696
rect 1104 25594 16836 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 16836 25594
rect 1104 25520 16836 25542
rect 10594 25440 10600 25492
rect 10652 25440 10658 25492
rect 11974 25440 11980 25492
rect 12032 25480 12038 25492
rect 12161 25483 12219 25489
rect 12161 25480 12173 25483
rect 12032 25452 12173 25480
rect 12032 25440 12038 25452
rect 12161 25449 12173 25452
rect 12207 25449 12219 25483
rect 12161 25443 12219 25449
rect 6914 25372 6920 25424
rect 6972 25412 6978 25424
rect 7837 25415 7895 25421
rect 7837 25412 7849 25415
rect 6972 25384 7849 25412
rect 6972 25372 6978 25384
rect 7837 25381 7849 25384
rect 7883 25381 7895 25415
rect 12434 25412 12440 25424
rect 7837 25375 7895 25381
rect 11532 25384 12440 25412
rect 5258 25344 5264 25356
rect 5092 25316 5264 25344
rect 4913 25279 4971 25285
rect 4913 25245 4925 25279
rect 4959 25276 4971 25279
rect 5092 25276 5120 25316
rect 5258 25304 5264 25316
rect 5316 25304 5322 25356
rect 7653 25347 7711 25353
rect 7653 25344 7665 25347
rect 7392 25316 7665 25344
rect 4959 25248 5120 25276
rect 5169 25279 5227 25285
rect 4959 25245 4971 25248
rect 4913 25239 4971 25245
rect 5169 25245 5181 25279
rect 5215 25276 5227 25279
rect 5721 25279 5779 25285
rect 5721 25276 5733 25279
rect 5215 25248 5733 25276
rect 5215 25245 5227 25248
rect 5169 25239 5227 25245
rect 5721 25245 5733 25248
rect 5767 25276 5779 25279
rect 5810 25276 5816 25288
rect 5767 25248 5816 25276
rect 5767 25245 5779 25248
rect 5721 25239 5779 25245
rect 5810 25236 5816 25248
rect 5868 25236 5874 25288
rect 5994 25285 6000 25288
rect 5988 25276 6000 25285
rect 5955 25248 6000 25276
rect 5988 25239 6000 25248
rect 5994 25236 6000 25239
rect 6052 25236 6058 25288
rect 6546 25276 6552 25288
rect 6196 25248 6552 25276
rect 4154 25168 4160 25220
rect 4212 25208 4218 25220
rect 5445 25211 5503 25217
rect 5445 25208 5457 25211
rect 4212 25180 5457 25208
rect 4212 25168 4218 25180
rect 5445 25177 5457 25180
rect 5491 25177 5503 25211
rect 5445 25171 5503 25177
rect 5629 25211 5687 25217
rect 5629 25177 5641 25211
rect 5675 25208 5687 25211
rect 6196 25208 6224 25248
rect 6546 25236 6552 25248
rect 6604 25236 6610 25288
rect 7098 25236 7104 25288
rect 7156 25276 7162 25288
rect 7285 25279 7343 25285
rect 7285 25276 7297 25279
rect 7156 25248 7297 25276
rect 7156 25236 7162 25248
rect 7285 25245 7297 25248
rect 7331 25245 7343 25279
rect 7285 25239 7343 25245
rect 7193 25211 7251 25217
rect 7193 25208 7205 25211
rect 5675 25180 6224 25208
rect 6288 25180 7205 25208
rect 5675 25177 5687 25180
rect 5629 25171 5687 25177
rect 3786 25100 3792 25152
rect 3844 25100 3850 25152
rect 5261 25143 5319 25149
rect 5261 25109 5273 25143
rect 5307 25140 5319 25143
rect 6288 25140 6316 25180
rect 7193 25177 7205 25180
rect 7239 25177 7251 25211
rect 7193 25171 7251 25177
rect 5307 25112 6316 25140
rect 5307 25109 5319 25112
rect 5261 25103 5319 25109
rect 6546 25100 6552 25152
rect 6604 25140 6610 25152
rect 7101 25143 7159 25149
rect 7101 25140 7113 25143
rect 6604 25112 7113 25140
rect 6604 25100 6610 25112
rect 7101 25109 7113 25112
rect 7147 25140 7159 25143
rect 7392 25140 7420 25316
rect 7653 25313 7665 25316
rect 7699 25313 7711 25347
rect 7653 25307 7711 25313
rect 7558 25236 7564 25288
rect 7616 25236 7622 25288
rect 7668 25276 7696 25307
rect 7926 25304 7932 25356
rect 7984 25344 7990 25356
rect 11532 25353 11560 25384
rect 12434 25372 12440 25384
rect 12492 25372 12498 25424
rect 11517 25347 11575 25353
rect 7984 25316 9168 25344
rect 7984 25304 7990 25316
rect 8294 25276 8300 25288
rect 7668 25248 8300 25276
rect 8294 25236 8300 25248
rect 8352 25276 8358 25288
rect 9140 25285 9168 25316
rect 11517 25313 11529 25347
rect 11563 25313 11575 25347
rect 11517 25307 11575 25313
rect 12002 25347 12060 25353
rect 12002 25313 12014 25347
rect 12048 25344 12060 25347
rect 12158 25344 12164 25356
rect 12048 25316 12164 25344
rect 12048 25313 12060 25316
rect 12002 25307 12060 25313
rect 12158 25304 12164 25316
rect 12216 25304 12222 25356
rect 8481 25279 8539 25285
rect 8481 25276 8493 25279
rect 8352 25248 8493 25276
rect 8352 25236 8358 25248
rect 8481 25245 8493 25248
rect 8527 25276 8539 25279
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8527 25248 8953 25276
rect 8527 25245 8539 25248
rect 8481 25239 8539 25245
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9125 25279 9183 25285
rect 9125 25245 9137 25279
rect 9171 25245 9183 25279
rect 9125 25239 9183 25245
rect 9217 25279 9275 25285
rect 9217 25245 9229 25279
rect 9263 25276 9275 25279
rect 10042 25276 10048 25288
rect 9263 25248 10048 25276
rect 9263 25245 9275 25248
rect 9217 25239 9275 25245
rect 10042 25236 10048 25248
rect 10100 25236 10106 25288
rect 11422 25236 11428 25288
rect 11480 25276 11486 25288
rect 11793 25279 11851 25285
rect 11793 25276 11805 25279
rect 11480 25248 11805 25276
rect 11480 25236 11486 25248
rect 11793 25245 11805 25248
rect 11839 25245 11851 25279
rect 11793 25239 11851 25245
rect 7466 25168 7472 25220
rect 7524 25208 7530 25220
rect 9490 25217 9496 25220
rect 7929 25211 7987 25217
rect 7929 25208 7941 25211
rect 7524 25180 7941 25208
rect 7524 25168 7530 25180
rect 7929 25177 7941 25180
rect 7975 25177 7987 25211
rect 9484 25208 9496 25217
rect 9451 25180 9496 25208
rect 7929 25171 7987 25177
rect 9484 25171 9496 25180
rect 9490 25168 9496 25171
rect 9548 25168 9554 25220
rect 7147 25112 7420 25140
rect 7147 25109 7159 25112
rect 7101 25103 7159 25109
rect 7650 25100 7656 25152
rect 7708 25140 7714 25152
rect 8386 25140 8392 25152
rect 7708 25112 8392 25140
rect 7708 25100 7714 25112
rect 8386 25100 8392 25112
rect 8444 25140 8450 25152
rect 8941 25143 8999 25149
rect 8941 25140 8953 25143
rect 8444 25112 8953 25140
rect 8444 25100 8450 25112
rect 8941 25109 8953 25112
rect 8987 25109 8999 25143
rect 8941 25103 8999 25109
rect 9306 25100 9312 25152
rect 9364 25140 9370 25152
rect 11885 25143 11943 25149
rect 11885 25140 11897 25143
rect 9364 25112 11897 25140
rect 9364 25100 9370 25112
rect 11885 25109 11897 25112
rect 11931 25109 11943 25143
rect 11885 25103 11943 25109
rect 1104 25050 16836 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 16836 25050
rect 1104 24976 16836 24998
rect 4154 24896 4160 24948
rect 4212 24896 4218 24948
rect 5626 24896 5632 24948
rect 5684 24896 5690 24948
rect 7929 24939 7987 24945
rect 7929 24905 7941 24939
rect 7975 24905 7987 24939
rect 7929 24899 7987 24905
rect 7558 24868 7564 24880
rect 5920 24840 7564 24868
rect 5281 24803 5339 24809
rect 5281 24769 5293 24803
rect 5327 24800 5339 24803
rect 5442 24800 5448 24812
rect 5327 24772 5448 24800
rect 5327 24769 5339 24772
rect 5281 24763 5339 24769
rect 5442 24760 5448 24772
rect 5500 24760 5506 24812
rect 5920 24744 5948 24840
rect 7558 24828 7564 24840
rect 7616 24828 7622 24880
rect 5997 24803 6055 24809
rect 5997 24769 6009 24803
rect 6043 24800 6055 24803
rect 7466 24800 7472 24812
rect 6043 24772 7472 24800
rect 6043 24769 6055 24772
rect 5997 24763 6055 24769
rect 7466 24760 7472 24772
rect 7524 24760 7530 24812
rect 7650 24760 7656 24812
rect 7708 24760 7714 24812
rect 7944 24800 7972 24899
rect 8277 24803 8335 24809
rect 8277 24800 8289 24803
rect 7944 24772 8289 24800
rect 8277 24769 8289 24772
rect 8323 24769 8335 24803
rect 8277 24763 8335 24769
rect 5537 24735 5595 24741
rect 5537 24701 5549 24735
rect 5583 24701 5595 24735
rect 5537 24695 5595 24701
rect 5552 24664 5580 24695
rect 5902 24692 5908 24744
rect 5960 24692 5966 24744
rect 6454 24692 6460 24744
rect 6512 24732 6518 24744
rect 6549 24735 6607 24741
rect 6549 24732 6561 24735
rect 6512 24704 6561 24732
rect 6512 24692 6518 24704
rect 6549 24701 6561 24704
rect 6595 24701 6607 24735
rect 6549 24695 6607 24701
rect 6822 24692 6828 24744
rect 6880 24732 6886 24744
rect 7282 24732 7288 24744
rect 6880 24704 7288 24732
rect 6880 24692 6886 24704
rect 7282 24692 7288 24704
rect 7340 24692 7346 24744
rect 7377 24735 7435 24741
rect 7377 24701 7389 24735
rect 7423 24732 7435 24735
rect 7558 24732 7564 24744
rect 7423 24704 7564 24732
rect 7423 24701 7435 24704
rect 7377 24695 7435 24701
rect 7558 24692 7564 24704
rect 7616 24692 7622 24744
rect 7742 24692 7748 24744
rect 7800 24692 7806 24744
rect 8021 24735 8079 24741
rect 8021 24701 8033 24735
rect 8067 24701 8079 24735
rect 8021 24695 8079 24701
rect 5810 24664 5816 24676
rect 5552 24636 5816 24664
rect 5810 24624 5816 24636
rect 5868 24664 5874 24676
rect 8036 24664 8064 24695
rect 5868 24636 8064 24664
rect 5868 24624 5874 24636
rect 7392 24608 7420 24636
rect 9122 24624 9128 24676
rect 9180 24664 9186 24676
rect 9401 24667 9459 24673
rect 9401 24664 9413 24667
rect 9180 24636 9413 24664
rect 9180 24624 9186 24636
rect 9401 24633 9413 24636
rect 9447 24633 9459 24667
rect 9401 24627 9459 24633
rect 6362 24556 6368 24608
rect 6420 24596 6426 24608
rect 6822 24596 6828 24608
rect 6420 24568 6828 24596
rect 6420 24556 6426 24568
rect 6822 24556 6828 24568
rect 6880 24556 6886 24608
rect 7190 24556 7196 24608
rect 7248 24556 7254 24608
rect 7374 24556 7380 24608
rect 7432 24556 7438 24608
rect 7558 24556 7564 24608
rect 7616 24596 7622 24608
rect 8202 24596 8208 24608
rect 7616 24568 8208 24596
rect 7616 24556 7622 24568
rect 8202 24556 8208 24568
rect 8260 24556 8266 24608
rect 1104 24506 16836 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 16836 24506
rect 1104 24432 16836 24454
rect 5442 24352 5448 24404
rect 5500 24352 5506 24404
rect 6454 24352 6460 24404
rect 6512 24352 6518 24404
rect 6549 24395 6607 24401
rect 6549 24361 6561 24395
rect 6595 24392 6607 24395
rect 7006 24392 7012 24404
rect 6595 24364 7012 24392
rect 6595 24361 6607 24364
rect 6549 24355 6607 24361
rect 7006 24352 7012 24364
rect 7064 24352 7070 24404
rect 7466 24352 7472 24404
rect 7524 24392 7530 24404
rect 7524 24364 7687 24392
rect 7524 24352 7530 24364
rect 5721 24327 5779 24333
rect 5721 24293 5733 24327
rect 5767 24324 5779 24327
rect 5902 24324 5908 24336
rect 5767 24296 5908 24324
rect 5767 24293 5779 24296
rect 5721 24287 5779 24293
rect 5902 24284 5908 24296
rect 5960 24284 5966 24336
rect 6730 24284 6736 24336
rect 6788 24284 6794 24336
rect 7659 24324 7687 24364
rect 7834 24352 7840 24404
rect 7892 24392 7898 24404
rect 8110 24392 8116 24404
rect 7892 24364 8116 24392
rect 7892 24352 7898 24364
rect 8110 24352 8116 24364
rect 8168 24392 8174 24404
rect 8205 24395 8263 24401
rect 8205 24392 8217 24395
rect 8168 24364 8217 24392
rect 8168 24352 8174 24364
rect 8205 24361 8217 24364
rect 8251 24361 8263 24395
rect 8205 24355 8263 24361
rect 9217 24327 9275 24333
rect 9217 24324 9229 24327
rect 7659 24296 9229 24324
rect 9217 24293 9229 24296
rect 9263 24293 9275 24327
rect 9217 24287 9275 24293
rect 3786 24216 3792 24268
rect 3844 24256 3850 24268
rect 4065 24259 4123 24265
rect 4065 24256 4077 24259
rect 3844 24228 4077 24256
rect 3844 24216 3850 24228
rect 4065 24225 4077 24228
rect 4111 24225 4123 24259
rect 4065 24219 4123 24225
rect 5810 24216 5816 24268
rect 5868 24216 5874 24268
rect 6748 24256 6776 24284
rect 6104 24228 6776 24256
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24157 5687 24191
rect 5629 24151 5687 24157
rect 5905 24191 5963 24197
rect 5905 24157 5917 24191
rect 5951 24188 5963 24191
rect 5994 24188 6000 24200
rect 5951 24160 6000 24188
rect 5951 24157 5963 24160
rect 5905 24151 5963 24157
rect 5644 24120 5672 24151
rect 5994 24148 6000 24160
rect 6052 24148 6058 24200
rect 6104 24197 6132 24228
rect 8294 24216 8300 24268
rect 8352 24216 8358 24268
rect 11609 24259 11667 24265
rect 11609 24225 11621 24259
rect 11655 24256 11667 24259
rect 11701 24259 11759 24265
rect 11701 24256 11713 24259
rect 11655 24228 11713 24256
rect 11655 24225 11667 24228
rect 11609 24219 11667 24225
rect 11701 24225 11713 24228
rect 11747 24225 11759 24259
rect 11701 24219 11759 24225
rect 6089 24191 6147 24197
rect 6089 24157 6101 24191
rect 6135 24157 6147 24191
rect 6089 24151 6147 24157
rect 6270 24148 6276 24200
rect 6328 24148 6334 24200
rect 6362 24148 6368 24200
rect 6420 24148 6426 24200
rect 6641 24191 6699 24197
rect 6641 24157 6653 24191
rect 6687 24157 6699 24191
rect 6641 24151 6699 24157
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24188 6791 24191
rect 7374 24188 7380 24200
rect 6779 24160 7380 24188
rect 6779 24157 6791 24160
rect 6733 24151 6791 24157
rect 6546 24120 6552 24132
rect 5644 24092 6552 24120
rect 6546 24080 6552 24092
rect 6604 24080 6610 24132
rect 4709 24055 4767 24061
rect 4709 24021 4721 24055
rect 4755 24052 4767 24055
rect 4798 24052 4804 24064
rect 4755 24024 4804 24052
rect 4755 24021 4767 24024
rect 4709 24015 4767 24021
rect 4798 24012 4804 24024
rect 4856 24012 4862 24064
rect 6656 24052 6684 24151
rect 7374 24148 7380 24160
rect 7432 24148 7438 24200
rect 8202 24148 8208 24200
rect 8260 24148 8266 24200
rect 10410 24148 10416 24200
rect 10468 24148 10474 24200
rect 11974 24148 11980 24200
rect 12032 24148 12038 24200
rect 12066 24148 12072 24200
rect 12124 24148 12130 24200
rect 12161 24191 12219 24197
rect 12161 24157 12173 24191
rect 12207 24157 12219 24191
rect 12161 24151 12219 24157
rect 7000 24123 7058 24129
rect 7000 24089 7012 24123
rect 7046 24120 7058 24123
rect 7190 24120 7196 24132
rect 7046 24092 7196 24120
rect 7046 24089 7058 24092
rect 7000 24083 7058 24089
rect 7190 24080 7196 24092
rect 7248 24080 7254 24132
rect 9033 24123 9091 24129
rect 9033 24089 9045 24123
rect 9079 24089 9091 24123
rect 9033 24083 9091 24089
rect 7742 24052 7748 24064
rect 6656 24024 7748 24052
rect 7742 24012 7748 24024
rect 7800 24012 7806 24064
rect 8573 24055 8631 24061
rect 8573 24021 8585 24055
rect 8619 24052 8631 24055
rect 8662 24052 8668 24064
rect 8619 24024 8668 24052
rect 8619 24021 8631 24024
rect 8573 24015 8631 24021
rect 8662 24012 8668 24024
rect 8720 24052 8726 24064
rect 9048 24052 9076 24083
rect 11606 24080 11612 24132
rect 11664 24120 11670 24132
rect 12176 24120 12204 24151
rect 12250 24148 12256 24200
rect 12308 24188 12314 24200
rect 12345 24191 12403 24197
rect 12345 24188 12357 24191
rect 12308 24160 12357 24188
rect 12308 24148 12314 24160
rect 12345 24157 12357 24160
rect 12391 24157 12403 24191
rect 12345 24151 12403 24157
rect 11664 24092 12204 24120
rect 11664 24080 11670 24092
rect 8720 24024 9076 24052
rect 8720 24012 8726 24024
rect 9766 24012 9772 24064
rect 9824 24052 9830 24064
rect 9861 24055 9919 24061
rect 9861 24052 9873 24055
rect 9824 24024 9873 24052
rect 9824 24012 9830 24024
rect 9861 24021 9873 24024
rect 9907 24021 9919 24055
rect 9861 24015 9919 24021
rect 10778 24012 10784 24064
rect 10836 24052 10842 24064
rect 10965 24055 11023 24061
rect 10965 24052 10977 24055
rect 10836 24024 10977 24052
rect 10836 24012 10842 24024
rect 10965 24021 10977 24024
rect 11011 24021 11023 24055
rect 10965 24015 11023 24021
rect 1104 23962 16836 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 16836 23962
rect 1104 23888 16836 23910
rect 4433 23851 4491 23857
rect 4433 23817 4445 23851
rect 4479 23848 4491 23851
rect 4614 23848 4620 23860
rect 4479 23820 4620 23848
rect 4479 23817 4491 23820
rect 4433 23811 4491 23817
rect 4614 23808 4620 23820
rect 4672 23808 4678 23860
rect 7742 23808 7748 23860
rect 7800 23848 7806 23860
rect 8021 23851 8079 23857
rect 8021 23848 8033 23851
rect 7800 23820 8033 23848
rect 7800 23808 7806 23820
rect 8021 23817 8033 23820
rect 8067 23817 8079 23851
rect 8021 23811 8079 23817
rect 8202 23808 8208 23860
rect 8260 23848 8266 23860
rect 11057 23851 11115 23857
rect 11057 23848 11069 23851
rect 8260 23820 11069 23848
rect 8260 23808 8266 23820
rect 11057 23817 11069 23820
rect 11103 23817 11115 23851
rect 11057 23811 11115 23817
rect 7653 23783 7711 23789
rect 7653 23749 7665 23783
rect 7699 23780 7711 23783
rect 10042 23780 10048 23792
rect 7699 23752 8156 23780
rect 7699 23749 7711 23752
rect 7653 23743 7711 23749
rect 8128 23724 8156 23752
rect 9508 23752 10048 23780
rect 3050 23672 3056 23724
rect 3108 23672 3114 23724
rect 3142 23672 3148 23724
rect 3200 23712 3206 23724
rect 3309 23715 3367 23721
rect 3309 23712 3321 23715
rect 3200 23684 3321 23712
rect 3200 23672 3206 23684
rect 3309 23681 3321 23684
rect 3355 23681 3367 23715
rect 3309 23675 3367 23681
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23681 7895 23715
rect 7837 23675 7895 23681
rect 7852 23644 7880 23675
rect 8110 23672 8116 23724
rect 8168 23712 8174 23724
rect 8205 23715 8263 23721
rect 8205 23712 8217 23715
rect 8168 23684 8217 23712
rect 8168 23672 8174 23684
rect 8205 23681 8217 23684
rect 8251 23681 8263 23715
rect 8205 23675 8263 23681
rect 8386 23672 8392 23724
rect 8444 23672 8450 23724
rect 9508 23721 9536 23752
rect 10042 23740 10048 23752
rect 10100 23740 10106 23792
rect 9766 23721 9772 23724
rect 9493 23715 9551 23721
rect 9493 23681 9505 23715
rect 9539 23681 9551 23715
rect 9760 23712 9772 23721
rect 9727 23684 9772 23712
rect 9493 23675 9551 23681
rect 9760 23675 9772 23684
rect 9766 23672 9772 23675
rect 9824 23672 9830 23724
rect 10965 23715 11023 23721
rect 10965 23712 10977 23715
rect 10888 23684 10977 23712
rect 8404 23644 8432 23672
rect 7852 23616 8432 23644
rect 6638 23536 6644 23588
rect 6696 23576 6702 23588
rect 10888 23585 10916 23684
rect 10965 23681 10977 23684
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23712 11207 23715
rect 11882 23712 11888 23724
rect 11195 23684 11888 23712
rect 11195 23681 11207 23684
rect 11149 23675 11207 23681
rect 11882 23672 11888 23684
rect 11940 23672 11946 23724
rect 13009 23715 13067 23721
rect 13009 23681 13021 23715
rect 13055 23712 13067 23715
rect 13170 23712 13176 23724
rect 13055 23684 13176 23712
rect 13055 23681 13067 23684
rect 13009 23675 13067 23681
rect 13170 23672 13176 23684
rect 13228 23672 13234 23724
rect 13262 23672 13268 23724
rect 13320 23712 13326 23724
rect 13814 23712 13820 23724
rect 13320 23684 13820 23712
rect 13320 23672 13326 23684
rect 13814 23672 13820 23684
rect 13872 23672 13878 23724
rect 8389 23579 8447 23585
rect 8389 23576 8401 23579
rect 6696 23548 8401 23576
rect 6696 23536 6702 23548
rect 8389 23545 8401 23548
rect 8435 23545 8447 23579
rect 8389 23539 8447 23545
rect 10873 23579 10931 23585
rect 10873 23545 10885 23579
rect 10919 23545 10931 23579
rect 10873 23539 10931 23545
rect 7466 23468 7472 23520
rect 7524 23468 7530 23520
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12158 23508 12164 23520
rect 11931 23480 12164 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12158 23468 12164 23480
rect 12216 23468 12222 23520
rect 1104 23418 16836 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 16836 23418
rect 1104 23344 16836 23366
rect 3142 23264 3148 23316
rect 3200 23264 3206 23316
rect 3326 23264 3332 23316
rect 3384 23304 3390 23316
rect 4706 23304 4712 23316
rect 3384 23276 4712 23304
rect 3384 23264 3390 23276
rect 4706 23264 4712 23276
rect 4764 23264 4770 23316
rect 11882 23264 11888 23316
rect 11940 23264 11946 23316
rect 11974 23264 11980 23316
rect 12032 23264 12038 23316
rect 13170 23264 13176 23316
rect 13228 23304 13234 23316
rect 13265 23307 13323 23313
rect 13265 23304 13277 23307
rect 13228 23276 13277 23304
rect 13228 23264 13234 23276
rect 13265 23273 13277 23276
rect 13311 23273 13323 23307
rect 13265 23267 13323 23273
rect 3068 23208 3832 23236
rect 3068 23180 3096 23208
rect 3050 23128 3056 23180
rect 3108 23128 3114 23180
rect 3804 23177 3832 23208
rect 3789 23171 3847 23177
rect 3789 23137 3801 23171
rect 3835 23137 3847 23171
rect 11900 23168 11928 23264
rect 12529 23171 12587 23177
rect 12529 23168 12541 23171
rect 11900 23140 12541 23168
rect 3789 23131 3847 23137
rect 12529 23137 12541 23140
rect 12575 23137 12587 23171
rect 12529 23131 12587 23137
rect 3326 23060 3332 23112
rect 3384 23060 3390 23112
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 3513 23103 3571 23109
rect 3513 23100 3525 23103
rect 3476 23072 3525 23100
rect 3476 23060 3482 23072
rect 3513 23069 3525 23072
rect 3559 23069 3571 23103
rect 3513 23063 3571 23069
rect 3605 23103 3663 23109
rect 3605 23069 3617 23103
rect 3651 23069 3663 23103
rect 5813 23103 5871 23109
rect 5813 23100 5825 23103
rect 3605 23063 3663 23069
rect 5184 23072 5825 23100
rect 2808 23035 2866 23041
rect 2808 23001 2820 23035
rect 2854 23032 2866 23035
rect 3234 23032 3240 23044
rect 2854 23004 3240 23032
rect 2854 23001 2866 23004
rect 2808 22995 2866 23001
rect 3234 22992 3240 23004
rect 3292 22992 3298 23044
rect 1673 22967 1731 22973
rect 1673 22933 1685 22967
rect 1719 22964 1731 22967
rect 2038 22964 2044 22976
rect 1719 22936 2044 22964
rect 1719 22933 1731 22936
rect 1673 22927 1731 22933
rect 2038 22924 2044 22936
rect 2096 22924 2102 22976
rect 3326 22924 3332 22976
rect 3384 22964 3390 22976
rect 3620 22964 3648 23063
rect 3694 22992 3700 23044
rect 3752 23032 3758 23044
rect 4034 23035 4092 23041
rect 4034 23032 4046 23035
rect 3752 23004 4046 23032
rect 3752 22992 3758 23004
rect 4034 23001 4046 23004
rect 4080 23001 4092 23035
rect 4034 22995 4092 23001
rect 3384 22936 3648 22964
rect 3384 22924 3390 22936
rect 4614 22924 4620 22976
rect 4672 22964 4678 22976
rect 5184 22973 5212 23072
rect 5813 23069 5825 23072
rect 5859 23069 5871 23103
rect 5813 23063 5871 23069
rect 6638 23060 6644 23112
rect 6696 23060 6702 23112
rect 8478 23060 8484 23112
rect 8536 23100 8542 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8536 23072 8953 23100
rect 8536 23060 8542 23072
rect 8941 23069 8953 23072
rect 8987 23100 8999 23103
rect 10042 23100 10048 23112
rect 8987 23072 10048 23100
rect 8987 23069 8999 23072
rect 8941 23063 8999 23069
rect 10042 23060 10048 23072
rect 10100 23100 10106 23112
rect 10778 23109 10784 23112
rect 10505 23103 10563 23109
rect 10505 23100 10517 23103
rect 10100 23072 10517 23100
rect 10100 23060 10106 23072
rect 10505 23069 10517 23072
rect 10551 23069 10563 23103
rect 10772 23100 10784 23109
rect 10739 23072 10784 23100
rect 10505 23063 10563 23069
rect 10772 23063 10784 23072
rect 10778 23060 10784 23063
rect 10836 23060 10842 23112
rect 12158 23060 12164 23112
rect 12216 23100 12222 23112
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 12216 23072 12725 23100
rect 12216 23060 12222 23072
rect 12713 23069 12725 23072
rect 12759 23100 12771 23103
rect 12802 23100 12808 23112
rect 12759 23072 12808 23100
rect 12759 23069 12771 23072
rect 12713 23063 12771 23069
rect 12802 23060 12808 23072
rect 12860 23060 12866 23112
rect 13078 23060 13084 23112
rect 13136 23060 13142 23112
rect 9214 23041 9220 23044
rect 9208 22995 9220 23041
rect 9214 22992 9220 22995
rect 9272 22992 9278 23044
rect 11698 22992 11704 23044
rect 11756 23032 11762 23044
rect 12897 23035 12955 23041
rect 12897 23032 12909 23035
rect 11756 23004 12909 23032
rect 11756 22992 11762 23004
rect 12897 23001 12909 23004
rect 12943 23001 12955 23035
rect 12897 22995 12955 23001
rect 12986 22992 12992 23044
rect 13044 22992 13050 23044
rect 5169 22967 5227 22973
rect 5169 22964 5181 22967
rect 4672 22936 5181 22964
rect 4672 22924 4678 22936
rect 5169 22933 5181 22936
rect 5215 22933 5227 22967
rect 5169 22927 5227 22933
rect 5258 22924 5264 22976
rect 5316 22924 5322 22976
rect 5994 22924 6000 22976
rect 6052 22964 6058 22976
rect 6089 22967 6147 22973
rect 6089 22964 6101 22967
rect 6052 22936 6101 22964
rect 6052 22924 6058 22936
rect 6089 22933 6101 22936
rect 6135 22933 6147 22967
rect 6089 22927 6147 22933
rect 9858 22924 9864 22976
rect 9916 22964 9922 22976
rect 10321 22967 10379 22973
rect 10321 22964 10333 22967
rect 9916 22936 10333 22964
rect 9916 22924 9922 22936
rect 10321 22933 10333 22936
rect 10367 22933 10379 22967
rect 10321 22927 10379 22933
rect 1104 22874 16836 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 16836 22874
rect 1104 22800 16836 22822
rect 3605 22763 3663 22769
rect 3605 22729 3617 22763
rect 3651 22729 3663 22763
rect 3605 22723 3663 22729
rect 3234 22652 3240 22704
rect 3292 22692 3298 22704
rect 3620 22692 3648 22723
rect 6270 22720 6276 22772
rect 6328 22760 6334 22772
rect 6457 22763 6515 22769
rect 6457 22760 6469 22763
rect 6328 22732 6469 22760
rect 6328 22720 6334 22732
rect 6457 22729 6469 22732
rect 6503 22729 6515 22763
rect 6457 22723 6515 22729
rect 9861 22763 9919 22769
rect 9861 22729 9873 22763
rect 9907 22760 9919 22763
rect 10410 22760 10416 22772
rect 9907 22732 10416 22760
rect 9907 22729 9919 22732
rect 9861 22723 9919 22729
rect 10410 22720 10416 22732
rect 10468 22720 10474 22772
rect 11698 22720 11704 22772
rect 11756 22720 11762 22772
rect 12066 22720 12072 22772
rect 12124 22760 12130 22772
rect 12253 22763 12311 22769
rect 12253 22760 12265 22763
rect 12124 22732 12265 22760
rect 12124 22720 12130 22732
rect 12253 22729 12265 22732
rect 12299 22729 12311 22763
rect 12253 22723 12311 22729
rect 3292 22664 3648 22692
rect 3773 22695 3831 22701
rect 3292 22652 3298 22664
rect 3773 22661 3785 22695
rect 3819 22692 3831 22695
rect 3878 22692 3884 22704
rect 3819 22664 3884 22692
rect 3819 22661 3831 22664
rect 3773 22655 3831 22661
rect 3878 22652 3884 22664
rect 3936 22652 3942 22704
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22692 4031 22695
rect 5258 22692 5264 22704
rect 4019 22664 5264 22692
rect 4019 22661 4031 22664
rect 3973 22655 4031 22661
rect 5258 22652 5264 22664
rect 5316 22652 5322 22704
rect 6288 22692 6316 22720
rect 5920 22664 6316 22692
rect 842 22584 848 22636
rect 900 22624 906 22636
rect 1489 22627 1547 22633
rect 1489 22624 1501 22627
rect 900 22596 1501 22624
rect 900 22584 906 22596
rect 1489 22593 1501 22596
rect 1535 22593 1547 22627
rect 1489 22587 1547 22593
rect 3418 22584 3424 22636
rect 3476 22584 3482 22636
rect 3513 22627 3571 22633
rect 3513 22593 3525 22627
rect 3559 22624 3571 22627
rect 4065 22627 4123 22633
rect 4065 22624 4077 22627
rect 3559 22596 4077 22624
rect 3559 22593 3571 22596
rect 3513 22587 3571 22593
rect 4065 22593 4077 22596
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 4798 22584 4804 22636
rect 4856 22584 4862 22636
rect 5920 22633 5948 22664
rect 4985 22627 5043 22633
rect 4985 22593 4997 22627
rect 5031 22593 5043 22627
rect 4985 22587 5043 22593
rect 5905 22627 5963 22633
rect 5905 22593 5917 22627
rect 5951 22593 5963 22627
rect 5905 22587 5963 22593
rect 3436 22556 3464 22584
rect 3878 22556 3884 22568
rect 3436 22528 3884 22556
rect 3878 22516 3884 22528
rect 3936 22516 3942 22568
rect 4709 22559 4767 22565
rect 4709 22525 4721 22559
rect 4755 22556 4767 22559
rect 4893 22559 4951 22565
rect 4893 22556 4905 22559
rect 4755 22528 4905 22556
rect 4755 22525 4767 22528
rect 4709 22519 4767 22525
rect 4893 22525 4905 22528
rect 4939 22525 4951 22559
rect 4893 22519 4951 22525
rect 1673 22491 1731 22497
rect 1673 22457 1685 22491
rect 1719 22488 1731 22491
rect 1762 22488 1768 22500
rect 1719 22460 1768 22488
rect 1719 22457 1731 22460
rect 1673 22451 1731 22457
rect 1762 22448 1768 22460
rect 1820 22448 1826 22500
rect 3237 22491 3295 22497
rect 3237 22457 3249 22491
rect 3283 22488 3295 22491
rect 3694 22488 3700 22500
rect 3283 22460 3700 22488
rect 3283 22457 3295 22460
rect 3237 22451 3295 22457
rect 3694 22448 3700 22460
rect 3752 22448 3758 22500
rect 4614 22448 4620 22500
rect 4672 22488 4678 22500
rect 5000 22488 5028 22587
rect 5810 22516 5816 22568
rect 5868 22516 5874 22568
rect 4672 22460 5028 22488
rect 4672 22448 4678 22460
rect 5920 22432 5948 22587
rect 5994 22584 6000 22636
rect 6052 22584 6058 22636
rect 6457 22627 6515 22633
rect 6457 22593 6469 22627
rect 6503 22593 6515 22627
rect 6457 22587 6515 22593
rect 6089 22559 6147 22565
rect 6089 22525 6101 22559
rect 6135 22525 6147 22559
rect 6472 22556 6500 22587
rect 6546 22584 6552 22636
rect 6604 22624 6610 22636
rect 6641 22627 6699 22633
rect 6641 22624 6653 22627
rect 6604 22596 6653 22624
rect 6604 22584 6610 22596
rect 6641 22593 6653 22596
rect 6687 22624 6699 22627
rect 6822 22624 6828 22636
rect 6687 22596 6828 22624
rect 6687 22593 6699 22596
rect 6641 22587 6699 22593
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 7282 22584 7288 22636
rect 7340 22624 7346 22636
rect 7466 22624 7472 22636
rect 7340 22596 7472 22624
rect 7340 22584 7346 22596
rect 7466 22584 7472 22596
rect 7524 22584 7530 22636
rect 7653 22627 7711 22633
rect 7653 22593 7665 22627
rect 7699 22593 7711 22627
rect 7653 22587 7711 22593
rect 6730 22556 6736 22568
rect 6472 22528 6736 22556
rect 6089 22519 6147 22525
rect 6104 22488 6132 22519
rect 6730 22516 6736 22528
rect 6788 22516 6794 22568
rect 7006 22488 7012 22500
rect 6104 22460 7012 22488
rect 7006 22448 7012 22460
rect 7064 22448 7070 22500
rect 7466 22448 7472 22500
rect 7524 22488 7530 22500
rect 7668 22488 7696 22587
rect 8478 22584 8484 22636
rect 8536 22584 8542 22636
rect 8754 22633 8760 22636
rect 8748 22587 8760 22633
rect 8754 22584 8760 22587
rect 8812 22584 8818 22636
rect 11606 22584 11612 22636
rect 11664 22584 11670 22636
rect 11793 22627 11851 22633
rect 11793 22593 11805 22627
rect 11839 22624 11851 22627
rect 12084 22624 12112 22720
rect 11839 22596 12112 22624
rect 11839 22593 11851 22596
rect 11793 22587 11851 22593
rect 8386 22516 8392 22568
rect 8444 22516 8450 22568
rect 7745 22491 7803 22497
rect 7745 22488 7757 22491
rect 7524 22460 7757 22488
rect 7524 22448 7530 22460
rect 7745 22457 7757 22460
rect 7791 22457 7803 22491
rect 12084 22488 12112 22596
rect 12158 22584 12164 22636
rect 12216 22584 12222 22636
rect 12345 22627 12403 22633
rect 12345 22593 12357 22627
rect 12391 22624 12403 22627
rect 12434 22624 12440 22636
rect 12391 22596 12440 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 12434 22584 12440 22596
rect 12492 22584 12498 22636
rect 16114 22584 16120 22636
rect 16172 22624 16178 22636
rect 16209 22627 16267 22633
rect 16209 22624 16221 22627
rect 16172 22596 16221 22624
rect 16172 22584 16178 22596
rect 16209 22593 16221 22596
rect 16255 22593 16267 22627
rect 16209 22587 16267 22593
rect 12802 22516 12808 22568
rect 12860 22556 12866 22568
rect 12897 22559 12955 22565
rect 12897 22556 12909 22559
rect 12860 22528 12909 22556
rect 12860 22516 12866 22528
rect 12897 22525 12909 22528
rect 12943 22525 12955 22559
rect 12897 22519 12955 22525
rect 13173 22491 13231 22497
rect 13173 22488 13185 22491
rect 12084 22460 13185 22488
rect 7745 22451 7803 22457
rect 13173 22457 13185 22460
rect 13219 22457 13231 22491
rect 13173 22451 13231 22457
rect 16390 22448 16396 22500
rect 16448 22448 16454 22500
rect 3789 22423 3847 22429
rect 3789 22389 3801 22423
rect 3835 22420 3847 22423
rect 4798 22420 4804 22432
rect 3835 22392 4804 22420
rect 3835 22389 3847 22392
rect 3789 22383 3847 22389
rect 4798 22380 4804 22392
rect 4856 22380 4862 22432
rect 5626 22380 5632 22432
rect 5684 22380 5690 22432
rect 5902 22380 5908 22432
rect 5960 22380 5966 22432
rect 7190 22380 7196 22432
rect 7248 22420 7254 22432
rect 7377 22423 7435 22429
rect 7377 22420 7389 22423
rect 7248 22392 7389 22420
rect 7248 22380 7254 22392
rect 7377 22389 7389 22392
rect 7423 22389 7435 22423
rect 7377 22383 7435 22389
rect 7558 22380 7564 22432
rect 7616 22380 7622 22432
rect 13357 22423 13415 22429
rect 13357 22389 13369 22423
rect 13403 22420 13415 22423
rect 14274 22420 14280 22432
rect 13403 22392 14280 22420
rect 13403 22389 13415 22392
rect 13357 22383 13415 22389
rect 14274 22380 14280 22392
rect 14332 22380 14338 22432
rect 1104 22330 16836 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 16836 22330
rect 1104 22256 16836 22278
rect 9861 22219 9919 22225
rect 9861 22185 9873 22219
rect 9907 22216 9919 22219
rect 9950 22216 9956 22228
rect 9907 22188 9956 22216
rect 9907 22185 9919 22188
rect 9861 22179 9919 22185
rect 9950 22176 9956 22188
rect 10008 22176 10014 22228
rect 16114 22176 16120 22228
rect 16172 22176 16178 22228
rect 8386 22108 8392 22160
rect 8444 22148 8450 22160
rect 8757 22151 8815 22157
rect 8757 22148 8769 22151
rect 8444 22120 8769 22148
rect 8444 22108 8450 22120
rect 8757 22117 8769 22120
rect 8803 22117 8815 22151
rect 8757 22111 8815 22117
rect 12434 22108 12440 22160
rect 12492 22108 12498 22160
rect 7374 22040 7380 22092
rect 7432 22040 7438 22092
rect 842 21972 848 22024
rect 900 22012 906 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 900 21984 1409 22012
rect 900 21972 906 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 22012 1731 22015
rect 1854 22012 1860 22024
rect 1719 21984 1860 22012
rect 1719 21981 1731 21984
rect 1673 21975 1731 21981
rect 1854 21972 1860 21984
rect 1912 22012 1918 22024
rect 1912 21984 2544 22012
rect 1912 21972 1918 21984
rect 106 21904 112 21956
rect 164 21944 170 21956
rect 2516 21944 2544 21984
rect 2774 21972 2780 22024
rect 2832 22012 2838 22024
rect 2869 22015 2927 22021
rect 2869 22012 2881 22015
rect 2832 21984 2881 22012
rect 2832 21972 2838 21984
rect 2869 21981 2881 21984
rect 2915 21981 2927 22015
rect 2869 21975 2927 21981
rect 3050 21972 3056 22024
rect 3108 22012 3114 22024
rect 4706 22012 4712 22024
rect 3108 21984 4712 22012
rect 3108 21972 3114 21984
rect 4706 21972 4712 21984
rect 4764 22012 4770 22024
rect 5353 22015 5411 22021
rect 5353 22012 5365 22015
rect 4764 21984 5365 22012
rect 4764 21972 4770 21984
rect 5353 21981 5365 21984
rect 5399 21981 5411 22015
rect 5353 21975 5411 21981
rect 5552 21984 6960 22012
rect 3786 21944 3792 21956
rect 164 21916 2452 21944
rect 2516 21916 3792 21944
rect 164 21904 170 21916
rect 2314 21836 2320 21888
rect 2372 21836 2378 21888
rect 2424 21876 2452 21916
rect 3786 21904 3792 21916
rect 3844 21944 3850 21956
rect 5552 21944 5580 21984
rect 3844 21916 5580 21944
rect 5620 21947 5678 21953
rect 3844 21904 3850 21916
rect 5620 21913 5632 21947
rect 5666 21944 5678 21947
rect 6825 21947 6883 21953
rect 6825 21944 6837 21947
rect 5666 21916 6837 21944
rect 5666 21913 5678 21916
rect 5620 21907 5678 21913
rect 6825 21913 6837 21916
rect 6871 21913 6883 21947
rect 6825 21907 6883 21913
rect 5810 21876 5816 21888
rect 2424 21848 5816 21876
rect 5810 21836 5816 21848
rect 5868 21836 5874 21888
rect 6546 21836 6552 21888
rect 6604 21876 6610 21888
rect 6730 21876 6736 21888
rect 6604 21848 6736 21876
rect 6604 21836 6610 21848
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 6932 21876 6960 21984
rect 7006 21972 7012 22024
rect 7064 21972 7070 22024
rect 7190 21972 7196 22024
rect 7248 21972 7254 22024
rect 7282 21972 7288 22024
rect 7340 22012 7346 22024
rect 8404 22012 8432 22108
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 10137 22083 10195 22089
rect 10137 22080 10149 22083
rect 10100 22052 10149 22080
rect 10100 22040 10106 22052
rect 10137 22049 10149 22052
rect 10183 22049 10195 22083
rect 10137 22043 10195 22049
rect 7340 21984 7382 22012
rect 7576 21984 8432 22012
rect 9493 22015 9551 22021
rect 7340 21972 7346 21984
rect 7374 21904 7380 21956
rect 7432 21944 7438 21956
rect 7576 21944 7604 21984
rect 9493 21981 9505 22015
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 7650 21953 7656 21956
rect 7432 21916 7604 21944
rect 7432 21904 7438 21916
rect 7644 21907 7656 21953
rect 7650 21904 7656 21907
rect 7708 21904 7714 21956
rect 9508 21876 9536 21975
rect 11330 21972 11336 22024
rect 11388 22012 11394 22024
rect 11609 22015 11667 22021
rect 11609 22012 11621 22015
rect 11388 21984 11621 22012
rect 11388 21972 11394 21984
rect 11609 21981 11621 21984
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 21981 11851 22015
rect 11793 21975 11851 21981
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 22012 12403 22015
rect 12526 22012 12532 22024
rect 12391 21984 12532 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 9858 21904 9864 21956
rect 9916 21904 9922 21956
rect 10404 21947 10462 21953
rect 10404 21913 10416 21947
rect 10450 21944 10462 21947
rect 11701 21947 11759 21953
rect 11701 21944 11713 21947
rect 10450 21916 11713 21944
rect 10450 21913 10462 21916
rect 10404 21907 10462 21913
rect 11701 21913 11713 21916
rect 11747 21913 11759 21947
rect 11808 21944 11836 21975
rect 12526 21972 12532 21984
rect 12584 22012 12590 22024
rect 12986 22012 12992 22024
rect 12584 21984 12992 22012
rect 12584 21972 12590 21984
rect 12986 21972 12992 21984
rect 13044 21972 13050 22024
rect 13814 21972 13820 22024
rect 13872 22012 13878 22024
rect 14366 22012 14372 22024
rect 13872 21984 14372 22012
rect 13872 21972 13878 21984
rect 14366 21972 14372 21984
rect 14424 21972 14430 22024
rect 15930 21972 15936 22024
rect 15988 21972 15994 22024
rect 16114 21972 16120 22024
rect 16172 22012 16178 22024
rect 16209 22015 16267 22021
rect 16209 22012 16221 22015
rect 16172 21984 16221 22012
rect 16172 21972 16178 21984
rect 16209 21981 16221 21984
rect 16255 21981 16267 22015
rect 16209 21975 16267 21981
rect 12618 21944 12624 21956
rect 11808 21916 12624 21944
rect 11701 21907 11759 21913
rect 12618 21904 12624 21916
rect 12676 21904 12682 21956
rect 13354 21904 13360 21956
rect 13412 21944 13418 21956
rect 13550 21947 13608 21953
rect 13550 21944 13562 21947
rect 13412 21916 13562 21944
rect 13412 21904 13418 21916
rect 13550 21913 13562 21916
rect 13596 21913 13608 21947
rect 13550 21907 13608 21913
rect 9674 21876 9680 21888
rect 6932 21848 9680 21876
rect 9674 21836 9680 21848
rect 9732 21836 9738 21888
rect 10045 21879 10103 21885
rect 10045 21845 10057 21879
rect 10091 21876 10103 21879
rect 11422 21876 11428 21888
rect 10091 21848 11428 21876
rect 10091 21845 10103 21848
rect 10045 21839 10103 21845
rect 11422 21836 11428 21848
rect 11480 21836 11486 21888
rect 11517 21879 11575 21885
rect 11517 21845 11529 21879
rect 11563 21876 11575 21879
rect 11790 21876 11796 21888
rect 11563 21848 11796 21876
rect 11563 21845 11575 21848
rect 11517 21839 11575 21845
rect 11790 21836 11796 21848
rect 11848 21876 11854 21888
rect 12158 21876 12164 21888
rect 11848 21848 12164 21876
rect 11848 21836 11854 21848
rect 12158 21836 12164 21848
rect 12216 21836 12222 21888
rect 12250 21836 12256 21888
rect 12308 21876 12314 21888
rect 13262 21876 13268 21888
rect 12308 21848 13268 21876
rect 12308 21836 12314 21848
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 16390 21836 16396 21888
rect 16448 21836 16454 21888
rect 1104 21786 16836 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 16836 21786
rect 1104 21712 16836 21734
rect 2685 21675 2743 21681
rect 2685 21641 2697 21675
rect 2731 21672 2743 21675
rect 2866 21672 2872 21684
rect 2731 21644 2872 21672
rect 2731 21641 2743 21644
rect 2685 21635 2743 21641
rect 2866 21632 2872 21644
rect 2924 21632 2930 21684
rect 3050 21632 3056 21684
rect 3108 21632 3114 21684
rect 6089 21675 6147 21681
rect 6089 21641 6101 21675
rect 6135 21672 6147 21675
rect 6135 21644 6592 21672
rect 6135 21641 6147 21644
rect 6089 21635 6147 21641
rect 3068 21604 3096 21632
rect 2792 21576 3096 21604
rect 4976 21607 5034 21613
rect 2792 21548 2820 21576
rect 4976 21573 4988 21607
rect 5022 21604 5034 21607
rect 5626 21604 5632 21616
rect 5022 21576 5632 21604
rect 5022 21573 5034 21576
rect 4976 21567 5034 21573
rect 5626 21564 5632 21576
rect 5684 21564 5690 21616
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21536 1731 21539
rect 1762 21536 1768 21548
rect 1719 21508 1768 21536
rect 1719 21505 1731 21508
rect 1673 21499 1731 21505
rect 1762 21496 1768 21508
rect 1820 21496 1826 21548
rect 2038 21496 2044 21548
rect 2096 21496 2102 21548
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 3050 21545 3056 21548
rect 3044 21499 3056 21545
rect 3050 21496 3056 21499
rect 3108 21496 3114 21548
rect 3878 21496 3884 21548
rect 3936 21536 3942 21548
rect 4249 21539 4307 21545
rect 4249 21536 4261 21539
rect 3936 21508 4261 21536
rect 3936 21496 3942 21508
rect 4249 21505 4261 21508
rect 4295 21505 4307 21539
rect 4249 21499 4307 21505
rect 4433 21539 4491 21545
rect 4433 21505 4445 21539
rect 4479 21536 4491 21539
rect 4614 21536 4620 21548
rect 4479 21508 4620 21536
rect 4479 21505 4491 21508
rect 4433 21499 4491 21505
rect 4614 21496 4620 21508
rect 4672 21496 4678 21548
rect 4706 21496 4712 21548
rect 4764 21496 4770 21548
rect 5718 21496 5724 21548
rect 5776 21536 5782 21548
rect 6564 21545 6592 21644
rect 7006 21632 7012 21684
rect 7064 21672 7070 21684
rect 7064 21644 7236 21672
rect 7064 21632 7070 21644
rect 6730 21564 6736 21616
rect 6788 21604 6794 21616
rect 7101 21607 7159 21613
rect 7101 21604 7113 21607
rect 6788 21576 7113 21604
rect 6788 21564 6794 21576
rect 7101 21573 7113 21576
rect 7147 21573 7159 21607
rect 7208 21604 7236 21644
rect 7650 21632 7656 21684
rect 7708 21632 7714 21684
rect 11330 21632 11336 21684
rect 11388 21632 11394 21684
rect 11422 21632 11428 21684
rect 11480 21672 11486 21684
rect 11885 21675 11943 21681
rect 11885 21672 11897 21675
rect 11480 21644 11897 21672
rect 11480 21632 11486 21644
rect 11885 21641 11897 21644
rect 11931 21641 11943 21675
rect 11885 21635 11943 21641
rect 12161 21675 12219 21681
rect 12161 21641 12173 21675
rect 12207 21641 12219 21675
rect 12161 21635 12219 21641
rect 12437 21675 12495 21681
rect 12437 21641 12449 21675
rect 12483 21672 12495 21675
rect 12526 21672 12532 21684
rect 12483 21644 12532 21672
rect 12483 21641 12495 21644
rect 12437 21635 12495 21641
rect 7837 21607 7895 21613
rect 7837 21604 7849 21607
rect 7208 21576 7849 21604
rect 7101 21567 7159 21573
rect 7837 21573 7849 21576
rect 7883 21573 7895 21607
rect 7837 21567 7895 21573
rect 6365 21539 6423 21545
rect 6365 21536 6377 21539
rect 5776 21508 6377 21536
rect 5776 21496 5782 21508
rect 6365 21505 6377 21508
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21536 6607 21539
rect 6638 21536 6644 21548
rect 6595 21508 6644 21536
rect 6595 21505 6607 21508
rect 6549 21499 6607 21505
rect 6638 21496 6644 21508
rect 6696 21496 6702 21548
rect 6914 21496 6920 21548
rect 6972 21536 6978 21548
rect 7282 21536 7288 21548
rect 6972 21508 7288 21536
rect 6972 21496 6978 21508
rect 7282 21496 7288 21508
rect 7340 21496 7346 21548
rect 7377 21539 7435 21545
rect 7377 21505 7389 21539
rect 7423 21536 7435 21539
rect 7466 21536 7472 21548
rect 7423 21508 7472 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 7466 21496 7472 21508
rect 7524 21496 7530 21548
rect 7745 21539 7803 21545
rect 7745 21505 7757 21539
rect 7791 21505 7803 21539
rect 7745 21499 7803 21505
rect 1946 21428 1952 21480
rect 2004 21428 2010 21480
rect 7558 21428 7564 21480
rect 7616 21468 7622 21480
rect 7653 21471 7711 21477
rect 7653 21468 7665 21471
rect 7616 21440 7665 21468
rect 7616 21428 7622 21440
rect 7653 21437 7665 21440
rect 7699 21437 7711 21471
rect 7653 21431 7711 21437
rect 1765 21403 1823 21409
rect 1765 21369 1777 21403
rect 1811 21400 1823 21403
rect 6733 21403 6791 21409
rect 1811 21372 2774 21400
rect 1811 21369 1823 21372
rect 1765 21363 1823 21369
rect 1857 21335 1915 21341
rect 1857 21301 1869 21335
rect 1903 21332 1915 21335
rect 2130 21332 2136 21344
rect 1903 21304 2136 21332
rect 1903 21301 1915 21304
rect 1857 21295 1915 21301
rect 2130 21292 2136 21304
rect 2188 21292 2194 21344
rect 2746 21332 2774 21372
rect 6733 21369 6745 21403
rect 6779 21400 6791 21403
rect 7760 21400 7788 21499
rect 9674 21496 9680 21548
rect 9732 21496 9738 21548
rect 9858 21496 9864 21548
rect 9916 21496 9922 21548
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 11146 21496 11152 21548
rect 11204 21496 11210 21548
rect 11900 21536 11928 21635
rect 12176 21604 12204 21635
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 12618 21604 12624 21616
rect 12176 21576 12624 21604
rect 12618 21564 12624 21576
rect 12676 21604 12682 21616
rect 13078 21604 13084 21616
rect 12676 21576 13084 21604
rect 12676 21564 12682 21576
rect 13078 21564 13084 21576
rect 13136 21604 13142 21616
rect 13173 21607 13231 21613
rect 13173 21604 13185 21607
rect 13136 21576 13185 21604
rect 13136 21564 13142 21576
rect 13173 21573 13185 21576
rect 13219 21573 13231 21607
rect 13173 21567 13231 21573
rect 12342 21536 12348 21548
rect 11900 21508 12348 21536
rect 12342 21496 12348 21508
rect 12400 21496 12406 21548
rect 13446 21496 13452 21548
rect 13504 21536 13510 21548
rect 13541 21539 13599 21545
rect 13541 21536 13553 21539
rect 13504 21508 13553 21536
rect 13504 21496 13510 21508
rect 13541 21505 13553 21508
rect 13587 21505 13599 21539
rect 13541 21499 13599 21505
rect 14366 21496 14372 21548
rect 14424 21496 14430 21548
rect 14642 21545 14648 21548
rect 14636 21499 14648 21545
rect 14642 21496 14648 21499
rect 14700 21496 14706 21548
rect 9766 21428 9772 21480
rect 9824 21468 9830 21480
rect 9968 21468 9996 21496
rect 9824 21440 9996 21468
rect 10873 21471 10931 21477
rect 9824 21428 9830 21440
rect 10873 21437 10885 21471
rect 10919 21468 10931 21471
rect 11517 21471 11575 21477
rect 11517 21468 11529 21471
rect 10919 21440 11529 21468
rect 10919 21437 10931 21440
rect 10873 21431 10931 21437
rect 11517 21437 11529 21440
rect 11563 21437 11575 21471
rect 11517 21431 11575 21437
rect 6779 21372 7788 21400
rect 10321 21403 10379 21409
rect 6779 21369 6791 21372
rect 6733 21363 6791 21369
rect 10321 21369 10333 21403
rect 10367 21400 10379 21403
rect 10965 21403 11023 21409
rect 10965 21400 10977 21403
rect 10367 21372 10977 21400
rect 10367 21369 10379 21372
rect 10321 21363 10379 21369
rect 10965 21369 10977 21372
rect 11011 21400 11023 21403
rect 11238 21400 11244 21412
rect 11011 21372 11244 21400
rect 11011 21369 11023 21372
rect 10965 21363 11023 21369
rect 11238 21360 11244 21372
rect 11296 21360 11302 21412
rect 11532 21400 11560 21431
rect 11790 21428 11796 21480
rect 11848 21428 11854 21480
rect 11974 21428 11980 21480
rect 12032 21477 12038 21480
rect 12032 21471 12060 21477
rect 12048 21437 12060 21471
rect 12032 21431 12060 21437
rect 12989 21471 13047 21477
rect 12989 21437 13001 21471
rect 13035 21437 13047 21471
rect 12989 21431 13047 21437
rect 12032 21428 12038 21431
rect 12158 21400 12164 21412
rect 11532 21372 12164 21400
rect 12158 21360 12164 21372
rect 12216 21360 12222 21412
rect 12526 21360 12532 21412
rect 12584 21400 12590 21412
rect 12894 21400 12900 21412
rect 12584 21372 12900 21400
rect 12584 21360 12590 21372
rect 12894 21360 12900 21372
rect 12952 21400 12958 21412
rect 13004 21400 13032 21431
rect 13262 21428 13268 21480
rect 13320 21468 13326 21480
rect 13357 21471 13415 21477
rect 13357 21468 13369 21471
rect 13320 21440 13369 21468
rect 13320 21428 13326 21440
rect 13357 21437 13369 21440
rect 13403 21437 13415 21471
rect 15930 21468 15936 21480
rect 13357 21431 13415 21437
rect 15764 21440 15936 21468
rect 13449 21403 13507 21409
rect 13449 21400 13461 21403
rect 12952 21372 13032 21400
rect 13280 21372 13461 21400
rect 12952 21360 12958 21372
rect 3970 21332 3976 21344
rect 2746 21304 3976 21332
rect 3970 21292 3976 21304
rect 4028 21292 4034 21344
rect 4062 21292 4068 21344
rect 4120 21332 4126 21344
rect 4157 21335 4215 21341
rect 4157 21332 4169 21335
rect 4120 21304 4169 21332
rect 4120 21292 4126 21304
rect 4157 21301 4169 21304
rect 4203 21301 4215 21335
rect 4157 21295 4215 21301
rect 4249 21335 4307 21341
rect 4249 21301 4261 21335
rect 4295 21332 4307 21335
rect 6454 21332 6460 21344
rect 4295 21304 6460 21332
rect 4295 21301 4307 21304
rect 4249 21295 4307 21301
rect 6454 21292 6460 21304
rect 6512 21292 6518 21344
rect 6546 21292 6552 21344
rect 6604 21292 6610 21344
rect 7285 21335 7343 21341
rect 7285 21301 7297 21335
rect 7331 21332 7343 21335
rect 7374 21332 7380 21344
rect 7331 21304 7380 21332
rect 7331 21301 7343 21304
rect 7285 21295 7343 21301
rect 7374 21292 7380 21304
rect 7432 21332 7438 21344
rect 7469 21335 7527 21341
rect 7469 21332 7481 21335
rect 7432 21304 7481 21332
rect 7432 21292 7438 21304
rect 7469 21301 7481 21304
rect 7515 21301 7527 21335
rect 7469 21295 7527 21301
rect 11606 21292 11612 21344
rect 11664 21332 11670 21344
rect 13280 21332 13308 21372
rect 13449 21369 13461 21372
rect 13495 21400 13507 21403
rect 14182 21400 14188 21412
rect 13495 21372 14188 21400
rect 13495 21369 13507 21372
rect 13449 21363 13507 21369
rect 14182 21360 14188 21372
rect 14240 21360 14246 21412
rect 15764 21409 15792 21440
rect 15930 21428 15936 21440
rect 15988 21468 15994 21480
rect 16393 21471 16451 21477
rect 16393 21468 16405 21471
rect 15988 21440 16405 21468
rect 15988 21428 15994 21440
rect 16393 21437 16405 21440
rect 16439 21437 16451 21471
rect 16393 21431 16451 21437
rect 15749 21403 15807 21409
rect 15749 21369 15761 21403
rect 15795 21369 15807 21403
rect 15749 21363 15807 21369
rect 11664 21304 13308 21332
rect 11664 21292 11670 21304
rect 13354 21292 13360 21344
rect 13412 21292 13418 21344
rect 15838 21292 15844 21344
rect 15896 21292 15902 21344
rect 1104 21242 16836 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 16836 21242
rect 1104 21168 16836 21190
rect 2682 21088 2688 21140
rect 2740 21128 2746 21140
rect 2777 21131 2835 21137
rect 2777 21128 2789 21131
rect 2740 21100 2789 21128
rect 2740 21088 2746 21100
rect 2777 21097 2789 21100
rect 2823 21097 2835 21131
rect 2777 21091 2835 21097
rect 3050 21088 3056 21140
rect 3108 21088 3114 21140
rect 3237 21131 3295 21137
rect 3237 21097 3249 21131
rect 3283 21128 3295 21131
rect 3878 21128 3884 21140
rect 3283 21100 3884 21128
rect 3283 21097 3295 21100
rect 3237 21091 3295 21097
rect 2961 21063 3019 21069
rect 2961 21029 2973 21063
rect 3007 21060 3019 21063
rect 3252 21060 3280 21091
rect 3878 21088 3884 21100
rect 3936 21088 3942 21140
rect 3970 21088 3976 21140
rect 4028 21128 4034 21140
rect 4617 21131 4675 21137
rect 4617 21128 4629 21131
rect 4028 21100 4629 21128
rect 4028 21088 4034 21100
rect 4617 21097 4629 21100
rect 4663 21097 4675 21131
rect 4617 21091 4675 21097
rect 4801 21131 4859 21137
rect 4801 21097 4813 21131
rect 4847 21097 4859 21131
rect 4801 21091 4859 21097
rect 3694 21060 3700 21072
rect 3007 21032 3280 21060
rect 3528 21032 3700 21060
rect 3007 21029 3019 21032
rect 2961 21023 3019 21029
rect 3142 20952 3148 21004
rect 3200 20952 3206 21004
rect 1397 20927 1455 20933
rect 1397 20893 1409 20927
rect 1443 20924 1455 20927
rect 2774 20924 2780 20936
rect 1443 20896 2780 20924
rect 1443 20893 1455 20896
rect 1397 20887 1455 20893
rect 2774 20884 2780 20896
rect 2832 20884 2838 20936
rect 2869 20927 2927 20933
rect 2869 20893 2881 20927
rect 2915 20924 2927 20927
rect 2958 20924 2964 20936
rect 2915 20896 2964 20924
rect 2915 20893 2927 20896
rect 2869 20887 2927 20893
rect 2958 20884 2964 20896
rect 3016 20924 3022 20936
rect 3326 20924 3332 20936
rect 3016 20896 3332 20924
rect 3016 20884 3022 20896
rect 3326 20884 3332 20896
rect 3384 20884 3390 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20926 3479 20927
rect 3528 20926 3556 21032
rect 3694 21020 3700 21032
rect 3752 21060 3758 21072
rect 4062 21060 4068 21072
rect 3752 21032 4068 21060
rect 3752 21020 3758 21032
rect 4062 21020 4068 21032
rect 4120 21060 4126 21072
rect 4816 21060 4844 21091
rect 5718 21088 5724 21140
rect 5776 21128 5782 21140
rect 5813 21131 5871 21137
rect 5813 21128 5825 21131
rect 5776 21100 5825 21128
rect 5776 21088 5782 21100
rect 5813 21097 5825 21100
rect 5859 21097 5871 21131
rect 5813 21091 5871 21097
rect 6273 21131 6331 21137
rect 6273 21097 6285 21131
rect 6319 21128 6331 21131
rect 6914 21128 6920 21140
rect 6319 21100 6920 21128
rect 6319 21097 6331 21100
rect 6273 21091 6331 21097
rect 6914 21088 6920 21100
rect 6972 21088 6978 21140
rect 8573 21131 8631 21137
rect 8573 21097 8585 21131
rect 8619 21097 8631 21131
rect 8573 21091 8631 21097
rect 4120 21032 4844 21060
rect 4120 21020 4126 21032
rect 5736 20992 5764 21088
rect 6362 21020 6368 21072
rect 6420 21060 6426 21072
rect 6457 21063 6515 21069
rect 6457 21060 6469 21063
rect 6420 21032 6469 21060
rect 6420 21020 6426 21032
rect 6457 21029 6469 21032
rect 6503 21029 6515 21063
rect 6457 21023 6515 21029
rect 6546 21020 6552 21072
rect 6604 21060 6610 21072
rect 8588 21060 8616 21091
rect 10226 21088 10232 21140
rect 10284 21088 10290 21140
rect 11146 21088 11152 21140
rect 11204 21128 11210 21140
rect 11514 21128 11520 21140
rect 11204 21100 11520 21128
rect 11204 21088 11210 21100
rect 11514 21088 11520 21100
rect 11572 21128 11578 21140
rect 11793 21131 11851 21137
rect 11793 21128 11805 21131
rect 11572 21100 11805 21128
rect 11572 21088 11578 21100
rect 11793 21097 11805 21100
rect 11839 21097 11851 21131
rect 11793 21091 11851 21097
rect 9858 21060 9864 21072
rect 6604 21032 9864 21060
rect 6604 21020 6610 21032
rect 9858 21020 9864 21032
rect 9916 21020 9922 21072
rect 3620 20964 5028 20992
rect 3620 20936 3648 20964
rect 3467 20898 3556 20926
rect 3467 20893 3479 20898
rect 3421 20887 3479 20893
rect 3602 20884 3608 20936
rect 3660 20884 3666 20936
rect 4157 20927 4215 20933
rect 4157 20924 4169 20927
rect 3712 20896 4169 20924
rect 1486 20816 1492 20868
rect 1544 20856 1550 20868
rect 1642 20859 1700 20865
rect 1642 20856 1654 20859
rect 1544 20828 1654 20856
rect 1544 20816 1550 20828
rect 1642 20825 1654 20828
rect 1688 20825 1700 20859
rect 1642 20819 1700 20825
rect 1762 20816 1768 20868
rect 1820 20856 1826 20868
rect 3712 20856 3740 20896
rect 4157 20893 4169 20896
rect 4203 20893 4215 20927
rect 4525 20927 4583 20933
rect 4525 20924 4537 20927
rect 4157 20887 4215 20893
rect 4264 20896 4537 20924
rect 1820 20828 3740 20856
rect 1820 20816 1826 20828
rect 3712 20788 3740 20828
rect 3786 20816 3792 20868
rect 3844 20856 3850 20868
rect 4264 20856 4292 20896
rect 4525 20893 4537 20896
rect 4571 20893 4583 20927
rect 4525 20887 4583 20893
rect 4614 20884 4620 20936
rect 4672 20924 4678 20936
rect 5000 20933 5028 20964
rect 5552 20964 5764 20992
rect 5552 20933 5580 20964
rect 5810 20952 5816 21004
rect 5868 20992 5874 21004
rect 11808 20992 11836 21091
rect 12250 21088 12256 21140
rect 12308 21128 12314 21140
rect 12437 21131 12495 21137
rect 12437 21128 12449 21131
rect 12308 21100 12449 21128
rect 12308 21088 12314 21100
rect 12437 21097 12449 21100
rect 12483 21097 12495 21131
rect 12437 21091 12495 21097
rect 12894 21088 12900 21140
rect 12952 21088 12958 21140
rect 13078 21088 13084 21140
rect 13136 21128 13142 21140
rect 13446 21128 13452 21140
rect 13136 21100 13452 21128
rect 13136 21088 13142 21100
rect 13446 21088 13452 21100
rect 13504 21088 13510 21140
rect 14642 21088 14648 21140
rect 14700 21128 14706 21140
rect 14829 21131 14887 21137
rect 14829 21128 14841 21131
rect 14700 21100 14841 21128
rect 14700 21088 14706 21100
rect 14829 21097 14841 21100
rect 14875 21097 14887 21131
rect 14829 21091 14887 21097
rect 16114 21088 16120 21140
rect 16172 21088 16178 21140
rect 12158 21020 12164 21072
rect 12216 21060 12222 21072
rect 12802 21060 12808 21072
rect 12216 21032 12808 21060
rect 12216 21020 12222 21032
rect 12802 21020 12808 21032
rect 12860 21060 12866 21072
rect 13265 21063 13323 21069
rect 12860 21032 13032 21060
rect 12860 21020 12866 21032
rect 13004 21001 13032 21032
rect 13265 21029 13277 21063
rect 13311 21060 13323 21063
rect 13538 21060 13544 21072
rect 13311 21032 13544 21060
rect 13311 21029 13323 21032
rect 13265 21023 13323 21029
rect 13538 21020 13544 21032
rect 13596 21060 13602 21072
rect 13596 21032 14136 21060
rect 13596 21020 13602 21032
rect 12989 20995 13047 21001
rect 5868 20964 8984 20992
rect 11808 20964 12940 20992
rect 5868 20952 5874 20964
rect 4801 20927 4859 20933
rect 4801 20924 4813 20927
rect 4672 20896 4813 20924
rect 4672 20884 4678 20896
rect 4801 20893 4813 20896
rect 4847 20893 4859 20927
rect 4801 20887 4859 20893
rect 4985 20927 5043 20933
rect 4985 20893 4997 20927
rect 5031 20893 5043 20927
rect 4985 20887 5043 20893
rect 5537 20927 5595 20933
rect 5537 20893 5549 20927
rect 5583 20893 5595 20927
rect 5537 20887 5595 20893
rect 5721 20927 5779 20933
rect 5721 20893 5733 20927
rect 5767 20924 5779 20927
rect 5902 20924 5908 20936
rect 5767 20896 5908 20924
rect 5767 20893 5779 20896
rect 5721 20887 5779 20893
rect 5902 20884 5908 20896
rect 5960 20884 5966 20936
rect 6089 20927 6147 20933
rect 6089 20893 6101 20927
rect 6135 20893 6147 20927
rect 6089 20887 6147 20893
rect 6365 20927 6423 20933
rect 6365 20893 6377 20927
rect 6411 20924 6423 20927
rect 6822 20924 6828 20936
rect 6411 20896 6828 20924
rect 6411 20893 6423 20896
rect 6365 20887 6423 20893
rect 3844 20828 4292 20856
rect 4367 20859 4425 20865
rect 3844 20816 3850 20828
rect 4367 20825 4379 20859
rect 4413 20856 4425 20859
rect 4706 20856 4712 20868
rect 4413 20828 4712 20856
rect 4413 20825 4425 20828
rect 4367 20819 4425 20825
rect 4706 20816 4712 20828
rect 4764 20816 4770 20868
rect 6104 20856 6132 20887
rect 6822 20884 6828 20896
rect 6880 20884 6886 20936
rect 7009 20927 7067 20933
rect 7009 20893 7021 20927
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 6178 20856 6184 20868
rect 5644 20828 6040 20856
rect 6104 20828 6184 20856
rect 5644 20788 5672 20828
rect 3712 20760 5672 20788
rect 5718 20748 5724 20800
rect 5776 20748 5782 20800
rect 6012 20788 6040 20828
rect 6178 20816 6184 20828
rect 6236 20856 6242 20868
rect 7024 20856 7052 20887
rect 7282 20884 7288 20936
rect 7340 20884 7346 20936
rect 7377 20927 7435 20933
rect 7377 20893 7389 20927
rect 7423 20924 7435 20927
rect 7466 20924 7472 20936
rect 7423 20896 7472 20924
rect 7423 20893 7435 20896
rect 7377 20887 7435 20893
rect 7466 20884 7472 20896
rect 7524 20884 7530 20936
rect 7558 20884 7564 20936
rect 7616 20884 7622 20936
rect 8956 20933 8984 20964
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 11701 20927 11759 20933
rect 11701 20893 11713 20927
rect 11747 20924 11759 20927
rect 11790 20924 11796 20936
rect 11747 20896 11796 20924
rect 11747 20893 11759 20896
rect 11701 20887 11759 20893
rect 11790 20884 11796 20896
rect 11848 20924 11854 20936
rect 12158 20924 12164 20936
rect 11848 20896 12164 20924
rect 11848 20884 11854 20896
rect 12158 20884 12164 20896
rect 12216 20924 12222 20936
rect 12912 20933 12940 20964
rect 12989 20961 13001 20995
rect 13035 20961 13047 20995
rect 12989 20955 13047 20961
rect 13096 20964 13584 20992
rect 12897 20927 12955 20933
rect 12216 20896 12848 20924
rect 12216 20884 12222 20896
rect 7834 20856 7840 20868
rect 6236 20828 7840 20856
rect 6236 20816 6242 20828
rect 7834 20816 7840 20828
rect 7892 20816 7898 20868
rect 8386 20816 8392 20868
rect 8444 20816 8450 20868
rect 9766 20856 9772 20868
rect 8496 20828 9772 20856
rect 8496 20788 8524 20828
rect 9766 20816 9772 20828
rect 9824 20816 9830 20868
rect 12820 20856 12848 20896
rect 12897 20893 12909 20927
rect 12943 20893 12955 20927
rect 13096 20924 13124 20964
rect 13556 20933 13584 20964
rect 14108 20933 14136 21032
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 13357 20927 13415 20933
rect 13357 20924 13369 20927
rect 12897 20887 12955 20893
rect 13004 20896 13124 20924
rect 13188 20896 13369 20924
rect 13004 20856 13032 20896
rect 12268 20828 12756 20856
rect 12820 20828 13032 20856
rect 12268 20800 12296 20828
rect 6012 20760 8524 20788
rect 8570 20748 8576 20800
rect 8628 20797 8634 20800
rect 8628 20791 8647 20797
rect 8635 20757 8647 20791
rect 8628 20751 8647 20757
rect 8628 20748 8634 20751
rect 8754 20748 8760 20800
rect 8812 20748 8818 20800
rect 12250 20748 12256 20800
rect 12308 20748 12314 20800
rect 12434 20748 12440 20800
rect 12492 20748 12498 20800
rect 12728 20788 12756 20828
rect 13188 20788 13216 20896
rect 13357 20893 13369 20896
rect 13403 20893 13415 20927
rect 13357 20887 13415 20893
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20893 13599 20927
rect 13541 20887 13599 20893
rect 14093 20927 14151 20933
rect 14093 20893 14105 20927
rect 14139 20893 14151 20927
rect 14093 20887 14151 20893
rect 14182 20884 14188 20936
rect 14240 20924 14246 20936
rect 15197 20927 15255 20933
rect 14240 20896 14285 20924
rect 14240 20884 14246 20896
rect 15197 20893 15209 20927
rect 15243 20924 15255 20927
rect 15838 20924 15844 20936
rect 15243 20896 15844 20924
rect 15243 20893 15255 20896
rect 15197 20887 15255 20893
rect 15838 20884 15844 20896
rect 15896 20884 15902 20936
rect 15930 20884 15936 20936
rect 15988 20884 15994 20936
rect 12728 20760 13216 20788
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14461 20791 14519 20797
rect 14461 20788 14473 20791
rect 13872 20760 14473 20788
rect 13872 20748 13878 20760
rect 14461 20757 14473 20760
rect 14507 20757 14519 20791
rect 14461 20751 14519 20757
rect 15010 20748 15016 20800
rect 15068 20788 15074 20800
rect 15289 20791 15347 20797
rect 15289 20788 15301 20791
rect 15068 20760 15301 20788
rect 15068 20748 15074 20760
rect 15289 20757 15301 20760
rect 15335 20757 15347 20791
rect 15289 20751 15347 20757
rect 1104 20698 16836 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 16836 20698
rect 1104 20624 16836 20646
rect 1486 20544 1492 20596
rect 1544 20544 1550 20596
rect 3142 20544 3148 20596
rect 3200 20584 3206 20596
rect 3421 20587 3479 20593
rect 3421 20584 3433 20587
rect 3200 20556 3433 20584
rect 3200 20544 3206 20556
rect 3421 20553 3433 20556
rect 3467 20553 3479 20587
rect 3421 20547 3479 20553
rect 6178 20544 6184 20596
rect 6236 20544 6242 20596
rect 6362 20544 6368 20596
rect 6420 20584 6426 20596
rect 6457 20587 6515 20593
rect 6457 20584 6469 20587
rect 6420 20556 6469 20584
rect 6420 20544 6426 20556
rect 6457 20553 6469 20556
rect 6503 20553 6515 20587
rect 6457 20547 6515 20553
rect 6822 20544 6828 20596
rect 6880 20584 6886 20596
rect 7009 20587 7067 20593
rect 7009 20584 7021 20587
rect 6880 20556 7021 20584
rect 6880 20544 6886 20556
rect 7009 20553 7021 20556
rect 7055 20553 7067 20587
rect 7466 20584 7472 20596
rect 7009 20547 7067 20553
rect 7116 20556 7472 20584
rect 1762 20476 1768 20528
rect 1820 20476 1826 20528
rect 1854 20476 1860 20528
rect 1912 20476 1918 20528
rect 1995 20519 2053 20525
rect 1995 20485 2007 20519
rect 2041 20516 2053 20519
rect 2314 20516 2320 20528
rect 2041 20488 2320 20516
rect 2041 20485 2053 20488
rect 1995 20479 2053 20485
rect 2314 20476 2320 20488
rect 2372 20476 2378 20528
rect 2866 20516 2872 20528
rect 2792 20488 2872 20516
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20417 1731 20451
rect 1673 20411 1731 20417
rect 1688 20380 1716 20411
rect 2130 20408 2136 20460
rect 2188 20408 2194 20460
rect 2501 20451 2559 20457
rect 2501 20417 2513 20451
rect 2547 20448 2559 20451
rect 2682 20448 2688 20460
rect 2547 20420 2688 20448
rect 2547 20417 2559 20420
rect 2501 20411 2559 20417
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 2792 20457 2820 20488
rect 2866 20476 2872 20488
rect 2924 20476 2930 20528
rect 3510 20516 3516 20528
rect 2976 20488 3516 20516
rect 2976 20457 3004 20488
rect 3510 20476 3516 20488
rect 3568 20516 3574 20528
rect 3568 20488 3740 20516
rect 3568 20476 3574 20488
rect 3712 20460 3740 20488
rect 5718 20476 5724 20528
rect 5776 20516 5782 20528
rect 5776 20488 6684 20516
rect 5776 20476 5782 20488
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20417 2835 20451
rect 2777 20411 2835 20417
rect 2961 20451 3019 20457
rect 2961 20417 2973 20451
rect 3007 20417 3019 20451
rect 2961 20411 3019 20417
rect 3050 20408 3056 20460
rect 3108 20408 3114 20460
rect 3694 20408 3700 20460
rect 3752 20408 3758 20460
rect 3786 20408 3792 20460
rect 3844 20448 3850 20460
rect 4801 20451 4859 20457
rect 4801 20448 4813 20451
rect 3844 20420 4813 20448
rect 3844 20408 3850 20420
rect 4801 20417 4813 20420
rect 4847 20417 4859 20451
rect 4801 20411 4859 20417
rect 5068 20451 5126 20457
rect 5068 20417 5080 20451
rect 5114 20448 5126 20451
rect 5114 20420 5948 20448
rect 5114 20417 5126 20420
rect 5068 20411 5126 20417
rect 1946 20380 1952 20392
rect 1688 20352 1952 20380
rect 1946 20340 1952 20352
rect 2004 20380 2010 20392
rect 2869 20383 2927 20389
rect 2004 20352 2452 20380
rect 2004 20340 2010 20352
rect 1302 20272 1308 20324
rect 1360 20312 1366 20324
rect 2317 20315 2375 20321
rect 2317 20312 2329 20315
rect 1360 20284 2329 20312
rect 1360 20272 1366 20284
rect 2317 20281 2329 20284
rect 2363 20281 2375 20315
rect 2424 20312 2452 20352
rect 2869 20349 2881 20383
rect 2915 20380 2927 20383
rect 3142 20380 3148 20392
rect 2915 20352 3148 20380
rect 2915 20349 2927 20352
rect 2869 20343 2927 20349
rect 3142 20340 3148 20352
rect 3200 20380 3206 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3200 20352 3433 20380
rect 3200 20340 3206 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 3602 20340 3608 20392
rect 3660 20380 3666 20392
rect 4617 20383 4675 20389
rect 4617 20380 4629 20383
rect 3660 20352 4629 20380
rect 3660 20340 3666 20352
rect 4617 20349 4629 20352
rect 4663 20349 4675 20383
rect 5920 20380 5948 20420
rect 6362 20408 6368 20460
rect 6420 20408 6426 20460
rect 6656 20457 6684 20488
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 6917 20451 6975 20457
rect 6917 20417 6929 20451
rect 6963 20448 6975 20451
rect 7006 20448 7012 20460
rect 6963 20420 7012 20448
rect 6963 20417 6975 20420
rect 6917 20411 6975 20417
rect 7006 20408 7012 20420
rect 7064 20408 7070 20460
rect 7116 20457 7144 20556
rect 7466 20544 7472 20556
rect 7524 20584 7530 20596
rect 8573 20587 8631 20593
rect 8573 20584 8585 20587
rect 7524 20556 8585 20584
rect 7524 20544 7530 20556
rect 8573 20553 8585 20556
rect 8619 20553 8631 20587
rect 8573 20547 8631 20553
rect 9858 20544 9864 20596
rect 9916 20593 9922 20596
rect 9916 20587 9935 20593
rect 9923 20553 9935 20587
rect 9916 20547 9935 20553
rect 9916 20544 9922 20547
rect 11238 20544 11244 20596
rect 11296 20584 11302 20596
rect 11882 20584 11888 20596
rect 11296 20556 11888 20584
rect 11296 20544 11302 20556
rect 11882 20544 11888 20556
rect 11940 20584 11946 20596
rect 13630 20584 13636 20596
rect 11940 20556 13636 20584
rect 11940 20544 11946 20556
rect 13630 20544 13636 20556
rect 13688 20584 13694 20596
rect 14185 20587 14243 20593
rect 13688 20556 13952 20584
rect 13688 20544 13694 20556
rect 9674 20476 9680 20528
rect 9732 20476 9738 20528
rect 11790 20476 11796 20528
rect 11848 20516 11854 20528
rect 11974 20516 11980 20528
rect 11848 20488 11980 20516
rect 11848 20476 11854 20488
rect 11974 20476 11980 20488
rect 12032 20516 12038 20528
rect 12032 20488 13860 20516
rect 12032 20476 12038 20488
rect 13832 20460 13860 20488
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20417 7159 20451
rect 7101 20411 7159 20417
rect 7460 20451 7518 20457
rect 7460 20417 7472 20451
rect 7506 20448 7518 20451
rect 7742 20448 7748 20460
rect 7506 20420 7748 20448
rect 7506 20417 7518 20420
rect 7460 20411 7518 20417
rect 7742 20408 7748 20420
rect 7800 20408 7806 20460
rect 11514 20408 11520 20460
rect 11572 20408 11578 20460
rect 12250 20408 12256 20460
rect 12308 20448 12314 20460
rect 13081 20451 13139 20457
rect 13081 20448 13093 20451
rect 12308 20420 13093 20448
rect 12308 20408 12314 20420
rect 13081 20417 13093 20420
rect 13127 20417 13139 20451
rect 13081 20411 13139 20417
rect 13265 20451 13323 20457
rect 13265 20417 13277 20451
rect 13311 20448 13323 20451
rect 13446 20448 13452 20460
rect 13311 20420 13452 20448
rect 13311 20417 13323 20420
rect 13265 20411 13323 20417
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 13541 20451 13599 20457
rect 13541 20417 13553 20451
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 5920 20352 6837 20380
rect 4617 20343 4675 20349
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7190 20340 7196 20392
rect 7248 20340 7254 20392
rect 9214 20340 9220 20392
rect 9272 20380 9278 20392
rect 9401 20383 9459 20389
rect 9401 20380 9413 20383
rect 9272 20352 9413 20380
rect 9272 20340 9278 20352
rect 9401 20349 9413 20352
rect 9447 20349 9459 20383
rect 9401 20343 9459 20349
rect 9490 20340 9496 20392
rect 9548 20380 9554 20392
rect 10137 20383 10195 20389
rect 10137 20380 10149 20383
rect 9548 20352 10149 20380
rect 9548 20340 9554 20352
rect 10137 20349 10149 20352
rect 10183 20349 10195 20383
rect 10137 20343 10195 20349
rect 11793 20383 11851 20389
rect 11793 20349 11805 20383
rect 11839 20380 11851 20383
rect 12268 20380 12296 20408
rect 11839 20352 12296 20380
rect 11839 20349 11851 20352
rect 11793 20343 11851 20349
rect 13170 20340 13176 20392
rect 13228 20380 13234 20392
rect 13556 20380 13584 20411
rect 13722 20408 13728 20460
rect 13780 20408 13786 20460
rect 13814 20408 13820 20460
rect 13872 20408 13878 20460
rect 13924 20457 13952 20556
rect 14185 20553 14197 20587
rect 14231 20584 14243 20587
rect 15378 20584 15384 20596
rect 14231 20556 15384 20584
rect 14231 20553 14243 20556
rect 14185 20547 14243 20553
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 13909 20451 13967 20457
rect 13909 20417 13921 20451
rect 13955 20417 13967 20451
rect 13909 20411 13967 20417
rect 14553 20451 14611 20457
rect 14553 20417 14565 20451
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 13228 20352 13584 20380
rect 13228 20340 13234 20352
rect 3237 20315 3295 20321
rect 3237 20312 3249 20315
rect 2424 20284 3249 20312
rect 2317 20275 2375 20281
rect 3237 20281 3249 20284
rect 3283 20312 3295 20315
rect 3326 20312 3332 20324
rect 3283 20284 3332 20312
rect 3283 20281 3295 20284
rect 3237 20275 3295 20281
rect 3326 20272 3332 20284
rect 3384 20312 3390 20324
rect 10045 20315 10103 20321
rect 3384 20284 4200 20312
rect 3384 20272 3390 20284
rect 3602 20204 3608 20256
rect 3660 20204 3666 20256
rect 3694 20204 3700 20256
rect 3752 20244 3758 20256
rect 4065 20247 4123 20253
rect 4065 20244 4077 20247
rect 3752 20216 4077 20244
rect 3752 20204 3758 20216
rect 4065 20213 4077 20216
rect 4111 20213 4123 20247
rect 4172 20244 4200 20284
rect 10045 20281 10057 20315
rect 10091 20312 10103 20315
rect 14458 20312 14464 20324
rect 10091 20284 14464 20312
rect 10091 20281 10103 20284
rect 10045 20275 10103 20281
rect 14458 20272 14464 20284
rect 14516 20312 14522 20324
rect 14568 20312 14596 20411
rect 15930 20340 15936 20392
rect 15988 20380 15994 20392
rect 16209 20383 16267 20389
rect 16209 20380 16221 20383
rect 15988 20352 16221 20380
rect 15988 20340 15994 20352
rect 16209 20349 16221 20352
rect 16255 20349 16267 20383
rect 16209 20343 16267 20349
rect 14516 20284 14596 20312
rect 14516 20272 14522 20284
rect 8386 20244 8392 20256
rect 4172 20216 8392 20244
rect 4065 20207 4123 20213
rect 8386 20204 8392 20216
rect 8444 20204 8450 20256
rect 8846 20204 8852 20256
rect 8904 20204 8910 20256
rect 9766 20204 9772 20256
rect 9824 20244 9830 20256
rect 9861 20247 9919 20253
rect 9861 20244 9873 20247
rect 9824 20216 9873 20244
rect 9824 20204 9830 20216
rect 9861 20213 9873 20216
rect 9907 20213 9919 20247
rect 9861 20207 9919 20213
rect 10778 20204 10784 20256
rect 10836 20204 10842 20256
rect 11514 20204 11520 20256
rect 11572 20244 11578 20256
rect 11609 20247 11667 20253
rect 11609 20244 11621 20247
rect 11572 20216 11621 20244
rect 11572 20204 11578 20216
rect 11609 20213 11621 20216
rect 11655 20213 11667 20247
rect 11609 20207 11667 20213
rect 11701 20247 11759 20253
rect 11701 20213 11713 20247
rect 11747 20244 11759 20247
rect 11974 20244 11980 20256
rect 11747 20216 11980 20244
rect 11747 20213 11759 20216
rect 11701 20207 11759 20213
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 13170 20204 13176 20256
rect 13228 20244 13234 20256
rect 13357 20247 13415 20253
rect 13357 20244 13369 20247
rect 13228 20216 13369 20244
rect 13228 20204 13234 20216
rect 13357 20213 13369 20216
rect 13403 20213 13415 20247
rect 13357 20207 13415 20213
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 13814 20244 13820 20256
rect 13504 20216 13820 20244
rect 13504 20204 13510 20216
rect 13814 20204 13820 20216
rect 13872 20244 13878 20256
rect 14369 20247 14427 20253
rect 14369 20244 14381 20247
rect 13872 20216 14381 20244
rect 13872 20204 13878 20216
rect 14369 20213 14381 20216
rect 14415 20213 14427 20247
rect 14369 20207 14427 20213
rect 15286 20204 15292 20256
rect 15344 20244 15350 20256
rect 15657 20247 15715 20253
rect 15657 20244 15669 20247
rect 15344 20216 15669 20244
rect 15344 20204 15350 20216
rect 15657 20213 15669 20216
rect 15703 20213 15715 20247
rect 15657 20207 15715 20213
rect 1104 20154 16836 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 16836 20154
rect 1104 20080 16836 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 2774 20040 2780 20052
rect 1627 20012 2780 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 2774 20000 2780 20012
rect 2832 20040 2838 20052
rect 2958 20040 2964 20052
rect 2832 20012 2964 20040
rect 2832 20000 2838 20012
rect 2958 20000 2964 20012
rect 3016 20000 3022 20052
rect 5169 20043 5227 20049
rect 5169 20040 5181 20043
rect 3252 20012 5181 20040
rect 3252 19984 3280 20012
rect 5169 20009 5181 20012
rect 5215 20009 5227 20043
rect 5169 20003 5227 20009
rect 6181 20043 6239 20049
rect 6181 20009 6193 20043
rect 6227 20040 6239 20043
rect 6362 20040 6368 20052
rect 6227 20012 6368 20040
rect 6227 20009 6239 20012
rect 6181 20003 6239 20009
rect 6362 20000 6368 20012
rect 6420 20000 6426 20052
rect 6457 20043 6515 20049
rect 6457 20009 6469 20043
rect 6503 20040 6515 20043
rect 7098 20040 7104 20052
rect 6503 20012 7104 20040
rect 6503 20009 6515 20012
rect 6457 20003 6515 20009
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7742 20000 7748 20052
rect 7800 20000 7806 20052
rect 8570 20000 8576 20052
rect 8628 20040 8634 20052
rect 8665 20043 8723 20049
rect 8665 20040 8677 20043
rect 8628 20012 8677 20040
rect 8628 20000 8634 20012
rect 8665 20009 8677 20012
rect 8711 20009 8723 20043
rect 8665 20003 8723 20009
rect 9125 20043 9183 20049
rect 9125 20009 9137 20043
rect 9171 20040 9183 20043
rect 9490 20040 9496 20052
rect 9171 20012 9496 20040
rect 9171 20009 9183 20012
rect 9125 20003 9183 20009
rect 9490 20000 9496 20012
rect 9548 20000 9554 20052
rect 15930 20000 15936 20052
rect 15988 20000 15994 20052
rect 3234 19972 3240 19984
rect 2148 19944 3240 19972
rect 842 19796 848 19848
rect 900 19836 906 19848
rect 1489 19839 1547 19845
rect 1489 19836 1501 19839
rect 900 19808 1501 19836
rect 900 19796 906 19808
rect 1489 19805 1501 19808
rect 1535 19805 1547 19839
rect 1489 19799 1547 19805
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19836 2007 19839
rect 2038 19836 2044 19848
rect 1995 19808 2044 19836
rect 1995 19805 2007 19808
rect 1949 19799 2007 19805
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 2148 19845 2176 19944
rect 3234 19932 3240 19944
rect 3292 19932 3298 19984
rect 7469 19975 7527 19981
rect 7469 19972 7481 19975
rect 6748 19944 7481 19972
rect 3142 19864 3148 19916
rect 3200 19864 3206 19916
rect 3786 19864 3792 19916
rect 3844 19864 3850 19916
rect 6748 19904 6776 19944
rect 7469 19941 7481 19944
rect 7515 19941 7527 19975
rect 7469 19935 7527 19941
rect 11609 19975 11667 19981
rect 11609 19941 11621 19975
rect 11655 19972 11667 19975
rect 12066 19972 12072 19984
rect 11655 19944 12072 19972
rect 11655 19941 11667 19944
rect 11609 19935 11667 19941
rect 12066 19932 12072 19944
rect 12124 19932 12130 19984
rect 13906 19972 13912 19984
rect 13280 19944 13912 19972
rect 7374 19904 7380 19916
rect 6288 19876 6776 19904
rect 2133 19839 2191 19845
rect 2133 19805 2145 19839
rect 2179 19805 2191 19839
rect 2133 19799 2191 19805
rect 2314 19796 2320 19848
rect 2372 19796 2378 19848
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 3694 19836 3700 19848
rect 3283 19808 3700 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 6288 19845 6316 19876
rect 6089 19839 6147 19845
rect 6089 19805 6101 19839
rect 6135 19805 6147 19839
rect 6089 19799 6147 19805
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19805 6331 19839
rect 6273 19799 6331 19805
rect 2056 19768 2084 19796
rect 3142 19768 3148 19780
rect 2056 19740 3148 19768
rect 3142 19728 3148 19740
rect 3200 19728 3206 19780
rect 4034 19771 4092 19777
rect 4034 19768 4046 19771
rect 3620 19740 4046 19768
rect 2130 19660 2136 19712
rect 2188 19660 2194 19712
rect 2866 19660 2872 19712
rect 2924 19660 2930 19712
rect 3620 19709 3648 19740
rect 4034 19737 4046 19740
rect 4080 19737 4092 19771
rect 6104 19768 6132 19799
rect 6638 19796 6644 19848
rect 6696 19796 6702 19848
rect 6748 19845 6776 19876
rect 6932 19876 7380 19904
rect 6733 19839 6791 19845
rect 6733 19805 6745 19839
rect 6779 19836 6791 19839
rect 6822 19836 6828 19848
rect 6779 19808 6828 19836
rect 6779 19805 6791 19808
rect 6733 19799 6791 19805
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 6932 19845 6960 19876
rect 7374 19864 7380 19876
rect 7432 19864 7438 19916
rect 10778 19864 10784 19916
rect 10836 19904 10842 19916
rect 11057 19907 11115 19913
rect 11057 19904 11069 19907
rect 10836 19876 11069 19904
rect 10836 19864 10842 19876
rect 11057 19873 11069 19876
rect 11103 19873 11115 19907
rect 11057 19867 11115 19873
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19904 11299 19907
rect 13081 19907 13139 19913
rect 13081 19904 13093 19907
rect 11287 19876 13093 19904
rect 11287 19873 11299 19876
rect 11241 19867 11299 19873
rect 13081 19873 13093 19876
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 7006 19796 7012 19848
rect 7064 19796 7070 19848
rect 7101 19839 7159 19845
rect 7101 19805 7113 19839
rect 7147 19805 7159 19839
rect 7101 19799 7159 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7466 19836 7472 19848
rect 7331 19808 7472 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 7116 19768 7144 19799
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 7558 19796 7564 19848
rect 7616 19796 7622 19848
rect 8757 19839 8815 19845
rect 8757 19805 8769 19839
rect 8803 19836 8815 19839
rect 8803 19808 9628 19836
rect 8803 19805 8815 19808
rect 8757 19799 8815 19805
rect 9600 19780 9628 19808
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 10505 19839 10563 19845
rect 10505 19836 10517 19839
rect 9916 19808 10517 19836
rect 9916 19796 9922 19808
rect 10505 19805 10517 19808
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 11790 19796 11796 19848
rect 11848 19796 11854 19848
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 13280 19845 13308 19944
rect 13906 19932 13912 19944
rect 13964 19932 13970 19984
rect 13357 19907 13415 19913
rect 13357 19873 13369 19907
rect 13403 19904 13415 19907
rect 13446 19904 13452 19916
rect 13403 19876 13452 19904
rect 13403 19873 13415 19876
rect 13357 19867 13415 19873
rect 13446 19864 13452 19876
rect 13504 19864 13510 19916
rect 13814 19904 13820 19916
rect 13556 19876 13820 19904
rect 13556 19845 13584 19876
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 11977 19839 12035 19845
rect 11977 19836 11989 19839
rect 11940 19808 11989 19836
rect 11940 19796 11946 19808
rect 11977 19805 11989 19808
rect 12023 19805 12035 19839
rect 11977 19799 12035 19805
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19805 13047 19839
rect 12989 19799 13047 19805
rect 13173 19839 13231 19845
rect 13173 19805 13185 19839
rect 13219 19805 13231 19839
rect 13173 19799 13231 19805
rect 13265 19839 13323 19845
rect 13265 19805 13277 19839
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 6104 19740 7144 19768
rect 4034 19731 4092 19737
rect 6748 19712 6776 19740
rect 9582 19728 9588 19780
rect 9640 19728 9646 19780
rect 10260 19771 10318 19777
rect 10260 19737 10272 19771
rect 10306 19768 10318 19771
rect 10965 19771 11023 19777
rect 10306 19740 10640 19768
rect 10306 19737 10318 19740
rect 10260 19731 10318 19737
rect 3605 19703 3663 19709
rect 3605 19669 3617 19703
rect 3651 19669 3663 19703
rect 3605 19663 3663 19669
rect 6730 19660 6736 19712
rect 6788 19660 6794 19712
rect 10612 19709 10640 19740
rect 10965 19737 10977 19771
rect 11011 19768 11023 19771
rect 11808 19768 11836 19796
rect 11011 19740 11836 19768
rect 11011 19737 11023 19740
rect 10965 19731 11023 19737
rect 10597 19703 10655 19709
rect 10597 19669 10609 19703
rect 10643 19669 10655 19703
rect 10597 19663 10655 19669
rect 11698 19660 11704 19712
rect 11756 19700 11762 19712
rect 11885 19703 11943 19709
rect 11885 19700 11897 19703
rect 11756 19672 11897 19700
rect 11756 19660 11762 19672
rect 11885 19669 11897 19672
rect 11931 19669 11943 19703
rect 13004 19700 13032 19799
rect 13188 19768 13216 19799
rect 13354 19768 13360 19780
rect 13188 19740 13360 19768
rect 13354 19728 13360 19740
rect 13412 19768 13418 19780
rect 13648 19768 13676 19799
rect 14550 19796 14556 19848
rect 14608 19796 14614 19848
rect 13412 19740 13676 19768
rect 14820 19771 14878 19777
rect 13412 19728 13418 19740
rect 14820 19737 14832 19771
rect 14866 19768 14878 19771
rect 14918 19768 14924 19780
rect 14866 19740 14924 19768
rect 14866 19737 14878 19740
rect 14820 19731 14878 19737
rect 14918 19728 14924 19740
rect 14976 19728 14982 19780
rect 13446 19700 13452 19712
rect 13004 19672 13452 19700
rect 11885 19663 11943 19669
rect 13446 19660 13452 19672
rect 13504 19660 13510 19712
rect 13817 19703 13875 19709
rect 13817 19669 13829 19703
rect 13863 19700 13875 19703
rect 15470 19700 15476 19712
rect 13863 19672 15476 19700
rect 13863 19669 13875 19672
rect 13817 19663 13875 19669
rect 15470 19660 15476 19672
rect 15528 19660 15534 19712
rect 1104 19610 16836 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 16836 19610
rect 1104 19536 16836 19558
rect 3142 19456 3148 19508
rect 3200 19456 3206 19508
rect 3234 19456 3240 19508
rect 3292 19456 3298 19508
rect 6638 19456 6644 19508
rect 6696 19496 6702 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 6696 19468 7021 19496
rect 6696 19456 6702 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 7377 19499 7435 19505
rect 7377 19465 7389 19499
rect 7423 19496 7435 19499
rect 9214 19496 9220 19508
rect 7423 19468 9220 19496
rect 7423 19465 7435 19468
rect 7377 19459 7435 19465
rect 9214 19456 9220 19468
rect 9272 19456 9278 19508
rect 11333 19499 11391 19505
rect 11333 19465 11345 19499
rect 11379 19496 11391 19499
rect 11422 19496 11428 19508
rect 11379 19468 11428 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 11422 19456 11428 19468
rect 11480 19456 11486 19508
rect 11517 19499 11575 19505
rect 11517 19465 11529 19499
rect 11563 19465 11575 19499
rect 11517 19459 11575 19465
rect 1664 19431 1722 19437
rect 1664 19397 1676 19431
rect 1710 19428 1722 19431
rect 3697 19431 3755 19437
rect 3697 19428 3709 19431
rect 1710 19400 3709 19428
rect 1710 19397 1722 19400
rect 1664 19391 1722 19397
rect 3697 19397 3709 19400
rect 3743 19397 3755 19431
rect 3697 19391 3755 19397
rect 7190 19388 7196 19440
rect 7248 19428 7254 19440
rect 8202 19428 8208 19440
rect 7248 19400 8208 19428
rect 7248 19388 7254 19400
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 2866 19320 2872 19372
rect 2924 19360 2930 19372
rect 3605 19363 3663 19369
rect 3605 19360 3617 19363
rect 2924 19332 3617 19360
rect 2924 19320 2930 19332
rect 3605 19329 3617 19332
rect 3651 19329 3663 19363
rect 3605 19323 3663 19329
rect 3789 19363 3847 19369
rect 3789 19329 3801 19363
rect 3835 19329 3847 19363
rect 3789 19323 3847 19329
rect 7469 19363 7527 19369
rect 7469 19329 7481 19363
rect 7515 19360 7527 19363
rect 7650 19360 7656 19372
rect 7515 19332 7656 19360
rect 7515 19329 7527 19332
rect 7469 19323 7527 19329
rect 3028 19295 3086 19301
rect 3028 19292 3040 19295
rect 2792 19264 3040 19292
rect 2792 19168 2820 19264
rect 3028 19261 3040 19264
rect 3074 19261 3086 19295
rect 3028 19255 3086 19261
rect 3510 19252 3516 19304
rect 3568 19252 3574 19304
rect 3694 19252 3700 19304
rect 3752 19292 3758 19304
rect 3804 19292 3832 19323
rect 7650 19320 7656 19332
rect 7708 19320 7714 19372
rect 7852 19369 7880 19400
rect 8202 19388 8208 19400
rect 8260 19388 8266 19440
rect 9766 19388 9772 19440
rect 9824 19428 9830 19440
rect 9861 19431 9919 19437
rect 9861 19428 9873 19431
rect 9824 19400 9873 19428
rect 9824 19388 9830 19400
rect 9861 19397 9873 19400
rect 9907 19397 9919 19431
rect 9861 19391 9919 19397
rect 10220 19431 10278 19437
rect 10220 19397 10232 19431
rect 10266 19428 10278 19431
rect 11532 19428 11560 19459
rect 11606 19456 11612 19508
rect 11664 19496 11670 19508
rect 11974 19496 11980 19508
rect 11664 19468 11980 19496
rect 11664 19456 11670 19468
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 13354 19456 13360 19508
rect 13412 19456 13418 19508
rect 13722 19456 13728 19508
rect 13780 19496 13786 19508
rect 13909 19499 13967 19505
rect 13909 19496 13921 19499
rect 13780 19468 13921 19496
rect 13780 19456 13786 19468
rect 13909 19465 13921 19468
rect 13955 19465 13967 19499
rect 13909 19459 13967 19465
rect 14918 19456 14924 19508
rect 14976 19456 14982 19508
rect 15286 19456 15292 19508
rect 15344 19456 15350 19508
rect 14553 19431 14611 19437
rect 14553 19428 14565 19431
rect 10266 19400 11560 19428
rect 13740 19400 14565 19428
rect 10266 19397 10278 19400
rect 10220 19391 10278 19397
rect 8110 19369 8116 19372
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 8104 19323 8116 19369
rect 8110 19320 8116 19323
rect 8168 19320 8174 19372
rect 9674 19320 9680 19372
rect 9732 19320 9738 19372
rect 11698 19320 11704 19372
rect 11756 19360 11762 19372
rect 11885 19363 11943 19369
rect 11885 19360 11897 19363
rect 11756 19332 11897 19360
rect 11756 19320 11762 19332
rect 11885 19329 11897 19332
rect 11931 19329 11943 19363
rect 11885 19323 11943 19329
rect 12250 19320 12256 19372
rect 12308 19360 12314 19372
rect 12897 19363 12955 19369
rect 12897 19360 12909 19363
rect 12308 19332 12909 19360
rect 12308 19320 12314 19332
rect 12897 19329 12909 19332
rect 12943 19329 12955 19363
rect 12897 19323 12955 19329
rect 13173 19363 13231 19369
rect 13173 19329 13185 19363
rect 13219 19360 13231 19363
rect 13262 19360 13268 19372
rect 13219 19332 13268 19360
rect 13219 19329 13231 19332
rect 13173 19323 13231 19329
rect 13262 19320 13268 19332
rect 13320 19320 13326 19372
rect 13538 19320 13544 19372
rect 13596 19320 13602 19372
rect 13630 19320 13636 19372
rect 13688 19360 13694 19372
rect 13740 19369 13768 19400
rect 14553 19397 14565 19400
rect 14599 19397 14611 19431
rect 14553 19391 14611 19397
rect 13725 19363 13783 19369
rect 13725 19360 13737 19363
rect 13688 19332 13737 19360
rect 13688 19320 13694 19332
rect 13725 19329 13737 19332
rect 13771 19329 13783 19363
rect 14277 19363 14335 19369
rect 14277 19360 14289 19363
rect 13725 19323 13783 19329
rect 13832 19332 14289 19360
rect 3752 19264 3832 19292
rect 7561 19295 7619 19301
rect 3752 19252 3758 19264
rect 7561 19261 7573 19295
rect 7607 19261 7619 19295
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 7561 19255 7619 19261
rect 9876 19264 9965 19292
rect 7576 19224 7604 19255
rect 9876 19236 9904 19264
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 9953 19255 10011 19261
rect 12066 19252 12072 19304
rect 12124 19292 12130 19304
rect 12526 19292 12532 19304
rect 12124 19264 12532 19292
rect 12124 19252 12130 19264
rect 12526 19252 12532 19264
rect 12584 19252 12590 19304
rect 13081 19295 13139 19301
rect 13081 19261 13093 19295
rect 13127 19292 13139 19295
rect 13354 19292 13360 19304
rect 13127 19264 13360 19292
rect 13127 19261 13139 19264
rect 13081 19255 13139 19261
rect 13354 19252 13360 19264
rect 13412 19292 13418 19304
rect 13556 19292 13584 19320
rect 13412 19264 13584 19292
rect 13412 19252 13418 19264
rect 7834 19224 7840 19236
rect 7576 19196 7840 19224
rect 7834 19184 7840 19196
rect 7892 19184 7898 19236
rect 8772 19196 9720 19224
rect 2774 19116 2780 19168
rect 2832 19116 2838 19168
rect 2866 19116 2872 19168
rect 2924 19116 2930 19168
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 8772 19156 8800 19196
rect 5316 19128 8800 19156
rect 5316 19116 5322 19128
rect 9582 19116 9588 19168
rect 9640 19116 9646 19168
rect 9692 19156 9720 19196
rect 9858 19184 9864 19236
rect 9916 19184 9922 19236
rect 12986 19184 12992 19236
rect 13044 19184 13050 19236
rect 13538 19184 13544 19236
rect 13596 19184 13602 19236
rect 13722 19184 13728 19236
rect 13780 19224 13786 19236
rect 13832 19224 13860 19332
rect 14277 19329 14289 19332
rect 14323 19329 14335 19363
rect 14277 19323 14335 19329
rect 14366 19320 14372 19372
rect 14424 19320 14430 19372
rect 14090 19252 14096 19304
rect 14148 19292 14154 19304
rect 14185 19295 14243 19301
rect 14185 19292 14197 19295
rect 14148 19264 14197 19292
rect 14148 19252 14154 19264
rect 14185 19261 14197 19264
rect 14231 19261 14243 19295
rect 14185 19255 14243 19261
rect 15378 19252 15384 19304
rect 15436 19252 15442 19304
rect 15470 19252 15476 19304
rect 15528 19252 15534 19304
rect 13780 19196 13860 19224
rect 13780 19184 13786 19196
rect 13906 19184 13912 19236
rect 13964 19224 13970 19236
rect 14734 19224 14740 19236
rect 13964 19196 14740 19224
rect 13964 19184 13970 19196
rect 14734 19184 14740 19196
rect 14792 19184 14798 19236
rect 13998 19156 14004 19168
rect 9692 19128 14004 19156
rect 13998 19116 14004 19128
rect 14056 19116 14062 19168
rect 14274 19116 14280 19168
rect 14332 19116 14338 19168
rect 1104 19066 16836 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 16836 19066
rect 1104 18992 16836 19014
rect 2130 18912 2136 18964
rect 2188 18952 2194 18964
rect 2225 18955 2283 18961
rect 2225 18952 2237 18955
rect 2188 18924 2237 18952
rect 2188 18912 2194 18924
rect 2225 18921 2237 18924
rect 2271 18921 2283 18955
rect 2225 18915 2283 18921
rect 2314 18912 2320 18964
rect 2372 18912 2378 18964
rect 5994 18912 6000 18964
rect 6052 18952 6058 18964
rect 6733 18955 6791 18961
rect 6733 18952 6745 18955
rect 6052 18924 6745 18952
rect 6052 18912 6058 18924
rect 6733 18921 6745 18924
rect 6779 18921 6791 18955
rect 6733 18915 6791 18921
rect 8021 18955 8079 18961
rect 8021 18921 8033 18955
rect 8067 18952 8079 18955
rect 8110 18952 8116 18964
rect 8067 18924 8116 18952
rect 8067 18921 8079 18924
rect 8021 18915 8079 18921
rect 8110 18912 8116 18924
rect 8168 18912 8174 18964
rect 12069 18955 12127 18961
rect 12069 18921 12081 18955
rect 12115 18952 12127 18955
rect 12250 18952 12256 18964
rect 12115 18924 12256 18952
rect 12115 18921 12127 18924
rect 12069 18915 12127 18921
rect 12250 18912 12256 18924
rect 12308 18912 12314 18964
rect 13354 18912 13360 18964
rect 13412 18912 13418 18964
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 13633 18955 13691 18961
rect 13633 18952 13645 18955
rect 13504 18924 13645 18952
rect 13504 18912 13510 18924
rect 13633 18921 13645 18924
rect 13679 18921 13691 18955
rect 14090 18952 14096 18964
rect 13633 18915 13691 18921
rect 13924 18924 14096 18952
rect 6641 18887 6699 18893
rect 6641 18853 6653 18887
rect 6687 18884 6699 18887
rect 6687 18856 7328 18884
rect 6687 18853 6699 18856
rect 6641 18847 6699 18853
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18816 2467 18819
rect 2501 18819 2559 18825
rect 2501 18816 2513 18819
rect 2455 18788 2513 18816
rect 2455 18785 2467 18788
rect 2409 18779 2467 18785
rect 2501 18785 2513 18788
rect 2547 18785 2559 18819
rect 2501 18779 2559 18785
rect 3786 18776 3792 18828
rect 3844 18816 3850 18828
rect 7300 18825 7328 18856
rect 8570 18844 8576 18896
rect 8628 18884 8634 18896
rect 8628 18856 9352 18884
rect 8628 18844 8634 18856
rect 5261 18819 5319 18825
rect 5261 18816 5273 18819
rect 3844 18788 5273 18816
rect 3844 18776 3850 18788
rect 5261 18785 5273 18788
rect 5307 18785 5319 18819
rect 5261 18779 5319 18785
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18816 7343 18819
rect 7466 18816 7472 18828
rect 7331 18788 7472 18816
rect 7331 18785 7343 18788
rect 7285 18779 7343 18785
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 8662 18776 8668 18828
rect 8720 18776 8726 18828
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 2148 18680 2176 18711
rect 2774 18708 2780 18760
rect 2832 18748 2838 18760
rect 3053 18751 3111 18757
rect 3053 18748 3065 18751
rect 2832 18720 3065 18748
rect 2832 18708 2838 18720
rect 3053 18717 3065 18720
rect 3099 18717 3111 18751
rect 3053 18711 3111 18717
rect 8481 18751 8539 18757
rect 8481 18717 8493 18751
rect 8527 18748 8539 18751
rect 8846 18748 8852 18760
rect 8527 18720 8852 18748
rect 8527 18717 8539 18720
rect 8481 18711 8539 18717
rect 8846 18708 8852 18720
rect 8904 18708 8910 18760
rect 9324 18757 9352 18856
rect 13262 18844 13268 18896
rect 13320 18884 13326 18896
rect 13924 18884 13952 18924
rect 14090 18912 14096 18924
rect 14148 18912 14154 18964
rect 15013 18955 15071 18961
rect 15013 18921 15025 18955
rect 15059 18952 15071 18955
rect 15378 18952 15384 18964
rect 15059 18924 15384 18952
rect 15059 18921 15071 18924
rect 15013 18915 15071 18921
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 13320 18856 13952 18884
rect 13320 18844 13326 18856
rect 13998 18844 14004 18896
rect 14056 18884 14062 18896
rect 14056 18856 14596 18884
rect 14056 18844 14062 18856
rect 9582 18776 9588 18828
rect 9640 18816 9646 18828
rect 10134 18816 10140 18828
rect 9640 18788 10140 18816
rect 9640 18776 9646 18788
rect 10134 18776 10140 18788
rect 10192 18776 10198 18828
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 11572 18788 12388 18816
rect 11572 18776 11578 18788
rect 12360 18760 12388 18788
rect 14458 18776 14464 18828
rect 14516 18776 14522 18828
rect 14568 18825 14596 18856
rect 14553 18819 14611 18825
rect 14553 18785 14565 18819
rect 14599 18785 14611 18819
rect 14553 18779 14611 18785
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 10778 18708 10784 18760
rect 10836 18708 10842 18760
rect 11425 18751 11483 18757
rect 11425 18717 11437 18751
rect 11471 18748 11483 18751
rect 12066 18748 12072 18760
rect 11471 18720 12072 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12342 18708 12348 18760
rect 12400 18708 12406 18760
rect 12526 18708 12532 18760
rect 12584 18708 12590 18760
rect 12986 18708 12992 18760
rect 13044 18748 13050 18760
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 13044 18720 13277 18748
rect 13044 18708 13050 18720
rect 13265 18717 13277 18720
rect 13311 18717 13323 18751
rect 13265 18711 13323 18717
rect 13354 18708 13360 18760
rect 13412 18708 13418 18760
rect 2958 18680 2964 18692
rect 2148 18652 2964 18680
rect 2958 18640 2964 18652
rect 3016 18680 3022 18692
rect 3510 18680 3516 18692
rect 3016 18652 3516 18680
rect 3016 18640 3022 18652
rect 3510 18640 3516 18652
rect 3568 18640 3574 18692
rect 5534 18689 5540 18692
rect 5528 18643 5540 18689
rect 5534 18640 5540 18643
rect 5592 18640 5598 18692
rect 8389 18683 8447 18689
rect 8389 18649 8401 18683
rect 8435 18680 8447 18683
rect 9401 18683 9459 18689
rect 8435 18652 8984 18680
rect 8435 18649 8447 18652
rect 8389 18643 8447 18649
rect 8956 18621 8984 18652
rect 9401 18649 9413 18683
rect 9447 18680 9459 18683
rect 9490 18680 9496 18692
rect 9447 18652 9496 18680
rect 9447 18649 9459 18652
rect 9401 18643 9459 18649
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 12158 18640 12164 18692
rect 12216 18680 12222 18692
rect 12253 18683 12311 18689
rect 12253 18680 12265 18683
rect 12216 18652 12265 18680
rect 12216 18640 12222 18652
rect 12253 18649 12265 18652
rect 12299 18649 12311 18683
rect 12894 18680 12900 18692
rect 12253 18643 12311 18649
rect 12360 18652 12900 18680
rect 8941 18615 8999 18621
rect 8941 18581 8953 18615
rect 8987 18581 8999 18615
rect 8941 18575 8999 18581
rect 11882 18572 11888 18624
rect 11940 18572 11946 18624
rect 12053 18615 12111 18621
rect 12053 18581 12065 18615
rect 12099 18612 12111 18615
rect 12360 18612 12388 18652
rect 12894 18640 12900 18652
rect 12952 18640 12958 18692
rect 12099 18584 12388 18612
rect 12099 18581 12111 18584
rect 12053 18575 12111 18581
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 13722 18612 13728 18624
rect 12492 18584 13728 18612
rect 12492 18572 12498 18584
rect 13722 18572 13728 18584
rect 13780 18572 13786 18624
rect 14642 18572 14648 18624
rect 14700 18572 14706 18624
rect 1104 18522 16836 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 16836 18522
rect 1104 18448 16836 18470
rect 2961 18411 3019 18417
rect 2961 18377 2973 18411
rect 3007 18408 3019 18411
rect 3050 18408 3056 18420
rect 3007 18380 3056 18408
rect 3007 18377 3019 18380
rect 2961 18371 3019 18377
rect 3050 18368 3056 18380
rect 3108 18408 3114 18420
rect 3694 18408 3700 18420
rect 3108 18380 3700 18408
rect 3108 18368 3114 18380
rect 3694 18368 3700 18380
rect 3752 18368 3758 18420
rect 5077 18411 5135 18417
rect 5077 18377 5089 18411
rect 5123 18408 5135 18411
rect 5258 18408 5264 18420
rect 5123 18380 5264 18408
rect 5123 18377 5135 18380
rect 5077 18371 5135 18377
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 5445 18411 5503 18417
rect 5445 18377 5457 18411
rect 5491 18408 5503 18411
rect 5534 18408 5540 18420
rect 5491 18380 5540 18408
rect 5491 18377 5503 18380
rect 5445 18371 5503 18377
rect 5534 18368 5540 18380
rect 5592 18368 5598 18420
rect 5813 18411 5871 18417
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 6457 18411 6515 18417
rect 6457 18408 6469 18411
rect 5859 18380 6469 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 6457 18377 6469 18380
rect 6503 18377 6515 18411
rect 6457 18371 6515 18377
rect 7466 18368 7472 18420
rect 7524 18417 7530 18420
rect 7524 18411 7543 18417
rect 7531 18377 7543 18411
rect 7524 18371 7543 18377
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 10778 18408 10784 18420
rect 9539 18380 10784 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 7524 18368 7530 18371
rect 2130 18300 2136 18352
rect 2188 18340 2194 18352
rect 5905 18343 5963 18349
rect 2188 18312 2636 18340
rect 2188 18300 2194 18312
rect 2608 18281 2636 18312
rect 5905 18309 5917 18343
rect 5951 18340 5963 18343
rect 5994 18340 6000 18352
rect 5951 18312 6000 18340
rect 5951 18309 5963 18312
rect 5905 18303 5963 18309
rect 5994 18300 6000 18312
rect 6052 18300 6058 18352
rect 7282 18300 7288 18352
rect 7340 18300 7346 18352
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18272 2099 18275
rect 2593 18275 2651 18281
rect 2087 18244 2544 18272
rect 2087 18241 2099 18244
rect 2041 18235 2099 18241
rect 2133 18207 2191 18213
rect 2133 18173 2145 18207
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 2148 18136 2176 18167
rect 2222 18164 2228 18216
rect 2280 18164 2286 18216
rect 2516 18204 2544 18244
rect 2593 18241 2605 18275
rect 2639 18241 2651 18275
rect 2593 18235 2651 18241
rect 2777 18275 2835 18281
rect 2777 18241 2789 18275
rect 2823 18272 2835 18275
rect 2958 18272 2964 18284
rect 2823 18244 2964 18272
rect 2823 18241 2835 18244
rect 2777 18235 2835 18241
rect 2958 18232 2964 18244
rect 3016 18232 3022 18284
rect 3697 18275 3755 18281
rect 3697 18241 3709 18275
rect 3743 18272 3755 18275
rect 3786 18272 3792 18284
rect 3743 18244 3792 18272
rect 3743 18241 3755 18244
rect 3697 18235 3755 18241
rect 3786 18232 3792 18244
rect 3844 18232 3850 18284
rect 3970 18281 3976 18284
rect 3964 18235 3976 18281
rect 3970 18232 3976 18235
rect 4028 18232 4034 18284
rect 6822 18232 6828 18284
rect 6880 18232 6886 18284
rect 6917 18275 6975 18281
rect 6917 18241 6929 18275
rect 6963 18272 6975 18275
rect 9508 18272 9536 18371
rect 10778 18368 10784 18380
rect 10836 18368 10842 18420
rect 11517 18411 11575 18417
rect 11517 18377 11529 18411
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 13633 18411 13691 18417
rect 13633 18377 13645 18411
rect 13679 18408 13691 18411
rect 14642 18408 14648 18420
rect 13679 18380 14648 18408
rect 13679 18377 13691 18380
rect 13633 18371 13691 18377
rect 10628 18343 10686 18349
rect 10628 18309 10640 18343
rect 10674 18340 10686 18343
rect 11532 18340 11560 18371
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 14921 18411 14979 18417
rect 14921 18377 14933 18411
rect 14967 18408 14979 18411
rect 15010 18408 15016 18420
rect 14967 18380 15016 18408
rect 14967 18377 14979 18380
rect 14921 18371 14979 18377
rect 15010 18368 15016 18380
rect 15068 18368 15074 18420
rect 10674 18312 11560 18340
rect 10674 18309 10686 18312
rect 10628 18303 10686 18309
rect 11790 18300 11796 18352
rect 11848 18300 11854 18352
rect 11885 18343 11943 18349
rect 11885 18309 11897 18343
rect 11931 18340 11943 18343
rect 12253 18343 12311 18349
rect 12253 18340 12265 18343
rect 11931 18312 12265 18340
rect 11931 18309 11943 18312
rect 11885 18303 11943 18309
rect 12253 18309 12265 18312
rect 12299 18309 12311 18343
rect 12253 18303 12311 18309
rect 12636 18312 14688 18340
rect 11701 18275 11759 18281
rect 6963 18244 9536 18272
rect 9692 18244 11008 18272
rect 6963 18241 6975 18244
rect 6917 18235 6975 18241
rect 2682 18204 2688 18216
rect 2516 18176 2688 18204
rect 2682 18164 2688 18176
rect 2740 18204 2746 18216
rect 3510 18204 3516 18216
rect 2740 18176 3516 18204
rect 2740 18164 2746 18176
rect 3510 18164 3516 18176
rect 3568 18164 3574 18216
rect 6086 18164 6092 18216
rect 6144 18164 6150 18216
rect 7101 18207 7159 18213
rect 7101 18173 7113 18207
rect 7147 18204 7159 18207
rect 9582 18204 9588 18216
rect 7147 18176 9588 18204
rect 7147 18173 7159 18176
rect 7101 18167 7159 18173
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 2958 18136 2964 18148
rect 2148 18108 2964 18136
rect 2958 18096 2964 18108
rect 3016 18136 3022 18148
rect 3418 18136 3424 18148
rect 3016 18108 3424 18136
rect 3016 18096 3022 18108
rect 3418 18096 3424 18108
rect 3476 18136 3482 18148
rect 9692 18136 9720 18244
rect 10873 18207 10931 18213
rect 10873 18173 10885 18207
rect 10919 18173 10931 18207
rect 10873 18167 10931 18173
rect 3476 18108 3740 18136
rect 3476 18096 3482 18108
rect 1670 18028 1676 18080
rect 1728 18028 1734 18080
rect 2774 18028 2780 18080
rect 2832 18028 2838 18080
rect 3712 18068 3740 18108
rect 4724 18108 9720 18136
rect 4724 18068 4752 18108
rect 3712 18040 4752 18068
rect 7466 18028 7472 18080
rect 7524 18028 7530 18080
rect 7653 18071 7711 18077
rect 7653 18037 7665 18071
rect 7699 18068 7711 18071
rect 8110 18068 8116 18080
rect 7699 18040 8116 18068
rect 7699 18037 7711 18040
rect 7653 18031 7711 18037
rect 8110 18028 8116 18040
rect 8168 18028 8174 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 10888 18068 10916 18167
rect 10980 18136 11008 18244
rect 11701 18241 11713 18275
rect 11747 18241 11759 18275
rect 11701 18235 11759 18241
rect 11716 18204 11744 18235
rect 12066 18232 12072 18284
rect 12124 18232 12130 18284
rect 12434 18232 12440 18284
rect 12492 18232 12498 18284
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 12250 18204 12256 18216
rect 11716 18176 12256 18204
rect 12250 18164 12256 18176
rect 12308 18164 12314 18216
rect 12636 18136 12664 18312
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18241 12771 18275
rect 12713 18235 12771 18241
rect 12728 18204 12756 18235
rect 12802 18232 12808 18284
rect 12860 18232 12866 18284
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13265 18275 13323 18281
rect 13265 18272 13277 18275
rect 13044 18244 13277 18272
rect 13044 18232 13050 18244
rect 13265 18241 13277 18244
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 13722 18232 13728 18284
rect 13780 18232 13786 18284
rect 13909 18275 13967 18281
rect 13909 18241 13921 18275
rect 13955 18272 13967 18275
rect 13998 18272 14004 18284
rect 13955 18244 14004 18272
rect 13955 18241 13967 18244
rect 13909 18235 13967 18241
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 14093 18275 14151 18281
rect 14093 18241 14105 18275
rect 14139 18272 14151 18275
rect 14369 18275 14427 18281
rect 14369 18272 14381 18275
rect 14139 18244 14381 18272
rect 14139 18241 14151 18244
rect 14093 18235 14151 18241
rect 14369 18241 14381 18244
rect 14415 18241 14427 18275
rect 14369 18235 14427 18241
rect 14458 18232 14464 18284
rect 14516 18272 14522 18284
rect 14660 18281 14688 18312
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14516 18244 14565 18272
rect 14516 18232 14522 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 14737 18275 14795 18281
rect 14737 18241 14749 18275
rect 14783 18241 14795 18275
rect 14737 18235 14795 18241
rect 13078 18204 13084 18216
rect 12728 18176 13084 18204
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 13357 18207 13415 18213
rect 13357 18173 13369 18207
rect 13403 18173 13415 18207
rect 13357 18167 13415 18173
rect 10980 18108 12664 18136
rect 13372 18136 13400 18167
rect 13814 18164 13820 18216
rect 13872 18204 13878 18216
rect 14274 18204 14280 18216
rect 13872 18176 14280 18204
rect 13872 18164 13878 18176
rect 14274 18164 14280 18176
rect 14332 18204 14338 18216
rect 14752 18204 14780 18235
rect 14332 18176 14780 18204
rect 14332 18164 14338 18176
rect 13998 18136 14004 18148
rect 13372 18108 14004 18136
rect 13998 18096 14004 18108
rect 14056 18096 14062 18148
rect 9916 18040 10916 18068
rect 9916 18028 9922 18040
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 12342 18068 12348 18080
rect 11940 18040 12348 18068
rect 11940 18028 11946 18040
rect 12342 18028 12348 18040
rect 12400 18068 12406 18080
rect 12802 18068 12808 18080
rect 12400 18040 12808 18068
rect 12400 18028 12406 18040
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 13449 18071 13507 18077
rect 13449 18037 13461 18071
rect 13495 18068 13507 18071
rect 14182 18068 14188 18080
rect 13495 18040 14188 18068
rect 13495 18037 13507 18040
rect 13449 18031 13507 18037
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 1104 17978 16836 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 16836 17978
rect 1104 17904 16836 17926
rect 2777 17867 2835 17873
rect 2777 17833 2789 17867
rect 2823 17864 2835 17867
rect 2958 17864 2964 17876
rect 2823 17836 2964 17864
rect 2823 17833 2835 17836
rect 2777 17827 2835 17833
rect 2958 17824 2964 17836
rect 3016 17824 3022 17876
rect 3326 17824 3332 17876
rect 3384 17824 3390 17876
rect 3513 17867 3571 17873
rect 3513 17833 3525 17867
rect 3559 17864 3571 17867
rect 3602 17864 3608 17876
rect 3559 17836 3608 17864
rect 3559 17833 3571 17836
rect 3513 17827 3571 17833
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 3881 17867 3939 17873
rect 3881 17833 3893 17867
rect 3927 17864 3939 17867
rect 3970 17864 3976 17876
rect 3927 17836 3976 17864
rect 3927 17833 3939 17836
rect 3881 17827 3939 17833
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 8205 17867 8263 17873
rect 8205 17833 8217 17867
rect 8251 17864 8263 17867
rect 8294 17864 8300 17876
rect 8251 17836 8300 17864
rect 8251 17833 8263 17836
rect 8205 17827 8263 17833
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 12897 17867 12955 17873
rect 12897 17833 12909 17867
rect 12943 17833 12955 17867
rect 12897 17827 12955 17833
rect 1394 17688 1400 17740
rect 1452 17688 1458 17740
rect 3050 17728 3056 17740
rect 2884 17700 3056 17728
rect 1412 17660 1440 17688
rect 2774 17660 2780 17672
rect 1412 17632 2780 17660
rect 2774 17620 2780 17632
rect 2832 17620 2838 17672
rect 1670 17601 1676 17604
rect 1664 17592 1676 17601
rect 1631 17564 1676 17592
rect 1664 17555 1676 17564
rect 1670 17552 1676 17555
rect 1728 17552 1734 17604
rect 2222 17552 2228 17604
rect 2280 17592 2286 17604
rect 2884 17592 2912 17700
rect 3050 17688 3056 17700
rect 3108 17688 3114 17740
rect 3620 17728 3648 17824
rect 4433 17731 4491 17737
rect 4433 17728 4445 17731
rect 3620 17700 4445 17728
rect 4433 17697 4445 17700
rect 4479 17697 4491 17731
rect 4433 17691 4491 17697
rect 6178 17688 6184 17740
rect 6236 17728 6242 17740
rect 6641 17731 6699 17737
rect 6641 17728 6653 17731
rect 6236 17700 6653 17728
rect 6236 17688 6242 17700
rect 6641 17697 6653 17700
rect 6687 17728 6699 17731
rect 6822 17728 6828 17740
rect 6687 17700 6828 17728
rect 6687 17697 6699 17700
rect 6641 17691 6699 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 12158 17728 12164 17740
rect 12084 17700 12164 17728
rect 3510 17620 3516 17672
rect 3568 17660 3574 17672
rect 3970 17660 3976 17672
rect 3568 17632 3976 17660
rect 3568 17620 3574 17632
rect 3970 17620 3976 17632
rect 4028 17660 4034 17672
rect 4341 17663 4399 17669
rect 4341 17660 4353 17663
rect 4028 17632 4353 17660
rect 4028 17620 4034 17632
rect 4341 17629 4353 17632
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 8021 17663 8079 17669
rect 8021 17629 8033 17663
rect 8067 17629 8079 17663
rect 8021 17623 8079 17629
rect 2280 17564 2912 17592
rect 2280 17552 2286 17564
rect 3050 17552 3056 17604
rect 3108 17592 3114 17604
rect 3145 17595 3203 17601
rect 3145 17592 3157 17595
rect 3108 17564 3157 17592
rect 3108 17552 3114 17564
rect 3145 17561 3157 17564
rect 3191 17561 3203 17595
rect 3145 17555 3203 17561
rect 4249 17595 4307 17601
rect 4249 17561 4261 17595
rect 4295 17592 4307 17595
rect 5258 17592 5264 17604
rect 4295 17564 5264 17592
rect 4295 17561 4307 17564
rect 4249 17555 4307 17561
rect 5258 17552 5264 17564
rect 5316 17552 5322 17604
rect 7745 17595 7803 17601
rect 7745 17561 7757 17595
rect 7791 17592 7803 17595
rect 7834 17592 7840 17604
rect 7791 17564 7840 17592
rect 7791 17561 7803 17564
rect 7745 17555 7803 17561
rect 7834 17552 7840 17564
rect 7892 17552 7898 17604
rect 8036 17592 8064 17623
rect 8110 17620 8116 17672
rect 8168 17660 8174 17672
rect 12084 17669 12112 17700
rect 12158 17688 12164 17700
rect 12216 17728 12222 17740
rect 12912 17728 12940 17827
rect 12986 17824 12992 17876
rect 13044 17864 13050 17876
rect 13081 17867 13139 17873
rect 13081 17864 13093 17867
rect 13044 17836 13093 17864
rect 13044 17824 13050 17836
rect 13081 17833 13093 17836
rect 13127 17833 13139 17867
rect 13081 17827 13139 17833
rect 12216 17700 12940 17728
rect 12216 17688 12222 17700
rect 14458 17688 14464 17740
rect 14516 17688 14522 17740
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 8168 17632 8217 17660
rect 8168 17620 8174 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 12069 17663 12127 17669
rect 12069 17629 12081 17663
rect 12115 17629 12127 17663
rect 12069 17623 12127 17629
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17660 12311 17663
rect 12986 17660 12992 17672
rect 12299 17632 12992 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 12928 17629 12992 17632
rect 8938 17592 8944 17604
rect 8036 17564 8944 17592
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 11882 17552 11888 17604
rect 11940 17552 11946 17604
rect 12526 17552 12532 17604
rect 12584 17592 12590 17604
rect 12713 17595 12771 17601
rect 12928 17598 12955 17629
rect 12713 17592 12725 17595
rect 12584 17564 12725 17592
rect 12584 17552 12590 17564
rect 12713 17561 12725 17564
rect 12759 17561 12771 17595
rect 12943 17595 12955 17598
rect 12989 17620 12992 17629
rect 13044 17620 13050 17672
rect 14182 17620 14188 17672
rect 14240 17620 14246 17672
rect 14274 17620 14280 17672
rect 14332 17620 14338 17672
rect 14737 17663 14795 17669
rect 14737 17629 14749 17663
rect 14783 17660 14795 17663
rect 14826 17660 14832 17672
rect 14783 17632 14832 17660
rect 14783 17629 14795 17632
rect 14737 17623 14795 17629
rect 14826 17620 14832 17632
rect 14884 17620 14890 17672
rect 16390 17620 16396 17672
rect 16448 17620 16454 17672
rect 12989 17595 13001 17620
rect 12943 17589 13001 17595
rect 12713 17555 12771 17561
rect 2866 17484 2872 17536
rect 2924 17524 2930 17536
rect 3345 17527 3403 17533
rect 3345 17524 3357 17527
rect 2924 17496 3357 17524
rect 2924 17484 2930 17496
rect 3345 17493 3357 17496
rect 3391 17493 3403 17527
rect 3345 17487 3403 17493
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 7193 17527 7251 17533
rect 7193 17524 7205 17527
rect 6788 17496 7205 17524
rect 6788 17484 6794 17496
rect 7193 17493 7205 17496
rect 7239 17493 7251 17527
rect 7193 17487 7251 17493
rect 8386 17484 8392 17536
rect 8444 17484 8450 17536
rect 12434 17484 12440 17536
rect 12492 17524 12498 17536
rect 13998 17524 14004 17536
rect 12492 17496 14004 17524
rect 12492 17484 12498 17496
rect 13998 17484 14004 17496
rect 14056 17524 14062 17536
rect 14645 17527 14703 17533
rect 14645 17524 14657 17527
rect 14056 17496 14657 17524
rect 14056 17484 14062 17496
rect 14645 17493 14657 17496
rect 14691 17493 14703 17527
rect 14645 17487 14703 17493
rect 15838 17484 15844 17536
rect 15896 17484 15902 17536
rect 1104 17434 16836 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 16836 17434
rect 1104 17360 16836 17382
rect 1857 17323 1915 17329
rect 1857 17289 1869 17323
rect 1903 17320 1915 17323
rect 2130 17320 2136 17332
rect 1903 17292 2136 17320
rect 1903 17289 1915 17292
rect 1857 17283 1915 17289
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 3326 17320 3332 17332
rect 2240 17292 3332 17320
rect 2240 17252 2268 17292
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 3694 17280 3700 17332
rect 3752 17320 3758 17332
rect 3752 17292 3832 17320
rect 3752 17280 3758 17292
rect 2774 17252 2780 17264
rect 2056 17224 2268 17252
rect 2332 17224 2780 17252
rect 2056 16989 2084 17224
rect 2222 17144 2228 17196
rect 2280 17144 2286 17196
rect 2332 17193 2360 17224
rect 2774 17212 2780 17224
rect 2832 17252 2838 17264
rect 3804 17261 3832 17292
rect 6178 17280 6184 17332
rect 6236 17280 6242 17332
rect 6365 17323 6423 17329
rect 6365 17289 6377 17323
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 3789 17255 3847 17261
rect 2832 17224 3740 17252
rect 2832 17212 2838 17224
rect 2317 17187 2375 17193
rect 2317 17153 2329 17187
rect 2363 17153 2375 17187
rect 2317 17147 2375 17153
rect 2584 17187 2642 17193
rect 2584 17153 2596 17187
rect 2630 17184 2642 17187
rect 2866 17184 2872 17196
rect 2630 17156 2872 17184
rect 2630 17153 2642 17156
rect 2584 17147 2642 17153
rect 2866 17144 2872 17156
rect 2924 17144 2930 17196
rect 3712 17184 3740 17224
rect 3789 17221 3801 17255
rect 3835 17221 3847 17255
rect 3789 17215 3847 17221
rect 3878 17212 3884 17264
rect 3936 17252 3942 17264
rect 3989 17255 4047 17261
rect 3989 17252 4001 17255
rect 3936 17224 4001 17252
rect 3936 17212 3942 17224
rect 3989 17221 4001 17224
rect 4035 17221 4047 17255
rect 3989 17215 4047 17221
rect 5068 17255 5126 17261
rect 5068 17221 5080 17255
rect 5114 17252 5126 17255
rect 6380 17252 6408 17283
rect 6730 17280 6736 17332
rect 6788 17280 6794 17332
rect 7006 17280 7012 17332
rect 7064 17320 7070 17332
rect 7561 17323 7619 17329
rect 7561 17320 7573 17323
rect 7064 17292 7573 17320
rect 7064 17280 7070 17292
rect 7561 17289 7573 17292
rect 7607 17289 7619 17323
rect 7561 17283 7619 17289
rect 8294 17280 8300 17332
rect 8352 17280 8358 17332
rect 8846 17320 8852 17332
rect 8404 17292 8852 17320
rect 8404 17252 8432 17292
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 8938 17280 8944 17332
rect 8996 17280 9002 17332
rect 11241 17323 11299 17329
rect 11241 17289 11253 17323
rect 11287 17320 11299 17323
rect 12158 17320 12164 17332
rect 11287 17292 12164 17320
rect 11287 17289 11299 17292
rect 11241 17283 11299 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12894 17280 12900 17332
rect 12952 17280 12958 17332
rect 13265 17323 13323 17329
rect 13265 17289 13277 17323
rect 13311 17320 13323 17323
rect 13354 17320 13360 17332
rect 13311 17292 13360 17320
rect 13311 17289 13323 17292
rect 13265 17283 13323 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 15930 17280 15936 17332
rect 15988 17320 15994 17332
rect 16117 17323 16175 17329
rect 16117 17320 16129 17323
rect 15988 17292 16129 17320
rect 15988 17280 15994 17292
rect 16117 17289 16129 17292
rect 16163 17320 16175 17323
rect 16390 17320 16396 17332
rect 16163 17292 16396 17320
rect 16163 17289 16175 17292
rect 16117 17283 16175 17289
rect 16390 17280 16396 17292
rect 16448 17280 16454 17332
rect 5114 17224 6408 17252
rect 7852 17224 8432 17252
rect 8481 17255 8539 17261
rect 5114 17221 5126 17224
rect 5068 17215 5126 17221
rect 3712 17156 3832 17184
rect 3804 17128 3832 17156
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7852 17193 7880 17224
rect 8481 17221 8493 17255
rect 8527 17252 8539 17255
rect 9766 17252 9772 17264
rect 8527 17224 9772 17252
rect 8527 17221 8539 17224
rect 8481 17215 8539 17221
rect 9766 17212 9772 17224
rect 9824 17212 9830 17264
rect 11885 17255 11943 17261
rect 11885 17221 11897 17255
rect 11931 17252 11943 17255
rect 12342 17252 12348 17264
rect 11931 17224 12348 17252
rect 11931 17221 11943 17224
rect 11885 17215 11943 17221
rect 12342 17212 12348 17224
rect 12400 17252 12406 17264
rect 12400 17224 13124 17252
rect 12400 17212 12406 17224
rect 7837 17187 7895 17193
rect 7837 17184 7849 17187
rect 7340 17156 7849 17184
rect 7340 17144 7346 17156
rect 7837 17153 7849 17156
rect 7883 17153 7895 17187
rect 7837 17147 7895 17153
rect 7929 17187 7987 17193
rect 7929 17153 7941 17187
rect 7975 17153 7987 17187
rect 7929 17147 7987 17153
rect 2133 17119 2191 17125
rect 2133 17085 2145 17119
rect 2179 17085 2191 17119
rect 2133 17079 2191 17085
rect 2041 16983 2099 16989
rect 2041 16949 2053 16983
rect 2087 16949 2099 16983
rect 2148 16980 2176 17079
rect 3786 17076 3792 17128
rect 3844 17116 3850 17128
rect 4801 17119 4859 17125
rect 4801 17116 4813 17119
rect 3844 17088 4813 17116
rect 3844 17076 3850 17088
rect 4801 17085 4813 17088
rect 4847 17085 4859 17119
rect 4801 17079 4859 17085
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 5868 17088 6837 17116
rect 5868 17076 5874 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 7009 17119 7067 17125
rect 7009 17085 7021 17119
rect 7055 17085 7067 17119
rect 7944 17116 7972 17147
rect 8018 17144 8024 17196
rect 8076 17144 8082 17196
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17184 8263 17187
rect 8386 17184 8392 17196
rect 8251 17156 8392 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 8386 17144 8392 17156
rect 8444 17144 8450 17196
rect 8846 17144 8852 17196
rect 8904 17144 8910 17196
rect 10128 17187 10186 17193
rect 10128 17153 10140 17187
rect 10174 17184 10186 17187
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 10174 17156 11529 17184
rect 10174 17153 10186 17156
rect 10128 17147 10186 17153
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 11790 17144 11796 17196
rect 11848 17144 11854 17196
rect 12003 17187 12061 17193
rect 12003 17184 12015 17187
rect 11900 17156 12015 17184
rect 9401 17119 9459 17125
rect 9401 17116 9413 17119
rect 7944 17088 9413 17116
rect 7009 17079 7067 17085
rect 3326 17008 3332 17060
rect 3384 17048 3390 17060
rect 7024 17048 7052 17079
rect 8294 17048 8300 17060
rect 3384 17020 4016 17048
rect 7024 17020 8300 17048
rect 3384 17008 3390 17020
rect 3050 16980 3056 16992
rect 2148 16952 3056 16980
rect 2041 16943 2099 16949
rect 3050 16940 3056 16952
rect 3108 16980 3114 16992
rect 3694 16980 3700 16992
rect 3108 16952 3700 16980
rect 3108 16940 3114 16952
rect 3694 16940 3700 16952
rect 3752 16940 3758 16992
rect 3988 16989 4016 17020
rect 8294 17008 8300 17020
rect 8352 17008 8358 17060
rect 8496 16992 8524 17088
rect 9401 17085 9413 17088
rect 9447 17085 9459 17119
rect 9401 17079 9459 17085
rect 9858 17076 9864 17128
rect 9916 17076 9922 17128
rect 11606 17076 11612 17128
rect 11664 17116 11670 17128
rect 11900 17116 11928 17156
rect 12003 17153 12015 17156
rect 12049 17153 12061 17187
rect 12003 17147 12061 17153
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12216 17156 12449 17184
rect 12216 17144 12222 17156
rect 12437 17153 12449 17156
rect 12483 17184 12495 17187
rect 12526 17184 12532 17196
rect 12483 17156 12532 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 12986 17144 12992 17196
rect 13044 17144 13050 17196
rect 13096 17193 13124 17224
rect 13081 17187 13139 17193
rect 13081 17153 13093 17187
rect 13127 17153 13139 17187
rect 13372 17184 13400 17280
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 14458 17252 14464 17264
rect 14240 17224 14464 17252
rect 14240 17212 14246 17224
rect 14458 17212 14464 17224
rect 14516 17212 14522 17264
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13372 17156 14013 17184
rect 13081 17147 13139 17153
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 14274 17144 14280 17196
rect 14332 17144 14338 17196
rect 14366 17144 14372 17196
rect 14424 17144 14430 17196
rect 14550 17144 14556 17196
rect 14608 17184 14614 17196
rect 15010 17193 15016 17196
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14608 17156 14749 17184
rect 14608 17144 14614 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 15004 17147 15016 17193
rect 15010 17144 15016 17147
rect 15068 17144 15074 17196
rect 16206 17144 16212 17196
rect 16264 17144 16270 17196
rect 11664 17088 11928 17116
rect 11664 17076 11670 17088
rect 9122 17008 9128 17060
rect 9180 17008 9186 17060
rect 12805 17051 12863 17057
rect 12805 17017 12817 17051
rect 12851 17048 12863 17051
rect 13004 17048 13032 17144
rect 13262 17076 13268 17128
rect 13320 17116 13326 17128
rect 13446 17116 13452 17128
rect 13320 17088 13452 17116
rect 13320 17076 13326 17088
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 12851 17020 13032 17048
rect 12851 17017 12863 17020
rect 12805 17011 12863 17017
rect 16390 17008 16396 17060
rect 16448 17008 16454 17060
rect 3973 16983 4031 16989
rect 3973 16949 3985 16983
rect 4019 16949 4031 16983
rect 3973 16943 4031 16949
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 4614 16980 4620 16992
rect 4203 16952 4620 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 8478 16940 8484 16992
rect 8536 16940 8542 16992
rect 11422 16940 11428 16992
rect 11480 16980 11486 16992
rect 12158 16980 12164 16992
rect 11480 16952 12164 16980
rect 11480 16940 11486 16952
rect 12158 16940 12164 16952
rect 12216 16940 12222 16992
rect 13262 16940 13268 16992
rect 13320 16980 13326 16992
rect 13538 16980 13544 16992
rect 13320 16952 13544 16980
rect 13320 16940 13326 16952
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 14553 16983 14611 16989
rect 14553 16949 14565 16983
rect 14599 16980 14611 16983
rect 15378 16980 15384 16992
rect 14599 16952 15384 16980
rect 14599 16949 14611 16952
rect 14553 16943 14611 16949
rect 15378 16940 15384 16952
rect 15436 16940 15442 16992
rect 1104 16890 16836 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 16836 16890
rect 1104 16816 16836 16838
rect 2866 16736 2872 16788
rect 2924 16736 2930 16788
rect 3513 16779 3571 16785
rect 3513 16745 3525 16779
rect 3559 16776 3571 16779
rect 3878 16776 3884 16788
rect 3559 16748 3884 16776
rect 3559 16745 3571 16748
rect 3513 16739 3571 16745
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 7561 16779 7619 16785
rect 7561 16776 7573 16779
rect 7524 16748 7573 16776
rect 7524 16736 7530 16748
rect 7561 16745 7573 16748
rect 7607 16776 7619 16779
rect 8478 16776 8484 16788
rect 7607 16748 8484 16776
rect 7607 16745 7619 16748
rect 7561 16739 7619 16745
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 11977 16779 12035 16785
rect 11977 16745 11989 16779
rect 12023 16776 12035 16779
rect 12066 16776 12072 16788
rect 12023 16748 12072 16776
rect 12023 16745 12035 16748
rect 11977 16739 12035 16745
rect 12066 16736 12072 16748
rect 12124 16776 12130 16788
rect 12342 16776 12348 16788
rect 12124 16748 12348 16776
rect 12124 16736 12130 16748
rect 12342 16736 12348 16748
rect 12400 16776 12406 16788
rect 13081 16779 13139 16785
rect 13081 16776 13093 16779
rect 12400 16748 13093 16776
rect 12400 16736 12406 16748
rect 13081 16745 13093 16748
rect 13127 16745 13139 16779
rect 13538 16776 13544 16788
rect 13081 16739 13139 16745
rect 13208 16748 13544 16776
rect 3142 16668 3148 16720
rect 3200 16668 3206 16720
rect 7193 16711 7251 16717
rect 7193 16677 7205 16711
rect 7239 16708 7251 16711
rect 7282 16708 7288 16720
rect 7239 16680 7288 16708
rect 7239 16677 7251 16680
rect 7193 16671 7251 16677
rect 7282 16668 7288 16680
rect 7340 16668 7346 16720
rect 8110 16668 8116 16720
rect 8168 16668 8174 16720
rect 8294 16668 8300 16720
rect 8352 16708 8358 16720
rect 8662 16708 8668 16720
rect 8352 16680 8668 16708
rect 8352 16668 8358 16680
rect 8662 16668 8668 16680
rect 8720 16668 8726 16720
rect 11241 16711 11299 16717
rect 11241 16677 11253 16711
rect 11287 16708 11299 16711
rect 13208 16708 13236 16748
rect 13538 16736 13544 16748
rect 13596 16776 13602 16788
rect 13596 16748 14596 16776
rect 13596 16736 13602 16748
rect 13998 16708 14004 16720
rect 11287 16680 11652 16708
rect 11287 16677 11299 16680
rect 11241 16671 11299 16677
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16640 2835 16643
rect 3160 16640 3188 16668
rect 3510 16640 3516 16652
rect 2823 16612 3096 16640
rect 3160 16612 3516 16640
rect 2823 16609 2835 16612
rect 2777 16603 2835 16609
rect 3068 16581 3096 16612
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3142 16532 3148 16584
rect 3200 16532 3206 16584
rect 3436 16581 3464 16612
rect 3510 16600 3516 16612
rect 3568 16600 3574 16652
rect 3786 16600 3792 16652
rect 3844 16640 3850 16652
rect 3973 16643 4031 16649
rect 3973 16640 3985 16643
rect 3844 16612 3985 16640
rect 3844 16600 3850 16612
rect 3973 16609 3985 16612
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 9582 16600 9588 16652
rect 9640 16600 9646 16652
rect 9858 16600 9864 16652
rect 9916 16600 9922 16652
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 10888 16612 11345 16640
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16541 7159 16575
rect 7101 16535 7159 16541
rect 10128 16575 10186 16581
rect 10128 16541 10140 16575
rect 10174 16572 10186 16575
rect 10888 16572 10916 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11333 16603 11391 16609
rect 10174 16544 10916 16572
rect 10174 16541 10186 16544
rect 10128 16535 10186 16541
rect 2409 16507 2467 16513
rect 2409 16473 2421 16507
rect 2455 16504 2467 16507
rect 2593 16507 2651 16513
rect 2455 16476 2544 16504
rect 2455 16473 2467 16476
rect 2409 16467 2467 16473
rect 2516 16448 2544 16476
rect 2593 16473 2605 16507
rect 2639 16504 2651 16507
rect 2866 16504 2872 16516
rect 2639 16476 2872 16504
rect 2639 16473 2651 16476
rect 2593 16467 2651 16473
rect 2866 16464 2872 16476
rect 2924 16464 2930 16516
rect 4062 16464 4068 16516
rect 4120 16504 4126 16516
rect 4218 16507 4276 16513
rect 4218 16504 4230 16507
rect 4120 16476 4230 16504
rect 4120 16464 4126 16476
rect 4218 16473 4230 16476
rect 4264 16473 4276 16507
rect 7116 16504 7144 16535
rect 11514 16532 11520 16584
rect 11572 16532 11578 16584
rect 11624 16581 11652 16680
rect 13096 16680 13236 16708
rect 13280 16680 14004 16708
rect 13096 16652 13124 16680
rect 12360 16612 12572 16640
rect 11609 16575 11667 16581
rect 11609 16541 11621 16575
rect 11655 16572 11667 16575
rect 11698 16572 11704 16584
rect 11655 16544 11704 16572
rect 11655 16541 11667 16544
rect 11609 16535 11667 16541
rect 11698 16532 11704 16544
rect 11756 16532 11762 16584
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 11885 16575 11943 16581
rect 11885 16541 11897 16575
rect 11931 16572 11943 16575
rect 11974 16572 11980 16584
rect 11931 16544 11980 16572
rect 11931 16541 11943 16544
rect 11885 16535 11943 16541
rect 7558 16504 7564 16516
rect 7116 16476 7564 16504
rect 4218 16467 4276 16473
rect 7558 16464 7564 16476
rect 7616 16464 7622 16516
rect 8478 16464 8484 16516
rect 8536 16504 8542 16516
rect 9030 16504 9036 16516
rect 8536 16476 9036 16504
rect 8536 16464 8542 16476
rect 9030 16464 9036 16476
rect 9088 16464 9094 16516
rect 2498 16396 2504 16448
rect 2556 16436 2562 16448
rect 2958 16436 2964 16448
rect 2556 16408 2964 16436
rect 2556 16396 2562 16408
rect 2958 16396 2964 16408
rect 3016 16396 3022 16448
rect 5350 16396 5356 16448
rect 5408 16396 5414 16448
rect 6454 16396 6460 16448
rect 6512 16396 6518 16448
rect 7742 16396 7748 16448
rect 7800 16396 7806 16448
rect 8021 16439 8079 16445
rect 8021 16405 8033 16439
rect 8067 16436 8079 16439
rect 8294 16436 8300 16448
rect 8067 16408 8300 16436
rect 8067 16405 8079 16408
rect 8021 16399 8079 16405
rect 8294 16396 8300 16408
rect 8352 16396 8358 16448
rect 8938 16396 8944 16448
rect 8996 16396 9002 16448
rect 9306 16396 9312 16448
rect 9364 16396 9370 16448
rect 9401 16439 9459 16445
rect 9401 16405 9413 16439
rect 9447 16436 9459 16439
rect 9950 16436 9956 16448
rect 9447 16408 9956 16436
rect 9447 16405 9459 16408
rect 9401 16399 9459 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 11606 16396 11612 16448
rect 11664 16436 11670 16448
rect 11808 16436 11836 16535
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12158 16532 12164 16584
rect 12216 16532 12222 16584
rect 12360 16581 12388 16612
rect 12544 16584 12572 16612
rect 13078 16600 13084 16652
rect 13136 16600 13142 16652
rect 13280 16649 13308 16680
rect 13998 16668 14004 16680
rect 14056 16668 14062 16720
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16609 13323 16643
rect 13265 16603 13323 16609
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13872 16612 13921 16640
rect 13872 16600 13878 16612
rect 13909 16609 13921 16612
rect 13955 16640 13967 16643
rect 14461 16643 14519 16649
rect 14461 16640 14473 16643
rect 13955 16612 14473 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 14461 16609 14473 16612
rect 14507 16609 14519 16643
rect 14461 16603 14519 16609
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16541 12495 16575
rect 12437 16535 12495 16541
rect 11664 16408 11836 16436
rect 12176 16436 12204 16532
rect 12452 16436 12480 16535
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 12621 16575 12679 16581
rect 12621 16572 12633 16575
rect 12584 16544 12633 16572
rect 12584 16532 12590 16544
rect 12621 16541 12633 16544
rect 12667 16541 12679 16575
rect 12621 16535 12679 16541
rect 12986 16532 12992 16584
rect 13044 16532 13050 16584
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 13412 16544 13553 16572
rect 13412 16532 13418 16544
rect 13541 16541 13553 16544
rect 13587 16541 13599 16575
rect 13541 16535 13599 16541
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14277 16575 14335 16581
rect 14277 16541 14289 16575
rect 14323 16541 14335 16575
rect 14277 16535 14335 16541
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16572 14427 16575
rect 14568 16572 14596 16748
rect 15010 16736 15016 16788
rect 15068 16776 15074 16788
rect 15105 16779 15163 16785
rect 15105 16776 15117 16779
rect 15068 16748 15117 16776
rect 15068 16736 15074 16748
rect 15105 16745 15117 16748
rect 15151 16745 15163 16779
rect 15105 16739 15163 16745
rect 16117 16779 16175 16785
rect 16117 16745 16129 16779
rect 16163 16776 16175 16779
rect 16206 16776 16212 16788
rect 16163 16748 16212 16776
rect 16163 16745 16175 16748
rect 16117 16739 16175 16745
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 14829 16643 14887 16649
rect 14829 16609 14841 16643
rect 14875 16640 14887 16643
rect 15657 16643 15715 16649
rect 15657 16640 15669 16643
rect 14875 16612 15669 16640
rect 14875 16609 14887 16612
rect 14829 16603 14887 16609
rect 15657 16609 15669 16612
rect 15703 16609 15715 16643
rect 15657 16603 15715 16609
rect 14415 16544 14596 16572
rect 14645 16575 14703 16581
rect 14415 16541 14427 16544
rect 14369 16535 14427 16541
rect 14645 16541 14657 16575
rect 14691 16572 14703 16575
rect 14734 16572 14740 16584
rect 14691 16544 14740 16572
rect 14691 16541 14703 16544
rect 14645 16535 14703 16541
rect 13722 16464 13728 16516
rect 13780 16464 13786 16516
rect 13906 16464 13912 16516
rect 13964 16504 13970 16516
rect 14108 16504 14136 16535
rect 13964 16476 14136 16504
rect 13964 16464 13970 16476
rect 12176 16408 12480 16436
rect 11664 16396 11670 16408
rect 12526 16396 12532 16448
rect 12584 16396 12590 16448
rect 13265 16439 13323 16445
rect 13265 16405 13277 16439
rect 13311 16436 13323 16439
rect 13630 16436 13636 16448
rect 13311 16408 13636 16436
rect 13311 16405 13323 16408
rect 13265 16399 13323 16405
rect 13630 16396 13636 16408
rect 13688 16436 13694 16448
rect 14292 16436 14320 16535
rect 14734 16532 14740 16544
rect 14792 16532 14798 16584
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15838 16572 15844 16584
rect 15519 16544 15844 16572
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 15930 16532 15936 16584
rect 15988 16532 15994 16584
rect 15378 16464 15384 16516
rect 15436 16504 15442 16516
rect 15565 16507 15623 16513
rect 15565 16504 15577 16507
rect 15436 16476 15577 16504
rect 15436 16464 15442 16476
rect 15565 16473 15577 16476
rect 15611 16473 15623 16507
rect 15565 16467 15623 16473
rect 13688 16408 14320 16436
rect 13688 16396 13694 16408
rect 1104 16346 16836 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 16836 16346
rect 1104 16272 16836 16294
rect 4062 16192 4068 16244
rect 4120 16192 4126 16244
rect 7558 16192 7564 16244
rect 7616 16232 7622 16244
rect 7745 16235 7803 16241
rect 7745 16232 7757 16235
rect 7616 16204 7757 16232
rect 7616 16192 7622 16204
rect 7745 16201 7757 16204
rect 7791 16201 7803 16235
rect 7745 16195 7803 16201
rect 7837 16235 7895 16241
rect 7837 16201 7849 16235
rect 7883 16232 7895 16235
rect 8018 16232 8024 16244
rect 7883 16204 8024 16232
rect 7883 16201 7895 16204
rect 7837 16195 7895 16201
rect 8018 16192 8024 16204
rect 8076 16192 8082 16244
rect 9766 16192 9772 16244
rect 9824 16232 9830 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9824 16204 9873 16232
rect 9824 16192 9830 16204
rect 9861 16201 9873 16204
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 4525 16167 4583 16173
rect 4525 16164 4537 16167
rect 4028 16136 4537 16164
rect 4028 16124 4034 16136
rect 4525 16133 4537 16136
rect 4571 16133 4583 16167
rect 6914 16164 6920 16176
rect 4525 16127 4583 16133
rect 6380 16136 6920 16164
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 4706 16096 4712 16108
rect 4479 16068 4712 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 4706 16056 4712 16068
rect 4764 16096 4770 16108
rect 5350 16096 5356 16108
rect 4764 16068 5356 16096
rect 4764 16056 4770 16068
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 6380 16105 6408 16136
rect 6914 16124 6920 16136
rect 6972 16164 6978 16176
rect 8202 16164 8208 16176
rect 6972 16136 8208 16164
rect 6972 16124 6978 16136
rect 8202 16124 8208 16136
rect 8260 16124 8266 16176
rect 8294 16124 8300 16176
rect 8352 16124 8358 16176
rect 8748 16167 8806 16173
rect 8748 16133 8760 16167
rect 8794 16164 8806 16167
rect 8938 16164 8944 16176
rect 8794 16136 8944 16164
rect 8794 16133 8806 16136
rect 8748 16127 8806 16133
rect 8938 16124 8944 16136
rect 8996 16124 9002 16176
rect 6638 16105 6644 16108
rect 6365 16099 6423 16105
rect 6365 16065 6377 16099
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 6632 16059 6644 16105
rect 6638 16056 6644 16059
rect 6696 16056 6702 16108
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 7892 16068 8033 16096
rect 7892 16056 7898 16068
rect 8021 16065 8033 16068
rect 8067 16065 8079 16099
rect 9876 16096 9904 16195
rect 9950 16192 9956 16244
rect 10008 16192 10014 16244
rect 11790 16192 11796 16244
rect 11848 16232 11854 16244
rect 12069 16235 12127 16241
rect 12069 16232 12081 16235
rect 11848 16204 12081 16232
rect 11848 16192 11854 16204
rect 12069 16201 12081 16204
rect 12115 16232 12127 16235
rect 12250 16232 12256 16244
rect 12115 16204 12256 16232
rect 12115 16201 12127 16204
rect 12069 16195 12127 16201
rect 12250 16192 12256 16204
rect 12308 16232 12314 16244
rect 12526 16232 12532 16244
rect 12308 16204 12532 16232
rect 12308 16192 12314 16204
rect 12526 16192 12532 16204
rect 12584 16192 12590 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 13262 16232 13268 16244
rect 12768 16204 13268 16232
rect 12768 16192 12774 16204
rect 13262 16192 13268 16204
rect 13320 16232 13326 16244
rect 13607 16235 13665 16241
rect 13607 16232 13619 16235
rect 13320 16204 13619 16232
rect 13320 16192 13326 16204
rect 13607 16201 13619 16204
rect 13653 16201 13665 16235
rect 13607 16195 13665 16201
rect 12805 16167 12863 16173
rect 12805 16164 12817 16167
rect 11725 16136 12817 16164
rect 11725 16108 11753 16136
rect 12805 16133 12817 16136
rect 12851 16164 12863 16167
rect 12986 16164 12992 16176
rect 12851 16136 12992 16164
rect 12851 16133 12863 16136
rect 12805 16127 12863 16133
rect 12986 16124 12992 16136
rect 13044 16124 13050 16176
rect 13814 16124 13820 16176
rect 13872 16124 13878 16176
rect 10505 16099 10563 16105
rect 10505 16096 10517 16099
rect 9876 16068 10517 16096
rect 8021 16059 8079 16065
rect 10505 16065 10517 16068
rect 10551 16065 10563 16099
rect 10505 16059 10563 16065
rect 11698 16056 11704 16108
rect 11756 16056 11762 16108
rect 14274 16096 14280 16108
rect 11808 16068 14280 16096
rect 4614 15988 4620 16040
rect 4672 15988 4678 16040
rect 7742 15988 7748 16040
rect 7800 16028 7806 16040
rect 8113 16031 8171 16037
rect 8113 16028 8125 16031
rect 7800 16000 8125 16028
rect 7800 15988 7806 16000
rect 8113 15997 8125 16000
rect 8159 15997 8171 16031
rect 8113 15991 8171 15997
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 8260 16000 8493 16028
rect 8260 15988 8266 16000
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 7300 15932 8423 15960
rect 5350 15852 5356 15904
rect 5408 15892 5414 15904
rect 7300 15892 7328 15932
rect 5408 15864 7328 15892
rect 5408 15852 5414 15864
rect 8294 15852 8300 15904
rect 8352 15852 8358 15904
rect 8395 15892 8423 15932
rect 11808 15892 11836 16068
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 15565 16099 15623 16105
rect 15565 16065 15577 16099
rect 15611 16096 15623 16099
rect 16114 16096 16120 16108
rect 15611 16068 16120 16096
rect 15611 16065 15623 16068
rect 15565 16059 15623 16065
rect 16114 16056 16120 16068
rect 16172 16096 16178 16108
rect 16393 16099 16451 16105
rect 16393 16096 16405 16099
rect 16172 16068 16405 16096
rect 16172 16056 16178 16068
rect 16393 16065 16405 16068
rect 16439 16065 16451 16099
rect 16393 16059 16451 16065
rect 12894 16028 12900 16040
rect 12268 16000 12900 16028
rect 12268 15969 12296 16000
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 12253 15963 12311 15969
rect 12253 15929 12265 15963
rect 12299 15929 12311 15963
rect 12253 15923 12311 15929
rect 12434 15920 12440 15972
rect 12492 15920 12498 15972
rect 13354 15960 13360 15972
rect 12928 15932 13360 15960
rect 8395 15864 11836 15892
rect 12066 15852 12072 15904
rect 12124 15852 12130 15904
rect 12345 15895 12403 15901
rect 12345 15861 12357 15895
rect 12391 15892 12403 15895
rect 12928 15892 12956 15932
rect 13354 15920 13360 15932
rect 13412 15920 13418 15972
rect 12391 15864 12956 15892
rect 12391 15861 12403 15864
rect 12345 15855 12403 15861
rect 12986 15852 12992 15904
rect 13044 15892 13050 15904
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 13044 15864 13461 15892
rect 13044 15852 13050 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 13630 15852 13636 15904
rect 13688 15852 13694 15904
rect 15746 15852 15752 15904
rect 15804 15852 15810 15904
rect 15838 15852 15844 15904
rect 15896 15852 15902 15904
rect 1104 15802 16836 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 16836 15802
rect 1104 15728 16836 15750
rect 2958 15688 2964 15700
rect 2240 15660 2964 15688
rect 2240 15561 2268 15660
rect 2958 15648 2964 15660
rect 3016 15688 3022 15700
rect 3145 15691 3203 15697
rect 3145 15688 3157 15691
rect 3016 15660 3157 15688
rect 3016 15648 3022 15660
rect 3145 15657 3157 15660
rect 3191 15688 3203 15691
rect 3326 15688 3332 15700
rect 3191 15660 3332 15688
rect 3191 15657 3203 15660
rect 3145 15651 3203 15657
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 6638 15648 6644 15700
rect 6696 15688 6702 15700
rect 6917 15691 6975 15697
rect 6917 15688 6929 15691
rect 6696 15660 6929 15688
rect 6696 15648 6702 15660
rect 6917 15657 6929 15660
rect 6963 15657 6975 15691
rect 6917 15651 6975 15657
rect 8294 15648 8300 15700
rect 8352 15688 8358 15700
rect 8941 15691 8999 15697
rect 8941 15688 8953 15691
rect 8352 15660 8953 15688
rect 8352 15648 8358 15660
rect 8941 15657 8953 15660
rect 8987 15657 8999 15691
rect 8941 15651 8999 15657
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 9088 15660 9137 15688
rect 9088 15648 9094 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 9401 15691 9459 15697
rect 9401 15688 9413 15691
rect 9364 15660 9413 15688
rect 9364 15648 9370 15660
rect 9401 15657 9413 15660
rect 9447 15657 9459 15691
rect 9401 15651 9459 15657
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12253 15691 12311 15697
rect 12253 15688 12265 15691
rect 12124 15660 12265 15688
rect 12124 15648 12130 15660
rect 12253 15657 12265 15660
rect 12299 15657 12311 15691
rect 12253 15651 12311 15657
rect 13909 15691 13967 15697
rect 13909 15657 13921 15691
rect 13955 15688 13967 15691
rect 15654 15688 15660 15700
rect 13955 15660 15660 15688
rect 13955 15657 13967 15660
rect 13909 15651 13967 15657
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 16114 15648 16120 15700
rect 16172 15648 16178 15700
rect 16390 15648 16396 15700
rect 16448 15648 16454 15700
rect 2866 15620 2872 15632
rect 2332 15592 2872 15620
rect 2225 15555 2283 15561
rect 2225 15521 2237 15555
rect 2271 15521 2283 15555
rect 2225 15515 2283 15521
rect 2332 15493 2360 15592
rect 2866 15580 2872 15592
rect 2924 15620 2930 15632
rect 3605 15623 3663 15629
rect 2924 15592 3372 15620
rect 2924 15580 2930 15592
rect 2409 15555 2467 15561
rect 2409 15521 2421 15555
rect 2455 15552 2467 15555
rect 3142 15552 3148 15564
rect 2455 15524 3148 15552
rect 2455 15521 2467 15524
rect 2409 15515 2467 15521
rect 2041 15487 2099 15493
rect 2041 15453 2053 15487
rect 2087 15453 2099 15487
rect 2041 15447 2099 15453
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15453 2375 15487
rect 2317 15447 2375 15453
rect 2056 15416 2084 15447
rect 2498 15444 2504 15496
rect 2556 15444 2562 15496
rect 2608 15493 2636 15524
rect 3142 15512 3148 15524
rect 3200 15512 3206 15564
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 2777 15487 2835 15493
rect 2777 15453 2789 15487
rect 2823 15484 2835 15487
rect 2958 15484 2964 15496
rect 2823 15456 2964 15484
rect 2823 15453 2835 15456
rect 2777 15447 2835 15453
rect 2608 15416 2636 15447
rect 2958 15444 2964 15456
rect 3016 15444 3022 15496
rect 3344 15493 3372 15592
rect 3605 15589 3617 15623
rect 3651 15620 3663 15623
rect 3651 15592 4660 15620
rect 3651 15589 3663 15592
rect 3605 15583 3663 15589
rect 4632 15561 4660 15592
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 5592 15592 12434 15620
rect 5592 15580 5598 15592
rect 4617 15555 4675 15561
rect 4617 15521 4629 15555
rect 4663 15521 4675 15555
rect 4617 15515 4675 15521
rect 6086 15512 6092 15564
rect 6144 15552 6150 15564
rect 6273 15555 6331 15561
rect 6273 15552 6285 15555
rect 6144 15524 6285 15552
rect 6144 15512 6150 15524
rect 6273 15521 6285 15524
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15453 3111 15487
rect 3053 15447 3111 15453
rect 3329 15487 3387 15493
rect 3329 15453 3341 15487
rect 3375 15453 3387 15487
rect 3329 15447 3387 15453
rect 2056 15388 2636 15416
rect 2682 15376 2688 15428
rect 2740 15376 2746 15428
rect 1857 15351 1915 15357
rect 1857 15317 1869 15351
rect 1903 15348 1915 15351
rect 2130 15348 2136 15360
rect 1903 15320 2136 15348
rect 1903 15317 1915 15320
rect 1857 15311 1915 15317
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 2590 15308 2596 15360
rect 2648 15348 2654 15360
rect 3068 15348 3096 15447
rect 3142 15376 3148 15428
rect 3200 15416 3206 15428
rect 3344 15416 3372 15447
rect 3970 15444 3976 15496
rect 4028 15484 4034 15496
rect 4433 15487 4491 15493
rect 4433 15484 4445 15487
rect 4028 15456 4445 15484
rect 4028 15444 4034 15456
rect 4433 15453 4445 15456
rect 4479 15453 4491 15487
rect 6288 15484 6316 15515
rect 6454 15512 6460 15564
rect 6512 15512 6518 15564
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 7929 15555 7987 15561
rect 7929 15552 7941 15555
rect 7708 15524 7941 15552
rect 7708 15512 7714 15524
rect 7929 15521 7941 15524
rect 7975 15521 7987 15555
rect 7929 15515 7987 15521
rect 8110 15512 8116 15564
rect 8168 15512 8174 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10134 15552 10140 15564
rect 9999 15524 10140 15552
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 10134 15512 10140 15524
rect 10192 15512 10198 15564
rect 12406 15552 12434 15592
rect 13170 15580 13176 15632
rect 13228 15620 13234 15632
rect 13814 15620 13820 15632
rect 13228 15592 13820 15620
rect 13228 15580 13234 15592
rect 13814 15580 13820 15592
rect 13872 15580 13878 15632
rect 12406 15524 14412 15552
rect 6822 15484 6828 15496
rect 6288 15456 6828 15484
rect 4433 15447 4491 15453
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15484 9919 15487
rect 10042 15484 10048 15496
rect 9907 15456 10048 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 10042 15444 10048 15456
rect 10100 15484 10106 15496
rect 11333 15487 11391 15493
rect 11333 15484 11345 15487
rect 10100 15456 11345 15484
rect 10100 15444 10106 15456
rect 11333 15453 11345 15456
rect 11379 15453 11391 15487
rect 11333 15447 11391 15453
rect 11977 15487 12035 15493
rect 11977 15453 11989 15487
rect 12023 15484 12035 15487
rect 12618 15484 12624 15496
rect 12023 15456 12624 15484
rect 12023 15453 12035 15456
rect 11977 15447 12035 15453
rect 12618 15444 12624 15456
rect 12676 15444 12682 15496
rect 13170 15444 13176 15496
rect 13228 15444 13234 15496
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 13449 15487 13507 15493
rect 13449 15453 13461 15487
rect 13495 15453 13507 15487
rect 13449 15447 13507 15453
rect 3200 15388 3372 15416
rect 3200 15376 3206 15388
rect 8846 15376 8852 15428
rect 8904 15416 8910 15428
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 8904 15388 9321 15416
rect 8904 15376 8910 15388
rect 9309 15385 9321 15388
rect 9355 15385 9367 15419
rect 9309 15379 9367 15385
rect 11698 15376 11704 15428
rect 11756 15416 11762 15428
rect 12069 15419 12127 15425
rect 12069 15416 12081 15419
rect 11756 15388 12081 15416
rect 11756 15376 11762 15388
rect 12069 15385 12081 15388
rect 12115 15385 12127 15419
rect 12069 15379 12127 15385
rect 12250 15376 12256 15428
rect 12308 15425 12314 15428
rect 12308 15419 12327 15425
rect 12315 15385 12327 15419
rect 12308 15379 12327 15385
rect 12308 15376 12314 15379
rect 2648 15320 3096 15348
rect 4065 15351 4123 15357
rect 2648 15308 2654 15320
rect 4065 15317 4077 15351
rect 4111 15348 4123 15351
rect 4246 15348 4252 15360
rect 4111 15320 4252 15348
rect 4111 15317 4123 15320
rect 4065 15311 4123 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 4525 15351 4583 15357
rect 4525 15317 4537 15351
rect 4571 15348 4583 15351
rect 5534 15348 5540 15360
rect 4571 15320 5540 15348
rect 4571 15317 4583 15320
rect 4525 15311 4583 15317
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 6549 15351 6607 15357
rect 6549 15317 6561 15351
rect 6595 15348 6607 15351
rect 7006 15348 7012 15360
rect 6595 15320 7012 15348
rect 6595 15317 6607 15320
rect 6549 15311 6607 15317
rect 7006 15308 7012 15320
rect 7064 15308 7070 15360
rect 7374 15308 7380 15360
rect 7432 15308 7438 15360
rect 8754 15308 8760 15360
rect 8812 15308 8818 15360
rect 9109 15351 9167 15357
rect 9109 15317 9121 15351
rect 9155 15348 9167 15351
rect 9490 15348 9496 15360
rect 9155 15320 9496 15348
rect 9155 15317 9167 15320
rect 9109 15311 9167 15317
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 9769 15351 9827 15357
rect 9769 15317 9781 15351
rect 9815 15348 9827 15351
rect 10318 15348 10324 15360
rect 9815 15320 10324 15348
rect 9815 15317 9827 15320
rect 9769 15311 9827 15317
rect 10318 15308 10324 15320
rect 10376 15308 10382 15360
rect 12434 15308 12440 15360
rect 12492 15348 12498 15360
rect 13372 15348 13400 15447
rect 13464 15416 13492 15447
rect 13538 15444 13544 15496
rect 13596 15444 13602 15496
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13688 15456 13737 15484
rect 13688 15444 13694 15456
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 14182 15444 14188 15496
rect 14240 15484 14246 15496
rect 14384 15493 14412 15524
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 14737 15555 14795 15561
rect 14737 15552 14749 15555
rect 14608 15524 14749 15552
rect 14608 15512 14614 15524
rect 14737 15521 14749 15524
rect 14783 15521 14795 15555
rect 14737 15515 14795 15521
rect 14277 15487 14335 15493
rect 14277 15484 14289 15487
rect 14240 15456 14289 15484
rect 14240 15444 14246 15456
rect 14277 15453 14289 15456
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15453 14427 15487
rect 14369 15447 14427 15453
rect 14458 15444 14464 15496
rect 14516 15444 14522 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 15804 15456 16221 15484
rect 15804 15444 15810 15456
rect 16209 15453 16221 15456
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 14734 15416 14740 15428
rect 13464 15388 14740 15416
rect 14292 15360 14320 15388
rect 14734 15376 14740 15388
rect 14792 15376 14798 15428
rect 15004 15419 15062 15425
rect 15004 15385 15016 15419
rect 15050 15416 15062 15419
rect 15102 15416 15108 15428
rect 15050 15388 15108 15416
rect 15050 15385 15062 15388
rect 15004 15379 15062 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 12492 15320 13400 15348
rect 12492 15308 12498 15320
rect 14274 15308 14280 15360
rect 14332 15308 14338 15360
rect 14645 15351 14703 15357
rect 14645 15317 14657 15351
rect 14691 15348 14703 15351
rect 15562 15348 15568 15360
rect 14691 15320 15568 15348
rect 14691 15317 14703 15320
rect 14645 15311 14703 15317
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 1104 15258 16836 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 16836 15258
rect 1104 15184 16836 15206
rect 2958 15104 2964 15156
rect 3016 15104 3022 15156
rect 5534 15104 5540 15156
rect 5592 15104 5598 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7745 15147 7803 15153
rect 7745 15144 7757 15147
rect 7708 15116 7757 15144
rect 7708 15104 7714 15116
rect 7745 15113 7757 15116
rect 7791 15113 7803 15147
rect 7745 15107 7803 15113
rect 7929 15147 7987 15153
rect 7929 15113 7941 15147
rect 7975 15144 7987 15147
rect 8110 15144 8116 15156
rect 7975 15116 8116 15144
rect 7975 15113 7987 15116
rect 7929 15107 7987 15113
rect 8110 15104 8116 15116
rect 8168 15104 8174 15156
rect 9953 15147 10011 15153
rect 9953 15113 9965 15147
rect 9999 15144 10011 15147
rect 10042 15144 10048 15156
rect 9999 15116 10048 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 12526 15144 12532 15156
rect 11716 15116 12532 15144
rect 2774 15076 2780 15088
rect 1596 15048 2780 15076
rect 1596 15017 1624 15048
rect 2774 15036 2780 15048
rect 2832 15036 2838 15088
rect 2976 15076 3004 15104
rect 6914 15076 6920 15088
rect 2976 15048 3740 15076
rect 1854 15017 1860 15020
rect 1581 15011 1639 15017
rect 1581 14977 1593 15011
rect 1627 14977 1639 15011
rect 1581 14971 1639 14977
rect 1848 14971 1860 15017
rect 1854 14968 1860 14971
rect 1912 14968 1918 15020
rect 3142 14968 3148 15020
rect 3200 15008 3206 15020
rect 3712 15017 3740 15048
rect 4172 15048 6920 15076
rect 4172 15017 4200 15048
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 3200 14980 3433 15008
rect 3200 14968 3206 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3697 15011 3755 15017
rect 3697 14977 3709 15011
rect 3743 14977 3755 15011
rect 3697 14971 3755 14977
rect 4157 15011 4215 15017
rect 4157 14977 4169 15011
rect 4203 14977 4215 15011
rect 4157 14971 4215 14977
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 6380 15017 6408 15048
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 8846 15036 8852 15088
rect 8904 15076 8910 15088
rect 9582 15076 9588 15088
rect 8904 15048 9588 15076
rect 8904 15036 8910 15048
rect 9582 15036 9588 15048
rect 9640 15036 9646 15088
rect 11088 15079 11146 15085
rect 11088 15045 11100 15079
rect 11134 15076 11146 15079
rect 11517 15079 11575 15085
rect 11517 15076 11529 15079
rect 11134 15048 11529 15076
rect 11134 15045 11146 15048
rect 11088 15039 11146 15045
rect 11517 15045 11529 15048
rect 11563 15045 11575 15079
rect 11517 15039 11575 15045
rect 6638 15017 6644 15020
rect 4413 15011 4471 15017
rect 4413 15008 4425 15011
rect 4304 14980 4425 15008
rect 4304 14968 4310 14980
rect 4413 14977 4425 14980
rect 4459 14977 4471 15011
rect 4413 14971 4471 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 14977 6423 15011
rect 6365 14971 6423 14977
rect 6632 14971 6644 15017
rect 6638 14968 6644 14971
rect 6696 14968 6702 15020
rect 9030 14968 9036 15020
rect 9088 15017 9094 15020
rect 9088 14971 9100 15017
rect 9088 14968 9094 14971
rect 11238 14968 11244 15020
rect 11296 15008 11302 15020
rect 11716 15017 11744 15116
rect 12526 15104 12532 15116
rect 12584 15144 12590 15156
rect 13078 15144 13084 15156
rect 12584 15116 13084 15144
rect 12584 15104 12590 15116
rect 13078 15104 13084 15116
rect 13136 15144 13142 15156
rect 14001 15147 14059 15153
rect 13136 15116 13584 15144
rect 13136 15104 13142 15116
rect 12434 15076 12440 15088
rect 12360 15048 12440 15076
rect 11333 15011 11391 15017
rect 11333 15008 11345 15011
rect 11296 14980 11345 15008
rect 11296 14968 11302 14980
rect 11333 14977 11345 14980
rect 11379 14977 11391 15011
rect 11333 14971 11391 14977
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 14977 11759 15011
rect 11701 14971 11759 14977
rect 11793 15011 11851 15017
rect 11793 14977 11805 15011
rect 11839 15008 11851 15011
rect 11882 15008 11888 15020
rect 11839 14980 11888 15008
rect 11839 14977 11851 14980
rect 11793 14971 11851 14977
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 12360 15017 12388 15048
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 13170 15076 13176 15088
rect 12544 15048 13176 15076
rect 11977 15011 12035 15017
rect 11977 14977 11989 15011
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12544 15008 12572 15048
rect 13170 15036 13176 15048
rect 13228 15076 13234 15088
rect 13449 15079 13507 15085
rect 13449 15076 13461 15079
rect 13228 15048 13461 15076
rect 13228 15036 13234 15048
rect 13449 15045 13461 15048
rect 13495 15045 13507 15079
rect 13556 15076 13584 15116
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14090 15144 14096 15156
rect 14047 15116 14096 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 15102 15104 15108 15156
rect 15160 15104 15166 15156
rect 15473 15147 15531 15153
rect 15473 15113 15485 15147
rect 15519 15144 15531 15147
rect 15838 15144 15844 15156
rect 15519 15116 15844 15144
rect 15519 15113 15531 15116
rect 15473 15107 15531 15113
rect 15838 15104 15844 15116
rect 15896 15104 15902 15156
rect 13633 15079 13691 15085
rect 13633 15076 13645 15079
rect 13556 15048 13645 15076
rect 13449 15039 13507 15045
rect 13633 15045 13645 15048
rect 13679 15045 13691 15079
rect 13633 15039 13691 15045
rect 15562 15036 15568 15088
rect 15620 15036 15626 15088
rect 12345 14971 12403 14977
rect 12452 14980 12572 15008
rect 9309 14943 9367 14949
rect 9309 14909 9321 14943
rect 9355 14909 9367 14943
rect 11992 14940 12020 14971
rect 12452 14949 12480 14980
rect 12618 14968 12624 15020
rect 12676 14968 12682 15020
rect 12802 14968 12808 15020
rect 12860 15008 12866 15020
rect 12989 15011 13047 15017
rect 12989 15008 13001 15011
rect 12860 14980 13001 15008
rect 12860 14968 12866 14980
rect 12989 14977 13001 14980
rect 13035 14977 13047 15011
rect 12989 14971 13047 14977
rect 12161 14943 12219 14949
rect 12161 14940 12173 14943
rect 11992 14912 12173 14940
rect 9309 14903 9367 14909
rect 12161 14909 12173 14912
rect 12207 14909 12219 14943
rect 12161 14903 12219 14909
rect 12437 14943 12495 14949
rect 12437 14909 12449 14943
rect 12483 14909 12495 14943
rect 12437 14903 12495 14909
rect 3418 14832 3424 14884
rect 3476 14872 3482 14884
rect 3973 14875 4031 14881
rect 3973 14872 3985 14875
rect 3476 14844 3985 14872
rect 3476 14832 3482 14844
rect 3973 14841 3985 14844
rect 4019 14841 4031 14875
rect 3973 14835 4031 14841
rect 3510 14764 3516 14816
rect 3568 14764 3574 14816
rect 8938 14764 8944 14816
rect 8996 14804 9002 14816
rect 9324 14804 9352 14903
rect 12526 14900 12532 14952
rect 12584 14940 12590 14952
rect 12710 14940 12716 14952
rect 12584 14912 12716 14940
rect 12584 14900 12590 14912
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 13004 14940 13032 14971
rect 13262 14968 13268 15020
rect 13320 14968 13326 15020
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 13817 15011 13875 15017
rect 13817 14977 13829 15011
rect 13863 15008 13875 15011
rect 14090 15008 14096 15020
rect 13863 14980 14096 15008
rect 13863 14977 13875 14980
rect 13817 14971 13875 14977
rect 13556 14940 13584 14971
rect 14090 14968 14096 14980
rect 14148 14968 14154 15020
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 15008 15991 15011
rect 16114 15008 16120 15020
rect 15979 14980 16120 15008
rect 15979 14977 15991 14980
rect 15933 14971 15991 14977
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 14366 14940 14372 14952
rect 13004 14912 14372 14940
rect 14366 14900 14372 14912
rect 14424 14900 14430 14952
rect 15654 14900 15660 14952
rect 15712 14900 15718 14952
rect 11882 14832 11888 14884
rect 11940 14832 11946 14884
rect 13262 14832 13268 14884
rect 13320 14872 13326 14884
rect 13538 14872 13544 14884
rect 13320 14844 13544 14872
rect 13320 14832 13326 14844
rect 13538 14832 13544 14844
rect 13596 14832 13602 14884
rect 8996 14776 9352 14804
rect 16117 14807 16175 14813
rect 8996 14764 9002 14776
rect 16117 14773 16129 14807
rect 16163 14804 16175 14807
rect 16206 14804 16212 14816
rect 16163 14776 16212 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 16206 14764 16212 14776
rect 16264 14764 16270 14816
rect 1104 14714 16836 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 16836 14714
rect 1104 14640 16836 14662
rect 1765 14603 1823 14609
rect 1765 14569 1777 14603
rect 1811 14600 1823 14603
rect 1854 14600 1860 14612
rect 1811 14572 1860 14600
rect 1811 14569 1823 14572
rect 1765 14563 1823 14569
rect 1854 14560 1860 14572
rect 1912 14560 1918 14612
rect 2685 14603 2743 14609
rect 2685 14569 2697 14603
rect 2731 14600 2743 14603
rect 2958 14600 2964 14612
rect 2731 14572 2964 14600
rect 2731 14569 2743 14572
rect 2685 14563 2743 14569
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 3142 14560 3148 14612
rect 3200 14560 3206 14612
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 6917 14603 6975 14609
rect 6917 14600 6929 14603
rect 6696 14572 6929 14600
rect 6696 14560 6702 14572
rect 6917 14569 6929 14572
rect 6963 14569 6975 14603
rect 8846 14600 8852 14612
rect 6917 14563 6975 14569
rect 7484 14572 8852 14600
rect 2317 14535 2375 14541
rect 2317 14501 2329 14535
rect 2363 14532 2375 14535
rect 3160 14532 3188 14560
rect 2363 14504 3188 14532
rect 2363 14501 2375 14504
rect 2317 14495 2375 14501
rect 6822 14492 6828 14544
rect 6880 14532 6886 14544
rect 7484 14532 7512 14572
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 8941 14603 8999 14609
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9030 14600 9036 14612
rect 8987 14572 9036 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 9030 14560 9036 14572
rect 9088 14560 9094 14612
rect 9861 14603 9919 14609
rect 9861 14569 9873 14603
rect 9907 14600 9919 14603
rect 9907 14572 11376 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 9876 14532 9904 14563
rect 6880 14504 7512 14532
rect 6880 14492 6886 14504
rect 2038 14464 2044 14476
rect 1964 14436 2044 14464
rect 1964 14405 1992 14436
rect 2038 14424 2044 14436
rect 2096 14464 2102 14476
rect 2682 14464 2688 14476
rect 2096 14436 2688 14464
rect 2096 14424 2102 14436
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 7374 14424 7380 14476
rect 7432 14424 7438 14476
rect 7484 14473 7512 14504
rect 8220 14504 9904 14532
rect 8220 14473 8248 14504
rect 7469 14467 7527 14473
rect 7469 14433 7481 14467
rect 7515 14433 7527 14467
rect 7469 14427 7527 14433
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14433 8263 14467
rect 8205 14427 8263 14433
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 1949 14399 2007 14405
rect 1949 14365 1961 14399
rect 1995 14365 2007 14399
rect 1949 14359 2007 14365
rect 2130 14356 2136 14408
rect 2188 14356 2194 14408
rect 2958 14356 2964 14408
rect 3016 14396 3022 14408
rect 3053 14399 3111 14405
rect 3053 14396 3065 14399
rect 3016 14368 3065 14396
rect 3016 14356 3022 14368
rect 3053 14365 3065 14368
rect 3099 14365 3111 14399
rect 3053 14359 3111 14365
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 3510 14396 3516 14408
rect 3467 14368 3516 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3510 14356 3516 14368
rect 3568 14356 3574 14408
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 4295 14368 6745 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 6733 14365 6745 14368
rect 6779 14396 6791 14399
rect 6914 14396 6920 14408
rect 6779 14368 6920 14396
rect 6779 14365 6791 14368
rect 6733 14359 6791 14365
rect 6914 14356 6920 14368
rect 6972 14356 6978 14408
rect 7926 14356 7932 14408
rect 7984 14396 7990 14408
rect 8312 14396 8340 14427
rect 8754 14424 8760 14476
rect 8812 14464 8818 14476
rect 9401 14467 9459 14473
rect 9401 14464 9413 14467
rect 8812 14436 9413 14464
rect 8812 14424 8818 14436
rect 9401 14433 9413 14436
rect 9447 14433 9459 14467
rect 9401 14427 9459 14433
rect 9582 14424 9588 14476
rect 9640 14424 9646 14476
rect 11348 14473 11376 14572
rect 12986 14560 12992 14612
rect 13044 14600 13050 14612
rect 13081 14603 13139 14609
rect 13081 14600 13093 14603
rect 13044 14572 13093 14600
rect 13044 14560 13050 14572
rect 13081 14569 13093 14572
rect 13127 14600 13139 14603
rect 13722 14600 13728 14612
rect 13127 14572 13728 14600
rect 13127 14569 13139 14572
rect 13081 14563 13139 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 16114 14560 16120 14612
rect 16172 14560 16178 14612
rect 11882 14492 11888 14544
rect 11940 14532 11946 14544
rect 11940 14504 12664 14532
rect 11940 14492 11946 14504
rect 11333 14467 11391 14473
rect 11333 14433 11345 14467
rect 11379 14433 11391 14467
rect 11333 14427 11391 14433
rect 11977 14467 12035 14473
rect 11977 14433 11989 14467
rect 12023 14464 12035 14467
rect 12023 14436 12388 14464
rect 12023 14433 12035 14436
rect 11977 14427 12035 14433
rect 7984 14368 8340 14396
rect 7984 14356 7990 14368
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9858 14396 9864 14408
rect 8996 14368 9864 14396
rect 8996 14356 9002 14368
rect 9858 14356 9864 14368
rect 9916 14396 9922 14408
rect 11238 14396 11244 14408
rect 9916 14368 11244 14396
rect 9916 14356 9922 14368
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11606 14356 11612 14408
rect 11664 14396 11670 14408
rect 12250 14396 12256 14408
rect 11664 14368 12256 14396
rect 11664 14356 11670 14368
rect 12250 14356 12256 14368
rect 12308 14356 12314 14408
rect 12360 14405 12388 14436
rect 12526 14424 12532 14476
rect 12584 14424 12590 14476
rect 12636 14405 12664 14504
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 13078 14464 13084 14476
rect 12768 14436 13084 14464
rect 12768 14424 12774 14436
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13814 14424 13820 14476
rect 13872 14464 13878 14476
rect 14182 14464 14188 14476
rect 13872 14436 14188 14464
rect 13872 14424 13878 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14550 14424 14556 14476
rect 14608 14464 14614 14476
rect 14734 14464 14740 14476
rect 14608 14436 14740 14464
rect 14608 14424 14614 14436
rect 14734 14424 14740 14436
rect 14792 14424 14798 14476
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14365 12403 14399
rect 12345 14359 12403 14365
rect 12621 14399 12679 14405
rect 12621 14365 12633 14399
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 12894 14356 12900 14408
rect 12952 14356 12958 14408
rect 13096 14396 13124 14424
rect 13173 14399 13231 14405
rect 13173 14396 13185 14399
rect 13096 14368 13185 14396
rect 13173 14365 13185 14368
rect 13219 14365 13231 14399
rect 13173 14359 13231 14365
rect 13354 14356 13360 14408
rect 13412 14356 13418 14408
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 13541 14399 13599 14405
rect 13541 14396 13553 14399
rect 13504 14368 13553 14396
rect 13504 14356 13510 14368
rect 13541 14365 13553 14368
rect 13587 14396 13599 14399
rect 16022 14396 16028 14408
rect 13587 14368 16028 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16206 14356 16212 14408
rect 16264 14356 16270 14408
rect 2590 14288 2596 14340
rect 2648 14328 2654 14340
rect 2685 14331 2743 14337
rect 2685 14328 2697 14331
rect 2648 14300 2697 14328
rect 2648 14288 2654 14300
rect 2685 14297 2697 14300
rect 2731 14297 2743 14331
rect 2685 14291 2743 14297
rect 4062 14288 4068 14340
rect 4120 14328 4126 14340
rect 4494 14331 4552 14337
rect 4494 14328 4506 14331
rect 4120 14300 4506 14328
rect 4120 14288 4126 14300
rect 4494 14297 4506 14300
rect 4540 14297 4552 14331
rect 5994 14328 6000 14340
rect 4494 14291 4552 14297
rect 5644 14300 6000 14328
rect 2866 14220 2872 14272
rect 2924 14220 2930 14272
rect 3602 14220 3608 14272
rect 3660 14220 3666 14272
rect 5644 14269 5672 14300
rect 5994 14288 6000 14300
rect 6052 14328 6058 14340
rect 10996 14331 11054 14337
rect 6052 14300 9674 14328
rect 6052 14288 6058 14300
rect 5629 14263 5687 14269
rect 5629 14229 5641 14263
rect 5675 14229 5687 14263
rect 5629 14223 5687 14229
rect 7285 14263 7343 14269
rect 7285 14229 7297 14263
rect 7331 14260 7343 14263
rect 7745 14263 7803 14269
rect 7745 14260 7757 14263
rect 7331 14232 7757 14260
rect 7331 14229 7343 14232
rect 7285 14223 7343 14229
rect 7745 14229 7757 14232
rect 7791 14229 7803 14263
rect 7745 14223 7803 14229
rect 8110 14220 8116 14272
rect 8168 14220 8174 14272
rect 9306 14220 9312 14272
rect 9364 14220 9370 14272
rect 9646 14260 9674 14300
rect 10996 14297 11008 14331
rect 11042 14328 11054 14331
rect 12069 14331 12127 14337
rect 12069 14328 12081 14331
rect 11042 14300 12081 14328
rect 11042 14297 11054 14300
rect 10996 14291 11054 14297
rect 12069 14297 12081 14300
rect 12115 14297 12127 14331
rect 12069 14291 12127 14297
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 13078 14328 13084 14340
rect 12584 14300 13084 14328
rect 12584 14288 12590 14300
rect 13078 14288 13084 14300
rect 13136 14288 13142 14340
rect 14642 14328 14648 14340
rect 13280 14300 14648 14328
rect 13280 14272 13308 14300
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 15010 14337 15016 14340
rect 15004 14291 15016 14337
rect 15010 14288 15016 14291
rect 15068 14288 15074 14340
rect 13170 14260 13176 14272
rect 9646 14232 13176 14260
rect 13170 14220 13176 14232
rect 13228 14220 13234 14272
rect 13262 14220 13268 14272
rect 13320 14220 13326 14272
rect 13538 14220 13544 14272
rect 13596 14260 13602 14272
rect 13725 14263 13783 14269
rect 13725 14260 13737 14263
rect 13596 14232 13737 14260
rect 13596 14220 13602 14232
rect 13725 14229 13737 14232
rect 13771 14260 13783 14263
rect 14826 14260 14832 14272
rect 13771 14232 14832 14260
rect 13771 14229 13783 14232
rect 13725 14223 13783 14229
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 1104 14170 16836 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 16836 14170
rect 1104 14096 16836 14118
rect 1949 14059 2007 14065
rect 1949 14025 1961 14059
rect 1995 14056 2007 14059
rect 2958 14056 2964 14068
rect 1995 14028 2964 14056
rect 1995 14025 2007 14028
rect 1949 14019 2007 14025
rect 2958 14016 2964 14028
rect 3016 14056 3022 14068
rect 3697 14059 3755 14065
rect 3697 14056 3709 14059
rect 3016 14028 3709 14056
rect 3016 14016 3022 14028
rect 3697 14025 3709 14028
rect 3743 14056 3755 14059
rect 3970 14056 3976 14068
rect 3743 14028 3976 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4062 14016 4068 14068
rect 4120 14016 4126 14068
rect 10226 14056 10232 14068
rect 6564 14028 10232 14056
rect 2774 13948 2780 14000
rect 2832 13988 2838 14000
rect 3786 13988 3792 14000
rect 2832 13960 3792 13988
rect 2832 13948 2838 13960
rect 3786 13948 3792 13960
rect 3844 13988 3850 14000
rect 4893 13991 4951 13997
rect 4893 13988 4905 13991
rect 3844 13960 4905 13988
rect 3844 13948 3850 13960
rect 4893 13957 4905 13960
rect 4939 13957 4951 13991
rect 4893 13951 4951 13957
rect 6362 13948 6368 14000
rect 6420 13988 6426 14000
rect 6564 13997 6592 14028
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11940 14028 12173 14056
rect 11940 14016 11946 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 12434 14016 12440 14068
rect 12492 14016 12498 14068
rect 12526 14016 12532 14068
rect 12584 14016 12590 14068
rect 12618 14016 12624 14068
rect 12676 14016 12682 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13725 14059 13783 14065
rect 13228 14028 13308 14056
rect 13228 14016 13234 14028
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6420 13960 6561 13988
rect 6420 13948 6426 13960
rect 6549 13957 6561 13960
rect 6595 13957 6607 13991
rect 6549 13951 6607 13957
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 6914 13988 6920 14000
rect 6696 13960 6920 13988
rect 6696 13948 6702 13960
rect 6914 13948 6920 13960
rect 6972 13988 6978 14000
rect 7285 13991 7343 13997
rect 7285 13988 7297 13991
rect 6972 13960 7297 13988
rect 6972 13948 6978 13960
rect 7285 13957 7297 13960
rect 7331 13957 7343 13991
rect 7285 13951 7343 13957
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13889 1915 13923
rect 1857 13883 1915 13889
rect 1872 13784 1900 13883
rect 2682 13880 2688 13932
rect 2740 13880 2746 13932
rect 2958 13920 2964 13932
rect 2792 13892 2964 13920
rect 2038 13812 2044 13864
rect 2096 13812 2102 13864
rect 2792 13861 2820 13892
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 4157 13923 4215 13929
rect 4157 13889 4169 13923
rect 4203 13920 4215 13923
rect 6380 13920 6408 13948
rect 4203 13892 6408 13920
rect 7300 13920 7328 13951
rect 9122 13948 9128 14000
rect 9180 13988 9186 14000
rect 9180 13960 11100 13988
rect 9180 13948 9186 13960
rect 8113 13923 8171 13929
rect 8113 13920 8125 13923
rect 7300 13892 8125 13920
rect 4203 13889 4215 13892
rect 4157 13883 4215 13889
rect 8113 13889 8125 13892
rect 8159 13889 8171 13923
rect 8113 13883 8171 13889
rect 8380 13923 8438 13929
rect 8380 13889 8392 13923
rect 8426 13920 8438 13923
rect 8426 13892 9628 13920
rect 8426 13889 8438 13892
rect 8380 13883 8438 13889
rect 2777 13855 2835 13861
rect 2777 13821 2789 13855
rect 2823 13821 2835 13855
rect 2777 13815 2835 13821
rect 2866 13812 2872 13864
rect 2924 13812 2930 13864
rect 3418 13812 3424 13864
rect 3476 13812 3482 13864
rect 3605 13855 3663 13861
rect 3605 13821 3617 13855
rect 3651 13852 3663 13855
rect 5994 13852 6000 13864
rect 3651 13824 6000 13852
rect 3651 13821 3663 13824
rect 3605 13815 3663 13821
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9180 13824 9536 13852
rect 9180 13812 9186 13824
rect 2590 13784 2596 13796
rect 1872 13756 2596 13784
rect 2590 13744 2596 13756
rect 2648 13784 2654 13796
rect 9508 13793 9536 13824
rect 9600 13793 9628 13892
rect 9950 13880 9956 13932
rect 10008 13880 10014 13932
rect 11072 13929 11100 13960
rect 11698 13948 11704 14000
rect 11756 13988 11762 14000
rect 12452 13988 12480 14016
rect 11756 13960 12480 13988
rect 11756 13948 11762 13960
rect 10045 13923 10103 13929
rect 10045 13889 10057 13923
rect 10091 13920 10103 13923
rect 10413 13923 10471 13929
rect 10413 13920 10425 13923
rect 10091 13892 10425 13920
rect 10091 13889 10103 13892
rect 10045 13883 10103 13889
rect 10413 13889 10425 13892
rect 10459 13889 10471 13923
rect 10413 13883 10471 13889
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13889 11115 13923
rect 11057 13883 11115 13889
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 11609 13923 11667 13929
rect 11609 13920 11621 13923
rect 11296 13892 11621 13920
rect 11296 13880 11302 13892
rect 11609 13889 11621 13892
rect 11655 13889 11667 13923
rect 11609 13883 11667 13889
rect 12158 13880 12164 13932
rect 12216 13880 12222 13932
rect 12360 13929 12388 13960
rect 12345 13923 12403 13929
rect 12345 13889 12357 13923
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 12636 13929 12664 14016
rect 12906 13960 13032 13988
rect 12906 13929 12934 13960
rect 12621 13923 12679 13929
rect 12621 13920 12633 13923
rect 12544 13892 12633 13920
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 9493 13787 9551 13793
rect 2648 13756 2774 13784
rect 2648 13744 2654 13756
rect 1486 13676 1492 13728
rect 1544 13676 1550 13728
rect 2222 13676 2228 13728
rect 2280 13716 2286 13728
rect 2317 13719 2375 13725
rect 2317 13716 2329 13719
rect 2280 13688 2329 13716
rect 2280 13676 2286 13688
rect 2317 13685 2329 13688
rect 2363 13685 2375 13719
rect 2746 13716 2774 13756
rect 9493 13753 9505 13787
rect 9539 13753 9551 13787
rect 9493 13747 9551 13753
rect 9585 13787 9643 13793
rect 9585 13753 9597 13787
rect 9631 13753 9643 13787
rect 9585 13747 9643 13753
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 10152 13784 10180 13815
rect 12544 13796 12572 13892
rect 12621 13889 12633 13892
rect 12667 13889 12679 13923
rect 12621 13883 12679 13889
rect 12719 13923 12777 13929
rect 12719 13889 12731 13923
rect 12765 13889 12777 13923
rect 12719 13883 12777 13889
rect 12891 13923 12949 13929
rect 12891 13889 12903 13923
rect 12937 13889 12949 13923
rect 12891 13883 12949 13889
rect 9732 13756 10180 13784
rect 9732 13744 9738 13756
rect 12526 13744 12532 13796
rect 12584 13744 12590 13796
rect 12729 13784 12757 13883
rect 13004 13852 13032 13960
rect 13170 13880 13176 13932
rect 13228 13880 13234 13932
rect 13280 13923 13308 14028
rect 13725 14025 13737 14059
rect 13771 14025 13783 14059
rect 13725 14019 13783 14025
rect 13357 13991 13415 13997
rect 13357 13957 13369 13991
rect 13403 13988 13415 13991
rect 13630 13988 13636 14000
rect 13403 13960 13636 13988
rect 13403 13957 13415 13960
rect 13357 13951 13415 13957
rect 13630 13948 13636 13960
rect 13688 13948 13694 14000
rect 13740 13988 13768 14019
rect 13814 14016 13820 14068
rect 13872 14056 13878 14068
rect 14458 14056 14464 14068
rect 13872 14028 14464 14056
rect 13872 14016 13878 14028
rect 14458 14016 14464 14028
rect 14516 14016 14522 14068
rect 15010 14016 15016 14068
rect 15068 14016 15074 14068
rect 15473 13991 15531 13997
rect 15473 13988 15485 13991
rect 13740 13960 15485 13988
rect 15473 13957 15485 13960
rect 15519 13957 15531 13991
rect 15473 13951 15531 13957
rect 13449 13923 13507 13929
rect 13280 13920 13400 13923
rect 13449 13920 13461 13923
rect 13280 13895 13461 13920
rect 13372 13892 13461 13895
rect 13449 13889 13461 13892
rect 13495 13889 13507 13923
rect 13449 13883 13507 13889
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13817 13923 13875 13929
rect 13817 13889 13829 13923
rect 13863 13920 13875 13923
rect 13906 13920 13912 13932
rect 13863 13892 13912 13920
rect 13863 13889 13875 13892
rect 13817 13883 13875 13889
rect 13262 13852 13268 13864
rect 13004 13824 13268 13852
rect 13262 13812 13268 13824
rect 13320 13812 13326 13864
rect 13556 13852 13584 13883
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 13998 13880 14004 13932
rect 14056 13880 14062 13932
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13889 14151 13923
rect 14093 13883 14151 13889
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 14274 13920 14280 13932
rect 14231 13892 14280 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 13630 13852 13636 13864
rect 13556 13824 13636 13852
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 14108 13852 14136 13883
rect 14274 13880 14280 13892
rect 14332 13880 14338 13932
rect 15381 13923 15439 13929
rect 15381 13889 15393 13923
rect 15427 13920 15439 13923
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15427 13892 15853 13920
rect 15427 13889 15439 13892
rect 15381 13883 15439 13889
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 15841 13883 15899 13889
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 16393 13923 16451 13929
rect 16393 13920 16405 13923
rect 16172 13892 16405 13920
rect 16172 13880 16178 13892
rect 16393 13889 16405 13892
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 14366 13852 14372 13864
rect 14108 13824 14372 13852
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 14461 13787 14519 13793
rect 12729 13756 13032 13784
rect 11790 13716 11796 13728
rect 2746 13688 11796 13716
rect 2317 13679 2375 13685
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12894 13676 12900 13728
rect 12952 13676 12958 13728
rect 13004 13716 13032 13756
rect 14461 13753 14473 13787
rect 14507 13784 14519 13787
rect 15580 13784 15608 13815
rect 14507 13756 15608 13784
rect 14507 13753 14519 13756
rect 14461 13747 14519 13753
rect 13538 13716 13544 13728
rect 13004 13688 13544 13716
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 1104 13626 16836 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 16836 13626
rect 1104 13552 16836 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2590 13512 2596 13524
rect 2372 13484 2596 13512
rect 2372 13472 2378 13484
rect 2590 13472 2596 13484
rect 2648 13512 2654 13524
rect 2777 13515 2835 13521
rect 2777 13512 2789 13515
rect 2648 13484 2789 13512
rect 2648 13472 2654 13484
rect 2777 13481 2789 13484
rect 2823 13481 2835 13515
rect 2777 13475 2835 13481
rect 13170 13472 13176 13524
rect 13228 13472 13234 13524
rect 13538 13472 13544 13524
rect 13596 13472 13602 13524
rect 13725 13515 13783 13521
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 13998 13512 14004 13524
rect 13771 13484 14004 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 2682 13404 2688 13456
rect 2740 13444 2746 13456
rect 3418 13444 3424 13456
rect 2740 13416 3424 13444
rect 2740 13404 2746 13416
rect 3418 13404 3424 13416
rect 3476 13404 3482 13456
rect 7929 13447 7987 13453
rect 7929 13413 7941 13447
rect 7975 13444 7987 13447
rect 7975 13416 9536 13444
rect 7975 13413 7987 13416
rect 7929 13407 7987 13413
rect 9508 13388 9536 13416
rect 12894 13404 12900 13456
rect 12952 13444 12958 13456
rect 13262 13444 13268 13456
rect 12952 13416 13268 13444
rect 12952 13404 12958 13416
rect 13262 13404 13268 13416
rect 13320 13444 13326 13456
rect 13556 13444 13584 13472
rect 13320 13416 13584 13444
rect 13320 13404 13326 13416
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 14274 13444 14280 13456
rect 13872 13416 14280 13444
rect 13872 13404 13878 13416
rect 14274 13404 14280 13416
rect 14332 13404 14338 13456
rect 3786 13336 3792 13388
rect 3844 13336 3850 13388
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 8665 13379 8723 13385
rect 6411 13348 6500 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 1397 13311 1455 13317
rect 1397 13277 1409 13311
rect 1443 13308 1455 13311
rect 2774 13308 2780 13320
rect 1443 13280 2780 13308
rect 1443 13277 1455 13280
rect 1397 13271 1455 13277
rect 2774 13268 2780 13280
rect 2832 13268 2838 13320
rect 1486 13200 1492 13252
rect 1544 13240 1550 13252
rect 1642 13243 1700 13249
rect 1642 13240 1654 13243
rect 1544 13212 1654 13240
rect 1544 13200 1550 13212
rect 1642 13209 1654 13212
rect 1688 13209 1700 13243
rect 1642 13203 1700 13209
rect 4056 13243 4114 13249
rect 4056 13209 4068 13243
rect 4102 13240 4114 13243
rect 4246 13240 4252 13252
rect 4102 13212 4252 13240
rect 4102 13209 4114 13212
rect 4056 13203 4114 13209
rect 4246 13200 4252 13212
rect 4304 13200 4310 13252
rect 6472 13240 6500 13348
rect 8665 13345 8677 13379
rect 8711 13376 8723 13379
rect 8846 13376 8852 13388
rect 8711 13348 8852 13376
rect 8711 13345 8723 13348
rect 8665 13339 8723 13345
rect 8846 13336 8852 13348
rect 8904 13336 8910 13388
rect 9490 13336 9496 13388
rect 9548 13336 9554 13388
rect 11238 13336 11244 13388
rect 11296 13376 11302 13388
rect 11333 13379 11391 13385
rect 11333 13376 11345 13379
rect 11296 13348 11345 13376
rect 11296 13336 11302 13348
rect 11333 13345 11345 13348
rect 11379 13345 11391 13379
rect 11333 13339 11391 13345
rect 12066 13336 12072 13388
rect 12124 13376 12130 13388
rect 12345 13379 12403 13385
rect 12345 13376 12357 13379
rect 12124 13348 12357 13376
rect 12124 13336 12130 13348
rect 12345 13345 12357 13348
rect 12391 13376 12403 13379
rect 12391 13348 13400 13376
rect 12391 13345 12403 13348
rect 12345 13339 12403 13345
rect 6549 13311 6607 13317
rect 6549 13277 6561 13311
rect 6595 13308 6607 13311
rect 6638 13308 6644 13320
rect 6595 13280 6644 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 8202 13308 8208 13320
rect 6748 13280 8208 13308
rect 6748 13240 6776 13280
rect 8202 13268 8208 13280
rect 8260 13268 8266 13320
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 10597 13311 10655 13317
rect 10597 13308 10609 13311
rect 10284 13280 10609 13308
rect 10284 13268 10290 13280
rect 10597 13277 10609 13280
rect 10643 13308 10655 13311
rect 11514 13308 11520 13320
rect 10643 13280 11520 13308
rect 10643 13277 10655 13280
rect 10597 13271 10655 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 6472 13212 6776 13240
rect 6816 13243 6874 13249
rect 6816 13209 6828 13243
rect 6862 13240 6874 13243
rect 6862 13212 8064 13240
rect 6862 13209 6874 13212
rect 6816 13203 6874 13209
rect 5169 13175 5227 13181
rect 5169 13141 5181 13175
rect 5215 13172 5227 13175
rect 5258 13172 5264 13184
rect 5215 13144 5264 13172
rect 5215 13141 5227 13144
rect 5169 13135 5227 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5718 13132 5724 13184
rect 5776 13132 5782 13184
rect 6086 13132 6092 13184
rect 6144 13132 6150 13184
rect 6178 13132 6184 13184
rect 6236 13132 6242 13184
rect 8036 13181 8064 13212
rect 9858 13200 9864 13252
rect 9916 13240 9922 13252
rect 11624 13240 11652 13271
rect 12526 13268 12532 13320
rect 12584 13268 12590 13320
rect 12618 13268 12624 13320
rect 12676 13308 12682 13320
rect 12897 13311 12955 13317
rect 12897 13308 12909 13311
rect 12676 13280 12909 13308
rect 12676 13268 12682 13280
rect 12897 13277 12909 13280
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 12989 13311 13047 13317
rect 12989 13277 13001 13311
rect 13035 13277 13047 13311
rect 12989 13271 13047 13277
rect 9916 13212 11652 13240
rect 9916 13200 9922 13212
rect 11790 13200 11796 13252
rect 11848 13240 11854 13252
rect 11848 13212 12434 13240
rect 11848 13200 11854 13212
rect 8021 13175 8079 13181
rect 8021 13141 8033 13175
rect 8067 13141 8079 13175
rect 8021 13135 8079 13141
rect 8386 13132 8392 13184
rect 8444 13132 8450 13184
rect 8481 13175 8539 13181
rect 8481 13141 8493 13175
rect 8527 13172 8539 13175
rect 8941 13175 8999 13181
rect 8941 13172 8953 13175
rect 8527 13144 8953 13172
rect 8527 13141 8539 13144
rect 8481 13135 8539 13141
rect 8941 13141 8953 13144
rect 8987 13141 8999 13175
rect 8941 13135 8999 13141
rect 11882 13132 11888 13184
rect 11940 13172 11946 13184
rect 12253 13175 12311 13181
rect 12253 13172 12265 13175
rect 11940 13144 12265 13172
rect 11940 13132 11946 13144
rect 12253 13141 12265 13144
rect 12299 13141 12311 13175
rect 12406 13172 12434 13212
rect 12710 13200 12716 13252
rect 12768 13240 12774 13252
rect 13004 13240 13032 13271
rect 13078 13268 13084 13320
rect 13136 13268 13142 13320
rect 13372 13317 13400 13348
rect 13446 13336 13452 13388
rect 13504 13336 13510 13388
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 14516 13348 14688 13376
rect 14516 13336 14522 13348
rect 13265 13311 13323 13317
rect 13265 13277 13277 13311
rect 13311 13277 13323 13311
rect 13265 13271 13323 13277
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 12768 13212 13032 13240
rect 12768 13200 12774 13212
rect 13170 13200 13176 13252
rect 13228 13240 13234 13252
rect 13280 13240 13308 13271
rect 13464 13240 13492 13336
rect 14274 13268 14280 13320
rect 14332 13268 14338 13320
rect 14660 13317 14688 13348
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13277 14703 13311
rect 14645 13271 14703 13277
rect 15749 13311 15807 13317
rect 15749 13277 15761 13311
rect 15795 13308 15807 13311
rect 15930 13308 15936 13320
rect 15795 13280 15936 13308
rect 15795 13277 15807 13280
rect 15749 13271 15807 13277
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 16390 13268 16396 13320
rect 16448 13268 16454 13320
rect 13228 13212 13492 13240
rect 13228 13200 13234 13212
rect 14182 13200 14188 13252
rect 14240 13240 14246 13252
rect 14366 13240 14372 13252
rect 14240 13212 14372 13240
rect 14240 13200 14246 13212
rect 14366 13200 14372 13212
rect 14424 13240 14430 13252
rect 14461 13243 14519 13249
rect 14461 13240 14473 13243
rect 14424 13212 14473 13240
rect 14424 13200 14430 13212
rect 14461 13209 14473 13212
rect 14507 13209 14519 13243
rect 14461 13203 14519 13209
rect 14553 13243 14611 13249
rect 14553 13209 14565 13243
rect 14599 13240 14611 13243
rect 15010 13240 15016 13252
rect 14599 13212 15016 13240
rect 14599 13209 14611 13212
rect 14553 13203 14611 13209
rect 14568 13172 14596 13203
rect 15010 13200 15016 13212
rect 15068 13200 15074 13252
rect 12406 13144 14596 13172
rect 14829 13175 14887 13181
rect 12253 13135 12311 13141
rect 14829 13141 14841 13175
rect 14875 13172 14887 13175
rect 15378 13172 15384 13184
rect 14875 13144 15384 13172
rect 14875 13141 14887 13144
rect 14829 13135 14887 13141
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15562 13132 15568 13184
rect 15620 13132 15626 13184
rect 15838 13132 15844 13184
rect 15896 13132 15902 13184
rect 1104 13082 16836 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 16836 13082
rect 1104 13008 16836 13030
rect 1302 12928 1308 12980
rect 1360 12968 1366 12980
rect 1489 12971 1547 12977
rect 1489 12968 1501 12971
rect 1360 12940 1501 12968
rect 1360 12928 1366 12940
rect 1489 12937 1501 12940
rect 1535 12937 1547 12971
rect 3329 12971 3387 12977
rect 1489 12931 1547 12937
rect 1688 12940 3188 12968
rect 1688 12841 1716 12940
rect 2774 12900 2780 12912
rect 1964 12872 2780 12900
rect 1964 12841 1992 12872
rect 2774 12860 2780 12872
rect 2832 12860 2838 12912
rect 2222 12841 2228 12844
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12801 2007 12835
rect 2216 12832 2228 12841
rect 2183 12804 2228 12832
rect 1949 12795 2007 12801
rect 2216 12795 2228 12804
rect 2222 12792 2228 12795
rect 2280 12792 2286 12844
rect 3160 12832 3188 12940
rect 3329 12937 3341 12971
rect 3375 12937 3387 12971
rect 3329 12931 3387 12937
rect 3881 12971 3939 12977
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 3970 12968 3976 12980
rect 3927 12940 3976 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 3344 12900 3372 12931
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4246 12928 4252 12980
rect 4304 12928 4310 12980
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6457 12971 6515 12977
rect 6457 12968 6469 12971
rect 6144 12940 6469 12968
rect 6144 12928 6150 12940
rect 6457 12937 6469 12940
rect 6503 12937 6515 12971
rect 6457 12931 6515 12937
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 8110 12968 8116 12980
rect 7156 12940 8116 12968
rect 7156 12928 7162 12940
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 9033 12971 9091 12977
rect 9033 12937 9045 12971
rect 9079 12968 9091 12971
rect 9306 12968 9312 12980
rect 9079 12940 9312 12968
rect 9079 12937 9091 12940
rect 9033 12931 9091 12937
rect 9306 12928 9312 12940
rect 9364 12928 9370 12980
rect 9493 12971 9551 12977
rect 9493 12937 9505 12971
rect 9539 12968 9551 12971
rect 9858 12968 9864 12980
rect 9539 12940 9864 12968
rect 9539 12937 9551 12940
rect 9493 12931 9551 12937
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 11517 12971 11575 12977
rect 11517 12937 11529 12971
rect 11563 12937 11575 12971
rect 11517 12931 11575 12937
rect 3418 12900 3424 12912
rect 3344 12872 3424 12900
rect 3418 12860 3424 12872
rect 3476 12900 3482 12912
rect 10996 12903 11054 12909
rect 3476 12872 10364 12900
rect 3476 12860 3482 12872
rect 3160 12804 4660 12832
rect 3602 12724 3608 12776
rect 3660 12724 3666 12776
rect 3789 12767 3847 12773
rect 3789 12733 3801 12767
rect 3835 12764 3847 12767
rect 4062 12764 4068 12776
rect 3835 12736 4068 12764
rect 3835 12733 3847 12736
rect 3789 12727 3847 12733
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 4632 12764 4660 12804
rect 7098 12792 7104 12844
rect 7156 12792 7162 12844
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12832 7343 12835
rect 7374 12832 7380 12844
rect 7331 12804 7380 12832
rect 7331 12801 7343 12804
rect 7285 12795 7343 12801
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 7469 12835 7527 12841
rect 7469 12801 7481 12835
rect 7515 12801 7527 12835
rect 7469 12795 7527 12801
rect 7561 12835 7619 12841
rect 7561 12801 7573 12835
rect 7607 12832 7619 12835
rect 8294 12832 8300 12844
rect 7607 12804 8300 12832
rect 7607 12801 7619 12804
rect 7561 12795 7619 12801
rect 4706 12764 4712 12776
rect 4632 12736 4712 12764
rect 4706 12724 4712 12736
rect 4764 12764 4770 12776
rect 7484 12764 7512 12795
rect 8294 12792 8300 12804
rect 8352 12792 8358 12844
rect 9401 12835 9459 12841
rect 9401 12801 9413 12835
rect 9447 12832 9459 12835
rect 10226 12832 10232 12844
rect 9447 12804 10232 12832
rect 9447 12801 9459 12804
rect 9401 12795 9459 12801
rect 10226 12792 10232 12804
rect 10284 12792 10290 12844
rect 10336 12832 10364 12872
rect 10996 12869 11008 12903
rect 11042 12900 11054 12903
rect 11532 12900 11560 12931
rect 11882 12928 11888 12980
rect 11940 12928 11946 12980
rect 13357 12971 13415 12977
rect 13357 12937 13369 12971
rect 13403 12937 13415 12971
rect 13357 12931 13415 12937
rect 14093 12971 14151 12977
rect 14093 12937 14105 12971
rect 14139 12968 14151 12971
rect 15746 12968 15752 12980
rect 14139 12940 15752 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 11042 12872 11560 12900
rect 11624 12872 13308 12900
rect 11042 12869 11054 12872
rect 10996 12863 11054 12869
rect 11624 12832 11652 12872
rect 10336 12804 11652 12832
rect 11977 12835 12035 12841
rect 11977 12801 11989 12835
rect 12023 12832 12035 12835
rect 12158 12832 12164 12844
rect 12023 12804 12164 12832
rect 12023 12801 12035 12804
rect 11977 12795 12035 12801
rect 12158 12792 12164 12804
rect 12216 12832 12222 12844
rect 12618 12832 12624 12844
rect 12216 12804 12624 12832
rect 12216 12792 12222 12804
rect 12618 12792 12624 12804
rect 12676 12792 12682 12844
rect 12894 12792 12900 12844
rect 12952 12832 12958 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12952 12804 13001 12832
rect 12952 12792 12958 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13170 12792 13176 12844
rect 13228 12792 13234 12844
rect 4764 12736 7512 12764
rect 4764 12724 4770 12736
rect 8110 12724 8116 12776
rect 8168 12724 8174 12776
rect 8662 12724 8668 12776
rect 8720 12724 8726 12776
rect 9585 12767 9643 12773
rect 9585 12733 9597 12767
rect 9631 12733 9643 12767
rect 9585 12727 9643 12733
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 11330 12764 11336 12776
rect 11287 12736 11336 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 7745 12699 7803 12705
rect 7745 12665 7757 12699
rect 7791 12696 7803 12699
rect 9030 12696 9036 12708
rect 7791 12668 9036 12696
rect 7791 12665 7803 12668
rect 7745 12659 7803 12665
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 2314 12588 2320 12640
rect 2372 12628 2378 12640
rect 2682 12628 2688 12640
rect 2372 12600 2688 12628
rect 2372 12588 2378 12600
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 7926 12588 7932 12640
rect 7984 12628 7990 12640
rect 9600 12628 9628 12727
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 12069 12767 12127 12773
rect 12069 12733 12081 12767
rect 12115 12764 12127 12767
rect 12342 12764 12348 12776
rect 12115 12736 12348 12764
rect 12115 12733 12127 12736
rect 12069 12727 12127 12733
rect 12342 12724 12348 12736
rect 12400 12724 12406 12776
rect 13280 12764 13308 12872
rect 13372 12832 13400 12931
rect 15746 12928 15752 12940
rect 15804 12928 15810 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 16172 12940 16221 12968
rect 16172 12928 16178 12940
rect 16209 12937 16221 12940
rect 16255 12968 16267 12971
rect 16390 12968 16396 12980
rect 16255 12940 16396 12968
rect 16255 12937 16267 12940
rect 16209 12931 16267 12937
rect 16390 12928 16396 12940
rect 16448 12928 16454 12980
rect 13906 12900 13912 12912
rect 13648 12872 13912 12900
rect 13648 12841 13676 12872
rect 13906 12860 13912 12872
rect 13964 12860 13970 12912
rect 14366 12860 14372 12912
rect 14424 12860 14430 12912
rect 15096 12903 15154 12909
rect 15096 12869 15108 12903
rect 15142 12900 15154 12903
rect 15194 12900 15200 12912
rect 15142 12872 15200 12900
rect 15142 12869 15154 12872
rect 15096 12863 15154 12869
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13372 12804 13461 12832
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13633 12835 13691 12841
rect 13633 12801 13645 12835
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 13722 12792 13728 12844
rect 13780 12792 13786 12844
rect 13814 12792 13820 12844
rect 13872 12792 13878 12844
rect 14182 12792 14188 12844
rect 14240 12792 14246 12844
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 14476 12764 14504 12795
rect 14550 12792 14556 12844
rect 14608 12792 14614 12844
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14792 12804 14841 12832
rect 14792 12792 14798 12804
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 16482 12792 16488 12844
rect 16540 12792 16546 12844
rect 14936 12764 14964 12792
rect 13280 12736 14964 12764
rect 12802 12656 12808 12708
rect 12860 12696 12866 12708
rect 13722 12696 13728 12708
rect 12860 12668 13728 12696
rect 12860 12656 12866 12668
rect 13722 12656 13728 12668
rect 13780 12656 13786 12708
rect 13906 12656 13912 12708
rect 13964 12696 13970 12708
rect 14550 12696 14556 12708
rect 13964 12668 14556 12696
rect 13964 12656 13970 12668
rect 14550 12656 14556 12668
rect 14608 12656 14614 12708
rect 16022 12656 16028 12708
rect 16080 12696 16086 12708
rect 16301 12699 16359 12705
rect 16301 12696 16313 12699
rect 16080 12668 16313 12696
rect 16080 12656 16086 12668
rect 16301 12665 16313 12668
rect 16347 12665 16359 12699
rect 16301 12659 16359 12665
rect 10134 12628 10140 12640
rect 7984 12600 10140 12628
rect 7984 12588 7990 12600
rect 10134 12588 10140 12600
rect 10192 12628 10198 12640
rect 10502 12628 10508 12640
rect 10192 12600 10508 12628
rect 10192 12588 10198 12600
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 12986 12588 12992 12640
rect 13044 12588 13050 12640
rect 14737 12631 14795 12637
rect 14737 12597 14749 12631
rect 14783 12628 14795 12631
rect 15562 12628 15568 12640
rect 14783 12600 15568 12628
rect 14783 12597 14795 12600
rect 14737 12591 14795 12597
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 1104 12538 16836 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 16836 12538
rect 1104 12464 16836 12486
rect 4062 12384 4068 12436
rect 4120 12424 4126 12436
rect 5258 12424 5264 12436
rect 4120 12396 5264 12424
rect 4120 12384 4126 12396
rect 5258 12384 5264 12396
rect 5316 12424 5322 12436
rect 6546 12424 6552 12436
rect 5316 12396 6552 12424
rect 5316 12384 5322 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 6733 12427 6791 12433
rect 6733 12393 6745 12427
rect 6779 12424 6791 12427
rect 7098 12424 7104 12436
rect 6779 12396 7104 12424
rect 6779 12393 6791 12396
rect 6733 12387 6791 12393
rect 7098 12384 7104 12396
rect 7156 12384 7162 12436
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 8478 12424 8484 12436
rect 8352 12396 8484 12424
rect 8352 12384 8358 12396
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 10318 12384 10324 12436
rect 10376 12384 10382 12436
rect 13909 12427 13967 12433
rect 13909 12393 13921 12427
rect 13955 12424 13967 12427
rect 14182 12424 14188 12436
rect 13955 12396 14188 12424
rect 13955 12393 13967 12396
rect 13909 12387 13967 12393
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 15194 12384 15200 12436
rect 15252 12384 15258 12436
rect 5350 12356 5356 12368
rect 2056 12328 5356 12356
rect 1670 12180 1676 12232
rect 1728 12180 1734 12232
rect 2056 12229 2084 12328
rect 5350 12316 5356 12328
rect 5408 12316 5414 12368
rect 3878 12248 3884 12300
rect 3936 12288 3942 12300
rect 8021 12291 8079 12297
rect 3936 12260 4108 12288
rect 3936 12248 3942 12260
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2685 12223 2743 12229
rect 2685 12189 2697 12223
rect 2731 12220 2743 12223
rect 2958 12220 2964 12232
rect 2731 12192 2964 12220
rect 2731 12189 2743 12192
rect 2685 12183 2743 12189
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 4080 12229 4108 12260
rect 8021 12257 8033 12291
rect 8067 12288 8079 12291
rect 8202 12288 8208 12300
rect 8067 12260 8208 12288
rect 8067 12257 8079 12260
rect 8021 12251 8079 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8938 12248 8944 12300
rect 8996 12248 9002 12300
rect 10336 12288 10364 12384
rect 16390 12316 16396 12368
rect 16448 12316 16454 12368
rect 10965 12291 11023 12297
rect 10965 12288 10977 12291
rect 10336 12260 10977 12288
rect 10965 12257 10977 12260
rect 11011 12257 11023 12291
rect 10965 12251 11023 12257
rect 11885 12291 11943 12297
rect 11885 12257 11897 12291
rect 11931 12288 11943 12291
rect 11974 12288 11980 12300
rect 11931 12260 11980 12288
rect 11931 12257 11943 12260
rect 11885 12251 11943 12257
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 12526 12288 12532 12300
rect 12176 12260 12532 12288
rect 4065 12223 4123 12229
rect 4065 12189 4077 12223
rect 4111 12189 4123 12223
rect 4065 12183 4123 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12189 4215 12223
rect 4157 12183 4215 12189
rect 4249 12223 4307 12229
rect 4249 12189 4261 12223
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 3878 12112 3884 12164
rect 3936 12152 3942 12164
rect 4172 12152 4200 12183
rect 3936 12124 4200 12152
rect 3936 12112 3942 12124
rect 842 12044 848 12096
rect 900 12084 906 12096
rect 1489 12087 1547 12093
rect 1489 12084 1501 12087
rect 900 12056 1501 12084
rect 900 12044 906 12056
rect 1489 12053 1501 12056
rect 1535 12053 1547 12087
rect 1489 12047 1547 12053
rect 1854 12044 1860 12096
rect 1912 12044 1918 12096
rect 2501 12087 2559 12093
rect 2501 12053 2513 12087
rect 2547 12084 2559 12087
rect 3050 12084 3056 12096
rect 2547 12056 3056 12084
rect 2547 12053 2559 12056
rect 2501 12047 2559 12053
rect 3050 12044 3056 12056
rect 3108 12044 3114 12096
rect 3602 12044 3608 12096
rect 3660 12084 3666 12096
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 3660 12056 3801 12084
rect 3660 12044 3666 12056
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 4264 12084 4292 12183
rect 4430 12180 4436 12232
rect 4488 12180 4494 12232
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12220 5411 12223
rect 6638 12220 6644 12232
rect 5399 12192 6644 12220
rect 5399 12189 5411 12192
rect 5353 12183 5411 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8110 12220 8116 12232
rect 7791 12192 8116 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 8665 12223 8723 12229
rect 8665 12189 8677 12223
rect 8711 12220 8723 12223
rect 8754 12220 8760 12232
rect 8711 12192 8760 12220
rect 8711 12189 8723 12192
rect 8665 12183 8723 12189
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 10100 12192 11161 12220
rect 10100 12180 10106 12192
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 11606 12180 11612 12232
rect 11664 12220 11670 12232
rect 12066 12220 12072 12232
rect 11664 12192 12072 12220
rect 11664 12180 11670 12192
rect 12066 12180 12072 12192
rect 12124 12180 12130 12232
rect 12176 12229 12204 12260
rect 12526 12248 12532 12260
rect 12584 12288 12590 12300
rect 13170 12288 13176 12300
rect 12584 12260 13176 12288
rect 12584 12248 12590 12260
rect 13170 12248 13176 12260
rect 13228 12248 13234 12300
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12288 13323 12291
rect 13814 12288 13820 12300
rect 13311 12260 13820 12288
rect 13311 12257 13323 12260
rect 13265 12251 13323 12257
rect 13814 12248 13820 12260
rect 13872 12288 13878 12300
rect 14734 12288 14740 12300
rect 13872 12260 14740 12288
rect 13872 12248 13878 12260
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15562 12248 15568 12300
rect 15620 12288 15626 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15620 12260 15669 12288
rect 15620 12248 15626 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15746 12248 15752 12300
rect 15804 12248 15810 12300
rect 12161 12223 12219 12229
rect 12161 12189 12173 12223
rect 12207 12189 12219 12223
rect 12161 12183 12219 12189
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 13541 12223 13599 12229
rect 13541 12220 13553 12223
rect 13044 12192 13553 12220
rect 13044 12180 13050 12192
rect 13541 12189 13553 12192
rect 13587 12189 13599 12223
rect 13541 12183 13599 12189
rect 13725 12223 13783 12229
rect 13725 12189 13737 12223
rect 13771 12220 13783 12223
rect 13998 12220 14004 12232
rect 13771 12192 14004 12220
rect 13771 12189 13783 12192
rect 13725 12183 13783 12189
rect 13998 12180 14004 12192
rect 14056 12220 14062 12232
rect 14366 12220 14372 12232
rect 14056 12192 14372 12220
rect 14056 12180 14062 12192
rect 14366 12180 14372 12192
rect 14424 12180 14430 12232
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12220 14611 12223
rect 16022 12220 16028 12232
rect 14599 12192 16028 12220
rect 14599 12189 14611 12192
rect 14553 12183 14611 12189
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 16209 12223 16267 12229
rect 16209 12189 16221 12223
rect 16255 12220 16267 12223
rect 16298 12220 16304 12232
rect 16255 12192 16304 12220
rect 16255 12189 16267 12192
rect 16209 12183 16267 12189
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 4525 12155 4583 12161
rect 4525 12121 4537 12155
rect 4571 12121 4583 12155
rect 4525 12115 4583 12121
rect 5620 12155 5678 12161
rect 5620 12121 5632 12155
rect 5666 12152 5678 12155
rect 5718 12152 5724 12164
rect 5666 12124 5724 12152
rect 5666 12121 5678 12124
rect 5620 12115 5678 12121
rect 4120 12056 4292 12084
rect 4120 12044 4126 12056
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4540 12084 4568 12115
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 9208 12155 9266 12161
rect 9208 12121 9220 12155
rect 9254 12152 9266 12155
rect 9490 12152 9496 12164
rect 9254 12124 9496 12152
rect 9254 12121 9266 12124
rect 9208 12115 9266 12121
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 11514 12112 11520 12164
rect 11572 12152 11578 12164
rect 11974 12152 11980 12164
rect 11572 12124 11980 12152
rect 11572 12112 11578 12124
rect 11974 12112 11980 12124
rect 12032 12152 12038 12164
rect 12437 12155 12495 12161
rect 12437 12152 12449 12155
rect 12032 12124 12449 12152
rect 12032 12112 12038 12124
rect 12437 12121 12449 12124
rect 12483 12121 12495 12155
rect 12437 12115 12495 12121
rect 15565 12155 15623 12161
rect 15565 12121 15577 12155
rect 15611 12152 15623 12155
rect 15838 12152 15844 12164
rect 15611 12124 15844 12152
rect 15611 12121 15623 12124
rect 15565 12115 15623 12121
rect 15838 12112 15844 12124
rect 15896 12112 15902 12164
rect 4396 12056 4568 12084
rect 4396 12044 4402 12056
rect 4798 12044 4804 12096
rect 4856 12084 4862 12096
rect 4893 12087 4951 12093
rect 4893 12084 4905 12087
rect 4856 12056 4905 12084
rect 4856 12044 4862 12056
rect 4893 12053 4905 12056
rect 4939 12053 4951 12087
rect 4893 12047 4951 12053
rect 7374 12044 7380 12096
rect 7432 12044 7438 12096
rect 7834 12044 7840 12096
rect 7892 12044 7898 12096
rect 8294 12044 8300 12096
rect 8352 12084 8358 12096
rect 8573 12087 8631 12093
rect 8573 12084 8585 12087
rect 8352 12056 8585 12084
rect 8352 12044 8358 12056
rect 8573 12053 8585 12056
rect 8619 12084 8631 12087
rect 8938 12084 8944 12096
rect 8619 12056 8944 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 8938 12044 8944 12056
rect 8996 12044 9002 12096
rect 10410 12044 10416 12096
rect 10468 12044 10474 12096
rect 11790 12044 11796 12096
rect 11848 12044 11854 12096
rect 11882 12044 11888 12096
rect 11940 12044 11946 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15470 12084 15476 12096
rect 15151 12056 15476 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 1104 11994 16836 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 16836 11994
rect 1104 11920 16836 11942
rect 3786 11880 3792 11892
rect 1688 11852 3792 11880
rect 1688 11821 1716 11852
rect 3786 11840 3792 11852
rect 3844 11880 3850 11892
rect 4338 11880 4344 11892
rect 3844 11852 4344 11880
rect 3844 11840 3850 11852
rect 4338 11840 4344 11852
rect 4396 11840 4402 11892
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 6181 11883 6239 11889
rect 6181 11880 6193 11883
rect 4764 11852 6193 11880
rect 4764 11840 4770 11852
rect 6181 11849 6193 11852
rect 6227 11849 6239 11883
rect 6181 11843 6239 11849
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8662 11880 8668 11892
rect 8343 11852 8668 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 9030 11840 9036 11892
rect 9088 11840 9094 11892
rect 9490 11840 9496 11892
rect 9548 11840 9554 11892
rect 9953 11883 10011 11889
rect 9953 11849 9965 11883
rect 9999 11880 10011 11883
rect 10042 11880 10048 11892
rect 9999 11852 10048 11880
rect 9999 11849 10011 11852
rect 9953 11843 10011 11849
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11849 11575 11883
rect 11517 11843 11575 11849
rect 1673 11815 1731 11821
rect 1673 11781 1685 11815
rect 1719 11781 1731 11815
rect 1673 11775 1731 11781
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 2866 11812 2872 11824
rect 1903 11784 2872 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 2866 11772 2872 11784
rect 2924 11772 2930 11824
rect 3344 11784 4844 11812
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3344 11753 3372 11784
rect 3602 11753 3608 11756
rect 3329 11747 3387 11753
rect 3329 11744 3341 11747
rect 2832 11716 3341 11744
rect 2832 11704 2838 11716
rect 3329 11713 3341 11716
rect 3375 11713 3387 11747
rect 3596 11744 3608 11753
rect 3563 11716 3608 11744
rect 3329 11707 3387 11713
rect 3596 11707 3608 11716
rect 3602 11704 3608 11707
rect 3660 11704 3666 11756
rect 4816 11753 4844 11784
rect 4890 11772 4896 11824
rect 4948 11812 4954 11824
rect 5534 11812 5540 11824
rect 4948 11784 5540 11812
rect 4948 11772 4954 11784
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 7184 11815 7242 11821
rect 7184 11781 7196 11815
rect 7230 11812 7242 11815
rect 7374 11812 7380 11824
rect 7230 11784 7380 11812
rect 7230 11781 7242 11784
rect 7184 11775 7242 11781
rect 7374 11772 7380 11784
rect 7432 11772 7438 11824
rect 9125 11815 9183 11821
rect 9125 11781 9137 11815
rect 9171 11812 9183 11815
rect 10410 11812 10416 11824
rect 9171 11784 10416 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 10410 11772 10416 11784
rect 10468 11772 10474 11824
rect 11088 11815 11146 11821
rect 11088 11781 11100 11815
rect 11134 11812 11146 11815
rect 11532 11812 11560 11843
rect 11790 11840 11796 11892
rect 11848 11880 11854 11892
rect 11848 11852 12112 11880
rect 11848 11840 11854 11852
rect 11134 11784 11560 11812
rect 11134 11781 11146 11784
rect 11088 11775 11146 11781
rect 11882 11772 11888 11824
rect 11940 11772 11946 11824
rect 5074 11753 5080 11756
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 5068 11707 5080 11753
rect 5074 11704 5080 11707
rect 5132 11704 5138 11756
rect 6638 11704 6644 11756
rect 6696 11744 6702 11756
rect 6917 11747 6975 11753
rect 6917 11744 6929 11747
rect 6696 11716 6929 11744
rect 6696 11704 6702 11716
rect 6917 11713 6929 11716
rect 6963 11713 6975 11747
rect 6917 11707 6975 11713
rect 11330 11704 11336 11756
rect 11388 11704 11394 11756
rect 11606 11704 11612 11756
rect 11664 11744 11670 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11664 11716 11713 11744
rect 11664 11704 11670 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11790 11704 11796 11756
rect 11848 11704 11854 11756
rect 12084 11753 12112 11852
rect 12618 11840 12624 11892
rect 12676 11840 12682 11892
rect 14274 11840 14280 11892
rect 14332 11880 14338 11892
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 14332 11852 14749 11880
rect 14332 11840 14338 11852
rect 14737 11849 14749 11852
rect 14783 11849 14795 11883
rect 14737 11843 14795 11849
rect 15470 11840 15476 11892
rect 15528 11840 15534 11892
rect 15930 11840 15936 11892
rect 15988 11840 15994 11892
rect 12636 11812 12664 11840
rect 13354 11812 13360 11824
rect 12360 11784 13360 11812
rect 12069 11747 12127 11753
rect 12069 11713 12081 11747
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 12158 11704 12164 11756
rect 12216 11704 12222 11756
rect 12360 11753 12388 11784
rect 13354 11772 13360 11784
rect 13412 11772 13418 11824
rect 12345 11747 12403 11753
rect 12345 11713 12357 11747
rect 12391 11713 12403 11747
rect 12345 11707 12403 11713
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 13814 11744 13820 11756
rect 12667 11716 13820 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 2958 11636 2964 11688
rect 3016 11636 3022 11688
rect 3234 11636 3240 11688
rect 3292 11636 3298 11688
rect 8938 11636 8944 11688
rect 8996 11676 9002 11688
rect 9582 11676 9588 11688
rect 8996 11648 9588 11676
rect 8996 11636 9002 11648
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 11348 11676 11376 11704
rect 12636 11676 12664 11707
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 13998 11704 14004 11756
rect 14056 11744 14062 11756
rect 14642 11744 14648 11756
rect 14056 11716 14648 11744
rect 14056 11704 14062 11716
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 11348 11648 12664 11676
rect 13170 11636 13176 11688
rect 13228 11676 13234 11688
rect 14844 11676 14872 11707
rect 16114 11704 16120 11756
rect 16172 11704 16178 11756
rect 16206 11704 16212 11756
rect 16264 11704 16270 11756
rect 13228 11648 14872 11676
rect 13228 11636 13234 11648
rect 15562 11636 15568 11688
rect 15620 11636 15626 11688
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 1670 11568 1676 11620
rect 1728 11608 1734 11620
rect 1728 11580 2774 11608
rect 1728 11568 1734 11580
rect 2041 11543 2099 11549
rect 2041 11509 2053 11543
rect 2087 11540 2099 11543
rect 2130 11540 2136 11552
rect 2087 11512 2136 11540
rect 2087 11509 2099 11512
rect 2041 11503 2099 11509
rect 2130 11500 2136 11512
rect 2188 11500 2194 11552
rect 2746 11540 2774 11580
rect 13906 11568 13912 11620
rect 13964 11608 13970 11620
rect 15672 11608 15700 11639
rect 13964 11580 15700 11608
rect 13964 11568 13970 11580
rect 16390 11568 16396 11620
rect 16448 11568 16454 11620
rect 3970 11540 3976 11552
rect 2746 11512 3976 11540
rect 3970 11500 3976 11512
rect 4028 11540 4034 11552
rect 4709 11543 4767 11549
rect 4709 11540 4721 11543
rect 4028 11512 4721 11540
rect 4028 11500 4034 11512
rect 4709 11509 4721 11512
rect 4755 11540 4767 11543
rect 5534 11540 5540 11552
rect 4755 11512 5540 11540
rect 4755 11509 4767 11512
rect 4709 11503 4767 11509
rect 5534 11500 5540 11512
rect 5592 11500 5598 11552
rect 12253 11543 12311 11549
rect 12253 11509 12265 11543
rect 12299 11540 12311 11543
rect 12434 11540 12440 11552
rect 12299 11512 12440 11540
rect 12299 11509 12311 11512
rect 12253 11503 12311 11509
rect 12434 11500 12440 11512
rect 12492 11500 12498 11552
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 14550 11540 14556 11552
rect 13228 11512 14556 11540
rect 13228 11500 13234 11512
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 15102 11500 15108 11552
rect 15160 11500 15166 11552
rect 1104 11450 16836 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 16836 11450
rect 1104 11376 16836 11398
rect 1118 11296 1124 11348
rect 1176 11336 1182 11348
rect 1489 11339 1547 11345
rect 1489 11336 1501 11339
rect 1176 11308 1501 11336
rect 1176 11296 1182 11308
rect 1489 11305 1501 11308
rect 1535 11305 1547 11339
rect 1489 11299 1547 11305
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 3694 11336 3700 11348
rect 3016 11308 3700 11336
rect 3016 11296 3022 11308
rect 3694 11296 3700 11308
rect 3752 11296 3758 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4157 11339 4215 11345
rect 4157 11336 4169 11339
rect 4120 11308 4169 11336
rect 4120 11296 4126 11308
rect 4157 11305 4169 11308
rect 4203 11305 4215 11339
rect 4157 11299 4215 11305
rect 4985 11339 5043 11345
rect 4985 11305 4997 11339
rect 5031 11336 5043 11339
rect 5074 11336 5080 11348
rect 5031 11308 5080 11336
rect 5031 11305 5043 11308
rect 4985 11299 5043 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 6917 11339 6975 11345
rect 6917 11305 6929 11339
rect 6963 11336 6975 11339
rect 7006 11336 7012 11348
rect 6963 11308 7012 11336
rect 6963 11305 6975 11308
rect 6917 11299 6975 11305
rect 7006 11296 7012 11308
rect 7064 11296 7070 11348
rect 8386 11296 8392 11348
rect 8444 11336 8450 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8444 11308 8585 11336
rect 8444 11296 8450 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 9677 11339 9735 11345
rect 9677 11305 9689 11339
rect 9723 11336 9735 11339
rect 9950 11336 9956 11348
rect 9723 11308 9956 11336
rect 9723 11305 9735 11308
rect 9677 11299 9735 11305
rect 9950 11296 9956 11308
rect 10008 11296 10014 11348
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 12894 11336 12900 11348
rect 11848 11308 12900 11336
rect 11848 11296 11854 11308
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13814 11336 13820 11348
rect 13044 11308 13820 11336
rect 13044 11296 13050 11308
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 13906 11296 13912 11348
rect 13964 11296 13970 11348
rect 14645 11339 14703 11345
rect 14645 11305 14657 11339
rect 14691 11336 14703 11339
rect 15562 11336 15568 11348
rect 14691 11308 15568 11336
rect 14691 11305 14703 11308
rect 14645 11299 14703 11305
rect 15562 11296 15568 11308
rect 15620 11296 15626 11348
rect 16022 11296 16028 11348
rect 16080 11336 16086 11348
rect 16209 11339 16267 11345
rect 16209 11336 16221 11339
rect 16080 11308 16221 11336
rect 16080 11296 16086 11308
rect 16209 11305 16221 11308
rect 16255 11305 16267 11339
rect 16209 11299 16267 11305
rect 2866 11228 2872 11280
rect 2924 11268 2930 11280
rect 3145 11271 3203 11277
rect 3145 11268 3157 11271
rect 2924 11240 3157 11268
rect 2924 11228 2930 11240
rect 3145 11237 3157 11240
rect 3191 11268 3203 11271
rect 3418 11268 3424 11280
rect 3191 11240 3424 11268
rect 3191 11237 3203 11240
rect 3145 11231 3203 11237
rect 3418 11228 3424 11240
rect 3476 11228 3482 11280
rect 4614 11268 4620 11280
rect 4428 11240 4620 11268
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1688 11064 1716 11095
rect 1762 11092 1768 11144
rect 1820 11092 1826 11144
rect 2866 11132 2872 11144
rect 1964 11104 2872 11132
rect 1964 11064 1992 11104
rect 2866 11092 2872 11104
rect 2924 11092 2930 11144
rect 3786 11092 3792 11144
rect 3844 11092 3850 11144
rect 3970 11092 3976 11144
rect 4028 11092 4034 11144
rect 4341 11135 4399 11141
rect 4341 11132 4353 11135
rect 4071 11104 4353 11132
rect 2038 11073 2044 11076
rect 1688 11036 1992 11064
rect 2032 11027 2044 11073
rect 2038 11024 2044 11027
rect 2096 11024 2102 11076
rect 2222 11024 2228 11076
rect 2280 11064 2286 11076
rect 3050 11064 3056 11076
rect 2280 11036 3056 11064
rect 2280 11024 2286 11036
rect 3050 11024 3056 11036
rect 3108 11064 3114 11076
rect 4071 11064 4099 11104
rect 4341 11101 4353 11104
rect 4387 11132 4399 11135
rect 4428 11132 4456 11240
rect 4614 11228 4620 11240
rect 4672 11228 4678 11280
rect 6546 11228 6552 11280
rect 6604 11268 6610 11280
rect 11514 11268 11520 11280
rect 6604 11240 11520 11268
rect 6604 11228 6610 11240
rect 11514 11228 11520 11240
rect 11572 11268 11578 11280
rect 13078 11268 13084 11280
rect 11572 11240 12112 11268
rect 11572 11228 11578 11240
rect 4798 11200 4804 11212
rect 4540 11172 4804 11200
rect 4540 11141 4568 11172
rect 4798 11160 4804 11172
rect 4856 11160 4862 11212
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 7926 11200 7932 11212
rect 7607 11172 7932 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11200 8171 11203
rect 8159 11172 9996 11200
rect 8159 11169 8171 11172
rect 8113 11163 8171 11169
rect 4387 11104 4456 11132
rect 4525 11135 4583 11141
rect 4387 11101 4399 11104
rect 4341 11095 4399 11101
rect 4525 11101 4537 11135
rect 4571 11101 4583 11135
rect 4525 11095 4583 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11132 4767 11135
rect 4890 11132 4896 11144
rect 4755 11104 4896 11132
rect 4755 11101 4767 11104
rect 4709 11095 4767 11101
rect 3108 11036 4099 11064
rect 3108 11024 3114 11036
rect 4246 11024 4252 11076
rect 4304 11064 4310 11076
rect 4632 11064 4660 11095
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5445 11135 5503 11141
rect 5445 11101 5457 11135
rect 5491 11132 5503 11135
rect 6638 11132 6644 11144
rect 5491 11104 6644 11132
rect 5491 11101 5503 11104
rect 5445 11095 5503 11101
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 8205 11135 8263 11141
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 8662 11132 8668 11144
rect 8251 11104 8668 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 8662 11092 8668 11104
rect 8720 11092 8726 11144
rect 9968 11132 9996 11172
rect 10042 11160 10048 11212
rect 10100 11200 10106 11212
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 10100 11172 10149 11200
rect 10100 11160 10106 11172
rect 10137 11169 10149 11172
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10502 11200 10508 11212
rect 10367 11172 10508 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 11974 11200 11980 11212
rect 11900 11172 11980 11200
rect 11330 11132 11336 11144
rect 9968 11104 11336 11132
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 11790 11092 11796 11144
rect 11848 11092 11854 11144
rect 11900 11141 11928 11172
rect 11974 11160 11980 11172
rect 12032 11160 12038 11212
rect 12084 11200 12112 11240
rect 12268 11240 13084 11268
rect 12268 11200 12296 11240
rect 13078 11228 13084 11240
rect 13136 11228 13142 11280
rect 13188 11240 14136 11268
rect 12084 11172 12296 11200
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11200 12403 11203
rect 13188 11200 13216 11240
rect 12391 11172 13216 11200
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13449 11203 13507 11209
rect 13449 11200 13461 11203
rect 13320 11172 13461 11200
rect 13320 11160 13326 11172
rect 13449 11169 13461 11172
rect 13495 11169 13507 11203
rect 13449 11163 13507 11169
rect 13538 11160 13544 11212
rect 13596 11160 13602 11212
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11101 11943 11135
rect 11885 11095 11943 11101
rect 12158 11092 12164 11144
rect 12216 11092 12222 11144
rect 12250 11092 12256 11144
rect 12308 11092 12314 11144
rect 12437 11135 12495 11141
rect 12437 11101 12449 11135
rect 12483 11132 12495 11135
rect 12526 11132 12532 11144
rect 12483 11104 12532 11132
rect 12483 11101 12495 11104
rect 12437 11095 12495 11101
rect 4304 11036 4660 11064
rect 5712 11067 5770 11073
rect 4304 11024 4310 11036
rect 5712 11033 5724 11067
rect 5758 11064 5770 11067
rect 6270 11064 6276 11076
rect 5758 11036 6276 11064
rect 5758 11033 5770 11036
rect 5712 11027 5770 11033
rect 6270 11024 6276 11036
rect 6328 11024 6334 11076
rect 7377 11067 7435 11073
rect 7377 11033 7389 11067
rect 7423 11064 7435 11067
rect 9490 11064 9496 11076
rect 7423 11036 9496 11064
rect 7423 11033 7435 11036
rect 7377 11027 7435 11033
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 11974 11024 11980 11076
rect 12032 11024 12038 11076
rect 2314 10956 2320 11008
rect 2372 10996 2378 11008
rect 2682 10996 2688 11008
rect 2372 10968 2688 10996
rect 2372 10956 2378 10968
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 4154 10956 4160 11008
rect 4212 10996 4218 11008
rect 4706 10996 4712 11008
rect 4212 10968 4712 10996
rect 4212 10956 4218 10968
rect 4706 10956 4712 10968
rect 4764 10956 4770 11008
rect 6825 10999 6883 11005
rect 6825 10965 6837 10999
rect 6871 10996 6883 10999
rect 7282 10996 7288 11008
rect 6871 10968 7288 10996
rect 6871 10965 6883 10968
rect 6825 10959 6883 10965
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 10045 10999 10103 11005
rect 10045 10965 10057 10999
rect 10091 10996 10103 10999
rect 10502 10996 10508 11008
rect 10091 10968 10508 10996
rect 10091 10965 10103 10968
rect 10045 10959 10103 10965
rect 10502 10956 10508 10968
rect 10560 10956 10566 11008
rect 11609 10999 11667 11005
rect 11609 10965 11621 10999
rect 11655 10996 11667 10999
rect 11698 10996 11704 11008
rect 11655 10968 11704 10996
rect 11655 10965 11667 10968
rect 11609 10959 11667 10965
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 12452 10996 12480 11095
rect 12526 11092 12532 11104
rect 12584 11092 12590 11144
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 12710 11092 12716 11144
rect 12768 11092 12774 11144
rect 12805 11135 12863 11141
rect 12805 11101 12817 11135
rect 12851 11101 12863 11135
rect 12805 11095 12863 11101
rect 12636 11064 12664 11092
rect 12820 11064 12848 11095
rect 12894 11092 12900 11144
rect 12952 11092 12958 11144
rect 12986 11092 12992 11144
rect 13044 11092 13050 11144
rect 13170 11092 13176 11144
rect 13228 11092 13234 11144
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13630 11132 13636 11144
rect 13403 11104 13636 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 13630 11092 13636 11104
rect 13688 11092 13694 11144
rect 13722 11092 13728 11144
rect 13780 11092 13786 11144
rect 14108 11141 14136 11240
rect 14734 11160 14740 11212
rect 14792 11200 14798 11212
rect 14829 11203 14887 11209
rect 14829 11200 14841 11203
rect 14792 11172 14841 11200
rect 14792 11160 14798 11172
rect 14829 11169 14841 11172
rect 14875 11169 14887 11203
rect 14829 11163 14887 11169
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11101 14151 11135
rect 14093 11095 14151 11101
rect 14182 11092 14188 11144
rect 14240 11132 14246 11144
rect 14277 11135 14335 11141
rect 14277 11132 14289 11135
rect 14240 11104 14289 11132
rect 14240 11092 14246 11104
rect 14277 11101 14289 11104
rect 14323 11101 14335 11135
rect 14277 11095 14335 11101
rect 14458 11092 14464 11144
rect 14516 11092 14522 11144
rect 15102 11141 15108 11144
rect 15096 11132 15108 11141
rect 15063 11104 15108 11132
rect 15096 11095 15108 11104
rect 15102 11092 15108 11095
rect 15160 11092 15166 11144
rect 16224 11132 16252 11299
rect 16298 11296 16304 11348
rect 16356 11296 16362 11348
rect 16485 11135 16543 11141
rect 16485 11132 16497 11135
rect 16224 11104 16497 11132
rect 16485 11101 16497 11104
rect 16531 11101 16543 11135
rect 16485 11095 16543 11101
rect 12636 11036 12848 11064
rect 13078 11024 13084 11076
rect 13136 11064 13142 11076
rect 14369 11067 14427 11073
rect 14369 11064 14381 11067
rect 13136 11036 14381 11064
rect 13136 11024 13142 11036
rect 14369 11033 14381 11036
rect 14415 11033 14427 11067
rect 14369 11027 14427 11033
rect 12308 10968 12480 10996
rect 12529 10999 12587 11005
rect 12308 10956 12314 10968
rect 12529 10965 12541 10999
rect 12575 10996 12587 10999
rect 12618 10996 12624 11008
rect 12575 10968 12624 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12618 10956 12624 10968
rect 12676 10956 12682 11008
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 13630 10996 13636 11008
rect 12768 10968 13636 10996
rect 12768 10956 12774 10968
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 1104 10906 16836 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 16836 10906
rect 1104 10832 16836 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 2038 10792 2044 10804
rect 1719 10764 2044 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 3697 10795 3755 10801
rect 2832 10764 3648 10792
rect 2832 10752 2838 10764
rect 2590 10724 2596 10736
rect 2056 10696 2596 10724
rect 2056 10665 2084 10696
rect 2590 10684 2596 10696
rect 2648 10684 2654 10736
rect 3620 10724 3648 10764
rect 3697 10761 3709 10795
rect 3743 10792 3755 10795
rect 5810 10792 5816 10804
rect 3743 10764 5816 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 5810 10752 5816 10764
rect 5868 10752 5874 10804
rect 6270 10752 6276 10804
rect 6328 10792 6334 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6328 10764 6377 10792
rect 6328 10752 6334 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 7834 10752 7840 10804
rect 7892 10792 7898 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 7892 10764 7941 10792
rect 7892 10752 7898 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 7929 10755 7987 10761
rect 12158 10752 12164 10804
rect 12216 10752 12222 10804
rect 12894 10792 12900 10804
rect 12360 10764 12480 10792
rect 3878 10724 3884 10736
rect 3620 10696 3884 10724
rect 3878 10684 3884 10696
rect 3936 10724 3942 10736
rect 4246 10724 4252 10736
rect 3936 10696 4252 10724
rect 3936 10684 3942 10696
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 1964 10520 1992 10619
rect 2130 10616 2136 10668
rect 2188 10616 2194 10668
rect 2222 10616 2228 10668
rect 2280 10656 2286 10668
rect 2317 10659 2375 10665
rect 2317 10656 2329 10659
rect 2280 10628 2329 10656
rect 2280 10616 2286 10628
rect 2317 10625 2329 10628
rect 2363 10625 2375 10659
rect 2317 10619 2375 10625
rect 2406 10616 2412 10668
rect 2464 10656 2470 10668
rect 2685 10659 2743 10665
rect 2464 10646 2544 10656
rect 2685 10646 2697 10659
rect 2464 10628 2697 10646
rect 2464 10616 2470 10628
rect 2516 10625 2697 10628
rect 2731 10625 2743 10659
rect 2516 10619 2743 10625
rect 2516 10618 2728 10619
rect 2771 10616 2777 10668
rect 2829 10616 2835 10668
rect 2890 10665 2948 10671
rect 2890 10631 2902 10665
rect 2936 10662 2948 10665
rect 2936 10634 3004 10662
rect 2936 10631 2948 10634
rect 2890 10625 2948 10631
rect 2976 10532 3004 10634
rect 3050 10616 3056 10668
rect 3108 10616 3114 10668
rect 3145 10659 3203 10665
rect 3145 10625 3157 10659
rect 3191 10625 3203 10659
rect 3145 10619 3203 10625
rect 3237 10659 3295 10665
rect 3237 10625 3249 10659
rect 3283 10656 3295 10659
rect 3326 10656 3332 10668
rect 3283 10628 3332 10656
rect 3283 10625 3295 10628
rect 3237 10619 3295 10625
rect 1964 10492 2544 10520
rect 2516 10464 2544 10492
rect 2958 10480 2964 10532
rect 3016 10480 3022 10532
rect 3160 10520 3188 10619
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 3418 10616 3424 10668
rect 3476 10616 3482 10668
rect 3510 10616 3516 10668
rect 3568 10616 3574 10668
rect 3694 10616 3700 10668
rect 3752 10656 3758 10668
rect 4080 10665 4108 10696
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 4433 10727 4491 10733
rect 4433 10693 4445 10727
rect 4479 10724 4491 10727
rect 4770 10727 4828 10733
rect 4770 10724 4782 10727
rect 4479 10696 4782 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 4770 10693 4782 10696
rect 4816 10693 4828 10727
rect 4770 10687 4828 10693
rect 5534 10684 5540 10736
rect 5592 10724 5598 10736
rect 5592 10696 8248 10724
rect 5592 10684 5598 10696
rect 3789 10659 3847 10665
rect 3789 10656 3801 10659
rect 3752 10628 3801 10656
rect 3752 10616 3758 10628
rect 3789 10625 3801 10628
rect 3835 10625 3847 10659
rect 3789 10619 3847 10625
rect 3973 10659 4031 10665
rect 3973 10625 3985 10659
rect 4019 10625 4031 10659
rect 3973 10619 4031 10625
rect 4065 10659 4123 10665
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4065 10619 4123 10625
rect 3418 10520 3424 10532
rect 3160 10492 3424 10520
rect 3418 10480 3424 10492
rect 3476 10480 3482 10532
rect 2406 10412 2412 10464
rect 2464 10412 2470 10464
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 3234 10452 3240 10464
rect 2556 10424 3240 10452
rect 2556 10412 2562 10424
rect 3234 10412 3240 10424
rect 3292 10412 3298 10464
rect 3988 10452 4016 10619
rect 4154 10616 4160 10668
rect 4212 10616 4218 10668
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 4614 10656 4620 10668
rect 4571 10628 4620 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4614 10616 4620 10628
rect 4672 10616 4678 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10656 6791 10659
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6779 10628 7205 10656
rect 6779 10625 6791 10628
rect 6733 10619 6791 10625
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7340 10628 7757 10656
rect 7340 10616 7346 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 8110 10616 8116 10668
rect 8168 10616 8174 10668
rect 8220 10665 8248 10696
rect 9490 10684 9496 10736
rect 9548 10724 9554 10736
rect 12360 10733 12388 10764
rect 12345 10727 12403 10733
rect 9548 10696 11560 10724
rect 9548 10684 9554 10696
rect 8205 10659 8263 10665
rect 8205 10625 8217 10659
rect 8251 10625 8263 10659
rect 8205 10619 8263 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 6822 10548 6828 10600
rect 6880 10548 6886 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10588 7067 10591
rect 8294 10588 8300 10600
rect 7055 10560 8300 10588
rect 7055 10557 7067 10560
rect 7009 10551 7067 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 8404 10588 8432 10619
rect 8478 10616 8484 10668
rect 8536 10616 8542 10668
rect 11532 10665 11560 10696
rect 12345 10693 12357 10727
rect 12391 10693 12403 10727
rect 12345 10687 12403 10693
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10656 9367 10659
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9355 10628 9781 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 11517 10659 11575 10665
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 12250 10616 12256 10668
rect 12308 10616 12314 10668
rect 12452 10656 12480 10764
rect 12544 10764 12900 10792
rect 12544 10733 12572 10764
rect 12894 10752 12900 10764
rect 12952 10752 12958 10804
rect 13998 10752 14004 10804
rect 14056 10752 14062 10804
rect 12529 10727 12587 10733
rect 12529 10693 12541 10727
rect 12575 10693 12587 10727
rect 12529 10687 12587 10693
rect 12621 10727 12679 10733
rect 12621 10693 12633 10727
rect 12667 10724 12679 10727
rect 12710 10724 12716 10736
rect 12667 10696 12716 10724
rect 12667 10693 12679 10696
rect 12621 10687 12679 10693
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 13262 10724 13268 10736
rect 12912 10696 13268 10724
rect 12802 10656 12808 10668
rect 12452 10628 12808 10656
rect 12802 10616 12808 10628
rect 12860 10616 12866 10668
rect 12912 10665 12940 10696
rect 13262 10684 13268 10696
rect 13320 10684 13326 10736
rect 13814 10724 13820 10736
rect 13464 10696 13820 10724
rect 12897 10659 12955 10665
rect 12897 10625 12909 10659
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 12986 10616 12992 10668
rect 13044 10656 13050 10668
rect 13173 10659 13231 10665
rect 13173 10656 13185 10659
rect 13044 10628 13185 10656
rect 13044 10616 13050 10628
rect 13173 10625 13185 10628
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 9122 10588 9128 10600
rect 8404 10560 9128 10588
rect 9122 10548 9128 10560
rect 9180 10548 9186 10600
rect 9398 10548 9404 10600
rect 9456 10548 9462 10600
rect 9582 10548 9588 10600
rect 9640 10548 9646 10600
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 10321 10591 10379 10597
rect 10321 10588 10333 10591
rect 10284 10560 10333 10588
rect 10284 10548 10290 10560
rect 10321 10557 10333 10560
rect 10367 10557 10379 10591
rect 10321 10551 10379 10557
rect 10502 10548 10508 10600
rect 10560 10588 10566 10600
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10560 10560 11161 10588
rect 10560 10548 10566 10560
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 11606 10548 11612 10600
rect 11664 10588 11670 10600
rect 11664 10560 12434 10588
rect 11664 10548 11670 10560
rect 11974 10480 11980 10532
rect 12032 10520 12038 10532
rect 12253 10523 12311 10529
rect 12253 10520 12265 10523
rect 12032 10492 12265 10520
rect 12032 10480 12038 10492
rect 12253 10489 12265 10492
rect 12299 10489 12311 10523
rect 12406 10520 12434 10560
rect 12618 10548 12624 10600
rect 12676 10548 12682 10600
rect 13265 10591 13323 10597
rect 13265 10557 13277 10591
rect 13311 10588 13323 10591
rect 13464 10588 13492 10696
rect 13814 10684 13820 10696
rect 13872 10724 13878 10736
rect 14366 10724 14372 10736
rect 13872 10696 14372 10724
rect 13872 10684 13878 10696
rect 14366 10684 14372 10696
rect 14424 10684 14430 10736
rect 13541 10659 13599 10665
rect 13541 10625 13553 10659
rect 13587 10625 13599 10659
rect 13541 10619 13599 10625
rect 13633 10659 13691 10665
rect 13633 10625 13645 10659
rect 13679 10656 13691 10659
rect 13722 10656 13728 10668
rect 13679 10628 13728 10656
rect 13679 10625 13691 10628
rect 13633 10619 13691 10625
rect 13311 10560 13492 10588
rect 13311 10557 13323 10560
rect 13265 10551 13323 10557
rect 13556 10520 13584 10619
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 13909 10659 13967 10665
rect 13909 10656 13921 10659
rect 13832 10628 13921 10656
rect 13832 10529 13860 10628
rect 13909 10625 13921 10628
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10656 14611 10659
rect 14642 10656 14648 10668
rect 14599 10628 14648 10656
rect 14599 10625 14611 10628
rect 14553 10619 14611 10625
rect 14642 10616 14648 10628
rect 14700 10616 14706 10668
rect 14826 10665 14832 10668
rect 14820 10619 14832 10665
rect 14826 10616 14832 10619
rect 14884 10616 14890 10668
rect 15194 10616 15200 10668
rect 15252 10656 15258 10668
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 15252 10628 16221 10656
rect 15252 10616 15258 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10588 14427 10591
rect 14458 10588 14464 10600
rect 14415 10560 14464 10588
rect 14415 10557 14427 10560
rect 14369 10551 14427 10557
rect 14458 10548 14464 10560
rect 14516 10548 14522 10600
rect 12406 10492 13584 10520
rect 13817 10523 13875 10529
rect 12253 10483 12311 10489
rect 13817 10489 13829 10523
rect 13863 10489 13875 10523
rect 13817 10483 13875 10489
rect 4706 10452 4712 10464
rect 3988 10424 4712 10452
rect 4706 10412 4712 10424
rect 4764 10412 4770 10464
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5500 10424 5917 10452
rect 5500 10412 5506 10424
rect 5905 10421 5917 10424
rect 5951 10421 5963 10455
rect 5905 10415 5963 10421
rect 8938 10412 8944 10464
rect 8996 10412 9002 10464
rect 10594 10412 10600 10464
rect 10652 10412 10658 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12492 10424 12817 10452
rect 12492 10412 12498 10424
rect 12805 10421 12817 10424
rect 12851 10452 12863 10455
rect 13538 10452 13544 10464
rect 12851 10424 13544 10452
rect 12851 10421 12863 10424
rect 12805 10415 12863 10421
rect 13538 10412 13544 10424
rect 13596 10412 13602 10464
rect 14185 10455 14243 10461
rect 14185 10421 14197 10455
rect 14231 10452 14243 10455
rect 15470 10452 15476 10464
rect 14231 10424 15476 10452
rect 14231 10421 14243 10424
rect 14185 10415 14243 10421
rect 15470 10412 15476 10424
rect 15528 10412 15534 10464
rect 15930 10412 15936 10464
rect 15988 10412 15994 10464
rect 16390 10412 16396 10464
rect 16448 10412 16454 10464
rect 1104 10362 16836 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 16836 10362
rect 1104 10288 16836 10310
rect 1765 10251 1823 10257
rect 1765 10217 1777 10251
rect 1811 10248 1823 10251
rect 2958 10248 2964 10260
rect 1811 10220 2964 10248
rect 1811 10217 1823 10220
rect 1765 10211 1823 10217
rect 2958 10208 2964 10220
rect 3016 10208 3022 10260
rect 5353 10251 5411 10257
rect 4816 10220 5304 10248
rect 1762 10072 1768 10124
rect 1820 10112 1826 10124
rect 1857 10115 1915 10121
rect 1857 10112 1869 10115
rect 1820 10084 1869 10112
rect 1820 10072 1826 10084
rect 1857 10081 1869 10084
rect 1903 10081 1915 10115
rect 1857 10075 1915 10081
rect 1872 10044 1900 10075
rect 1872 10016 2774 10044
rect 1394 9936 1400 9988
rect 1452 9936 1458 9988
rect 1581 9979 1639 9985
rect 1581 9945 1593 9979
rect 1627 9945 1639 9979
rect 1581 9939 1639 9945
rect 2124 9979 2182 9985
rect 2124 9945 2136 9979
rect 2170 9976 2182 9979
rect 2406 9976 2412 9988
rect 2170 9948 2412 9976
rect 2170 9945 2182 9948
rect 2124 9939 2182 9945
rect 1596 9908 1624 9939
rect 2406 9936 2412 9948
rect 2464 9936 2470 9988
rect 2746 9976 2774 10016
rect 3510 10004 3516 10056
rect 3568 10044 3574 10056
rect 4816 10053 4844 10220
rect 5276 10112 5304 10220
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 6822 10248 6828 10260
rect 5399 10220 6828 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 8205 10251 8263 10257
rect 8205 10217 8217 10251
rect 8251 10248 8263 10251
rect 9398 10248 9404 10260
rect 8251 10220 9404 10248
rect 8251 10217 8263 10220
rect 8205 10211 8263 10217
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 9490 10208 9496 10260
rect 9548 10248 9554 10260
rect 9548 10220 10088 10248
rect 9548 10208 9554 10220
rect 10060 10180 10088 10220
rect 10502 10208 10508 10260
rect 10560 10208 10566 10260
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 11388 10220 12081 10248
rect 11388 10208 11394 10220
rect 12069 10217 12081 10220
rect 12115 10248 12127 10251
rect 12115 10220 14780 10248
rect 12115 10217 12127 10220
rect 12069 10211 12127 10217
rect 10597 10183 10655 10189
rect 10597 10180 10609 10183
rect 10060 10152 10609 10180
rect 10597 10149 10609 10152
rect 10643 10149 10655 10183
rect 10597 10143 10655 10149
rect 13630 10140 13636 10192
rect 13688 10140 13694 10192
rect 14642 10140 14648 10192
rect 14700 10140 14706 10192
rect 13449 10115 13507 10121
rect 5000 10084 5212 10112
rect 5276 10084 9260 10112
rect 4801 10047 4859 10053
rect 3568 10016 4752 10044
rect 3568 10004 3574 10016
rect 3789 9979 3847 9985
rect 3789 9976 3801 9979
rect 2746 9948 3801 9976
rect 3789 9945 3801 9948
rect 3835 9976 3847 9979
rect 4154 9976 4160 9988
rect 3835 9948 4160 9976
rect 3835 9945 3847 9948
rect 3789 9939 3847 9945
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 4724 9976 4752 10016
rect 4801 10013 4813 10047
rect 4847 10013 4859 10047
rect 4801 10007 4859 10013
rect 4890 10004 4896 10056
rect 4948 10004 4954 10056
rect 5000 9976 5028 10084
rect 5184 10053 5212 10084
rect 5077 10047 5135 10053
rect 5077 10013 5089 10047
rect 5123 10013 5135 10047
rect 5077 10007 5135 10013
rect 5169 10047 5227 10053
rect 5169 10013 5181 10047
rect 5215 10044 5227 10047
rect 8110 10044 8116 10056
rect 5215 10016 8116 10044
rect 5215 10013 5227 10016
rect 5169 10007 5227 10013
rect 4724 9948 5028 9976
rect 1670 9908 1676 9920
rect 1596 9880 1676 9908
rect 1670 9868 1676 9880
rect 1728 9908 1734 9920
rect 3237 9911 3295 9917
rect 3237 9908 3249 9911
rect 1728 9880 3249 9908
rect 1728 9868 1734 9880
rect 3237 9877 3249 9880
rect 3283 9908 3295 9911
rect 5092 9908 5120 10007
rect 8110 10004 8116 10016
rect 8168 10044 8174 10056
rect 8386 10044 8392 10056
rect 8168 10016 8392 10044
rect 8168 10004 8174 10016
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8481 10047 8539 10053
rect 8481 10013 8493 10047
rect 8527 10013 8539 10047
rect 8481 10007 8539 10013
rect 8665 10047 8723 10053
rect 8665 10013 8677 10047
rect 8711 10013 8723 10047
rect 8665 10007 8723 10013
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 8496 9976 8524 10007
rect 5408 9948 8524 9976
rect 5408 9936 5414 9948
rect 3283 9880 5120 9908
rect 8680 9908 8708 10007
rect 8754 10004 8760 10056
rect 8812 10004 8818 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9232 10044 9260 10084
rect 13449 10081 13461 10115
rect 13495 10112 13507 10115
rect 14660 10112 14688 10140
rect 14752 10121 14780 10220
rect 14826 10208 14832 10260
rect 14884 10248 14890 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14884 10220 14933 10248
rect 14884 10208 14890 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 14921 10211 14979 10217
rect 13495 10084 14688 10112
rect 14737 10115 14795 10121
rect 13495 10081 13507 10084
rect 13449 10075 13507 10081
rect 14737 10081 14749 10115
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 10686 10044 10692 10056
rect 9232 10016 10692 10044
rect 9125 10007 9183 10013
rect 9140 9976 9168 10007
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 11698 10004 11704 10056
rect 11756 10053 11762 10056
rect 11756 10044 11768 10053
rect 11977 10047 12035 10053
rect 11756 10016 11801 10044
rect 11756 10007 11768 10016
rect 11977 10013 11989 10047
rect 12023 10044 12035 10047
rect 13464 10044 13492 10075
rect 15378 10072 15384 10124
rect 15436 10072 15442 10124
rect 15470 10072 15476 10124
rect 15528 10072 15534 10124
rect 15930 10072 15936 10124
rect 15988 10112 15994 10124
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 15988 10084 16313 10112
rect 15988 10072 15994 10084
rect 16301 10081 16313 10084
rect 16347 10112 16359 10115
rect 16482 10112 16488 10124
rect 16347 10084 16488 10112
rect 16347 10081 16359 10084
rect 16301 10075 16359 10081
rect 16482 10072 16488 10084
rect 16540 10072 16546 10124
rect 12023 10016 13492 10044
rect 12023 10013 12035 10016
rect 11977 10007 12035 10013
rect 11756 10004 11762 10007
rect 13538 10004 13544 10056
rect 13596 10004 13602 10056
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10044 13783 10047
rect 13814 10044 13820 10056
rect 13771 10016 13820 10044
rect 13771 10013 13783 10016
rect 13725 10007 13783 10013
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 9214 9976 9220 9988
rect 9140 9948 9220 9976
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9392 9979 9450 9985
rect 9392 9945 9404 9979
rect 9438 9976 9450 9979
rect 10134 9976 10140 9988
rect 9438 9948 10140 9976
rect 9438 9945 9450 9948
rect 9392 9939 9450 9945
rect 10134 9936 10140 9948
rect 10192 9936 10198 9988
rect 12710 9936 12716 9988
rect 12768 9976 12774 9988
rect 13182 9979 13240 9985
rect 13182 9976 13194 9979
rect 12768 9948 13194 9976
rect 12768 9936 12774 9948
rect 13182 9945 13194 9948
rect 13228 9945 13240 9979
rect 13182 9939 13240 9945
rect 10870 9908 10876 9920
rect 8680 9880 10876 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 10870 9868 10876 9880
rect 10928 9868 10934 9920
rect 14090 9868 14096 9920
rect 14148 9868 14154 9920
rect 15289 9911 15347 9917
rect 15289 9877 15301 9911
rect 15335 9908 15347 9911
rect 15749 9911 15807 9917
rect 15749 9908 15761 9911
rect 15335 9880 15761 9908
rect 15335 9877 15347 9880
rect 15289 9871 15347 9877
rect 15749 9877 15761 9880
rect 15795 9877 15807 9911
rect 15749 9871 15807 9877
rect 1104 9818 16836 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 16836 9818
rect 1104 9744 16836 9766
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 5074 9704 5080 9716
rect 4120 9676 5080 9704
rect 4120 9664 4126 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 5166 9664 5172 9716
rect 5224 9704 5230 9716
rect 5626 9704 5632 9716
rect 5224 9676 5632 9704
rect 5224 9664 5230 9676
rect 5626 9664 5632 9676
rect 5684 9664 5690 9716
rect 10134 9664 10140 9716
rect 10192 9664 10198 9716
rect 10505 9707 10563 9713
rect 10505 9673 10517 9707
rect 10551 9704 10563 9707
rect 10594 9704 10600 9716
rect 10551 9676 10600 9704
rect 10551 9673 10563 9676
rect 10505 9667 10563 9673
rect 10594 9664 10600 9676
rect 10652 9664 10658 9716
rect 10686 9664 10692 9716
rect 10744 9704 10750 9716
rect 13998 9704 14004 9716
rect 10744 9676 14004 9704
rect 10744 9664 10750 9676
rect 13998 9664 14004 9676
rect 14056 9664 14062 9716
rect 3329 9639 3387 9645
rect 3329 9605 3341 9639
rect 3375 9636 3387 9639
rect 3786 9636 3792 9648
rect 3375 9608 3792 9636
rect 3375 9605 3387 9608
rect 3329 9599 3387 9605
rect 3786 9596 3792 9608
rect 3844 9596 3850 9648
rect 4709 9639 4767 9645
rect 4709 9605 4721 9639
rect 4755 9636 4767 9639
rect 6362 9636 6368 9648
rect 4755 9608 6368 9636
rect 4755 9605 4767 9608
rect 4709 9599 4767 9605
rect 6362 9596 6368 9608
rect 6420 9596 6426 9648
rect 8938 9645 8944 9648
rect 8932 9636 8944 9645
rect 8899 9608 8944 9636
rect 8932 9599 8944 9608
rect 8938 9596 8944 9599
rect 8996 9596 9002 9648
rect 13906 9596 13912 9648
rect 13964 9636 13970 9648
rect 14185 9639 14243 9645
rect 14185 9636 14197 9639
rect 13964 9608 14197 9636
rect 13964 9596 13970 9608
rect 14185 9605 14197 9608
rect 14231 9605 14243 9639
rect 14185 9599 14243 9605
rect 1670 9528 1676 9580
rect 1728 9528 1734 9580
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2498 9568 2504 9580
rect 2087 9540 2504 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3804 9568 3832 9596
rect 4801 9571 4859 9577
rect 4801 9568 4813 9571
rect 3804 9540 4813 9568
rect 3513 9531 3571 9537
rect 4801 9537 4813 9540
rect 4847 9537 4859 9571
rect 4801 9531 4859 9537
rect 4985 9571 5043 9577
rect 4985 9537 4997 9571
rect 5031 9568 5043 9571
rect 5350 9568 5356 9580
rect 5031 9540 5356 9568
rect 5031 9537 5043 9540
rect 4985 9531 5043 9537
rect 1026 9392 1032 9444
rect 1084 9432 1090 9444
rect 1857 9435 1915 9441
rect 1857 9432 1869 9435
rect 1084 9404 1869 9432
rect 1084 9392 1090 9404
rect 1857 9401 1869 9404
rect 1903 9401 1915 9435
rect 3528 9432 3556 9531
rect 5350 9528 5356 9540
rect 5408 9528 5414 9580
rect 6089 9571 6147 9577
rect 6089 9537 6101 9571
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9500 4031 9503
rect 4154 9500 4160 9512
rect 4019 9472 4160 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 4154 9460 4160 9472
rect 4212 9500 4218 9512
rect 4614 9500 4620 9512
rect 4212 9472 4620 9500
rect 4212 9460 4218 9472
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 5169 9503 5227 9509
rect 5169 9500 5181 9503
rect 4764 9472 5181 9500
rect 4764 9460 4770 9472
rect 5169 9469 5181 9472
rect 5215 9469 5227 9503
rect 6104 9500 6132 9531
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 6914 9528 6920 9580
rect 6972 9528 6978 9580
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9568 7067 9571
rect 7282 9568 7288 9580
rect 7055 9540 7288 9568
rect 7055 9537 7067 9540
rect 7009 9531 7067 9537
rect 7282 9528 7288 9540
rect 7340 9528 7346 9580
rect 7466 9577 7472 9580
rect 7460 9531 7472 9577
rect 7466 9528 7472 9531
rect 7524 9528 7530 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 9214 9568 9220 9580
rect 8711 9540 9220 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 9214 9528 9220 9540
rect 9272 9528 9278 9580
rect 14090 9528 14096 9580
rect 14148 9528 14154 9580
rect 16482 9528 16488 9580
rect 16540 9528 16546 9580
rect 7193 9503 7251 9509
rect 6104 9472 6960 9500
rect 5169 9463 5227 9469
rect 6932 9444 6960 9472
rect 7193 9469 7205 9503
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 6730 9432 6736 9444
rect 1857 9395 1915 9401
rect 2746 9404 6736 9432
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 1489 9367 1547 9373
rect 1489 9364 1501 9367
rect 1360 9336 1501 9364
rect 1360 9324 1366 9336
rect 1489 9333 1501 9336
rect 1535 9333 1547 9367
rect 1489 9327 1547 9333
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 2746 9364 2774 9404
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 6914 9392 6920 9444
rect 6972 9432 6978 9444
rect 7208 9432 7236 9463
rect 10594 9460 10600 9512
rect 10652 9460 10658 9512
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9469 10747 9503
rect 10689 9463 10747 9469
rect 6972 9404 7236 9432
rect 6972 9392 6978 9404
rect 8570 9392 8576 9444
rect 8628 9392 8634 9444
rect 10045 9435 10103 9441
rect 10045 9401 10057 9435
rect 10091 9432 10103 9435
rect 10226 9432 10232 9444
rect 10091 9404 10232 9432
rect 10091 9401 10103 9404
rect 10045 9395 10103 9401
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 1728 9336 2774 9364
rect 3697 9367 3755 9373
rect 1728 9324 1734 9336
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 4062 9364 4068 9376
rect 3743 9336 4068 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 4062 9324 4068 9336
rect 4120 9324 4126 9376
rect 6457 9367 6515 9373
rect 6457 9333 6469 9367
rect 6503 9364 6515 9367
rect 7926 9364 7932 9376
rect 6503 9336 7932 9364
rect 6503 9333 6515 9336
rect 6457 9327 6515 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 9582 9364 9588 9376
rect 8352 9336 9588 9364
rect 8352 9324 8358 9336
rect 9582 9324 9588 9336
rect 9640 9364 9646 9376
rect 10704 9364 10732 9463
rect 16206 9392 16212 9444
rect 16264 9432 16270 9444
rect 16301 9435 16359 9441
rect 16301 9432 16313 9435
rect 16264 9404 16313 9432
rect 16264 9392 16270 9404
rect 16301 9401 16313 9404
rect 16347 9401 16359 9435
rect 16301 9395 16359 9401
rect 9640 9336 10732 9364
rect 9640 9324 9646 9336
rect 1104 9274 16836 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 16836 9274
rect 1104 9200 16836 9222
rect 4430 9120 4436 9172
rect 4488 9160 4494 9172
rect 5902 9160 5908 9172
rect 4488 9132 5908 9160
rect 4488 9120 4494 9132
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 5997 9163 6055 9169
rect 5997 9129 6009 9163
rect 6043 9160 6055 9163
rect 6730 9160 6736 9172
rect 6043 9132 6736 9160
rect 6043 9129 6055 9132
rect 5997 9123 6055 9129
rect 6730 9120 6736 9132
rect 6788 9120 6794 9172
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 7524 9132 7573 9160
rect 7524 9120 7530 9132
rect 7561 9129 7573 9132
rect 7607 9129 7619 9163
rect 7561 9123 7619 9129
rect 9030 9120 9036 9172
rect 9088 9160 9094 9172
rect 9861 9163 9919 9169
rect 9861 9160 9873 9163
rect 9088 9132 9873 9160
rect 9088 9120 9094 9132
rect 9861 9129 9873 9132
rect 9907 9129 9919 9163
rect 9861 9123 9919 9129
rect 10870 9120 10876 9172
rect 10928 9120 10934 9172
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 12802 9160 12808 9172
rect 11112 9132 12808 9160
rect 11112 9120 11118 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 842 9052 848 9104
rect 900 9092 906 9104
rect 1489 9095 1547 9101
rect 1489 9092 1501 9095
rect 900 9064 1501 9092
rect 900 9052 906 9064
rect 1489 9061 1501 9064
rect 1535 9061 1547 9095
rect 2774 9092 2780 9104
rect 1489 9055 1547 9061
rect 1964 9064 2780 9092
rect 1670 8916 1676 8968
rect 1728 8916 1734 8968
rect 1964 8965 1992 9064
rect 2774 9052 2780 9064
rect 2832 9092 2838 9104
rect 3510 9092 3516 9104
rect 2832 9064 3516 9092
rect 2832 9052 2838 9064
rect 3510 9052 3516 9064
rect 3568 9052 3574 9104
rect 7282 9052 7288 9104
rect 7340 9092 7346 9104
rect 12989 9095 13047 9101
rect 12989 9092 13001 9095
rect 7340 9064 13001 9092
rect 7340 9052 7346 9064
rect 12989 9061 13001 9064
rect 13035 9061 13047 9095
rect 12989 9055 13047 9061
rect 2590 9024 2596 9036
rect 2240 8996 2596 9024
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 2240 8965 2268 8996
rect 2590 8984 2596 8996
rect 2648 9024 2654 9036
rect 4338 9024 4344 9036
rect 2648 8996 4344 9024
rect 2648 8984 2654 8996
rect 2133 8959 2191 8965
rect 2133 8956 2145 8959
rect 2096 8928 2145 8956
rect 2096 8916 2102 8928
rect 2133 8925 2145 8928
rect 2179 8925 2191 8959
rect 2133 8919 2191 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8925 2283 8959
rect 2225 8919 2283 8925
rect 2314 8916 2320 8968
rect 2372 8916 2378 8968
rect 2958 8916 2964 8968
rect 3016 8916 3022 8968
rect 3694 8916 3700 8968
rect 3752 8956 3758 8968
rect 3881 8959 3939 8965
rect 3881 8956 3893 8959
rect 3752 8928 3893 8956
rect 3752 8916 3758 8928
rect 3881 8925 3893 8928
rect 3927 8925 3939 8959
rect 3881 8919 3939 8925
rect 2590 8780 2596 8832
rect 2648 8780 2654 8832
rect 2774 8780 2780 8832
rect 2832 8780 2838 8832
rect 3896 8820 3924 8919
rect 4062 8916 4068 8968
rect 4120 8916 4126 8968
rect 4172 8965 4200 8996
rect 4338 8984 4344 8996
rect 4396 8984 4402 9036
rect 4614 8984 4620 9036
rect 4672 8984 4678 9036
rect 7926 8984 7932 9036
rect 7984 9024 7990 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 7984 8996 8033 9024
rect 7984 8984 7990 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8205 9027 8263 9033
rect 8205 8993 8217 9027
rect 8251 9024 8263 9027
rect 8294 9024 8300 9036
rect 8251 8996 8300 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 8294 8984 8300 8996
rect 8352 8984 8358 9036
rect 8570 8984 8576 9036
rect 8628 9024 8634 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8628 8996 9505 9024
rect 8628 8984 8634 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9493 8987 9551 8993
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 13262 9024 13268 9036
rect 9640 8996 10088 9024
rect 9640 8984 9646 8996
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8925 4215 8959
rect 4157 8919 4215 8925
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4706 8956 4712 8968
rect 4295 8928 4712 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4706 8916 4712 8928
rect 4764 8956 4770 8968
rect 5442 8956 5448 8968
rect 4764 8928 5448 8956
rect 4764 8916 4770 8928
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6089 8959 6147 8965
rect 6089 8925 6101 8959
rect 6135 8956 6147 8959
rect 6914 8956 6920 8968
rect 6135 8928 6920 8956
rect 6135 8925 6147 8928
rect 6089 8919 6147 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 7024 8928 9996 8956
rect 4525 8891 4583 8897
rect 4525 8857 4537 8891
rect 4571 8888 4583 8891
rect 4862 8891 4920 8897
rect 4862 8888 4874 8891
rect 4571 8860 4874 8888
rect 4571 8857 4583 8860
rect 4525 8851 4583 8857
rect 4862 8857 4874 8860
rect 4908 8857 4920 8891
rect 4862 8851 4920 8857
rect 5074 8848 5080 8900
rect 5132 8888 5138 8900
rect 5350 8888 5356 8900
rect 5132 8860 5356 8888
rect 5132 8848 5138 8860
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 6356 8891 6414 8897
rect 6356 8857 6368 8891
rect 6402 8888 6414 8891
rect 6454 8888 6460 8900
rect 6402 8860 6460 8888
rect 6402 8857 6414 8860
rect 6356 8851 6414 8857
rect 6454 8848 6460 8860
rect 6512 8848 6518 8900
rect 7024 8888 7052 8928
rect 6564 8860 7052 8888
rect 7929 8891 7987 8897
rect 6564 8820 6592 8860
rect 7929 8857 7941 8891
rect 7975 8888 7987 8891
rect 8941 8891 8999 8897
rect 8941 8888 8953 8891
rect 7975 8860 8953 8888
rect 7975 8857 7987 8860
rect 7929 8851 7987 8857
rect 8941 8857 8953 8860
rect 8987 8857 8999 8891
rect 8941 8851 8999 8857
rect 9674 8848 9680 8900
rect 9732 8848 9738 8900
rect 3896 8792 6592 8820
rect 6638 8780 6644 8832
rect 6696 8820 6702 8832
rect 7466 8820 7472 8832
rect 6696 8792 7472 8820
rect 6696 8780 6702 8792
rect 7466 8780 7472 8792
rect 7524 8780 7530 8832
rect 9858 8780 9864 8832
rect 9916 8780 9922 8832
rect 9968 8820 9996 8928
rect 10060 8888 10088 8996
rect 11164 8996 13268 9024
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 11054 8956 11060 8968
rect 10183 8928 11060 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 11054 8916 11060 8928
rect 11112 8916 11118 8968
rect 11164 8965 11192 8996
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 11149 8959 11207 8965
rect 11149 8925 11161 8959
rect 11195 8925 11207 8959
rect 11149 8919 11207 8925
rect 11422 8916 11428 8968
rect 11480 8916 11486 8968
rect 11517 8959 11575 8965
rect 11517 8925 11529 8959
rect 11563 8956 11575 8959
rect 11793 8959 11851 8965
rect 11563 8928 11652 8956
rect 11563 8925 11575 8928
rect 11517 8919 11575 8925
rect 10321 8891 10379 8897
rect 10321 8888 10333 8891
rect 10060 8860 10333 8888
rect 10321 8857 10333 8860
rect 10367 8857 10379 8891
rect 10321 8851 10379 8857
rect 10505 8891 10563 8897
rect 10505 8857 10517 8891
rect 10551 8888 10563 8891
rect 10962 8888 10968 8900
rect 10551 8860 10968 8888
rect 10551 8857 10563 8860
rect 10505 8851 10563 8857
rect 10962 8848 10968 8860
rect 11020 8888 11026 8900
rect 11241 8891 11299 8897
rect 11241 8888 11253 8891
rect 11020 8860 11253 8888
rect 11020 8848 11026 8860
rect 11241 8857 11253 8860
rect 11287 8857 11299 8891
rect 11241 8851 11299 8857
rect 11624 8820 11652 8928
rect 11793 8925 11805 8959
rect 11839 8956 11851 8959
rect 12158 8956 12164 8968
rect 11839 8928 12164 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 12437 8959 12495 8965
rect 12437 8925 12449 8959
rect 12483 8956 12495 8959
rect 12526 8956 12532 8968
rect 12483 8928 12532 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 12526 8916 12532 8928
rect 12584 8916 12590 8968
rect 12802 8916 12808 8968
rect 12860 8916 12866 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13096 8928 14105 8956
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 12621 8891 12679 8897
rect 12621 8888 12633 8891
rect 11756 8860 12633 8888
rect 11756 8848 11762 8860
rect 12621 8857 12633 8860
rect 12667 8857 12679 8891
rect 12621 8851 12679 8857
rect 12713 8891 12771 8897
rect 12713 8857 12725 8891
rect 12759 8888 12771 8891
rect 12894 8888 12900 8900
rect 12759 8860 12900 8888
rect 12759 8857 12771 8860
rect 12713 8851 12771 8857
rect 12894 8848 12900 8860
rect 12952 8848 12958 8900
rect 13096 8888 13124 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 13004 8860 13124 8888
rect 9968 8792 11652 8820
rect 12158 8780 12164 8832
rect 12216 8820 12222 8832
rect 13004 8820 13032 8860
rect 13262 8848 13268 8900
rect 13320 8848 13326 8900
rect 13446 8848 13452 8900
rect 13504 8848 13510 8900
rect 14108 8888 14136 8919
rect 14274 8916 14280 8968
rect 14332 8916 14338 8968
rect 14366 8916 14372 8968
rect 14424 8916 14430 8968
rect 14458 8916 14464 8968
rect 14516 8916 14522 8968
rect 15378 8888 15384 8900
rect 14108 8860 15384 8888
rect 15378 8848 15384 8860
rect 15436 8848 15442 8900
rect 12216 8792 13032 8820
rect 12216 8780 12222 8792
rect 13078 8780 13084 8832
rect 13136 8780 13142 8832
rect 14734 8780 14740 8832
rect 14792 8780 14798 8832
rect 1104 8730 16836 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 16836 8730
rect 1104 8656 16836 8678
rect 2038 8576 2044 8628
rect 2096 8576 2102 8628
rect 3142 8616 3148 8628
rect 2332 8588 3148 8616
rect 1394 8508 1400 8560
rect 1452 8548 1458 8560
rect 1673 8551 1731 8557
rect 1673 8548 1685 8551
rect 1452 8520 1685 8548
rect 1452 8508 1458 8520
rect 1673 8517 1685 8520
rect 1719 8517 1731 8551
rect 1673 8511 1731 8517
rect 1857 8551 1915 8557
rect 1857 8517 1869 8551
rect 1903 8548 1915 8551
rect 2332 8548 2360 8588
rect 3142 8576 3148 8588
rect 3200 8616 3206 8628
rect 3513 8619 3571 8625
rect 3513 8616 3525 8619
rect 3200 8588 3525 8616
rect 3200 8576 3206 8588
rect 3513 8585 3525 8588
rect 3559 8585 3571 8619
rect 6178 8616 6184 8628
rect 3513 8579 3571 8585
rect 3896 8588 6184 8616
rect 1903 8520 2360 8548
rect 2400 8551 2458 8557
rect 1903 8517 1915 8520
rect 1857 8511 1915 8517
rect 2400 8517 2412 8551
rect 2446 8548 2458 8551
rect 2590 8548 2596 8560
rect 2446 8520 2596 8548
rect 2446 8517 2458 8520
rect 2400 8511 2458 8517
rect 1688 8480 1716 8511
rect 2590 8508 2596 8520
rect 2648 8508 2654 8560
rect 2958 8508 2964 8560
rect 3016 8548 3022 8560
rect 3797 8551 3855 8557
rect 3797 8548 3809 8551
rect 3016 8520 3809 8548
rect 3016 8508 3022 8520
rect 3797 8517 3809 8520
rect 3843 8548 3855 8551
rect 3896 8548 3924 8588
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 13320 8588 14657 8616
rect 13320 8576 13326 8588
rect 14645 8585 14657 8588
rect 14691 8616 14703 8619
rect 15194 8616 15200 8628
rect 14691 8588 15200 8616
rect 14691 8585 14703 8588
rect 14645 8579 14703 8585
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 3843 8520 3924 8548
rect 3973 8551 4031 8557
rect 3843 8517 3855 8520
rect 3797 8511 3855 8517
rect 3973 8517 3985 8551
rect 4019 8548 4031 8551
rect 4019 8520 4292 8548
rect 4019 8517 4031 8520
rect 3973 8511 4031 8517
rect 3605 8483 3663 8489
rect 3605 8480 3617 8483
rect 1688 8452 3617 8480
rect 3605 8449 3617 8452
rect 3651 8480 3663 8483
rect 3878 8480 3884 8492
rect 3651 8452 3884 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4264 8489 4292 8520
rect 4816 8520 5212 8548
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 1762 8372 1768 8424
rect 1820 8412 1826 8424
rect 2133 8415 2191 8421
rect 2133 8412 2145 8415
rect 1820 8384 2145 8412
rect 1820 8372 1826 8384
rect 2133 8381 2145 8384
rect 2179 8381 2191 8415
rect 2133 8375 2191 8381
rect 3510 8372 3516 8424
rect 3568 8412 3574 8424
rect 3786 8412 3792 8424
rect 3568 8384 3792 8412
rect 3568 8372 3574 8384
rect 3786 8372 3792 8384
rect 3844 8412 3850 8424
rect 4080 8412 4108 8443
rect 4338 8440 4344 8492
rect 4396 8440 4402 8492
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4816 8489 4844 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 5057 8483 5115 8489
rect 5057 8480 5069 8483
rect 4801 8443 4859 8449
rect 4908 8452 5069 8480
rect 3844 8384 4108 8412
rect 4356 8412 4384 8440
rect 4614 8412 4620 8424
rect 4356 8384 4620 8412
rect 3844 8372 3850 8384
rect 4614 8372 4620 8384
rect 4672 8372 4678 8424
rect 4709 8415 4767 8421
rect 4709 8381 4721 8415
rect 4755 8412 4767 8415
rect 4908 8412 4936 8452
rect 5057 8449 5069 8452
rect 5103 8449 5115 8483
rect 5184 8480 5212 8520
rect 6362 8508 6368 8560
rect 6420 8508 6426 8560
rect 6730 8508 6736 8560
rect 6788 8548 6794 8560
rect 7377 8551 7435 8557
rect 7377 8548 7389 8551
rect 6788 8520 7389 8548
rect 6788 8508 6794 8520
rect 7377 8517 7389 8520
rect 7423 8517 7435 8551
rect 9309 8551 9367 8557
rect 9309 8548 9321 8551
rect 7377 8511 7435 8517
rect 8312 8520 9321 8548
rect 6914 8480 6920 8492
rect 5184 8452 6920 8480
rect 5057 8443 5115 8449
rect 6914 8440 6920 8452
rect 6972 8480 6978 8492
rect 6972 8452 7144 8480
rect 6972 8440 6978 8452
rect 7116 8421 7144 8452
rect 7466 8440 7472 8492
rect 7524 8480 7530 8492
rect 7929 8483 7987 8489
rect 7929 8480 7941 8483
rect 7524 8452 7941 8480
rect 7524 8440 7530 8452
rect 7929 8449 7941 8452
rect 7975 8480 7987 8483
rect 8205 8483 8263 8489
rect 8205 8480 8217 8483
rect 7975 8452 8217 8480
rect 7975 8449 7987 8452
rect 7929 8443 7987 8449
rect 8205 8449 8217 8452
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 4755 8384 4936 8412
rect 7101 8415 7159 8421
rect 4755 8381 4767 8384
rect 4709 8375 4767 8381
rect 7101 8381 7113 8415
rect 7147 8412 7159 8415
rect 7374 8412 7380 8424
rect 7147 8384 7380 8412
rect 7147 8381 7159 8384
rect 7101 8375 7159 8381
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 6178 8304 6184 8356
rect 6236 8304 6242 8356
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 8312 8276 8340 8520
rect 9309 8517 9321 8520
rect 9355 8548 9367 8551
rect 9582 8548 9588 8560
rect 9355 8520 9588 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 11882 8508 11888 8560
rect 11940 8548 11946 8560
rect 13081 8551 13139 8557
rect 11940 8520 12296 8548
rect 11940 8508 11946 8520
rect 12268 8492 12296 8520
rect 13081 8517 13093 8551
rect 13127 8548 13139 8551
rect 14090 8548 14096 8560
rect 13127 8520 14096 8548
rect 13127 8517 13139 8520
rect 13081 8511 13139 8517
rect 8386 8440 8392 8492
rect 8444 8480 8450 8492
rect 8573 8483 8631 8489
rect 8573 8480 8585 8483
rect 8444 8452 8585 8480
rect 8444 8440 8450 8452
rect 8573 8449 8585 8452
rect 8619 8480 8631 8483
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8619 8452 8769 8480
rect 8619 8449 8631 8452
rect 8573 8443 8631 8449
rect 8757 8449 8769 8452
rect 8803 8480 8815 8483
rect 8846 8480 8852 8492
rect 8803 8452 8852 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 9766 8480 9772 8492
rect 9272 8452 9772 8480
rect 9272 8440 9278 8452
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 10962 8480 10968 8492
rect 10919 8452 10968 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 10962 8440 10968 8452
rect 11020 8480 11026 8492
rect 11698 8480 11704 8492
rect 11020 8452 11704 8480
rect 11020 8440 11026 8452
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 12161 8483 12219 8489
rect 12161 8449 12173 8483
rect 12207 8449 12219 8483
rect 12161 8443 12219 8449
rect 9125 8415 9183 8421
rect 9125 8381 9137 8415
rect 9171 8381 9183 8415
rect 9125 8375 9183 8381
rect 9140 8344 9168 8375
rect 10502 8372 10508 8424
rect 10560 8372 10566 8424
rect 11882 8372 11888 8424
rect 11940 8412 11946 8424
rect 12176 8412 12204 8443
rect 12250 8440 12256 8492
rect 12308 8440 12314 8492
rect 13096 8412 13124 8511
rect 14090 8508 14096 8520
rect 14148 8508 14154 8560
rect 13170 8440 13176 8492
rect 13228 8480 13234 8492
rect 13521 8483 13579 8489
rect 13521 8480 13533 8483
rect 13228 8452 13533 8480
rect 13228 8440 13234 8452
rect 13521 8449 13533 8452
rect 13567 8449 13579 8483
rect 13521 8443 13579 8449
rect 16206 8440 16212 8492
rect 16264 8440 16270 8492
rect 13265 8415 13323 8421
rect 13265 8412 13277 8415
rect 11940 8384 13277 8412
rect 11940 8372 11946 8384
rect 13265 8381 13277 8384
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 9858 8344 9864 8356
rect 9140 8316 9864 8344
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 16393 8347 16451 8353
rect 16393 8313 16405 8347
rect 16439 8344 16451 8347
rect 16574 8344 16580 8356
rect 16439 8316 16580 8344
rect 16439 8313 16451 8316
rect 16393 8307 16451 8313
rect 16574 8304 16580 8316
rect 16632 8304 16638 8356
rect 3108 8248 8340 8276
rect 3108 8236 3114 8248
rect 1104 8186 16836 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 16836 8186
rect 1104 8112 16836 8134
rect 1762 8072 1768 8084
rect 1412 8044 1768 8072
rect 1412 7945 1440 8044
rect 1762 8032 1768 8044
rect 1820 8032 1826 8084
rect 2498 8032 2504 8084
rect 2556 8072 2562 8084
rect 2777 8075 2835 8081
rect 2777 8072 2789 8075
rect 2556 8044 2789 8072
rect 2556 8032 2562 8044
rect 2777 8041 2789 8044
rect 2823 8041 2835 8075
rect 2777 8035 2835 8041
rect 4525 8075 4583 8081
rect 4525 8041 4537 8075
rect 4571 8072 4583 8075
rect 4614 8072 4620 8084
rect 4571 8044 4620 8072
rect 4571 8041 4583 8044
rect 4525 8035 4583 8041
rect 4614 8032 4620 8044
rect 4672 8032 4678 8084
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6454 8072 6460 8084
rect 6411 8044 6460 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6454 8032 6460 8044
rect 6512 8032 6518 8084
rect 8757 8075 8815 8081
rect 6564 8044 8340 8072
rect 3602 7964 3608 8016
rect 3660 8004 3666 8016
rect 4341 8007 4399 8013
rect 3660 7976 4200 8004
rect 3660 7964 3666 7976
rect 1397 7939 1455 7945
rect 1397 7905 1409 7939
rect 1443 7905 1455 7939
rect 4172 7936 4200 7976
rect 4341 7973 4353 8007
rect 4387 8004 4399 8007
rect 6086 8004 6092 8016
rect 4387 7976 6092 8004
rect 4387 7973 4399 7976
rect 4341 7967 4399 7973
rect 6086 7964 6092 7976
rect 6144 7964 6150 8016
rect 4522 7936 4528 7948
rect 1397 7899 1455 7905
rect 3160 7908 4108 7936
rect 3160 7880 3188 7908
rect 3142 7828 3148 7880
rect 3200 7828 3206 7880
rect 3418 7828 3424 7880
rect 3476 7868 3482 7880
rect 3789 7871 3847 7877
rect 3789 7868 3801 7871
rect 3476 7840 3801 7868
rect 3476 7828 3482 7840
rect 3789 7837 3801 7840
rect 3835 7837 3847 7871
rect 3789 7831 3847 7837
rect 3881 7871 3939 7877
rect 3881 7837 3893 7871
rect 3927 7868 3939 7871
rect 3970 7868 3976 7880
rect 3927 7840 3976 7868
rect 3927 7837 3939 7840
rect 3881 7831 3939 7837
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4080 7877 4108 7908
rect 4172 7908 4528 7936
rect 4172 7877 4200 7908
rect 4522 7896 4528 7908
rect 4580 7896 4586 7948
rect 4985 7939 5043 7945
rect 4985 7905 4997 7939
rect 5031 7936 5043 7939
rect 5350 7936 5356 7948
rect 5031 7908 5356 7936
rect 5031 7905 5043 7908
rect 4985 7899 5043 7905
rect 5350 7896 5356 7908
rect 5408 7936 5414 7948
rect 6564 7936 6592 8044
rect 8312 8004 8340 8044
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9030 8072 9036 8084
rect 8803 8044 9036 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9030 8032 9036 8044
rect 9088 8032 9094 8084
rect 10686 8072 10692 8084
rect 9140 8044 10692 8072
rect 9140 8004 9168 8044
rect 10686 8032 10692 8044
rect 10744 8072 10750 8084
rect 12894 8072 12900 8084
rect 10744 8044 12900 8072
rect 10744 8032 10750 8044
rect 12894 8032 12900 8044
rect 12952 8032 12958 8084
rect 13170 8032 13176 8084
rect 13228 8032 13234 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 14274 8072 14280 8084
rect 13679 8044 14280 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 14274 8032 14280 8044
rect 14332 8032 14338 8084
rect 8312 7976 9168 8004
rect 6825 7939 6883 7945
rect 6825 7936 6837 7939
rect 5408 7908 6592 7936
rect 6656 7908 6837 7936
rect 5408 7896 5414 7908
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7837 4215 7871
rect 4157 7831 4215 7837
rect 4246 7828 4252 7880
rect 4304 7868 4310 7880
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4304 7840 4813 7868
rect 4304 7828 4310 7840
rect 4801 7837 4813 7840
rect 4847 7868 4859 7871
rect 4893 7871 4951 7877
rect 4893 7868 4905 7871
rect 4847 7840 4905 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 4893 7837 4905 7840
rect 4939 7868 4951 7871
rect 5258 7868 5264 7880
rect 4939 7840 5264 7868
rect 4939 7837 4951 7840
rect 4893 7831 4951 7837
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5994 7828 6000 7880
rect 6052 7868 6058 7880
rect 6656 7868 6684 7908
rect 6825 7905 6837 7908
rect 6871 7905 6883 7939
rect 6825 7899 6883 7905
rect 7009 7939 7067 7945
rect 7009 7905 7021 7939
rect 7055 7936 7067 7939
rect 13078 7936 13084 7948
rect 7055 7908 7512 7936
rect 7055 7905 7067 7908
rect 7009 7899 7067 7905
rect 6052 7840 6684 7868
rect 6052 7828 6058 7840
rect 6730 7828 6736 7880
rect 6788 7828 6794 7880
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 7484 7868 7512 7908
rect 12728 7908 13084 7936
rect 7484 7840 8340 7868
rect 8312 7812 8340 7840
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 8941 7871 8999 7877
rect 8941 7868 8953 7871
rect 8904 7840 8953 7868
rect 8904 7828 8910 7840
rect 8941 7837 8953 7840
rect 8987 7837 8999 7871
rect 8941 7831 8999 7837
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7868 9275 7871
rect 9766 7868 9772 7880
rect 9263 7840 9772 7868
rect 9263 7837 9275 7840
rect 9217 7831 9275 7837
rect 9766 7828 9772 7840
rect 9824 7868 9830 7880
rect 10873 7871 10931 7877
rect 9824 7840 10180 7868
rect 9824 7828 9830 7840
rect 10152 7812 10180 7840
rect 10873 7837 10885 7871
rect 10919 7868 10931 7871
rect 11882 7868 11888 7880
rect 10919 7840 11888 7868
rect 10919 7837 10931 7840
rect 10873 7831 10931 7837
rect 11882 7828 11888 7840
rect 11940 7828 11946 7880
rect 12158 7828 12164 7880
rect 12216 7868 12222 7880
rect 12728 7877 12756 7908
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 12529 7871 12587 7877
rect 12529 7868 12541 7871
rect 12216 7840 12541 7868
rect 12216 7828 12222 7840
rect 12529 7837 12541 7840
rect 12575 7837 12587 7871
rect 12529 7831 12587 7837
rect 12713 7871 12771 7877
rect 12713 7837 12725 7871
rect 12759 7837 12771 7871
rect 12713 7831 12771 7837
rect 12802 7828 12808 7880
rect 12860 7828 12866 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 1670 7809 1676 7812
rect 1664 7763 1676 7809
rect 1670 7760 1676 7763
rect 1728 7760 1734 7812
rect 4614 7760 4620 7812
rect 4672 7800 4678 7812
rect 7644 7803 7702 7809
rect 4672 7772 7420 7800
rect 4672 7760 4678 7772
rect 2958 7692 2964 7744
rect 3016 7692 3022 7744
rect 7392 7732 7420 7772
rect 7644 7769 7656 7803
rect 7690 7800 7702 7803
rect 8018 7800 8024 7812
rect 7690 7772 8024 7800
rect 7690 7769 7702 7772
rect 7644 7763 7702 7769
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 8294 7760 8300 7812
rect 8352 7800 8358 7812
rect 8662 7800 8668 7812
rect 8352 7772 8668 7800
rect 8352 7760 8358 7772
rect 8662 7760 8668 7772
rect 8720 7760 8726 7812
rect 9490 7809 9496 7812
rect 9484 7763 9496 7809
rect 9490 7760 9496 7763
rect 9548 7760 9554 7812
rect 10134 7760 10140 7812
rect 10192 7760 10198 7812
rect 11140 7803 11198 7809
rect 11140 7769 11152 7803
rect 11186 7800 11198 7803
rect 11514 7800 11520 7812
rect 11186 7772 11520 7800
rect 11186 7769 11198 7772
rect 11140 7763 11198 7769
rect 11514 7760 11520 7772
rect 11572 7760 11578 7812
rect 12434 7760 12440 7812
rect 12492 7800 12498 7812
rect 12912 7800 12940 7831
rect 12986 7828 12992 7880
rect 13044 7868 13050 7880
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 13044 7840 13461 7868
rect 13044 7828 13050 7840
rect 13449 7837 13461 7840
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 12492 7772 12940 7800
rect 13265 7803 13323 7809
rect 12492 7760 12498 7772
rect 13265 7769 13277 7803
rect 13311 7800 13323 7803
rect 13311 7772 13400 7800
rect 13311 7769 13323 7772
rect 13265 7763 13323 7769
rect 13372 7744 13400 7772
rect 9033 7735 9091 7741
rect 9033 7732 9045 7735
rect 7392 7704 9045 7732
rect 9033 7701 9045 7704
rect 9079 7732 9091 7735
rect 9306 7732 9312 7744
rect 9079 7704 9312 7732
rect 9079 7701 9091 7704
rect 9033 7695 9091 7701
rect 9306 7692 9312 7704
rect 9364 7732 9370 7744
rect 9674 7732 9680 7744
rect 9364 7704 9680 7732
rect 9364 7692 9370 7704
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10597 7735 10655 7741
rect 10597 7701 10609 7735
rect 10643 7732 10655 7735
rect 10870 7732 10876 7744
rect 10643 7704 10876 7732
rect 10643 7701 10655 7704
rect 10597 7695 10655 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 12253 7735 12311 7741
rect 12253 7701 12265 7735
rect 12299 7732 12311 7735
rect 12618 7732 12624 7744
rect 12299 7704 12624 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 12802 7692 12808 7744
rect 12860 7732 12866 7744
rect 13078 7732 13084 7744
rect 12860 7704 13084 7732
rect 12860 7692 12866 7704
rect 13078 7692 13084 7704
rect 13136 7692 13142 7744
rect 13354 7692 13360 7744
rect 13412 7692 13418 7744
rect 13464 7732 13492 7831
rect 14090 7828 14096 7880
rect 14148 7868 14154 7880
rect 15102 7868 15108 7880
rect 14148 7840 15108 7868
rect 14148 7828 14154 7840
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 14360 7803 14418 7809
rect 14360 7769 14372 7803
rect 14406 7800 14418 7803
rect 14734 7800 14740 7812
rect 14406 7772 14740 7800
rect 14406 7769 14418 7772
rect 14360 7763 14418 7769
rect 14734 7760 14740 7772
rect 14792 7760 14798 7812
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 13464 7704 15485 7732
rect 15473 7701 15485 7704
rect 15519 7732 15531 7735
rect 16206 7732 16212 7744
rect 15519 7704 16212 7732
rect 15519 7701 15531 7704
rect 15473 7695 15531 7701
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 1104 7642 16836 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 16836 7642
rect 1104 7568 16836 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1670 7528 1676 7540
rect 1627 7500 1676 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 4798 7528 4804 7540
rect 3375 7500 4804 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 8389 7531 8447 7537
rect 8389 7497 8401 7531
rect 8435 7528 8447 7531
rect 9030 7528 9036 7540
rect 8435 7500 9036 7528
rect 8435 7497 8447 7500
rect 8389 7491 8447 7497
rect 9030 7488 9036 7500
rect 9088 7488 9094 7540
rect 9125 7531 9183 7537
rect 9125 7497 9137 7531
rect 9171 7528 9183 7531
rect 9398 7528 9404 7540
rect 9171 7500 9404 7528
rect 9171 7497 9183 7500
rect 9125 7491 9183 7497
rect 9398 7488 9404 7500
rect 9456 7528 9462 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9456 7500 9597 7528
rect 9456 7488 9462 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 11330 7528 11336 7540
rect 9585 7491 9643 7497
rect 10612 7500 11336 7528
rect 2317 7463 2375 7469
rect 2317 7460 2329 7463
rect 2056 7432 2329 7460
rect 1857 7395 1915 7401
rect 1857 7361 1869 7395
rect 1903 7361 1915 7395
rect 1857 7355 1915 7361
rect 1872 7188 1900 7355
rect 1946 7352 1952 7404
rect 2004 7352 2010 7404
rect 2056 7401 2084 7432
rect 2317 7429 2329 7432
rect 2363 7429 2375 7463
rect 2317 7423 2375 7429
rect 2498 7420 2504 7472
rect 2556 7460 2562 7472
rect 2556 7432 2820 7460
rect 2556 7420 2562 7432
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2225 7355 2283 7361
rect 1964 7256 1992 7352
rect 2240 7324 2268 7355
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 2792 7401 2820 7432
rect 2866 7420 2872 7472
rect 2924 7460 2930 7472
rect 3053 7463 3111 7469
rect 3053 7460 3065 7463
rect 2924 7432 3065 7460
rect 2924 7420 2930 7432
rect 3053 7429 3065 7432
rect 3099 7429 3111 7463
rect 3053 7423 3111 7429
rect 3160 7432 3832 7460
rect 2685 7395 2743 7401
rect 2685 7392 2697 7395
rect 2648 7364 2697 7392
rect 2648 7352 2654 7364
rect 2685 7361 2697 7364
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7361 2835 7395
rect 2777 7355 2835 7361
rect 2958 7352 2964 7404
rect 3016 7352 3022 7404
rect 3160 7401 3188 7432
rect 3160 7395 3227 7401
rect 3160 7364 3181 7395
rect 3169 7361 3181 7364
rect 3215 7361 3227 7395
rect 3804 7392 3832 7432
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4341 7463 4399 7469
rect 4341 7460 4353 7463
rect 4212 7432 4353 7460
rect 4212 7420 4218 7432
rect 4341 7429 4353 7432
rect 4387 7429 4399 7463
rect 4341 7423 4399 7429
rect 4522 7420 4528 7472
rect 4580 7460 4586 7472
rect 4580 7432 5488 7460
rect 4580 7420 4586 7432
rect 3804 7364 4200 7392
rect 3169 7355 3227 7361
rect 3694 7324 3700 7336
rect 2240 7296 3700 7324
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 4172 7324 4200 7364
rect 4246 7352 4252 7404
rect 4304 7352 4310 7404
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 4614 7392 4620 7404
rect 4479 7364 4620 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4985 7395 5043 7401
rect 4985 7361 4997 7395
rect 5031 7361 5043 7395
rect 4985 7355 5043 7361
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5350 7392 5356 7404
rect 5215 7364 5356 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5000 7324 5028 7355
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 5460 7392 5488 7432
rect 6178 7420 6184 7472
rect 6236 7460 6242 7472
rect 6236 7432 7052 7460
rect 6236 7420 6242 7432
rect 7024 7401 7052 7432
rect 9306 7420 9312 7472
rect 9364 7420 9370 7472
rect 10612 7460 10640 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 11514 7488 11520 7540
rect 11572 7488 11578 7540
rect 15197 7531 15255 7537
rect 15197 7497 15209 7531
rect 15243 7497 15255 7531
rect 15197 7491 15255 7497
rect 9600 7432 10640 7460
rect 10689 7463 10747 7469
rect 6917 7395 6975 7401
rect 6917 7392 6929 7395
rect 5460 7364 6929 7392
rect 6917 7361 6929 7364
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 7190 7352 7196 7404
rect 7248 7352 7254 7404
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 9600 7392 9628 7432
rect 10689 7429 10701 7463
rect 10735 7460 10747 7463
rect 12250 7460 12256 7472
rect 10735 7432 12256 7460
rect 10735 7429 10747 7432
rect 10689 7423 10747 7429
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 12710 7420 12716 7472
rect 12768 7460 12774 7472
rect 15212 7460 15240 7491
rect 12768 7432 13492 7460
rect 12768 7420 12774 7432
rect 7331 7364 9628 7392
rect 9677 7395 9735 7401
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 9677 7361 9689 7395
rect 9723 7392 9735 7395
rect 9858 7392 9864 7404
rect 9723 7364 9864 7392
rect 9723 7361 9735 7364
rect 9677 7355 9735 7361
rect 9858 7352 9864 7364
rect 9916 7392 9922 7404
rect 10870 7392 10876 7404
rect 9916 7364 10876 7392
rect 9916 7352 9922 7364
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 11790 7352 11796 7404
rect 11848 7352 11854 7404
rect 11885 7395 11943 7401
rect 11885 7361 11897 7395
rect 11931 7361 11943 7395
rect 11885 7355 11943 7361
rect 11977 7395 12035 7401
rect 11977 7361 11989 7395
rect 12023 7361 12035 7395
rect 11977 7355 12035 7361
rect 5442 7324 5448 7336
rect 4172 7296 5448 7324
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 8386 7284 8392 7336
rect 8444 7324 8450 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8444 7296 8493 7324
rect 8444 7284 8450 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 8662 7284 8668 7336
rect 8720 7284 8726 7336
rect 9953 7327 10011 7333
rect 9953 7293 9965 7327
rect 9999 7324 10011 7327
rect 10134 7324 10140 7336
rect 9999 7296 10140 7324
rect 9999 7293 10011 7296
rect 9953 7287 10011 7293
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 10781 7327 10839 7333
rect 10781 7324 10793 7327
rect 10744 7296 10793 7324
rect 10744 7284 10750 7296
rect 10781 7293 10793 7296
rect 10827 7293 10839 7327
rect 11900 7324 11928 7355
rect 10781 7287 10839 7293
rect 10888 7296 11928 7324
rect 11992 7324 12020 7355
rect 12158 7352 12164 7404
rect 12216 7352 12222 7404
rect 12342 7352 12348 7404
rect 12400 7352 12406 7404
rect 12529 7395 12587 7401
rect 12529 7361 12541 7395
rect 12575 7392 12587 7395
rect 12618 7392 12624 7404
rect 12575 7364 12624 7392
rect 12575 7361 12587 7364
rect 12529 7355 12587 7361
rect 12618 7352 12624 7364
rect 12676 7352 12682 7404
rect 12820 7401 12848 7432
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7361 12863 7395
rect 12805 7355 12863 7361
rect 12894 7352 12900 7404
rect 12952 7392 12958 7404
rect 13464 7401 13492 7432
rect 14476 7432 15240 7460
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12952 7364 13001 7392
rect 12952 7352 12958 7364
rect 12989 7361 13001 7364
rect 13035 7392 13047 7395
rect 13265 7395 13323 7401
rect 13265 7392 13277 7395
rect 13035 7364 13277 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13265 7361 13277 7364
rect 13311 7361 13323 7395
rect 13265 7355 13323 7361
rect 13449 7395 13507 7401
rect 13449 7361 13461 7395
rect 13495 7392 13507 7395
rect 13538 7392 13544 7404
rect 13495 7364 13544 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14476 7401 14504 7432
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 14332 7364 14473 7392
rect 14332 7352 14338 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 14642 7352 14648 7404
rect 14700 7352 14706 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7361 14795 7395
rect 14737 7355 14795 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7392 14887 7395
rect 14918 7392 14924 7404
rect 14875 7364 14924 7392
rect 14875 7361 14887 7364
rect 14829 7355 14887 7361
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 11992 7296 12725 7324
rect 6733 7259 6791 7265
rect 1964 7228 6684 7256
rect 2682 7188 2688 7200
rect 1872 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7188 2746 7200
rect 2958 7188 2964 7200
rect 2740 7160 2964 7188
rect 2740 7148 2746 7160
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4672 7160 4813 7188
rect 4672 7148 4678 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 6656 7188 6684 7228
rect 6733 7225 6745 7259
rect 6779 7256 6791 7259
rect 10594 7256 10600 7268
rect 6779 7228 10600 7256
rect 6779 7225 6791 7228
rect 6733 7219 6791 7225
rect 10594 7216 10600 7228
rect 10652 7216 10658 7268
rect 8570 7188 8576 7200
rect 6656 7160 8576 7188
rect 4801 7151 4859 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 8938 7148 8944 7200
rect 8996 7148 9002 7200
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9125 7191 9183 7197
rect 9125 7188 9137 7191
rect 9088 7160 9137 7188
rect 9088 7148 9094 7160
rect 9125 7157 9137 7160
rect 9171 7157 9183 7191
rect 9125 7151 9183 7157
rect 10502 7148 10508 7200
rect 10560 7188 10566 7200
rect 10888 7188 10916 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 13078 7284 13084 7336
rect 13136 7324 13142 7336
rect 14366 7324 14372 7336
rect 13136 7296 14372 7324
rect 13136 7284 13142 7296
rect 14366 7284 14372 7296
rect 14424 7324 14430 7336
rect 14752 7324 14780 7355
rect 14918 7352 14924 7364
rect 14976 7352 14982 7404
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 14424 7296 14780 7324
rect 14424 7284 14430 7296
rect 12342 7256 12348 7268
rect 11164 7228 12348 7256
rect 10560 7160 10916 7188
rect 10560 7148 10566 7160
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11164 7197 11192 7228
rect 12342 7216 12348 7228
rect 12400 7216 12406 7268
rect 14458 7256 14464 7268
rect 12820 7228 14464 7256
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 11112 7160 11161 7188
rect 11112 7148 11118 7160
rect 11149 7157 11161 7160
rect 11195 7157 11207 7191
rect 11149 7151 11207 7157
rect 11790 7148 11796 7200
rect 11848 7188 11854 7200
rect 12820 7188 12848 7228
rect 14458 7216 14464 7228
rect 14516 7216 14522 7268
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7256 15163 7259
rect 15378 7256 15384 7268
rect 15151 7228 15384 7256
rect 15151 7225 15163 7228
rect 15105 7219 15163 7225
rect 15378 7216 15384 7228
rect 15436 7216 15442 7268
rect 11848 7160 12848 7188
rect 11848 7148 11854 7160
rect 12894 7148 12900 7200
rect 12952 7148 12958 7200
rect 13446 7148 13452 7200
rect 13504 7188 13510 7200
rect 13633 7191 13691 7197
rect 13633 7188 13645 7191
rect 13504 7160 13645 7188
rect 13504 7148 13510 7160
rect 13633 7157 13645 7160
rect 13679 7157 13691 7191
rect 13633 7151 13691 7157
rect 1104 7098 16836 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 16836 7098
rect 1104 7024 16836 7046
rect 2774 6944 2780 6996
rect 2832 6984 2838 6996
rect 3050 6984 3056 6996
rect 2832 6956 3056 6984
rect 2832 6944 2838 6956
rect 3050 6944 3056 6956
rect 3108 6944 3114 6996
rect 5445 6987 5503 6993
rect 5445 6984 5457 6987
rect 4632 6956 5457 6984
rect 1762 6808 1768 6860
rect 1820 6848 1826 6860
rect 2038 6848 2044 6860
rect 1820 6820 2044 6848
rect 1820 6808 1826 6820
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 4632 6848 4660 6956
rect 4632 6820 4752 6848
rect 3786 6740 3792 6792
rect 3844 6780 3850 6792
rect 4430 6780 4436 6792
rect 3844 6752 4436 6780
rect 3844 6740 3850 6752
rect 4430 6740 4436 6752
rect 4488 6740 4494 6792
rect 4522 6740 4528 6792
rect 4580 6780 4586 6792
rect 4724 6789 4752 6820
rect 5368 6792 5396 6956
rect 5445 6953 5457 6956
rect 5491 6953 5503 6987
rect 5445 6947 5503 6953
rect 9490 6944 9496 6996
rect 9548 6944 9554 6996
rect 13909 6987 13967 6993
rect 13909 6953 13921 6987
rect 13955 6984 13967 6987
rect 14642 6984 14648 6996
rect 13955 6956 14648 6984
rect 13955 6953 13967 6956
rect 13909 6947 13967 6953
rect 14642 6944 14648 6956
rect 14700 6944 14706 6996
rect 8386 6876 8392 6928
rect 8444 6916 8450 6928
rect 13354 6916 13360 6928
rect 8444 6888 13360 6916
rect 8444 6876 8450 6888
rect 13354 6876 13360 6888
rect 13412 6876 13418 6928
rect 8662 6808 8668 6860
rect 8720 6848 8726 6860
rect 10045 6851 10103 6857
rect 10045 6848 10057 6851
rect 8720 6820 10057 6848
rect 8720 6808 8726 6820
rect 10045 6817 10057 6820
rect 10091 6817 10103 6851
rect 10045 6811 10103 6817
rect 10870 6808 10876 6860
rect 10928 6808 10934 6860
rect 14918 6848 14924 6860
rect 14660 6820 14924 6848
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4580 6752 4629 6780
rect 4580 6740 4586 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 4709 6783 4767 6789
rect 4709 6749 4721 6783
rect 4755 6749 4767 6783
rect 4709 6743 4767 6749
rect 4798 6740 4804 6792
rect 4856 6740 4862 6792
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 5442 6740 5448 6792
rect 5500 6780 5506 6792
rect 5537 6783 5595 6789
rect 5537 6780 5549 6783
rect 5500 6752 5549 6780
rect 5500 6740 5506 6752
rect 5537 6749 5549 6752
rect 5583 6780 5595 6783
rect 6546 6780 6552 6792
rect 5583 6752 6552 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 6546 6740 6552 6752
rect 6604 6740 6610 6792
rect 7374 6780 7380 6792
rect 6932 6752 7380 6780
rect 2308 6715 2366 6721
rect 2308 6681 2320 6715
rect 2354 6712 2366 6715
rect 2682 6712 2688 6724
rect 2354 6684 2688 6712
rect 2354 6681 2366 6684
rect 2308 6675 2366 6681
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 3973 6715 4031 6721
rect 3973 6712 3985 6715
rect 3436 6684 3985 6712
rect 2866 6604 2872 6656
rect 2924 6644 2930 6656
rect 3436 6653 3464 6684
rect 3973 6681 3985 6684
rect 4019 6681 4031 6715
rect 3973 6675 4031 6681
rect 4154 6672 4160 6724
rect 4212 6672 4218 6724
rect 4816 6712 4844 6740
rect 6932 6724 6960 6752
rect 7374 6740 7380 6752
rect 7432 6740 7438 6792
rect 7745 6783 7803 6789
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 4816 6684 6132 6712
rect 3421 6647 3479 6653
rect 3421 6644 3433 6647
rect 2924 6616 3433 6644
rect 2924 6604 2930 6616
rect 3421 6613 3433 6616
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 3786 6604 3792 6656
rect 3844 6604 3850 6656
rect 4172 6644 4200 6672
rect 4614 6644 4620 6656
rect 4172 6616 4620 6644
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5077 6647 5135 6653
rect 5077 6644 5089 6647
rect 4764 6616 5089 6644
rect 4764 6604 4770 6616
rect 5077 6613 5089 6616
rect 5123 6613 5135 6647
rect 5077 6607 5135 6613
rect 5994 6604 6000 6656
rect 6052 6604 6058 6656
rect 6104 6644 6132 6684
rect 6914 6672 6920 6724
rect 6972 6672 6978 6724
rect 7132 6715 7190 6721
rect 7132 6681 7144 6715
rect 7178 6712 7190 6715
rect 7469 6715 7527 6721
rect 7469 6712 7481 6715
rect 7178 6684 7481 6712
rect 7178 6681 7190 6684
rect 7132 6675 7190 6681
rect 7469 6681 7481 6684
rect 7515 6681 7527 6715
rect 7469 6675 7527 6681
rect 7760 6712 7788 6743
rect 7834 6740 7840 6792
rect 7892 6740 7898 6792
rect 7926 6740 7932 6792
rect 7984 6740 7990 6792
rect 8018 6740 8024 6792
rect 8076 6780 8082 6792
rect 8113 6783 8171 6789
rect 8113 6780 8125 6783
rect 8076 6752 8125 6780
rect 8076 6740 8082 6752
rect 8113 6749 8125 6752
rect 8159 6749 8171 6783
rect 11790 6780 11796 6792
rect 8113 6743 8171 6749
rect 9784 6752 11796 6780
rect 9784 6712 9812 6752
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 14274 6740 14280 6792
rect 14332 6740 14338 6792
rect 14458 6740 14464 6792
rect 14516 6740 14522 6792
rect 14660 6789 14688 6820
rect 14918 6808 14924 6820
rect 14976 6808 14982 6860
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 14645 6783 14703 6789
rect 14645 6749 14657 6783
rect 14691 6749 14703 6783
rect 14645 6743 14703 6749
rect 15013 6783 15071 6789
rect 15013 6749 15025 6783
rect 15059 6780 15071 6783
rect 15102 6780 15108 6792
rect 15059 6752 15108 6780
rect 15059 6749 15071 6752
rect 15013 6743 15071 6749
rect 7760 6684 9812 6712
rect 9861 6715 9919 6721
rect 7760 6644 7788 6684
rect 9861 6681 9873 6715
rect 9907 6712 9919 6715
rect 10321 6715 10379 6721
rect 10321 6712 10333 6715
rect 9907 6684 10333 6712
rect 9907 6681 9919 6684
rect 9861 6675 9919 6681
rect 10321 6681 10333 6684
rect 10367 6681 10379 6715
rect 10321 6675 10379 6681
rect 11146 6672 11152 6724
rect 11204 6672 11210 6724
rect 13446 6672 13452 6724
rect 13504 6712 13510 6724
rect 13541 6715 13599 6721
rect 13541 6712 13553 6715
rect 13504 6684 13553 6712
rect 13504 6672 13510 6684
rect 13541 6681 13553 6684
rect 13587 6681 13599 6715
rect 13541 6675 13599 6681
rect 13725 6715 13783 6721
rect 13725 6681 13737 6715
rect 13771 6712 13783 6715
rect 14366 6712 14372 6724
rect 13771 6684 14372 6712
rect 13771 6681 13783 6684
rect 13725 6675 13783 6681
rect 14366 6672 14372 6684
rect 14424 6672 14430 6724
rect 6104 6616 7788 6644
rect 9953 6647 10011 6653
rect 9953 6613 9965 6647
rect 9999 6644 10011 6647
rect 10042 6644 10048 6656
rect 9999 6616 10048 6644
rect 9999 6613 10011 6616
rect 9953 6607 10011 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 11238 6604 11244 6656
rect 11296 6604 11302 6656
rect 13262 6604 13268 6656
rect 13320 6644 13326 6656
rect 14568 6644 14596 6743
rect 15102 6740 15108 6752
rect 15160 6740 15166 6792
rect 14921 6715 14979 6721
rect 14921 6681 14933 6715
rect 14967 6712 14979 6715
rect 15258 6715 15316 6721
rect 15258 6712 15270 6715
rect 14967 6684 15270 6712
rect 14967 6681 14979 6684
rect 14921 6675 14979 6681
rect 15258 6681 15270 6684
rect 15304 6681 15316 6715
rect 15258 6675 15316 6681
rect 13320 6616 14596 6644
rect 13320 6604 13326 6616
rect 15838 6604 15844 6656
rect 15896 6644 15902 6656
rect 16393 6647 16451 6653
rect 16393 6644 16405 6647
rect 15896 6616 16405 6644
rect 15896 6604 15902 6616
rect 16393 6613 16405 6616
rect 16439 6613 16451 6647
rect 16393 6607 16451 6613
rect 1104 6554 16836 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 16836 6554
rect 1104 6480 16836 6502
rect 2682 6400 2688 6452
rect 2740 6400 2746 6452
rect 4522 6400 4528 6452
rect 4580 6400 4586 6452
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 5258 6440 5264 6452
rect 4672 6412 5264 6440
rect 4672 6400 4678 6412
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 6917 6443 6975 6449
rect 6917 6409 6929 6443
rect 6963 6440 6975 6443
rect 7006 6440 7012 6452
rect 6963 6412 7012 6440
rect 6963 6409 6975 6412
rect 6917 6403 6975 6409
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7377 6443 7435 6449
rect 7377 6409 7389 6443
rect 7423 6440 7435 6443
rect 7926 6440 7932 6452
rect 7423 6412 7932 6440
rect 7423 6409 7435 6412
rect 7377 6403 7435 6409
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8662 6400 8668 6452
rect 8720 6440 8726 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8720 6412 9045 6440
rect 8720 6400 8726 6412
rect 9033 6409 9045 6412
rect 9079 6440 9091 6443
rect 11146 6440 11152 6452
rect 9079 6412 11152 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 11146 6400 11152 6412
rect 11204 6400 11210 6452
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 14185 6443 14243 6449
rect 11940 6412 13584 6440
rect 11940 6400 11946 6412
rect 13556 6384 13584 6412
rect 14185 6409 14197 6443
rect 14231 6440 14243 6443
rect 14458 6440 14464 6452
rect 14231 6412 14464 6440
rect 14231 6409 14243 6412
rect 14185 6403 14243 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 16206 6440 16212 6452
rect 14568 6412 16212 6440
rect 3786 6372 3792 6384
rect 3160 6344 3792 6372
rect 2958 6264 2964 6316
rect 3016 6264 3022 6316
rect 3050 6264 3056 6316
rect 3108 6264 3114 6316
rect 3160 6313 3188 6344
rect 3786 6332 3792 6344
rect 3844 6332 3850 6384
rect 4430 6372 4436 6384
rect 3896 6344 4436 6372
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6273 3203 6307
rect 3145 6267 3203 6273
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6304 3479 6307
rect 3896 6304 3924 6344
rect 4430 6332 4436 6344
rect 4488 6332 4494 6384
rect 5442 6372 5448 6384
rect 4632 6344 5448 6372
rect 3467 6276 3924 6304
rect 3467 6273 3479 6276
rect 3421 6267 3479 6273
rect 3344 6236 3372 6267
rect 4154 6264 4160 6316
rect 4212 6264 4218 6316
rect 4632 6313 4660 6344
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 5994 6332 6000 6384
rect 6052 6372 6058 6384
rect 6641 6375 6699 6381
rect 6641 6372 6653 6375
rect 6052 6344 6653 6372
rect 6052 6332 6058 6344
rect 6641 6341 6653 6344
rect 6687 6372 6699 6375
rect 7193 6375 7251 6381
rect 7193 6372 7205 6375
rect 6687 6344 7205 6372
rect 6687 6341 6699 6344
rect 6641 6335 6699 6341
rect 7193 6341 7205 6344
rect 7239 6341 7251 6375
rect 7193 6335 7251 6341
rect 9582 6332 9588 6384
rect 9640 6372 9646 6384
rect 12342 6372 12348 6384
rect 9640 6344 12348 6372
rect 9640 6332 9646 6344
rect 12342 6332 12348 6344
rect 12400 6332 12406 6384
rect 13538 6332 13544 6384
rect 13596 6372 13602 6384
rect 13596 6344 14136 6372
rect 13596 6332 13602 6344
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 4617 6307 4675 6313
rect 4387 6276 4568 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 3344 6208 3648 6236
rect 3620 6109 3648 6208
rect 3605 6103 3663 6109
rect 3605 6069 3617 6103
rect 3651 6100 3663 6103
rect 3878 6100 3884 6112
rect 3651 6072 3884 6100
rect 3651 6069 3663 6072
rect 3605 6063 3663 6069
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 4540 6100 4568 6276
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 4873 6307 4931 6313
rect 4873 6304 4885 6307
rect 4764 6276 4885 6304
rect 4764 6264 4770 6276
rect 4873 6273 4885 6276
rect 4919 6273 4931 6307
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 4873 6267 4931 6273
rect 6012 6276 6377 6304
rect 4798 6100 4804 6112
rect 4540 6072 4804 6100
rect 4798 6060 4804 6072
rect 4856 6100 4862 6112
rect 6012 6109 6040 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 6564 6168 6592 6264
rect 6748 6236 6776 6267
rect 7006 6264 7012 6316
rect 7064 6264 7070 6316
rect 8846 6264 8852 6316
rect 8904 6304 8910 6316
rect 8941 6307 8999 6313
rect 8941 6304 8953 6307
rect 8904 6276 8953 6304
rect 8904 6264 8910 6276
rect 8941 6273 8953 6276
rect 8987 6273 8999 6307
rect 8941 6267 8999 6273
rect 9030 6264 9036 6316
rect 9088 6304 9094 6316
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 9088 6276 9229 6304
rect 9088 6264 9094 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 9217 6267 9275 6273
rect 9398 6264 9404 6316
rect 9456 6264 9462 6316
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 10209 6307 10267 6313
rect 10209 6304 10221 6307
rect 9916 6276 10221 6304
rect 9916 6264 9922 6276
rect 10209 6273 10221 6276
rect 10255 6273 10267 6307
rect 10209 6267 10267 6273
rect 11238 6264 11244 6316
rect 11296 6304 11302 6316
rect 12621 6307 12679 6313
rect 12621 6304 12633 6307
rect 11296 6276 12633 6304
rect 11296 6264 11302 6276
rect 7098 6236 7104 6248
rect 6748 6208 7104 6236
rect 7098 6196 7104 6208
rect 7156 6196 7162 6248
rect 9953 6239 10011 6245
rect 9953 6205 9965 6239
rect 9999 6205 10011 6239
rect 9953 6199 10011 6205
rect 8938 6168 8944 6180
rect 6564 6140 8944 6168
rect 8938 6128 8944 6140
rect 8996 6128 9002 6180
rect 5997 6103 6055 6109
rect 5997 6100 6009 6103
rect 4856 6072 6009 6100
rect 4856 6060 4862 6072
rect 5997 6069 6009 6072
rect 6043 6069 6055 6103
rect 9968 6100 9996 6199
rect 10134 6100 10140 6112
rect 9968 6072 10140 6100
rect 5997 6063 6055 6069
rect 10134 6060 10140 6072
rect 10192 6060 10198 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 10284 6072 11345 6100
rect 10284 6060 10290 6072
rect 11333 6069 11345 6072
rect 11379 6100 11391 6103
rect 11422 6100 11428 6112
rect 11379 6072 11428 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 12360 6100 12388 6276
rect 12621 6273 12633 6276
rect 12667 6304 12679 6307
rect 12897 6307 12955 6313
rect 12897 6304 12909 6307
rect 12667 6276 12909 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 12897 6273 12909 6276
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 12802 6196 12808 6248
rect 12860 6236 12866 6248
rect 13096 6236 13124 6267
rect 12860 6208 13124 6236
rect 12860 6196 12866 6208
rect 13262 6196 13268 6248
rect 13320 6196 13326 6248
rect 13832 6180 13860 6267
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14001 6307 14059 6313
rect 14001 6304 14013 6307
rect 13964 6276 14013 6304
rect 13964 6264 13970 6276
rect 14001 6273 14013 6276
rect 14047 6273 14059 6307
rect 14108 6304 14136 6344
rect 14366 6332 14372 6384
rect 14424 6372 14430 6384
rect 14568 6381 14596 6412
rect 16206 6400 16212 6412
rect 16264 6440 16270 6452
rect 16485 6443 16543 6449
rect 16485 6440 16497 6443
rect 16264 6412 16497 6440
rect 16264 6400 16270 6412
rect 16485 6409 16497 6412
rect 16531 6409 16543 6443
rect 16485 6403 16543 6409
rect 15378 6381 15384 6384
rect 14553 6375 14611 6381
rect 14553 6372 14565 6375
rect 14424 6344 14565 6372
rect 14424 6332 14430 6344
rect 14553 6341 14565 6344
rect 14599 6341 14611 6375
rect 15372 6372 15384 6381
rect 15339 6344 15384 6372
rect 14553 6335 14611 6341
rect 15372 6335 15384 6344
rect 15378 6332 15384 6335
rect 15436 6332 15442 6384
rect 14458 6304 14464 6316
rect 14108 6276 14464 6304
rect 14001 6267 14059 6273
rect 14458 6264 14464 6276
rect 14516 6264 14522 6316
rect 14642 6264 14648 6316
rect 14700 6264 14706 6316
rect 14826 6264 14832 6316
rect 14884 6304 14890 6316
rect 15838 6304 15844 6316
rect 14884 6276 15844 6304
rect 14884 6264 14890 6276
rect 15838 6264 15844 6276
rect 15896 6264 15902 6316
rect 15102 6196 15108 6248
rect 15160 6196 15166 6248
rect 12437 6171 12495 6177
rect 12437 6137 12449 6171
rect 12483 6168 12495 6171
rect 13814 6168 13820 6180
rect 12483 6140 13820 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 13814 6128 13820 6140
rect 13872 6128 13878 6180
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 14277 6171 14335 6177
rect 14277 6168 14289 6171
rect 14056 6140 14289 6168
rect 14056 6128 14062 6140
rect 14277 6137 14289 6140
rect 14323 6137 14335 6171
rect 14277 6131 14335 6137
rect 14458 6128 14464 6180
rect 14516 6168 14522 6180
rect 14918 6168 14924 6180
rect 14516 6140 14924 6168
rect 14516 6128 14522 6140
rect 14918 6128 14924 6140
rect 14976 6128 14982 6180
rect 14642 6100 14648 6112
rect 12360 6072 14648 6100
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 1104 6010 16836 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 16836 6010
rect 1104 5936 16836 5958
rect 2746 5868 8708 5896
rect 2222 5788 2228 5840
rect 2280 5828 2286 5840
rect 2590 5828 2596 5840
rect 2280 5800 2596 5828
rect 2280 5788 2286 5800
rect 2590 5788 2596 5800
rect 2648 5828 2654 5840
rect 2746 5828 2774 5868
rect 2648 5800 2774 5828
rect 2648 5788 2654 5800
rect 3050 5788 3056 5840
rect 3108 5828 3114 5840
rect 3108 5800 3188 5828
rect 3108 5788 3114 5800
rect 2866 5760 2872 5772
rect 1688 5732 2872 5760
rect 1688 5701 1716 5732
rect 2866 5720 2872 5732
rect 2924 5720 2930 5772
rect 3160 5760 3188 5800
rect 7006 5788 7012 5840
rect 7064 5788 7070 5840
rect 8680 5828 8708 5868
rect 8754 5856 8760 5908
rect 8812 5856 8818 5908
rect 9858 5856 9864 5908
rect 9916 5856 9922 5908
rect 12176 5868 13768 5896
rect 8680 5800 10088 5828
rect 5350 5760 5356 5772
rect 3160 5732 5356 5760
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 2222 5692 2228 5704
rect 1820 5664 2228 5692
rect 1820 5652 1826 5664
rect 2222 5652 2228 5664
rect 2280 5652 2286 5704
rect 2314 5652 2320 5704
rect 2372 5692 2378 5704
rect 3160 5701 3188 5732
rect 5350 5720 5356 5732
rect 5408 5720 5414 5772
rect 7024 5760 7052 5788
rect 8386 5760 8392 5772
rect 6932 5732 8392 5760
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2372 5664 3065 5692
rect 2372 5652 2378 5664
rect 3053 5661 3065 5664
rect 3099 5661 3111 5695
rect 3053 5655 3111 5661
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 3234 5652 3240 5704
rect 3292 5652 3298 5704
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 3510 5692 3516 5704
rect 3467 5664 3516 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 3510 5652 3516 5664
rect 3568 5692 3574 5704
rect 3878 5692 3884 5704
rect 3568 5664 3884 5692
rect 3568 5652 3574 5664
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 2041 5627 2099 5633
rect 2041 5593 2053 5627
rect 2087 5624 2099 5627
rect 2130 5624 2136 5636
rect 2087 5596 2136 5624
rect 2087 5593 2099 5596
rect 2041 5587 2099 5593
rect 2130 5584 2136 5596
rect 2188 5584 2194 5636
rect 6932 5624 6960 5732
rect 8386 5720 8392 5732
rect 8444 5720 8450 5772
rect 8846 5760 8852 5772
rect 8496 5732 8852 5760
rect 7006 5652 7012 5704
rect 7064 5692 7070 5704
rect 8205 5695 8263 5701
rect 8205 5692 8217 5695
rect 7064 5664 8217 5692
rect 7064 5652 7070 5664
rect 8205 5661 8217 5664
rect 8251 5661 8263 5695
rect 8205 5655 8263 5661
rect 7285 5627 7343 5633
rect 7285 5624 7297 5627
rect 6932 5596 7297 5624
rect 7285 5593 7297 5596
rect 7331 5593 7343 5627
rect 7285 5587 7343 5593
rect 7469 5627 7527 5633
rect 7469 5593 7481 5627
rect 7515 5624 7527 5627
rect 7558 5624 7564 5636
rect 7515 5596 7564 5624
rect 7515 5593 7527 5596
rect 7469 5587 7527 5593
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 8496 5633 8524 5732
rect 8846 5720 8852 5732
rect 8904 5720 8910 5772
rect 9953 5763 10011 5769
rect 9953 5760 9965 5763
rect 9416 5732 9965 5760
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 8754 5692 8760 5704
rect 8619 5664 8760 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 9214 5652 9220 5704
rect 9272 5652 9278 5704
rect 9416 5701 9444 5732
rect 9953 5729 9965 5732
rect 9999 5729 10011 5763
rect 9953 5723 10011 5729
rect 9401 5695 9459 5701
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 9401 5655 9459 5661
rect 9493 5695 9551 5701
rect 9493 5661 9505 5695
rect 9539 5661 9551 5695
rect 9493 5655 9551 5661
rect 8389 5627 8447 5633
rect 8389 5593 8401 5627
rect 8435 5593 8447 5627
rect 8389 5587 8447 5593
rect 8481 5627 8539 5633
rect 8481 5593 8493 5627
rect 8527 5593 8539 5627
rect 8481 5587 8539 5593
rect 1489 5559 1547 5565
rect 1489 5525 1501 5559
rect 1535 5556 1547 5559
rect 1578 5556 1584 5568
rect 1535 5528 1584 5556
rect 1535 5525 1547 5528
rect 1489 5519 1547 5525
rect 1578 5516 1584 5528
rect 1636 5516 1642 5568
rect 1857 5559 1915 5565
rect 1857 5525 1869 5559
rect 1903 5556 1915 5559
rect 1946 5556 1952 5568
rect 1903 5528 1952 5556
rect 1903 5525 1915 5528
rect 1857 5519 1915 5525
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2774 5516 2780 5568
rect 2832 5516 2838 5568
rect 7650 5516 7656 5568
rect 7708 5516 7714 5568
rect 8404 5556 8432 5587
rect 8662 5584 8668 5636
rect 8720 5624 8726 5636
rect 9508 5624 9536 5655
rect 9582 5652 9588 5704
rect 9640 5652 9646 5704
rect 10060 5692 10088 5800
rect 10134 5720 10140 5772
rect 10192 5760 10198 5772
rect 10413 5763 10471 5769
rect 10413 5760 10425 5763
rect 10192 5732 10425 5760
rect 10192 5720 10198 5732
rect 10413 5729 10425 5732
rect 10459 5729 10471 5763
rect 10413 5723 10471 5729
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 10060 5664 10333 5692
rect 10321 5661 10333 5664
rect 10367 5692 10379 5695
rect 11054 5692 11060 5704
rect 10367 5664 11060 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 11054 5652 11060 5664
rect 11112 5692 11118 5704
rect 11238 5692 11244 5704
rect 11112 5664 11244 5692
rect 11112 5652 11118 5664
rect 11238 5652 11244 5664
rect 11296 5652 11302 5704
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12069 5695 12127 5701
rect 12069 5692 12081 5695
rect 12032 5664 12081 5692
rect 12032 5652 12038 5664
rect 12069 5661 12081 5664
rect 12115 5692 12127 5695
rect 12176 5692 12204 5868
rect 13740 5837 13768 5868
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5828 13783 5831
rect 15194 5828 15200 5840
rect 13771 5800 15200 5828
rect 13771 5797 13783 5800
rect 13725 5791 13783 5797
rect 15194 5788 15200 5800
rect 15252 5788 15258 5840
rect 12115 5664 12204 5692
rect 12345 5695 12403 5701
rect 12115 5661 12127 5664
rect 12069 5655 12127 5661
rect 12345 5661 12357 5695
rect 12391 5692 12403 5695
rect 13078 5692 13084 5704
rect 12391 5664 13084 5692
rect 12391 5661 12403 5664
rect 12345 5655 12403 5661
rect 13078 5652 13084 5664
rect 13136 5652 13142 5704
rect 16206 5652 16212 5704
rect 16264 5652 16270 5704
rect 8720 5596 9536 5624
rect 8720 5584 8726 5596
rect 8938 5556 8944 5568
rect 8404 5528 8944 5556
rect 8938 5516 8944 5528
rect 8996 5516 9002 5568
rect 9508 5556 9536 5596
rect 9950 5584 9956 5636
rect 10008 5624 10014 5636
rect 10137 5627 10195 5633
rect 10137 5624 10149 5627
rect 10008 5596 10149 5624
rect 10008 5584 10014 5596
rect 10137 5593 10149 5596
rect 10183 5624 10195 5627
rect 10226 5624 10232 5636
rect 10183 5596 10232 5624
rect 10183 5593 10195 5596
rect 10137 5587 10195 5593
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 10410 5584 10416 5636
rect 10468 5624 10474 5636
rect 10658 5627 10716 5633
rect 10658 5624 10670 5627
rect 10468 5596 10670 5624
rect 10468 5584 10474 5596
rect 10658 5593 10670 5596
rect 10704 5593 10716 5627
rect 10658 5587 10716 5593
rect 12253 5627 12311 5633
rect 12253 5593 12265 5627
rect 12299 5624 12311 5627
rect 12612 5627 12670 5633
rect 12299 5596 12572 5624
rect 12299 5593 12311 5596
rect 12253 5587 12311 5593
rect 10502 5556 10508 5568
rect 9508 5528 10508 5556
rect 10502 5516 10508 5528
rect 10560 5516 10566 5568
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 11793 5559 11851 5565
rect 11793 5556 11805 5559
rect 11112 5528 11805 5556
rect 11112 5516 11118 5528
rect 11793 5525 11805 5528
rect 11839 5525 11851 5559
rect 11793 5519 11851 5525
rect 11885 5559 11943 5565
rect 11885 5525 11897 5559
rect 11931 5556 11943 5559
rect 12434 5556 12440 5568
rect 11931 5528 12440 5556
rect 11931 5525 11943 5528
rect 11885 5519 11943 5525
rect 12434 5516 12440 5528
rect 12492 5516 12498 5568
rect 12544 5556 12572 5596
rect 12612 5593 12624 5627
rect 12658 5624 12670 5627
rect 12986 5624 12992 5636
rect 12658 5596 12992 5624
rect 12658 5593 12670 5596
rect 12612 5587 12670 5593
rect 12986 5584 12992 5596
rect 13044 5584 13050 5636
rect 13446 5584 13452 5636
rect 13504 5624 13510 5636
rect 14185 5627 14243 5633
rect 14185 5624 14197 5627
rect 13504 5596 14197 5624
rect 13504 5584 13510 5596
rect 14185 5593 14197 5596
rect 14231 5593 14243 5627
rect 14185 5587 14243 5593
rect 14366 5584 14372 5636
rect 14424 5584 14430 5636
rect 13464 5556 13492 5584
rect 12544 5528 13492 5556
rect 14550 5516 14556 5568
rect 14608 5516 14614 5568
rect 16393 5559 16451 5565
rect 16393 5525 16405 5559
rect 16439 5556 16451 5559
rect 16574 5556 16580 5568
rect 16439 5528 16580 5556
rect 16439 5525 16451 5528
rect 16393 5519 16451 5525
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 1104 5466 16836 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 16836 5466
rect 1104 5392 16836 5414
rect 2314 5352 2320 5364
rect 1872 5324 2320 5352
rect 1872 5284 1900 5324
rect 2314 5312 2320 5324
rect 2372 5312 2378 5364
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 3697 5355 3755 5361
rect 3697 5352 3709 5355
rect 3292 5324 3709 5352
rect 3292 5312 3298 5324
rect 3697 5321 3709 5324
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 3878 5312 3884 5364
rect 3936 5352 3942 5364
rect 8018 5352 8024 5364
rect 3936 5324 8024 5352
rect 3936 5312 3942 5324
rect 1780 5256 1900 5284
rect 2492 5287 2550 5293
rect 1780 5225 1808 5256
rect 2492 5253 2504 5287
rect 2538 5284 2550 5287
rect 2774 5284 2780 5296
rect 2538 5256 2780 5284
rect 2538 5253 2550 5256
rect 2492 5247 2550 5253
rect 2774 5244 2780 5256
rect 2832 5244 2838 5296
rect 1765 5219 1823 5225
rect 1765 5185 1777 5219
rect 1811 5185 1823 5219
rect 1765 5179 1823 5185
rect 1854 5176 1860 5228
rect 1912 5176 1918 5228
rect 1946 5176 1952 5228
rect 2004 5176 2010 5228
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2424 5216 2544 5219
rect 3510 5216 3516 5228
rect 2179 5191 3516 5216
rect 2179 5188 2452 5191
rect 2516 5188 3516 5191
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 3881 5219 3939 5225
rect 3881 5216 3893 5219
rect 3620 5188 3893 5216
rect 2038 5108 2044 5160
rect 2096 5148 2102 5160
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 2096 5120 2237 5148
rect 2096 5108 2102 5120
rect 2225 5117 2237 5120
rect 2271 5117 2283 5151
rect 2225 5111 2283 5117
rect 1486 4972 1492 5024
rect 1544 4972 1550 5024
rect 2958 4972 2964 5024
rect 3016 5012 3022 5024
rect 3620 5021 3648 5188
rect 3881 5185 3893 5188
rect 3927 5185 3939 5219
rect 3881 5179 3939 5185
rect 4062 5176 4068 5228
rect 4120 5176 4126 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5185 4583 5219
rect 4525 5179 4583 5185
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5185 4675 5219
rect 4617 5179 4675 5185
rect 4540 5080 4568 5179
rect 4632 5148 4660 5179
rect 4706 5176 4712 5228
rect 4764 5176 4770 5228
rect 4908 5225 4936 5324
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8588 5324 11284 5352
rect 6181 5287 6239 5293
rect 6181 5284 6193 5287
rect 5276 5256 6193 5284
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5185 4951 5219
rect 4893 5179 4951 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5216 5135 5219
rect 5166 5216 5172 5228
rect 5123 5188 5172 5216
rect 5123 5185 5135 5188
rect 5077 5179 5135 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 5276 5225 5304 5256
rect 6181 5253 6193 5256
rect 6227 5253 6239 5287
rect 6181 5247 6239 5253
rect 6822 5244 6828 5296
rect 6880 5284 6886 5296
rect 8588 5284 8616 5324
rect 10134 5284 10140 5296
rect 6880 5256 8616 5284
rect 8680 5256 10140 5284
rect 6880 5244 6886 5256
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5185 5319 5219
rect 5261 5179 5319 5185
rect 5350 5176 5356 5228
rect 5408 5176 5414 5228
rect 5445 5219 5503 5225
rect 5445 5185 5457 5219
rect 5491 5216 5503 5219
rect 5534 5216 5540 5228
rect 5491 5188 5540 5216
rect 5491 5185 5503 5188
rect 5445 5179 5503 5185
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 5810 5176 5816 5228
rect 5868 5176 5874 5228
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 7006 5216 7012 5228
rect 6043 5188 7012 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7190 5225 7196 5228
rect 7184 5179 7196 5225
rect 7190 5176 7196 5179
rect 7248 5176 7254 5228
rect 8680 5225 8708 5256
rect 10134 5244 10140 5256
rect 10192 5244 10198 5296
rect 8938 5225 8944 5228
rect 8665 5219 8723 5225
rect 8665 5185 8677 5219
rect 8711 5185 8723 5219
rect 8665 5179 8723 5185
rect 8932 5179 8944 5225
rect 8938 5176 8944 5179
rect 8996 5176 9002 5228
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 10520 5225 10548 5324
rect 10965 5287 11023 5293
rect 10965 5284 10977 5287
rect 10704 5256 10977 5284
rect 10505 5219 10563 5225
rect 9272 5188 9720 5216
rect 9272 5176 9278 5188
rect 5368 5148 5396 5176
rect 9692 5160 9720 5188
rect 10505 5185 10517 5219
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 10594 5176 10600 5228
rect 10652 5176 10658 5228
rect 10704 5225 10732 5256
rect 10965 5253 10977 5256
rect 11011 5253 11023 5287
rect 11256 5284 11284 5324
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 11701 5355 11759 5361
rect 11701 5352 11713 5355
rect 11388 5324 11713 5352
rect 11388 5312 11394 5324
rect 11701 5321 11713 5324
rect 11747 5321 11759 5355
rect 12342 5352 12348 5364
rect 11701 5315 11759 5321
rect 11900 5324 12348 5352
rect 11900 5284 11928 5324
rect 12342 5312 12348 5324
rect 12400 5312 12406 5364
rect 12986 5312 12992 5364
rect 13044 5312 13050 5364
rect 14366 5312 14372 5364
rect 14424 5352 14430 5364
rect 14921 5355 14979 5361
rect 14921 5352 14933 5355
rect 14424 5324 14933 5352
rect 14424 5312 14430 5324
rect 14921 5321 14933 5324
rect 14967 5352 14979 5355
rect 14967 5324 15332 5352
rect 14967 5321 14979 5324
rect 14921 5315 14979 5321
rect 11256 5256 11928 5284
rect 10965 5247 11023 5253
rect 11974 5244 11980 5296
rect 12032 5244 12038 5296
rect 12802 5284 12808 5296
rect 12636 5256 12808 5284
rect 10689 5219 10747 5225
rect 10689 5185 10701 5219
rect 10735 5185 10747 5219
rect 10689 5179 10747 5185
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 10873 5179 10931 5185
rect 6914 5148 6920 5160
rect 4632 5120 5396 5148
rect 5552 5120 6920 5148
rect 5552 5092 5580 5120
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10888 5148 10916 5179
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11149 5219 11207 5225
rect 11149 5216 11161 5219
rect 11112 5188 11161 5216
rect 11112 5176 11118 5188
rect 11149 5185 11161 5188
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 9732 5120 10916 5148
rect 11164 5148 11192 5179
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 11296 5188 11345 5216
rect 11296 5176 11302 5188
rect 11333 5185 11345 5188
rect 11379 5185 11391 5219
rect 11333 5179 11391 5185
rect 11882 5176 11888 5228
rect 11940 5176 11946 5228
rect 12066 5176 12072 5228
rect 12124 5176 12130 5228
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 12176 5188 12265 5216
rect 12176 5148 12204 5188
rect 12253 5185 12265 5188
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12360 5148 12388 5179
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12636 5225 12664 5256
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 13078 5244 13084 5296
rect 13136 5284 13142 5296
rect 15102 5284 15108 5296
rect 13136 5256 15108 5284
rect 13136 5244 13142 5256
rect 13556 5225 13584 5256
rect 15102 5244 15108 5256
rect 15160 5244 15166 5296
rect 15304 5293 15332 5324
rect 15289 5287 15347 5293
rect 15289 5253 15301 5287
rect 15335 5284 15347 5287
rect 15654 5284 15660 5296
rect 15335 5256 15660 5284
rect 15335 5253 15347 5256
rect 15289 5247 15347 5253
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 12529 5219 12587 5225
rect 12529 5216 12541 5219
rect 12492 5188 12541 5216
rect 12492 5176 12498 5188
rect 12529 5185 12541 5188
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 12621 5219 12679 5225
rect 12621 5185 12633 5219
rect 12667 5185 12679 5219
rect 12621 5179 12679 5185
rect 12713 5219 12771 5225
rect 12713 5185 12725 5219
rect 12759 5185 12771 5219
rect 12713 5179 12771 5185
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 13808 5219 13866 5225
rect 13808 5185 13820 5219
rect 13854 5216 13866 5219
rect 14090 5216 14096 5228
rect 13854 5188 14096 5216
rect 13854 5185 13866 5188
rect 13808 5179 13866 5185
rect 11164 5120 12204 5148
rect 12268 5120 12388 5148
rect 9732 5108 9738 5120
rect 4540 5052 4752 5080
rect 3605 5015 3663 5021
rect 3605 5012 3617 5015
rect 3016 4984 3617 5012
rect 3016 4972 3022 4984
rect 3605 4981 3617 4984
rect 3651 4981 3663 5015
rect 3605 4975 3663 4981
rect 4249 5015 4307 5021
rect 4249 4981 4261 5015
rect 4295 5012 4307 5015
rect 4614 5012 4620 5024
rect 4295 4984 4620 5012
rect 4295 4981 4307 4984
rect 4249 4975 4307 4981
rect 4614 4972 4620 4984
rect 4672 4972 4678 5024
rect 4724 5012 4752 5052
rect 5534 5040 5540 5092
rect 5592 5040 5598 5092
rect 5902 5080 5908 5092
rect 5644 5052 5908 5080
rect 5644 5012 5672 5052
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 10229 5083 10287 5089
rect 10229 5049 10241 5083
rect 10275 5080 10287 5083
rect 10410 5080 10416 5092
rect 10275 5052 10416 5080
rect 10275 5049 10287 5052
rect 10229 5043 10287 5049
rect 10410 5040 10416 5052
rect 10468 5040 10474 5092
rect 4724 4984 5672 5012
rect 5718 4972 5724 5024
rect 5776 4972 5782 5024
rect 7558 4972 7564 5024
rect 7616 5012 7622 5024
rect 8297 5015 8355 5021
rect 8297 5012 8309 5015
rect 7616 4984 8309 5012
rect 7616 4972 7622 4984
rect 8297 4981 8309 4984
rect 8343 4981 8355 5015
rect 8297 4975 8355 4981
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10045 5015 10103 5021
rect 10045 5012 10057 5015
rect 9640 4984 10057 5012
rect 9640 4972 9646 4984
rect 10045 4981 10057 4984
rect 10091 4981 10103 5015
rect 10888 5012 10916 5120
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 11882 5080 11888 5092
rect 11020 5052 11888 5080
rect 11020 5040 11026 5052
rect 11882 5040 11888 5052
rect 11940 5040 11946 5092
rect 12268 5012 12296 5120
rect 12342 5040 12348 5092
rect 12400 5080 12406 5092
rect 12728 5080 12756 5179
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 14182 5176 14188 5228
rect 14240 5216 14246 5228
rect 14240 5188 14688 5216
rect 14240 5176 14246 5188
rect 14660 5160 14688 5188
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 14976 5188 15209 5216
rect 14976 5176 14982 5188
rect 15197 5185 15209 5188
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 15381 5219 15439 5225
rect 15381 5185 15393 5219
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 15396 5148 15424 5179
rect 15562 5176 15568 5228
rect 15620 5176 15626 5228
rect 14700 5120 15424 5148
rect 14700 5108 14706 5120
rect 12400 5052 12756 5080
rect 12400 5040 12406 5052
rect 14734 5012 14740 5024
rect 10888 4984 14740 5012
rect 10045 4975 10103 4981
rect 14734 4972 14740 4984
rect 14792 4972 14798 5024
rect 15010 4972 15016 5024
rect 15068 4972 15074 5024
rect 1104 4922 16836 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 16836 4922
rect 1104 4848 16836 4870
rect 2130 4768 2136 4820
rect 2188 4808 2194 4820
rect 2777 4811 2835 4817
rect 2777 4808 2789 4811
rect 2188 4780 2789 4808
rect 2188 4768 2194 4780
rect 2777 4777 2789 4780
rect 2823 4777 2835 4811
rect 2777 4771 2835 4777
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 2038 4604 2044 4616
rect 1443 4576 2044 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 2792 4604 2820 4771
rect 3418 4768 3424 4820
rect 3476 4768 3482 4820
rect 3970 4768 3976 4820
rect 4028 4808 4034 4820
rect 6917 4811 6975 4817
rect 4028 4780 6868 4808
rect 4028 4768 4034 4780
rect 6840 4740 6868 4780
rect 6917 4777 6929 4811
rect 6963 4808 6975 4811
rect 7006 4808 7012 4820
rect 6963 4780 7012 4808
rect 6963 4777 6975 4780
rect 6917 4771 6975 4777
rect 7006 4768 7012 4780
rect 7064 4768 7070 4820
rect 7190 4768 7196 4820
rect 7248 4768 7254 4820
rect 7760 4780 12434 4808
rect 7760 4740 7788 4780
rect 6840 4712 7788 4740
rect 7834 4700 7840 4752
rect 7892 4700 7898 4752
rect 8938 4700 8944 4752
rect 8996 4700 9002 4752
rect 12406 4740 12434 4780
rect 14090 4768 14096 4820
rect 14148 4768 14154 4820
rect 15010 4740 15016 4752
rect 12406 4712 15016 4740
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 7852 4672 7880 4700
rect 8202 4672 8208 4684
rect 7576 4644 8208 4672
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2792 4576 2881 4604
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 2958 4564 2964 4616
rect 3016 4604 3022 4616
rect 3145 4607 3203 4613
rect 3145 4604 3157 4607
rect 3016 4576 3157 4604
rect 3016 4564 3022 4576
rect 3145 4573 3157 4576
rect 3191 4573 3203 4607
rect 3145 4567 3203 4573
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3510 4604 3516 4616
rect 3283 4576 3516 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3510 4564 3516 4576
rect 3568 4564 3574 4616
rect 4062 4564 4068 4616
rect 4120 4564 4126 4616
rect 4332 4607 4390 4613
rect 4332 4573 4344 4607
rect 4378 4604 4390 4607
rect 4614 4604 4620 4616
rect 4378 4576 4620 4604
rect 4378 4573 4390 4576
rect 4332 4567 4390 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5534 4564 5540 4616
rect 5592 4564 5598 4616
rect 7576 4613 7604 4644
rect 8202 4632 8208 4644
rect 8260 4672 8266 4684
rect 13262 4672 13268 4684
rect 8260 4644 13268 4672
rect 8260 4632 8266 4644
rect 5804 4607 5862 4613
rect 5804 4573 5816 4607
rect 5850 4573 5862 4607
rect 5804 4567 5862 4573
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7561 4607 7619 4613
rect 7561 4573 7573 4607
rect 7607 4573 7619 4607
rect 7561 4567 7619 4573
rect 1486 4496 1492 4548
rect 1544 4536 1550 4548
rect 1642 4539 1700 4545
rect 1642 4536 1654 4539
rect 1544 4508 1654 4536
rect 1544 4496 1550 4508
rect 1642 4505 1654 4508
rect 1688 4505 1700 4539
rect 3053 4539 3111 4545
rect 3053 4536 3065 4539
rect 1642 4499 1700 4505
rect 2884 4508 3065 4536
rect 2884 4480 2912 4508
rect 3053 4505 3065 4508
rect 3099 4505 3111 4539
rect 3053 4499 3111 4505
rect 5718 4496 5724 4548
rect 5776 4536 5782 4548
rect 5828 4536 5856 4567
rect 5776 4508 5856 4536
rect 5776 4496 5782 4508
rect 5902 4496 5908 4548
rect 5960 4536 5966 4548
rect 6822 4536 6828 4548
rect 5960 4508 6828 4536
rect 5960 4496 5966 4508
rect 6822 4496 6828 4508
rect 6880 4536 6886 4548
rect 7484 4536 7512 4567
rect 7650 4564 7656 4616
rect 7708 4564 7714 4616
rect 7837 4607 7895 4613
rect 7837 4573 7849 4607
rect 7883 4604 7895 4607
rect 8018 4604 8024 4616
rect 7883 4576 8024 4604
rect 7883 4573 7895 4576
rect 7837 4567 7895 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 9214 4604 9220 4616
rect 8496 4576 9220 4604
rect 6880 4508 7512 4536
rect 6880 4496 6886 4508
rect 8386 4496 8392 4548
rect 8444 4496 8450 4548
rect 2866 4428 2872 4480
rect 2924 4428 2930 4480
rect 4614 4428 4620 4480
rect 4672 4468 4678 4480
rect 5445 4471 5503 4477
rect 5445 4468 5457 4471
rect 4672 4440 5457 4468
rect 4672 4428 4678 4440
rect 5445 4437 5457 4440
rect 5491 4437 5503 4471
rect 5445 4431 5503 4437
rect 5626 4428 5632 4480
rect 5684 4468 5690 4480
rect 8496 4468 8524 4576
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9324 4613 9352 4644
rect 13262 4632 13268 4644
rect 13320 4672 13326 4684
rect 13320 4644 14044 4672
rect 13320 4632 13326 4644
rect 9309 4607 9367 4613
rect 9309 4573 9321 4607
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 9585 4607 9643 4613
rect 9585 4573 9597 4607
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 10321 4607 10379 4613
rect 10321 4573 10333 4607
rect 10367 4604 10379 4607
rect 12158 4604 12164 4616
rect 10367 4576 12164 4604
rect 10367 4573 10379 4576
rect 10321 4567 10379 4573
rect 8573 4539 8631 4545
rect 8573 4505 8585 4539
rect 8619 4505 8631 4539
rect 8573 4499 8631 4505
rect 8757 4539 8815 4545
rect 8757 4505 8769 4539
rect 8803 4536 8815 4539
rect 9416 4536 9444 4567
rect 8803 4508 9444 4536
rect 8803 4505 8815 4508
rect 8757 4499 8815 4505
rect 5684 4440 8524 4468
rect 8588 4468 8616 4499
rect 9600 4480 9628 4567
rect 12158 4564 12164 4576
rect 12216 4564 12222 4616
rect 13541 4607 13599 4613
rect 13541 4604 13553 4607
rect 12406 4576 13553 4604
rect 9674 4496 9680 4548
rect 9732 4536 9738 4548
rect 12406 4536 12434 4576
rect 13541 4573 13553 4576
rect 13587 4604 13599 4607
rect 13906 4604 13912 4616
rect 13587 4576 13912 4604
rect 13587 4573 13599 4576
rect 13541 4567 13599 4573
rect 13906 4564 13912 4576
rect 13964 4564 13970 4616
rect 14016 4604 14044 4644
rect 14090 4632 14096 4684
rect 14148 4672 14154 4684
rect 14148 4644 14504 4672
rect 14148 4632 14154 4644
rect 14274 4604 14280 4616
rect 14016 4576 14280 4604
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14366 4564 14372 4616
rect 14424 4564 14430 4616
rect 14476 4613 14504 4644
rect 14642 4632 14648 4684
rect 14700 4672 14706 4684
rect 15102 4672 15108 4684
rect 14700 4644 15108 4672
rect 14700 4632 14706 4644
rect 15102 4632 15108 4644
rect 15160 4632 15166 4684
rect 14461 4607 14519 4613
rect 14461 4573 14473 4607
rect 14507 4573 14519 4607
rect 14461 4567 14519 4573
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14734 4564 14740 4616
rect 14792 4564 14798 4616
rect 9732 4508 12434 4536
rect 13725 4539 13783 4545
rect 9732 4496 9738 4508
rect 13725 4505 13737 4539
rect 13771 4536 13783 4539
rect 13771 4508 15056 4536
rect 13771 4505 13783 4508
rect 13725 4499 13783 4505
rect 8846 4468 8852 4480
rect 8588 4440 8852 4468
rect 5684 4428 5690 4440
rect 8846 4428 8852 4440
rect 8904 4468 8910 4480
rect 9490 4468 9496 4480
rect 8904 4440 9496 4468
rect 8904 4428 8910 4440
rect 9490 4428 9496 4440
rect 9548 4428 9554 4480
rect 9582 4428 9588 4480
rect 9640 4468 9646 4480
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 9640 4440 10149 4468
rect 9640 4428 9646 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 13909 4471 13967 4477
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 14550 4468 14556 4480
rect 13955 4440 14556 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 14550 4428 14556 4440
rect 14608 4428 14614 4480
rect 15028 4468 15056 4508
rect 15102 4496 15108 4548
rect 15160 4536 15166 4548
rect 15350 4539 15408 4545
rect 15350 4536 15362 4539
rect 15160 4508 15362 4536
rect 15160 4496 15166 4508
rect 15350 4505 15362 4508
rect 15396 4505 15408 4539
rect 15350 4499 15408 4505
rect 15562 4468 15568 4480
rect 15028 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4468 15626 4480
rect 16482 4468 16488 4480
rect 15620 4440 16488 4468
rect 15620 4428 15626 4440
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 1104 4378 16836 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 16836 4378
rect 1104 4304 16836 4326
rect 4525 4267 4583 4273
rect 4525 4233 4537 4267
rect 4571 4264 4583 4267
rect 4706 4264 4712 4276
rect 4571 4236 4712 4264
rect 4571 4233 4583 4236
rect 4525 4227 4583 4233
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 7190 4224 7196 4276
rect 7248 4264 7254 4276
rect 7248 4236 7972 4264
rect 7248 4224 7254 4236
rect 2866 4156 2872 4208
rect 2924 4196 2930 4208
rect 3145 4199 3203 4205
rect 3145 4196 3157 4199
rect 2924 4168 3157 4196
rect 2924 4156 2930 4168
rect 3145 4165 3157 4168
rect 3191 4165 3203 4199
rect 3145 4159 3203 4165
rect 3970 4156 3976 4208
rect 4028 4196 4034 4208
rect 4157 4199 4215 4205
rect 4157 4196 4169 4199
rect 4028 4168 4169 4196
rect 4028 4156 4034 4168
rect 4157 4165 4169 4168
rect 4203 4165 4215 4199
rect 4157 4159 4215 4165
rect 4341 4199 4399 4205
rect 4341 4165 4353 4199
rect 4387 4196 4399 4199
rect 4614 4196 4620 4208
rect 4387 4168 4620 4196
rect 4387 4165 4399 4168
rect 4341 4159 4399 4165
rect 4614 4156 4620 4168
rect 4672 4156 4678 4208
rect 6546 4156 6552 4208
rect 6604 4196 6610 4208
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 6604 4168 6929 4196
rect 6604 4156 6610 4168
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 7558 4196 7564 4208
rect 6917 4159 6975 4165
rect 7024 4168 7564 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 1688 3992 1716 4091
rect 2130 4088 2136 4140
rect 2188 4128 2194 4140
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 2188 4100 2329 4128
rect 2188 4088 2194 4100
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2685 4131 2743 4137
rect 2685 4097 2697 4131
rect 2731 4128 2743 4131
rect 2774 4128 2780 4140
rect 2731 4100 2780 4128
rect 2731 4097 2743 4100
rect 2685 4091 2743 4097
rect 2774 4088 2780 4100
rect 2832 4128 2838 4140
rect 2961 4131 3019 4137
rect 2961 4128 2973 4131
rect 2832 4100 2973 4128
rect 2832 4088 2838 4100
rect 2961 4097 2973 4100
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4128 3387 4131
rect 3510 4128 3516 4140
rect 3375 4100 3516 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 3252 4060 3280 4091
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3605 4131 3663 4137
rect 3605 4097 3617 4131
rect 3651 4128 3663 4131
rect 3694 4128 3700 4140
rect 3651 4100 3700 4128
rect 3651 4097 3663 4100
rect 3605 4091 3663 4097
rect 3620 4060 3648 4091
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 4632 4128 4660 4156
rect 7024 4137 7052 4168
rect 7558 4156 7564 4168
rect 7616 4156 7622 4208
rect 7834 4156 7840 4208
rect 7892 4156 7898 4208
rect 7944 4196 7972 4236
rect 8386 4224 8392 4276
rect 8444 4264 8450 4276
rect 9674 4264 9680 4276
rect 8444 4236 9680 4264
rect 8444 4224 8450 4236
rect 9674 4224 9680 4236
rect 9732 4224 9738 4276
rect 11606 4224 11612 4276
rect 11664 4264 11670 4276
rect 12802 4264 12808 4276
rect 11664 4236 12112 4264
rect 11664 4224 11670 4236
rect 8754 4196 8760 4208
rect 7944 4168 8760 4196
rect 6733 4131 6791 4137
rect 6733 4128 6745 4131
rect 4632 4100 6745 4128
rect 6733 4097 6745 4100
rect 6779 4097 6791 4131
rect 6733 4091 6791 4097
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4097 7067 4131
rect 7009 4091 7067 4097
rect 7101 4131 7159 4137
rect 7101 4097 7113 4131
rect 7147 4128 7159 4131
rect 7190 4128 7196 4140
rect 7147 4100 7196 4128
rect 7147 4097 7159 4100
rect 7101 4091 7159 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 8036 4137 8064 4168
rect 8754 4156 8760 4168
rect 8812 4156 8818 4208
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 11149 4199 11207 4205
rect 9640 4168 10916 4196
rect 9640 4156 9646 4168
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7929 4131 7987 4137
rect 7929 4097 7941 4131
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 8021 4131 8079 4137
rect 8021 4097 8033 4131
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 3252 4032 3648 4060
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7668 4060 7696 4091
rect 6880 4032 7696 4060
rect 7944 4060 7972 4091
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10100 4100 10517 4128
rect 10100 4088 10106 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10594 4088 10600 4140
rect 10652 4088 10658 4140
rect 10888 4137 10916 4168
rect 11149 4165 11161 4199
rect 11195 4196 11207 4199
rect 12084 4196 12112 4236
rect 12544 4236 12808 4264
rect 11195 4168 12020 4196
rect 12084 4168 12204 4196
rect 11195 4165 11207 4168
rect 11149 4159 11207 4165
rect 11992 4140 12020 4168
rect 10689 4131 10747 4137
rect 10689 4097 10701 4131
rect 10735 4097 10747 4131
rect 10689 4091 10747 4097
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 8294 4060 8300 4072
rect 7944 4032 8300 4060
rect 6880 4020 6886 4032
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10612 4060 10640 4088
rect 9824 4032 10640 4060
rect 10704 4060 10732 4091
rect 11238 4088 11244 4140
rect 11296 4128 11302 4140
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 11296 4100 11345 4128
rect 11296 4088 11302 4100
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 11698 4088 11704 4140
rect 11756 4088 11762 4140
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4097 11851 4131
rect 11793 4091 11851 4097
rect 10965 4063 11023 4069
rect 10965 4060 10977 4063
rect 10704 4032 10977 4060
rect 9824 4020 9830 4032
rect 10965 4029 10977 4032
rect 11011 4029 11023 4063
rect 11606 4060 11612 4072
rect 10965 4023 11023 4029
rect 11072 4032 11612 4060
rect 3142 3992 3148 4004
rect 1688 3964 3148 3992
rect 3142 3952 3148 3964
rect 3200 3952 3206 4004
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 3789 3995 3847 4001
rect 3789 3992 3801 3995
rect 3384 3964 3801 3992
rect 3384 3952 3390 3964
rect 3789 3961 3801 3964
rect 3835 3961 3847 3995
rect 3789 3955 3847 3961
rect 7282 3952 7288 4004
rect 7340 3952 7346 4004
rect 8205 3995 8263 4001
rect 8205 3961 8217 3995
rect 8251 3992 8263 3995
rect 8478 3992 8484 4004
rect 8251 3964 8484 3992
rect 8251 3961 8263 3964
rect 8205 3955 8263 3961
rect 8478 3952 8484 3964
rect 8536 3952 8542 4004
rect 9674 3952 9680 4004
rect 9732 3992 9738 4004
rect 11072 3992 11100 4032
rect 11606 4020 11612 4032
rect 11664 4020 11670 4072
rect 11808 4060 11836 4091
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 11974 4088 11980 4140
rect 12032 4128 12038 4140
rect 12069 4131 12127 4137
rect 12069 4128 12081 4131
rect 12032 4100 12081 4128
rect 12032 4088 12038 4100
rect 12069 4097 12081 4100
rect 12115 4097 12127 4131
rect 12176 4128 12204 4168
rect 12544 4137 12572 4236
rect 12802 4224 12808 4236
rect 12860 4264 12866 4276
rect 14090 4264 14096 4276
rect 12860 4236 14096 4264
rect 12860 4224 12866 4236
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 14274 4224 14280 4276
rect 14332 4224 14338 4276
rect 14366 4224 14372 4276
rect 14424 4264 14430 4276
rect 14424 4236 14872 4264
rect 14424 4224 14430 4236
rect 13265 4199 13323 4205
rect 13265 4165 13277 4199
rect 13311 4196 13323 4199
rect 13446 4196 13452 4208
rect 13311 4168 13452 4196
rect 13311 4165 13323 4168
rect 13265 4159 13323 4165
rect 13446 4156 13452 4168
rect 13504 4156 13510 4208
rect 13538 4156 13544 4208
rect 13596 4196 13602 4208
rect 14292 4196 14320 4224
rect 14844 4196 14872 4236
rect 14918 4196 14924 4208
rect 13596 4168 14044 4196
rect 14292 4168 14780 4196
rect 13596 4156 13602 4168
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 12176 4100 12449 4128
rect 12069 4091 12127 4097
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 12437 4091 12495 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4128 12863 4131
rect 12851 4100 13032 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 12250 4060 12256 4072
rect 11808 4032 12256 4060
rect 12250 4020 12256 4032
rect 12308 4020 12314 4072
rect 12636 4060 12664 4091
rect 12897 4063 12955 4069
rect 12897 4060 12909 4063
rect 12636 4032 12909 4060
rect 12897 4029 12909 4032
rect 12943 4029 12955 4063
rect 13004 4060 13032 4100
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 13814 4128 13820 4140
rect 13188 4100 13820 4128
rect 13188 4060 13216 4100
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14016 4137 14044 4168
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4097 14059 4131
rect 14001 4091 14059 4097
rect 14093 4131 14151 4137
rect 14093 4097 14105 4131
rect 14139 4097 14151 4131
rect 14093 4091 14151 4097
rect 13004 4032 13216 4060
rect 14108 4060 14136 4091
rect 14182 4088 14188 4140
rect 14240 4088 14246 4140
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 14369 4131 14427 4137
rect 14369 4128 14381 4131
rect 14332 4100 14381 4128
rect 14332 4088 14338 4100
rect 14369 4097 14381 4100
rect 14415 4097 14427 4131
rect 14369 4091 14427 4097
rect 14458 4088 14464 4140
rect 14516 4088 14522 4140
rect 14550 4088 14556 4140
rect 14608 4128 14614 4140
rect 14752 4137 14780 4168
rect 14844 4168 14924 4196
rect 14844 4137 14872 4168
rect 14918 4156 14924 4168
rect 14976 4156 14982 4208
rect 14645 4131 14703 4137
rect 14645 4128 14657 4131
rect 14608 4100 14657 4128
rect 14608 4088 14614 4100
rect 14645 4097 14657 4100
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14737 4131 14795 4137
rect 14737 4097 14749 4131
rect 14783 4097 14795 4131
rect 14737 4091 14795 4097
rect 14829 4131 14887 4137
rect 14829 4097 14841 4131
rect 14875 4097 14887 4131
rect 15473 4131 15531 4137
rect 15473 4128 15485 4131
rect 14829 4091 14887 4097
rect 14927 4100 15485 4128
rect 14927 4060 14955 4100
rect 15473 4097 15485 4100
rect 15519 4128 15531 4131
rect 15562 4128 15568 4140
rect 15519 4100 15568 4128
rect 15519 4097 15531 4100
rect 15473 4091 15531 4097
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 15838 4088 15844 4140
rect 15896 4088 15902 4140
rect 16482 4088 16488 4140
rect 16540 4088 16546 4140
rect 14108 4032 14955 4060
rect 12897 4023 12955 4029
rect 15102 4020 15108 4072
rect 15160 4020 15166 4072
rect 17402 4060 17408 4072
rect 15672 4032 17408 4060
rect 9732 3964 11100 3992
rect 9732 3952 9738 3964
rect 11514 3952 11520 4004
rect 11572 3952 11578 4004
rect 12526 3952 12532 4004
rect 12584 3992 12590 4004
rect 15672 4001 15700 4032
rect 17402 4020 17408 4032
rect 17460 4020 17466 4072
rect 13817 3995 13875 4001
rect 13817 3992 13829 3995
rect 12584 3964 13829 3992
rect 12584 3952 12590 3964
rect 13817 3961 13829 3964
rect 13863 3961 13875 3995
rect 13817 3955 13875 3961
rect 15657 3995 15715 4001
rect 15657 3961 15669 3995
rect 15703 3961 15715 3995
rect 15657 3955 15715 3961
rect 16025 3995 16083 4001
rect 16025 3961 16037 3995
rect 16071 3992 16083 3995
rect 16758 3992 16764 4004
rect 16071 3964 16764 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16758 3952 16764 3964
rect 16816 3952 16822 4004
rect 1394 3884 1400 3936
rect 1452 3924 1458 3936
rect 1489 3927 1547 3933
rect 1489 3924 1501 3927
rect 1452 3896 1501 3924
rect 1452 3884 1458 3896
rect 1489 3893 1501 3896
rect 1535 3893 1547 3927
rect 1489 3887 1547 3893
rect 2130 3884 2136 3936
rect 2188 3884 2194 3936
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 2372 3896 2513 3924
rect 2372 3884 2378 3896
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 3418 3884 3424 3936
rect 3476 3924 3482 3936
rect 3513 3927 3571 3933
rect 3513 3924 3525 3927
rect 3476 3896 3525 3924
rect 3476 3884 3482 3896
rect 3513 3893 3525 3896
rect 3559 3893 3571 3927
rect 3513 3887 3571 3893
rect 10226 3884 10232 3936
rect 10284 3884 10290 3936
rect 11882 3884 11888 3936
rect 11940 3924 11946 3936
rect 12161 3927 12219 3933
rect 12161 3924 12173 3927
rect 11940 3896 12173 3924
rect 11940 3884 11946 3896
rect 12161 3893 12173 3896
rect 12207 3893 12219 3927
rect 12161 3887 12219 3893
rect 14090 3884 14096 3936
rect 14148 3924 14154 3936
rect 14458 3924 14464 3936
rect 14148 3896 14464 3924
rect 14148 3884 14154 3896
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16301 3927 16359 3933
rect 16301 3924 16313 3927
rect 16172 3896 16313 3924
rect 16172 3884 16178 3896
rect 16301 3893 16313 3896
rect 16347 3893 16359 3927
rect 16301 3887 16359 3893
rect 1104 3834 16836 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 16836 3834
rect 1104 3760 16836 3782
rect 3602 3680 3608 3732
rect 3660 3720 3666 3732
rect 6733 3723 6791 3729
rect 3660 3692 6684 3720
rect 3660 3680 3666 3692
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 3108 3624 3188 3652
rect 3108 3612 3114 3624
rect 2406 3584 2412 3596
rect 1780 3556 2412 3584
rect 1780 3525 1808 3556
rect 2406 3544 2412 3556
rect 2464 3584 2470 3596
rect 3160 3584 3188 3624
rect 6656 3584 6684 3692
rect 6733 3689 6745 3723
rect 6779 3720 6791 3723
rect 6822 3720 6828 3732
rect 6779 3692 6828 3720
rect 6779 3689 6791 3692
rect 6733 3683 6791 3689
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 10042 3720 10048 3732
rect 7340 3692 10048 3720
rect 7340 3680 7346 3692
rect 10042 3680 10048 3692
rect 10100 3680 10106 3732
rect 12342 3720 12348 3732
rect 10152 3692 12348 3720
rect 10152 3652 10180 3692
rect 12342 3680 12348 3692
rect 12400 3680 12406 3732
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13078 3720 13084 3732
rect 13035 3692 13084 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 13412 3692 15240 3720
rect 13412 3680 13418 3692
rect 7300 3624 10180 3652
rect 7300 3584 7328 3624
rect 14366 3612 14372 3664
rect 14424 3612 14430 3664
rect 15212 3652 15240 3692
rect 15212 3624 15332 3652
rect 8202 3584 8208 3596
rect 2464 3556 3096 3584
rect 2464 3544 2470 3556
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3485 1823 3519
rect 1765 3479 1823 3485
rect 1854 3476 1860 3528
rect 1912 3476 1918 3528
rect 1946 3476 1952 3528
rect 2004 3476 2010 3528
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3485 2191 3519
rect 2133 3479 2191 3485
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 2958 3516 2964 3528
rect 2731 3488 2964 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 2148 3448 2176 3479
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3068 3525 3096 3556
rect 3160 3556 4936 3584
rect 6656 3556 7328 3584
rect 7392 3556 8208 3584
rect 3160 3525 3188 3556
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3234 3476 3240 3528
rect 3292 3476 3298 3528
rect 3421 3519 3479 3525
rect 3421 3485 3433 3519
rect 3467 3516 3479 3519
rect 3878 3516 3884 3528
rect 3467 3488 3884 3516
rect 3467 3485 3479 3488
rect 3421 3479 3479 3485
rect 3436 3448 3464 3479
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 4172 3525 4200 3556
rect 4065 3519 4123 3525
rect 4065 3485 4077 3519
rect 4111 3485 4123 3519
rect 4065 3479 4123 3485
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 2148 3420 3464 3448
rect 1486 3340 1492 3392
rect 1544 3340 1550 3392
rect 2498 3340 2504 3392
rect 2556 3340 2562 3392
rect 2590 3340 2596 3392
rect 2648 3380 2654 3392
rect 2777 3383 2835 3389
rect 2777 3380 2789 3383
rect 2648 3352 2789 3380
rect 2648 3340 2654 3352
rect 2777 3349 2789 3352
rect 2823 3349 2835 3383
rect 4080 3380 4108 3479
rect 4246 3476 4252 3528
rect 4304 3476 4310 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 4632 3448 4660 3479
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 4908 3525 4936 3556
rect 4893 3519 4951 3525
rect 4893 3485 4905 3519
rect 4939 3485 4951 3519
rect 4893 3479 4951 3485
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3516 5411 3519
rect 5442 3516 5448 3528
rect 5399 3488 5448 3516
rect 5399 3485 5411 3488
rect 5353 3479 5411 3485
rect 5442 3476 5448 3488
rect 5500 3476 5506 3528
rect 7282 3476 7288 3528
rect 7340 3476 7346 3528
rect 7392 3525 7420 3556
rect 8202 3544 8208 3556
rect 8260 3584 8266 3596
rect 8260 3556 8524 3584
rect 8260 3544 8266 3556
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3485 7435 3519
rect 7377 3479 7435 3485
rect 7466 3476 7472 3528
rect 7524 3476 7530 3528
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3516 7711 3519
rect 8018 3516 8024 3528
rect 7699 3488 8024 3516
rect 7699 3485 7711 3488
rect 7653 3479 7711 3485
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 8496 3525 8524 3556
rect 8680 3556 9720 3584
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 5166 3448 5172 3460
rect 4632 3420 5172 3448
rect 5166 3408 5172 3420
rect 5224 3408 5230 3460
rect 5261 3451 5319 3457
rect 5261 3417 5273 3451
rect 5307 3448 5319 3451
rect 5598 3451 5656 3457
rect 5598 3448 5610 3451
rect 5307 3420 5610 3448
rect 5307 3417 5319 3420
rect 5261 3411 5319 3417
rect 5598 3417 5610 3420
rect 5644 3417 5656 3451
rect 8404 3448 8432 3479
rect 8570 3476 8576 3528
rect 8628 3476 8634 3528
rect 8680 3448 8708 3556
rect 9692 3528 9720 3556
rect 13262 3544 13268 3596
rect 13320 3584 13326 3596
rect 13814 3584 13820 3596
rect 13320 3556 13492 3584
rect 13320 3544 13326 3556
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 5598 3411 5656 3417
rect 5736 3420 8708 3448
rect 8772 3448 8800 3479
rect 9582 3476 9588 3528
rect 9640 3476 9646 3528
rect 9674 3476 9680 3528
rect 9732 3476 9738 3528
rect 9766 3476 9772 3528
rect 9824 3476 9830 3528
rect 9858 3476 9864 3528
rect 9916 3476 9922 3528
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 9600 3448 9628 3476
rect 10060 3448 10088 3479
rect 10134 3476 10140 3528
rect 10192 3476 10198 3528
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10393 3519 10451 3525
rect 10393 3516 10405 3519
rect 10284 3488 10405 3516
rect 10284 3476 10290 3488
rect 10393 3485 10405 3488
rect 10439 3485 10451 3519
rect 10393 3479 10451 3485
rect 11609 3519 11667 3525
rect 11609 3485 11621 3519
rect 11655 3516 11667 3519
rect 12434 3516 12440 3528
rect 11655 3488 12440 3516
rect 11655 3485 11667 3488
rect 11609 3479 11667 3485
rect 12434 3476 12440 3488
rect 12492 3476 12498 3528
rect 13354 3476 13360 3528
rect 13412 3476 13418 3528
rect 13464 3525 13492 3556
rect 13740 3556 13820 3584
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13538 3476 13544 3528
rect 13596 3476 13602 3528
rect 13740 3525 13768 3556
rect 13814 3544 13820 3556
rect 13872 3584 13878 3596
rect 14384 3584 14412 3612
rect 13872 3556 14412 3584
rect 14479 3556 15240 3584
rect 13872 3544 13878 3556
rect 14479 3528 14507 3556
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 14182 3476 14188 3528
rect 14240 3476 14246 3528
rect 14366 3476 14372 3528
rect 14424 3476 14430 3528
rect 14458 3476 14464 3528
rect 14516 3476 14522 3528
rect 14550 3476 14556 3528
rect 14608 3476 14614 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 15212 3525 15240 3556
rect 15304 3525 15332 3624
rect 15470 3612 15476 3664
rect 15528 3652 15534 3664
rect 16209 3655 16267 3661
rect 16209 3652 16221 3655
rect 15528 3624 16221 3652
rect 15528 3612 15534 3624
rect 16209 3621 16221 3624
rect 16255 3621 16267 3655
rect 16209 3615 16267 3621
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14792 3488 14933 3516
rect 14792 3476 14798 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 15105 3516 15163 3522
rect 15105 3482 15117 3516
rect 15151 3482 15163 3516
rect 15105 3476 15163 3482
rect 15197 3519 15255 3525
rect 15197 3485 15209 3519
rect 15243 3485 15255 3519
rect 15197 3479 15255 3485
rect 15289 3519 15347 3525
rect 15289 3485 15301 3519
rect 15335 3485 15347 3519
rect 15289 3479 15347 3485
rect 15654 3476 15660 3528
rect 15712 3476 15718 3528
rect 16022 3476 16028 3528
rect 16080 3476 16086 3528
rect 11882 3457 11888 3460
rect 11876 3448 11888 3457
rect 8772 3420 10088 3448
rect 11843 3420 11888 3448
rect 4154 3380 4160 3392
rect 4080 3352 4160 3380
rect 2777 3343 2835 3349
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4522 3340 4528 3392
rect 4580 3340 4586 3392
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 5736 3380 5764 3420
rect 11876 3411 11888 3420
rect 11882 3408 11888 3411
rect 11940 3408 11946 3460
rect 15120 3392 15148 3476
rect 5040 3352 5764 3380
rect 5040 3340 5046 3352
rect 7006 3340 7012 3392
rect 7064 3340 7070 3392
rect 8110 3340 8116 3392
rect 8168 3340 8174 3392
rect 9401 3383 9459 3389
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9582 3380 9588 3392
rect 9447 3352 9588 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 10042 3340 10048 3392
rect 10100 3380 10106 3392
rect 10962 3380 10968 3392
rect 10100 3352 10968 3380
rect 10100 3340 10106 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11517 3383 11575 3389
rect 11517 3349 11529 3383
rect 11563 3380 11575 3383
rect 11974 3380 11980 3392
rect 11563 3352 11980 3380
rect 11563 3349 11575 3352
rect 11517 3343 11575 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 13078 3340 13084 3392
rect 13136 3340 13142 3392
rect 14182 3340 14188 3392
rect 14240 3380 14246 3392
rect 14734 3380 14740 3392
rect 14240 3352 14740 3380
rect 14240 3340 14246 3352
rect 14734 3340 14740 3352
rect 14792 3340 14798 3392
rect 14829 3383 14887 3389
rect 14829 3349 14841 3383
rect 14875 3380 14887 3383
rect 14918 3380 14924 3392
rect 14875 3352 14924 3380
rect 14875 3349 14887 3352
rect 14829 3343 14887 3349
rect 14918 3340 14924 3352
rect 14976 3340 14982 3392
rect 15102 3340 15108 3392
rect 15160 3340 15166 3392
rect 15378 3340 15384 3392
rect 15436 3380 15442 3392
rect 15565 3383 15623 3389
rect 15565 3380 15577 3383
rect 15436 3352 15577 3380
rect 15436 3340 15442 3352
rect 15565 3349 15577 3352
rect 15611 3349 15623 3383
rect 15565 3343 15623 3349
rect 15838 3340 15844 3392
rect 15896 3340 15902 3392
rect 1104 3290 16836 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 16836 3290
rect 1104 3216 16836 3238
rect 1946 3136 1952 3188
rect 2004 3136 2010 3188
rect 2774 3176 2780 3188
rect 2056 3148 2780 3176
rect 1581 3111 1639 3117
rect 1581 3077 1593 3111
rect 1627 3108 1639 3111
rect 1670 3108 1676 3120
rect 1627 3080 1676 3108
rect 1627 3077 1639 3080
rect 1581 3071 1639 3077
rect 1670 3068 1676 3080
rect 1728 3068 1734 3120
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 2056 3108 2084 3148
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 4154 3136 4160 3188
rect 4212 3136 4218 3188
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 5721 3179 5779 3185
rect 5721 3176 5733 3179
rect 4856 3148 5733 3176
rect 4856 3136 4862 3148
rect 5721 3145 5733 3148
rect 5767 3145 5779 3179
rect 5721 3139 5779 3145
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 9401 3179 9459 3185
rect 9401 3176 9413 3179
rect 8352 3148 9413 3176
rect 8352 3136 8358 3148
rect 9401 3145 9413 3148
rect 9447 3145 9459 3179
rect 9401 3139 9459 3145
rect 9858 3136 9864 3188
rect 9916 3176 9922 3188
rect 10965 3179 11023 3185
rect 10965 3176 10977 3179
rect 9916 3148 10977 3176
rect 9916 3136 9922 3148
rect 10965 3145 10977 3148
rect 11011 3145 11023 3179
rect 12986 3176 12992 3188
rect 10965 3139 11023 3145
rect 11808 3148 12992 3176
rect 4522 3117 4528 3120
rect 4516 3108 4528 3117
rect 1811 3080 2084 3108
rect 2148 3080 4108 3108
rect 4483 3080 4528 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 2038 3000 2044 3052
rect 2096 3040 2102 3052
rect 2148 3040 2176 3080
rect 4080 3052 4108 3080
rect 4516 3071 4528 3080
rect 4522 3068 4528 3071
rect 4580 3068 4586 3120
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 5905 3111 5963 3117
rect 5905 3108 5917 3111
rect 5500 3080 5917 3108
rect 5500 3068 5506 3080
rect 5905 3077 5917 3080
rect 5951 3108 5963 3111
rect 6822 3108 6828 3120
rect 5951 3080 6828 3108
rect 5951 3077 5963 3080
rect 5905 3071 5963 3077
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 7006 3068 7012 3120
rect 7064 3108 7070 3120
rect 7570 3111 7628 3117
rect 7570 3108 7582 3111
rect 7064 3080 7582 3108
rect 7064 3068 7070 3080
rect 7570 3077 7582 3080
rect 7616 3077 7628 3111
rect 10134 3108 10140 3120
rect 7570 3071 7628 3077
rect 8036 3080 10140 3108
rect 2222 3040 2228 3052
rect 2096 3012 2228 3040
rect 2096 3000 2102 3012
rect 2222 3000 2228 3012
rect 2280 3040 2286 3052
rect 2590 3049 2596 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2280 3012 2329 3040
rect 2280 3000 2286 3012
rect 2317 3009 2329 3012
rect 2363 3009 2375 3043
rect 2584 3040 2596 3049
rect 2551 3012 2596 3040
rect 2317 3003 2375 3009
rect 2584 3003 2596 3012
rect 2590 3000 2596 3003
rect 2648 3000 2654 3052
rect 3142 3000 3148 3052
rect 3200 3040 3206 3052
rect 3789 3043 3847 3049
rect 3200 3012 3740 3040
rect 3200 3000 3206 3012
rect 3712 2972 3740 3012
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 3878 3040 3884 3052
rect 3835 3012 3884 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 3878 3000 3884 3012
rect 3936 3000 3942 3052
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 3988 2972 4016 3003
rect 4062 3000 4068 3052
rect 4120 3040 4126 3052
rect 8036 3049 8064 3080
rect 4249 3043 4307 3049
rect 4249 3040 4261 3043
rect 4120 3012 4261 3040
rect 4120 3000 4126 3012
rect 4249 3009 4261 3012
rect 4295 3009 4307 3043
rect 6089 3043 6147 3049
rect 4249 3003 4307 3009
rect 4356 3012 5580 3040
rect 4356 2972 4384 3012
rect 3712 2944 4016 2972
rect 3694 2796 3700 2848
rect 3752 2796 3758 2848
rect 3988 2836 4016 2944
rect 4080 2944 4384 2972
rect 5552 2972 5580 3012
rect 6089 3009 6101 3043
rect 6135 3009 6147 3043
rect 6089 3003 6147 3009
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7883 3012 8033 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8021 3009 8033 3012
rect 8067 3009 8079 3043
rect 8021 3003 8079 3009
rect 5810 2972 5816 2984
rect 5552 2944 5816 2972
rect 4080 2916 4108 2944
rect 5810 2932 5816 2944
rect 5868 2972 5874 2984
rect 6104 2972 6132 3003
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 9508 3049 9536 3080
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 11808 3117 11836 3148
rect 12986 3136 12992 3148
rect 13044 3136 13050 3188
rect 13538 3136 13544 3188
rect 13596 3176 13602 3188
rect 14277 3179 14335 3185
rect 14277 3176 14289 3179
rect 13596 3148 14289 3176
rect 13596 3136 13602 3148
rect 14277 3145 14289 3148
rect 14323 3145 14335 3179
rect 14277 3139 14335 3145
rect 14458 3136 14464 3188
rect 14516 3176 14522 3188
rect 16022 3176 16028 3188
rect 14516 3148 16028 3176
rect 14516 3136 14522 3148
rect 16022 3136 16028 3148
rect 16080 3136 16086 3188
rect 11333 3111 11391 3117
rect 11333 3108 11345 3111
rect 11296 3080 11345 3108
rect 11296 3068 11302 3080
rect 11333 3077 11345 3080
rect 11379 3077 11391 3111
rect 11333 3071 11391 3077
rect 11793 3111 11851 3117
rect 11793 3077 11805 3111
rect 11839 3077 11851 3111
rect 11793 3071 11851 3077
rect 11882 3068 11888 3120
rect 11940 3068 11946 3120
rect 14642 3108 14648 3120
rect 12636 3080 14648 3108
rect 8277 3043 8335 3049
rect 8277 3040 8289 3043
rect 8168 3012 8289 3040
rect 8168 3000 8174 3012
rect 8277 3009 8289 3012
rect 8323 3009 8335 3043
rect 8277 3003 8335 3009
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3009 9551 3043
rect 9493 3003 9551 3009
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 9749 3043 9807 3049
rect 9749 3040 9761 3043
rect 9640 3012 9761 3040
rect 9640 3000 9646 3012
rect 9749 3009 9761 3012
rect 9795 3009 9807 3043
rect 9749 3003 9807 3009
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11164 2972 11192 3003
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 12069 3043 12127 3049
rect 12069 3009 12081 3043
rect 12115 3009 12127 3043
rect 12636 3040 12664 3080
rect 14642 3068 14648 3080
rect 14700 3068 14706 3120
rect 12069 3003 12127 3009
rect 12544 3012 12664 3040
rect 12704 3043 12762 3049
rect 11422 2972 11428 2984
rect 5868 2944 6132 2972
rect 10888 2944 11428 2972
rect 5868 2932 5874 2944
rect 4062 2864 4068 2916
rect 4120 2864 4126 2916
rect 6546 2904 6552 2916
rect 5644 2876 6552 2904
rect 5644 2845 5672 2876
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 10888 2913 10916 2944
rect 11422 2932 11428 2944
rect 11480 2972 11486 2984
rect 12084 2972 12112 3003
rect 11480 2944 12112 2972
rect 11480 2932 11486 2944
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12544 2972 12572 3012
rect 12704 3009 12716 3043
rect 12750 3040 12762 3043
rect 13078 3040 13084 3052
rect 12750 3012 13084 3040
rect 12750 3009 12762 3012
rect 12704 3003 12762 3009
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13906 3000 13912 3052
rect 13964 3000 13970 3052
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3040 14151 3043
rect 14274 3040 14280 3052
rect 14139 3012 14280 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 12492 2944 12572 2972
rect 12492 2932 12498 2944
rect 10873 2907 10931 2913
rect 10873 2873 10885 2907
rect 10919 2873 10931 2907
rect 10873 2867 10931 2873
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 13817 2907 13875 2913
rect 11020 2876 12434 2904
rect 11020 2864 11026 2876
rect 5629 2839 5687 2845
rect 5629 2836 5641 2839
rect 3988 2808 5641 2836
rect 5629 2805 5641 2808
rect 5675 2805 5687 2839
rect 5629 2799 5687 2805
rect 6178 2796 6184 2848
rect 6236 2836 6242 2848
rect 6457 2839 6515 2845
rect 6457 2836 6469 2839
rect 6236 2808 6469 2836
rect 6236 2796 6242 2808
rect 6457 2805 6469 2808
rect 6503 2805 6515 2839
rect 6457 2799 6515 2805
rect 9122 2796 9128 2848
rect 9180 2836 9186 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 9180 2808 11529 2836
rect 9180 2796 9186 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 12406 2836 12434 2876
rect 13817 2873 13829 2907
rect 13863 2904 13875 2907
rect 13906 2904 13912 2916
rect 13863 2876 13912 2904
rect 13863 2873 13875 2876
rect 13817 2867 13875 2873
rect 13906 2864 13912 2876
rect 13964 2904 13970 2916
rect 14108 2904 14136 3003
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14918 3049 14924 3052
rect 14912 3040 14924 3049
rect 14879 3012 14924 3040
rect 14912 3003 14924 3012
rect 14918 3000 14924 3003
rect 14976 3000 14982 3052
rect 15194 3000 15200 3052
rect 15252 3040 15258 3052
rect 16117 3043 16175 3049
rect 16117 3040 16129 3043
rect 15252 3012 16129 3040
rect 15252 3000 15258 3012
rect 16117 3009 16129 3012
rect 16163 3009 16175 3043
rect 16117 3003 16175 3009
rect 14642 2932 14648 2984
rect 14700 2932 14706 2984
rect 13964 2876 14136 2904
rect 13964 2864 13970 2876
rect 14550 2836 14556 2848
rect 12406 2808 14556 2836
rect 11517 2799 11575 2805
rect 14550 2796 14556 2808
rect 14608 2796 14614 2848
rect 16298 2796 16304 2848
rect 16356 2796 16362 2848
rect 1104 2746 16836 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 16836 2746
rect 1104 2672 16836 2694
rect 2774 2592 2780 2644
rect 2832 2592 2838 2644
rect 3053 2635 3111 2641
rect 3053 2601 3065 2635
rect 3099 2632 3111 2635
rect 3234 2632 3240 2644
rect 3099 2604 3240 2632
rect 3099 2601 3111 2604
rect 3053 2595 3111 2601
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 6914 2632 6920 2644
rect 5092 2604 6920 2632
rect 1397 2431 1455 2437
rect 1397 2397 1409 2431
rect 1443 2428 1455 2431
rect 2222 2428 2228 2440
rect 1443 2400 2228 2428
rect 1443 2397 1455 2400
rect 1397 2391 1455 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3694 2428 3700 2440
rect 3283 2400 3700 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3694 2388 3700 2400
rect 3752 2388 3758 2440
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4614 2428 4620 2440
rect 4295 2400 4620 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4706 2388 4712 2440
rect 4764 2388 4770 2440
rect 5092 2437 5120 2604
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7524 2604 7573 2632
rect 7524 2592 7530 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 7561 2595 7619 2601
rect 8570 2592 8576 2644
rect 8628 2632 8634 2644
rect 8757 2635 8815 2641
rect 8757 2632 8769 2635
rect 8628 2604 8769 2632
rect 8628 2592 8634 2604
rect 8757 2601 8769 2604
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 14461 2635 14519 2641
rect 14461 2632 14473 2635
rect 14424 2604 14473 2632
rect 14424 2592 14430 2604
rect 14461 2601 14473 2604
rect 14507 2601 14519 2635
rect 14461 2595 14519 2601
rect 14921 2635 14979 2641
rect 14921 2601 14933 2635
rect 14967 2632 14979 2635
rect 15102 2632 15108 2644
rect 14967 2604 15108 2632
rect 14967 2601 14979 2604
rect 14921 2595 14979 2601
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 5261 2567 5319 2573
rect 5261 2533 5273 2567
rect 5307 2564 5319 2567
rect 5810 2564 5816 2576
rect 5307 2536 5816 2564
rect 5307 2533 5319 2536
rect 5261 2527 5319 2533
rect 5810 2524 5816 2536
rect 5868 2524 5874 2576
rect 7101 2567 7159 2573
rect 7101 2533 7113 2567
rect 7147 2564 7159 2567
rect 8018 2564 8024 2576
rect 7147 2536 8024 2564
rect 7147 2533 7159 2536
rect 7101 2527 7159 2533
rect 8018 2524 8024 2536
rect 8076 2524 8082 2576
rect 6196 2468 7420 2496
rect 6196 2440 6224 2468
rect 5077 2431 5135 2437
rect 5077 2397 5089 2431
rect 5123 2397 5135 2431
rect 5077 2391 5135 2397
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 5994 2428 6000 2440
rect 5859 2400 6000 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6178 2388 6184 2440
rect 6236 2388 6242 2440
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 6638 2388 6644 2440
rect 6696 2428 6702 2440
rect 6840 2437 6868 2468
rect 6733 2431 6791 2437
rect 6733 2428 6745 2431
rect 6696 2400 6745 2428
rect 6696 2388 6702 2400
rect 6733 2397 6745 2400
rect 6779 2397 6791 2431
rect 6733 2391 6791 2397
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 7282 2428 7288 2440
rect 6963 2400 7288 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7392 2437 7420 2468
rect 9490 2456 9496 2508
rect 9548 2496 9554 2508
rect 9548 2468 10456 2496
rect 9548 2456 9554 2468
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 7377 2391 7435 2397
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 7929 2431 7987 2437
rect 7929 2428 7941 2431
rect 7616 2400 7941 2428
rect 7616 2388 7622 2400
rect 7929 2397 7941 2400
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 8021 2431 8079 2437
rect 8021 2397 8033 2431
rect 8067 2428 8079 2431
rect 8294 2428 8300 2440
rect 8067 2400 8300 2428
rect 8067 2397 8079 2400
rect 8021 2391 8079 2397
rect 8294 2388 8300 2400
rect 8352 2428 8358 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 8352 2400 8585 2428
rect 8352 2388 8358 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2428 9459 2431
rect 9950 2428 9956 2440
rect 9447 2400 9956 2428
rect 9447 2397 9459 2400
rect 9401 2391 9459 2397
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10428 2437 10456 2468
rect 12250 2456 12256 2508
rect 12308 2496 12314 2508
rect 14458 2496 14464 2508
rect 12308 2468 14464 2496
rect 12308 2456 12314 2468
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2397 10103 2431
rect 10045 2391 10103 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2428 11391 2431
rect 11422 2428 11428 2440
rect 11379 2400 11428 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 1486 2320 1492 2372
rect 1544 2360 1550 2372
rect 1642 2363 1700 2369
rect 1642 2360 1654 2363
rect 1544 2332 1654 2360
rect 1544 2320 1550 2332
rect 1642 2329 1654 2332
rect 1688 2329 1700 2363
rect 1642 2323 1700 2329
rect 3421 2363 3479 2369
rect 3421 2329 3433 2363
rect 3467 2360 3479 2363
rect 3786 2360 3792 2372
rect 3467 2332 3792 2360
rect 3467 2329 3479 2332
rect 3421 2323 3479 2329
rect 3786 2320 3792 2332
rect 3844 2320 3850 2372
rect 6454 2360 6460 2372
rect 5644 2332 6460 2360
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 4522 2252 4528 2304
rect 4580 2252 4586 2304
rect 4893 2295 4951 2301
rect 4893 2261 4905 2295
rect 4939 2292 4951 2295
rect 5166 2292 5172 2304
rect 4939 2264 5172 2292
rect 4939 2261 4951 2264
rect 4893 2255 4951 2261
rect 5166 2252 5172 2264
rect 5224 2252 5230 2304
rect 5644 2301 5672 2332
rect 6454 2320 6460 2332
rect 6512 2320 6518 2372
rect 7193 2363 7251 2369
rect 7193 2329 7205 2363
rect 7239 2360 7251 2363
rect 8386 2360 8392 2372
rect 7239 2332 8392 2360
rect 7239 2329 7251 2332
rect 7193 2323 7251 2329
rect 8386 2320 8392 2332
rect 8444 2320 8450 2372
rect 10060 2360 10088 2391
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 11974 2388 11980 2440
rect 12032 2388 12038 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 12986 2388 12992 2440
rect 13044 2388 13050 2440
rect 13906 2388 13912 2440
rect 13964 2388 13970 2440
rect 14292 2437 14320 2468
rect 14458 2456 14464 2468
rect 14516 2456 14522 2508
rect 14642 2456 14648 2508
rect 14700 2496 14706 2508
rect 15105 2499 15163 2505
rect 15105 2496 15117 2499
rect 14700 2468 15117 2496
rect 14700 2456 14706 2468
rect 15105 2465 15117 2468
rect 15151 2465 15163 2499
rect 15105 2459 15163 2465
rect 15378 2437 15384 2440
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2397 14335 2431
rect 15372 2428 15384 2437
rect 15339 2400 15384 2428
rect 14277 2391 14335 2397
rect 15372 2391 15384 2400
rect 15378 2388 15384 2391
rect 15436 2388 15442 2440
rect 11054 2360 11060 2372
rect 10060 2332 11060 2360
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 14093 2363 14151 2369
rect 14093 2360 14105 2363
rect 13320 2332 14105 2360
rect 13320 2320 13326 2332
rect 14093 2329 14105 2332
rect 14139 2360 14151 2363
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14139 2332 14565 2360
rect 14139 2329 14151 2332
rect 14093 2323 14151 2329
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 14737 2363 14795 2369
rect 14737 2329 14749 2363
rect 14783 2360 14795 2363
rect 15562 2360 15568 2372
rect 14783 2332 15568 2360
rect 14783 2329 14795 2332
rect 14737 2323 14795 2329
rect 15562 2320 15568 2332
rect 15620 2360 15626 2372
rect 15620 2332 16528 2360
rect 15620 2320 15626 2332
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2261 5687 2295
rect 5629 2255 5687 2261
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 7006 2292 7012 2304
rect 6043 2264 7012 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7742 2252 7748 2304
rect 7800 2252 7806 2304
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2292 8263 2295
rect 8294 2292 8300 2304
rect 8251 2264 8300 2292
rect 8251 2261 8263 2264
rect 8205 2255 8263 2261
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 9030 2252 9036 2304
rect 9088 2292 9094 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 9088 2264 9229 2292
rect 9088 2252 9094 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9861 2295 9919 2301
rect 9861 2292 9873 2295
rect 9732 2264 9873 2292
rect 9732 2252 9738 2264
rect 9861 2261 9873 2264
rect 9907 2261 9919 2295
rect 9861 2255 9919 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 10376 2264 10609 2292
rect 10376 2252 10382 2264
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10597 2255 10655 2261
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 11149 2295 11207 2301
rect 11149 2292 11161 2295
rect 11020 2264 11161 2292
rect 11020 2252 11026 2264
rect 11149 2261 11161 2264
rect 11195 2261 11207 2295
rect 11149 2255 11207 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 11793 2255 11851 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 12437 2295 12495 2301
rect 12437 2292 12449 2295
rect 12308 2264 12449 2292
rect 12308 2252 12314 2264
rect 12437 2261 12449 2264
rect 12483 2261 12495 2295
rect 12437 2255 12495 2261
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 16500 2301 16528 2332
rect 13725 2295 13783 2301
rect 13725 2292 13737 2295
rect 13596 2264 13737 2292
rect 13596 2252 13602 2264
rect 13725 2261 13737 2264
rect 13771 2261 13783 2295
rect 13725 2255 13783 2261
rect 16485 2295 16543 2301
rect 16485 2261 16497 2295
rect 16531 2261 16543 2295
rect 16485 2255 16543 2261
rect 1104 2202 16836 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 16836 2202
rect 1104 2128 16836 2150
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 1578 1340 1584 1352
rect 72 1312 1584 1340
rect 72 1300 78 1312
rect 1578 1300 1584 1312
rect 1636 1300 1642 1352
rect 14182 1300 14188 1352
rect 14240 1340 14246 1352
rect 16298 1340 16304 1352
rect 14240 1312 16304 1340
rect 14240 1300 14246 1312
rect 16298 1300 16304 1312
rect 16356 1300 16362 1352
rect 658 1232 664 1284
rect 716 1272 722 1284
rect 2314 1272 2320 1284
rect 716 1244 2320 1272
rect 716 1232 722 1244
rect 2314 1232 2320 1244
rect 2372 1232 2378 1284
rect 14826 1096 14832 1148
rect 14884 1136 14890 1148
rect 15838 1136 15844 1148
rect 14884 1108 15844 1136
rect 14884 1096 14890 1108
rect 15838 1096 15844 1108
rect 15896 1096 15902 1148
<< via1 >>
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 8668 39584 8720 39636
rect 10968 39380 11020 39432
rect 12900 39380 12952 39432
rect 8208 39312 8260 39364
rect 10048 39287 10100 39296
rect 10048 39253 10057 39287
rect 10057 39253 10091 39287
rect 10091 39253 10100 39287
rect 10048 39244 10100 39253
rect 10784 39244 10836 39296
rect 11336 39244 11388 39296
rect 12624 39244 12676 39296
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 7012 38972 7064 39024
rect 6920 38947 6972 38956
rect 6920 38913 6929 38947
rect 6929 38913 6963 38947
rect 6963 38913 6972 38947
rect 6920 38904 6972 38913
rect 7104 38947 7156 38956
rect 7104 38913 7113 38947
rect 7113 38913 7147 38947
rect 7147 38913 7156 38947
rect 7104 38904 7156 38913
rect 7380 39015 7432 39024
rect 7380 38981 7405 39015
rect 7405 38981 7432 39015
rect 10048 39040 10100 39092
rect 7380 38972 7432 38981
rect 8208 38904 8260 38956
rect 12716 38904 12768 38956
rect 6092 38836 6144 38888
rect 9772 38836 9824 38888
rect 13912 38836 13964 38888
rect 7104 38743 7156 38752
rect 7104 38709 7113 38743
rect 7113 38709 7147 38743
rect 7147 38709 7156 38743
rect 7104 38700 7156 38709
rect 7932 38700 7984 38752
rect 8300 38700 8352 38752
rect 11060 38700 11112 38752
rect 12072 38700 12124 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 7748 38496 7800 38548
rect 7932 38496 7984 38548
rect 8668 38496 8720 38548
rect 10784 38539 10836 38548
rect 10784 38505 10793 38539
rect 10793 38505 10827 38539
rect 10827 38505 10836 38539
rect 10784 38496 10836 38505
rect 12164 38496 12216 38548
rect 12716 38496 12768 38548
rect 7380 38428 7432 38480
rect 6092 38403 6144 38412
rect 6092 38369 6101 38403
rect 6101 38369 6135 38403
rect 6135 38369 6144 38403
rect 6092 38360 6144 38369
rect 6644 38224 6696 38276
rect 8116 38335 8168 38344
rect 8116 38301 8125 38335
rect 8125 38301 8159 38335
rect 8159 38301 8168 38335
rect 8116 38292 8168 38301
rect 8484 38292 8536 38344
rect 9772 38292 9824 38344
rect 10600 38335 10652 38344
rect 10600 38301 10609 38335
rect 10609 38301 10643 38335
rect 10643 38301 10652 38335
rect 10600 38292 10652 38301
rect 13912 38403 13964 38412
rect 13912 38369 13921 38403
rect 13921 38369 13955 38403
rect 13955 38369 13964 38403
rect 13912 38360 13964 38369
rect 11060 38335 11112 38344
rect 11060 38301 11069 38335
rect 11069 38301 11103 38335
rect 11103 38301 11112 38335
rect 11060 38292 11112 38301
rect 11520 38292 11572 38344
rect 12164 38292 12216 38344
rect 7564 38156 7616 38208
rect 7656 38199 7708 38208
rect 7656 38165 7665 38199
rect 7665 38165 7699 38199
rect 7699 38165 7708 38199
rect 7656 38156 7708 38165
rect 7840 38199 7892 38208
rect 7840 38165 7867 38199
rect 7867 38165 7892 38199
rect 7840 38156 7892 38165
rect 8208 38224 8260 38276
rect 8300 38156 8352 38208
rect 8576 38199 8628 38208
rect 11888 38267 11940 38276
rect 11888 38233 11897 38267
rect 11897 38233 11931 38267
rect 11931 38233 11940 38267
rect 11888 38224 11940 38233
rect 13084 38224 13136 38276
rect 8576 38165 8601 38199
rect 8601 38165 8628 38199
rect 8576 38156 8628 38165
rect 10324 38199 10376 38208
rect 10324 38165 10333 38199
rect 10333 38165 10367 38199
rect 10367 38165 10376 38199
rect 10324 38156 10376 38165
rect 12348 38156 12400 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 6644 37995 6696 38004
rect 6644 37961 6653 37995
rect 6653 37961 6687 37995
rect 6687 37961 6696 37995
rect 6644 37952 6696 37961
rect 7104 37952 7156 38004
rect 7196 37995 7248 38004
rect 7196 37961 7205 37995
rect 7205 37961 7239 37995
rect 7239 37961 7248 37995
rect 7196 37952 7248 37961
rect 7656 37952 7708 38004
rect 8116 37995 8168 38004
rect 8116 37961 8131 37995
rect 8131 37961 8165 37995
rect 8165 37961 8168 37995
rect 8116 37952 8168 37961
rect 8760 37952 8812 38004
rect 9956 37952 10008 38004
rect 10324 37952 10376 38004
rect 10600 37952 10652 38004
rect 12256 37952 12308 38004
rect 13084 37995 13136 38004
rect 13084 37961 13093 37995
rect 13093 37961 13127 37995
rect 13127 37961 13136 37995
rect 13084 37952 13136 37961
rect 7012 37927 7064 37936
rect 7012 37893 7021 37927
rect 7021 37893 7055 37927
rect 7055 37893 7064 37927
rect 7012 37884 7064 37893
rect 7840 37884 7892 37936
rect 7564 37859 7616 37868
rect 7564 37825 7573 37859
rect 7573 37825 7607 37859
rect 7607 37825 7616 37859
rect 7564 37816 7616 37825
rect 7656 37859 7708 37868
rect 7656 37825 7665 37859
rect 7665 37825 7699 37859
rect 7699 37825 7708 37859
rect 7656 37816 7708 37825
rect 8576 37748 8628 37800
rect 8760 37859 8812 37868
rect 8760 37825 8776 37859
rect 8776 37825 8810 37859
rect 8810 37825 8812 37859
rect 8760 37816 8812 37825
rect 12624 37884 12676 37936
rect 11060 37816 11112 37868
rect 11244 37748 11296 37800
rect 12072 37816 12124 37868
rect 12348 37859 12400 37868
rect 12348 37825 12357 37859
rect 12357 37825 12391 37859
rect 12391 37825 12400 37859
rect 12348 37816 12400 37825
rect 12808 37859 12860 37868
rect 12808 37825 12817 37859
rect 12817 37825 12851 37859
rect 12851 37825 12860 37859
rect 12808 37816 12860 37825
rect 12624 37748 12676 37800
rect 13360 37859 13412 37868
rect 13360 37825 13369 37859
rect 13369 37825 13403 37859
rect 13403 37825 13412 37859
rect 13360 37816 13412 37825
rect 8300 37680 8352 37732
rect 11704 37680 11756 37732
rect 12164 37723 12216 37732
rect 12164 37689 12173 37723
rect 12173 37689 12207 37723
rect 12207 37689 12216 37723
rect 12164 37680 12216 37689
rect 6828 37655 6880 37664
rect 6828 37621 6837 37655
rect 6837 37621 6871 37655
rect 6871 37621 6880 37655
rect 6828 37612 6880 37621
rect 6920 37612 6972 37664
rect 10876 37612 10928 37664
rect 11152 37612 11204 37664
rect 11888 37612 11940 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 6828 37408 6880 37460
rect 8668 37408 8720 37460
rect 11520 37451 11572 37460
rect 11520 37417 11529 37451
rect 11529 37417 11563 37451
rect 11563 37417 11572 37451
rect 11520 37408 11572 37417
rect 11704 37451 11756 37460
rect 11704 37417 11713 37451
rect 11713 37417 11747 37451
rect 11747 37417 11756 37451
rect 11704 37408 11756 37417
rect 12808 37408 12860 37460
rect 10600 37340 10652 37392
rect 10876 37340 10928 37392
rect 7012 37204 7064 37256
rect 9864 37247 9916 37256
rect 9864 37213 9873 37247
rect 9873 37213 9907 37247
rect 9907 37213 9916 37247
rect 9864 37204 9916 37213
rect 9956 37247 10008 37256
rect 9956 37213 9965 37247
rect 9965 37213 9999 37247
rect 9999 37213 10008 37247
rect 9956 37204 10008 37213
rect 11704 37272 11756 37324
rect 12348 37272 12400 37324
rect 10784 37247 10836 37256
rect 10784 37213 10793 37247
rect 10793 37213 10827 37247
rect 10827 37213 10836 37247
rect 10784 37204 10836 37213
rect 11060 37247 11112 37256
rect 11060 37213 11069 37247
rect 11069 37213 11103 37247
rect 11103 37213 11112 37247
rect 11060 37204 11112 37213
rect 11244 37247 11296 37256
rect 11244 37213 11253 37247
rect 11253 37213 11287 37247
rect 11287 37213 11296 37247
rect 11244 37204 11296 37213
rect 12624 37247 12676 37256
rect 12624 37213 12633 37247
rect 12633 37213 12667 37247
rect 12667 37213 12676 37247
rect 12624 37204 12676 37213
rect 13360 37204 13412 37256
rect 6736 37111 6788 37120
rect 6736 37077 6745 37111
rect 6745 37077 6779 37111
rect 6779 37077 6788 37111
rect 6736 37068 6788 37077
rect 7012 37068 7064 37120
rect 10048 37068 10100 37120
rect 11244 37068 11296 37120
rect 12072 37136 12124 37188
rect 12992 37136 13044 37188
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 9956 36864 10008 36916
rect 2964 36839 3016 36848
rect 2964 36805 2991 36839
rect 2991 36805 3016 36839
rect 2964 36796 3016 36805
rect 2044 36660 2096 36712
rect 6736 36796 6788 36848
rect 9036 36796 9088 36848
rect 11152 36796 11204 36848
rect 4068 36728 4120 36780
rect 6092 36728 6144 36780
rect 3608 36660 3660 36712
rect 10048 36771 10100 36780
rect 10048 36737 10057 36771
rect 10057 36737 10091 36771
rect 10091 36737 10100 36771
rect 10048 36728 10100 36737
rect 10416 36728 10468 36780
rect 11244 36728 11296 36780
rect 9864 36660 9916 36712
rect 10232 36660 10284 36712
rect 11704 36660 11756 36712
rect 7932 36592 7984 36644
rect 8208 36592 8260 36644
rect 12164 36592 12216 36644
rect 2780 36567 2832 36576
rect 2780 36533 2789 36567
rect 2789 36533 2823 36567
rect 2823 36533 2832 36567
rect 2780 36524 2832 36533
rect 3976 36524 4028 36576
rect 5356 36567 5408 36576
rect 5356 36533 5365 36567
rect 5365 36533 5399 36567
rect 5399 36533 5408 36567
rect 5356 36524 5408 36533
rect 7288 36524 7340 36576
rect 10508 36524 10560 36576
rect 10784 36567 10836 36576
rect 10784 36533 10793 36567
rect 10793 36533 10827 36567
rect 10827 36533 10836 36567
rect 10784 36524 10836 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 2044 36363 2096 36372
rect 2044 36329 2053 36363
rect 2053 36329 2087 36363
rect 2087 36329 2096 36363
rect 2044 36320 2096 36329
rect 4068 36320 4120 36372
rect 4160 36363 4212 36372
rect 4160 36329 4169 36363
rect 4169 36329 4203 36363
rect 4203 36329 4212 36363
rect 4160 36320 4212 36329
rect 2136 36159 2188 36168
rect 2136 36125 2145 36159
rect 2145 36125 2179 36159
rect 2179 36125 2188 36159
rect 2136 36116 2188 36125
rect 2780 36116 2832 36168
rect 3608 36159 3660 36168
rect 3608 36125 3617 36159
rect 3617 36125 3651 36159
rect 3651 36125 3660 36159
rect 3608 36116 3660 36125
rect 7012 36363 7064 36372
rect 7012 36329 7021 36363
rect 7021 36329 7055 36363
rect 7055 36329 7064 36363
rect 7012 36320 7064 36329
rect 10048 36320 10100 36372
rect 4528 36116 4580 36168
rect 4712 36227 4764 36236
rect 4712 36193 4721 36227
rect 4721 36193 4755 36227
rect 4755 36193 4764 36227
rect 4712 36184 4764 36193
rect 4804 36159 4856 36168
rect 4804 36125 4813 36159
rect 4813 36125 4847 36159
rect 4847 36125 4856 36159
rect 4804 36116 4856 36125
rect 4896 36159 4948 36168
rect 4896 36125 4905 36159
rect 4905 36125 4939 36159
rect 4939 36125 4948 36159
rect 4896 36116 4948 36125
rect 5356 36116 5408 36168
rect 5632 36159 5684 36168
rect 5632 36125 5641 36159
rect 5641 36125 5675 36159
rect 5675 36125 5684 36159
rect 5632 36116 5684 36125
rect 5908 36159 5960 36168
rect 5908 36125 5917 36159
rect 5917 36125 5951 36159
rect 5951 36125 5960 36159
rect 5908 36116 5960 36125
rect 6920 36184 6972 36236
rect 5172 36048 5224 36100
rect 3240 35980 3292 36032
rect 4620 35980 4672 36032
rect 4988 35980 5040 36032
rect 5356 35980 5408 36032
rect 7196 36116 7248 36168
rect 9128 36159 9180 36168
rect 9128 36125 9137 36159
rect 9137 36125 9171 36159
rect 9171 36125 9180 36159
rect 9128 36116 9180 36125
rect 9956 36116 10008 36168
rect 11428 36320 11480 36372
rect 12164 36320 12216 36372
rect 10784 36252 10836 36304
rect 12072 36252 12124 36304
rect 10600 36116 10652 36168
rect 7104 36048 7156 36100
rect 8576 36048 8628 36100
rect 11152 36116 11204 36168
rect 11428 36227 11480 36236
rect 11428 36193 11437 36227
rect 11437 36193 11471 36227
rect 11471 36193 11480 36227
rect 11428 36184 11480 36193
rect 13912 36227 13964 36236
rect 13912 36193 13921 36227
rect 13921 36193 13955 36227
rect 13955 36193 13964 36227
rect 13912 36184 13964 36193
rect 11336 36048 11388 36100
rect 11520 36159 11572 36168
rect 11520 36125 11529 36159
rect 11529 36125 11563 36159
rect 11563 36125 11572 36159
rect 11520 36116 11572 36125
rect 13084 36116 13136 36168
rect 12808 36048 12860 36100
rect 7472 35980 7524 36032
rect 8208 35980 8260 36032
rect 9036 35980 9088 36032
rect 10600 35980 10652 36032
rect 11060 36023 11112 36032
rect 11060 35989 11069 36023
rect 11069 35989 11103 36023
rect 11103 35989 11112 36023
rect 11060 35980 11112 35989
rect 12256 36023 12308 36032
rect 12256 35989 12265 36023
rect 12265 35989 12299 36023
rect 12299 35989 12308 36023
rect 12256 35980 12308 35989
rect 12440 36023 12492 36032
rect 12440 35989 12449 36023
rect 12449 35989 12483 36023
rect 12483 35989 12492 36023
rect 12440 35980 12492 35989
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 2964 35776 3016 35828
rect 4804 35776 4856 35828
rect 3240 35751 3292 35760
rect 3240 35717 3249 35751
rect 3249 35717 3283 35751
rect 3283 35717 3292 35751
rect 3240 35708 3292 35717
rect 4528 35708 4580 35760
rect 5264 35776 5316 35828
rect 5540 35776 5592 35828
rect 8576 35819 8628 35828
rect 8576 35785 8585 35819
rect 8585 35785 8619 35819
rect 8619 35785 8628 35819
rect 8576 35776 8628 35785
rect 9128 35776 9180 35828
rect 9956 35819 10008 35828
rect 9956 35785 9965 35819
rect 9965 35785 9999 35819
rect 9999 35785 10008 35819
rect 9956 35776 10008 35785
rect 10232 35776 10284 35828
rect 2136 35640 2188 35692
rect 4804 35683 4856 35692
rect 4804 35649 4813 35683
rect 4813 35649 4847 35683
rect 4847 35649 4856 35683
rect 4804 35640 4856 35649
rect 5356 35572 5408 35624
rect 5540 35683 5592 35692
rect 5540 35649 5549 35683
rect 5549 35649 5583 35683
rect 5583 35649 5592 35683
rect 5540 35640 5592 35649
rect 5632 35683 5684 35692
rect 5632 35649 5641 35683
rect 5641 35649 5675 35683
rect 5675 35649 5684 35683
rect 5632 35640 5684 35649
rect 5724 35683 5776 35692
rect 5724 35649 5733 35683
rect 5733 35649 5767 35683
rect 5767 35649 5776 35683
rect 5724 35640 5776 35649
rect 6736 35683 6788 35692
rect 6736 35649 6745 35683
rect 6745 35649 6779 35683
rect 6779 35649 6788 35683
rect 6736 35640 6788 35649
rect 7196 35683 7248 35692
rect 7196 35649 7205 35683
rect 7205 35649 7239 35683
rect 7239 35649 7248 35683
rect 7196 35640 7248 35649
rect 7472 35683 7524 35692
rect 7472 35649 7481 35683
rect 7481 35649 7515 35683
rect 7515 35649 7524 35683
rect 7472 35640 7524 35649
rect 6000 35572 6052 35624
rect 4160 35436 4212 35488
rect 4712 35436 4764 35488
rect 5356 35436 5408 35488
rect 8024 35572 8076 35624
rect 7840 35504 7892 35556
rect 8944 35615 8996 35624
rect 8944 35581 8953 35615
rect 8953 35581 8987 35615
rect 8987 35581 8996 35615
rect 8944 35572 8996 35581
rect 9496 35640 9548 35692
rect 10324 35751 10376 35760
rect 10324 35717 10333 35751
rect 10333 35717 10367 35751
rect 10367 35717 10376 35751
rect 10324 35708 10376 35717
rect 11060 35708 11112 35760
rect 11520 35776 11572 35828
rect 13084 35776 13136 35828
rect 11428 35708 11480 35760
rect 12164 35751 12216 35760
rect 12164 35717 12173 35751
rect 12173 35717 12207 35751
rect 12207 35717 12216 35751
rect 12164 35708 12216 35717
rect 12348 35751 12400 35760
rect 12348 35717 12373 35751
rect 12373 35717 12400 35751
rect 12348 35708 12400 35717
rect 12532 35708 12584 35760
rect 9956 35640 10008 35692
rect 8116 35436 8168 35488
rect 8208 35436 8260 35488
rect 9680 35572 9732 35624
rect 9772 35572 9824 35624
rect 10232 35683 10284 35692
rect 10232 35649 10241 35683
rect 10241 35649 10275 35683
rect 10275 35649 10284 35683
rect 10232 35640 10284 35649
rect 10508 35683 10560 35692
rect 10508 35649 10517 35683
rect 10517 35649 10551 35683
rect 10551 35649 10560 35683
rect 10508 35640 10560 35649
rect 10600 35683 10652 35692
rect 10600 35649 10609 35683
rect 10609 35649 10643 35683
rect 10643 35649 10652 35683
rect 10600 35640 10652 35649
rect 12072 35683 12124 35692
rect 10968 35572 11020 35624
rect 10876 35504 10928 35556
rect 9864 35479 9916 35488
rect 9864 35445 9873 35479
rect 9873 35445 9907 35479
rect 9907 35445 9916 35479
rect 9864 35436 9916 35445
rect 12072 35649 12081 35683
rect 12081 35649 12115 35683
rect 12115 35649 12124 35683
rect 12072 35640 12124 35649
rect 11336 35504 11388 35556
rect 12440 35572 12492 35624
rect 12624 35615 12676 35624
rect 12624 35581 12633 35615
rect 12633 35581 12667 35615
rect 12667 35581 12676 35615
rect 12624 35572 12676 35581
rect 12256 35436 12308 35488
rect 12808 35436 12860 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 2136 35232 2188 35284
rect 4620 35232 4672 35284
rect 5724 35232 5776 35284
rect 6000 35275 6052 35284
rect 6000 35241 6009 35275
rect 6009 35241 6043 35275
rect 6043 35241 6052 35275
rect 6000 35232 6052 35241
rect 8024 35275 8076 35284
rect 8024 35241 8033 35275
rect 8033 35241 8067 35275
rect 8067 35241 8076 35275
rect 8024 35232 8076 35241
rect 8392 35275 8444 35284
rect 8392 35241 8401 35275
rect 8401 35241 8435 35275
rect 8435 35241 8444 35275
rect 8392 35232 8444 35241
rect 4068 35164 4120 35216
rect 5908 35164 5960 35216
rect 6828 35164 6880 35216
rect 3608 35071 3660 35080
rect 3608 35037 3617 35071
rect 3617 35037 3651 35071
rect 3651 35037 3660 35071
rect 3608 35028 3660 35037
rect 6092 35028 6144 35080
rect 7564 35028 7616 35080
rect 7840 35071 7892 35080
rect 7840 35037 7849 35071
rect 7849 35037 7883 35071
rect 7883 35037 7892 35071
rect 7840 35028 7892 35037
rect 8116 35096 8168 35148
rect 8944 35275 8996 35284
rect 8944 35241 8953 35275
rect 8953 35241 8987 35275
rect 8987 35241 8996 35275
rect 8944 35232 8996 35241
rect 9772 35275 9824 35284
rect 9772 35241 9781 35275
rect 9781 35241 9815 35275
rect 9815 35241 9824 35275
rect 9772 35232 9824 35241
rect 9956 35275 10008 35284
rect 9956 35241 9965 35275
rect 9965 35241 9999 35275
rect 9999 35241 10008 35275
rect 9956 35232 10008 35241
rect 10232 35232 10284 35284
rect 12348 35232 12400 35284
rect 9312 35164 9364 35216
rect 10416 35164 10468 35216
rect 10784 35164 10836 35216
rect 9956 35096 10008 35148
rect 12256 35096 12308 35148
rect 3056 34960 3108 35012
rect 4160 34935 4212 34944
rect 4160 34901 4169 34935
rect 4169 34901 4203 34935
rect 4203 34901 4212 34935
rect 4160 34892 4212 34901
rect 5540 34960 5592 35012
rect 6736 34960 6788 35012
rect 8300 34960 8352 35012
rect 9496 35071 9548 35080
rect 9496 35037 9505 35071
rect 9505 35037 9539 35071
rect 9539 35037 9548 35071
rect 9496 35028 9548 35037
rect 9680 35071 9732 35080
rect 9680 35037 9689 35071
rect 9689 35037 9723 35071
rect 9723 35037 9732 35071
rect 9680 35028 9732 35037
rect 10508 35028 10560 35080
rect 10232 34960 10284 35012
rect 10324 35003 10376 35012
rect 10324 34969 10333 35003
rect 10333 34969 10367 35003
rect 10367 34969 10376 35003
rect 10324 34960 10376 34969
rect 10416 35003 10468 35012
rect 10416 34969 10425 35003
rect 10425 34969 10459 35003
rect 10459 34969 10468 35003
rect 10416 34960 10468 34969
rect 11336 35071 11388 35080
rect 11336 35037 11345 35071
rect 11345 35037 11379 35071
rect 11379 35037 11388 35071
rect 11336 35028 11388 35037
rect 11520 35028 11572 35080
rect 11612 35071 11664 35080
rect 11612 35037 11621 35071
rect 11621 35037 11655 35071
rect 11655 35037 11664 35071
rect 11612 35028 11664 35037
rect 12072 34960 12124 35012
rect 12440 34892 12492 34944
rect 12992 35028 13044 35080
rect 12716 34892 12768 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 3056 34731 3108 34740
rect 3056 34697 3065 34731
rect 3065 34697 3099 34731
rect 3099 34697 3108 34731
rect 3056 34688 3108 34697
rect 8392 34688 8444 34740
rect 11152 34688 11204 34740
rect 2136 34620 2188 34672
rect 10692 34620 10744 34672
rect 11336 34620 11388 34672
rect 13176 34663 13228 34672
rect 7472 34552 7524 34604
rect 8208 34552 8260 34604
rect 12256 34595 12308 34604
rect 12256 34561 12265 34595
rect 12265 34561 12299 34595
rect 12299 34561 12308 34595
rect 12256 34552 12308 34561
rect 12532 34595 12584 34604
rect 12532 34561 12541 34595
rect 12541 34561 12575 34595
rect 12575 34561 12584 34595
rect 12532 34552 12584 34561
rect 12716 34595 12768 34604
rect 12716 34561 12725 34595
rect 12725 34561 12759 34595
rect 12759 34561 12768 34595
rect 12716 34552 12768 34561
rect 12808 34595 12860 34604
rect 12808 34561 12817 34595
rect 12817 34561 12851 34595
rect 12851 34561 12860 34595
rect 12808 34552 12860 34561
rect 13176 34629 13185 34663
rect 13185 34629 13219 34663
rect 13219 34629 13228 34663
rect 13176 34620 13228 34629
rect 13084 34595 13136 34604
rect 13084 34561 13093 34595
rect 13093 34561 13127 34595
rect 13127 34561 13136 34595
rect 13084 34552 13136 34561
rect 13360 34552 13412 34604
rect 2872 34459 2924 34468
rect 2872 34425 2881 34459
rect 2881 34425 2915 34459
rect 2915 34425 2924 34459
rect 2872 34416 2924 34425
rect 4160 34416 4212 34468
rect 7288 34416 7340 34468
rect 8668 34416 8720 34468
rect 9220 34416 9272 34468
rect 12440 34484 12492 34536
rect 12900 34484 12952 34536
rect 12808 34416 12860 34468
rect 7196 34348 7248 34400
rect 9036 34348 9088 34400
rect 12348 34348 12400 34400
rect 12716 34348 12768 34400
rect 12992 34348 13044 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 4528 34144 4580 34196
rect 4160 34076 4212 34128
rect 4436 34008 4488 34060
rect 5908 34144 5960 34196
rect 7288 34144 7340 34196
rect 7840 34144 7892 34196
rect 8208 34187 8260 34196
rect 8208 34153 8217 34187
rect 8217 34153 8251 34187
rect 8251 34153 8260 34187
rect 8208 34144 8260 34153
rect 10416 34144 10468 34196
rect 12532 34144 12584 34196
rect 13084 34144 13136 34196
rect 13728 34144 13780 34196
rect 7380 34076 7432 34128
rect 7932 34076 7984 34128
rect 6092 34051 6144 34060
rect 6092 34017 6101 34051
rect 6101 34017 6135 34051
rect 6135 34017 6144 34051
rect 6092 34008 6144 34017
rect 4344 33940 4396 33992
rect 4712 33940 4764 33992
rect 10048 34008 10100 34060
rect 12716 34076 12768 34128
rect 12992 34076 13044 34128
rect 13360 34076 13412 34128
rect 7012 33940 7064 33992
rect 3976 33872 4028 33924
rect 5448 33872 5500 33924
rect 7196 33915 7248 33924
rect 7196 33881 7223 33915
rect 7223 33881 7248 33915
rect 7196 33872 7248 33881
rect 7380 33915 7432 33924
rect 7380 33881 7389 33915
rect 7389 33881 7423 33915
rect 7423 33881 7432 33915
rect 7380 33872 7432 33881
rect 8024 33940 8076 33992
rect 9036 33983 9088 33992
rect 9036 33949 9045 33983
rect 9045 33949 9079 33983
rect 9079 33949 9088 33983
rect 9036 33940 9088 33949
rect 9864 33940 9916 33992
rect 9956 33983 10008 33992
rect 9956 33949 9965 33983
rect 9965 33949 9999 33983
rect 9999 33949 10008 33983
rect 9956 33940 10008 33949
rect 4620 33847 4672 33856
rect 4620 33813 4645 33847
rect 4645 33813 4672 33847
rect 4620 33804 4672 33813
rect 4804 33847 4856 33856
rect 4804 33813 4813 33847
rect 4813 33813 4847 33847
rect 4847 33813 4856 33847
rect 4804 33804 4856 33813
rect 6920 33804 6972 33856
rect 7472 33847 7524 33856
rect 7472 33813 7481 33847
rect 7481 33813 7515 33847
rect 7515 33813 7524 33847
rect 7472 33804 7524 33813
rect 9220 33872 9272 33924
rect 10416 33983 10468 33992
rect 10416 33949 10425 33983
rect 10425 33949 10459 33983
rect 10459 33949 10468 33983
rect 10416 33940 10468 33949
rect 12440 34008 12492 34060
rect 11152 33983 11204 33992
rect 11152 33949 11160 33983
rect 11160 33949 11194 33983
rect 11194 33949 11204 33983
rect 11152 33940 11204 33949
rect 11244 33983 11296 33992
rect 11244 33949 11253 33983
rect 11253 33949 11287 33983
rect 11287 33949 11296 33983
rect 11244 33940 11296 33949
rect 12256 33940 12308 33992
rect 13912 34008 13964 34060
rect 12808 33983 12860 33992
rect 12808 33949 12817 33983
rect 12817 33949 12851 33983
rect 12851 33949 12860 33983
rect 12808 33940 12860 33949
rect 13176 33983 13228 33992
rect 13176 33949 13185 33983
rect 13185 33949 13219 33983
rect 13219 33949 13228 33983
rect 13176 33940 13228 33949
rect 8116 33804 8168 33856
rect 12072 33804 12124 33856
rect 12348 33872 12400 33924
rect 13728 33915 13780 33924
rect 13728 33881 13737 33915
rect 13737 33881 13771 33915
rect 13771 33881 13780 33915
rect 13728 33872 13780 33881
rect 12992 33804 13044 33856
rect 13084 33847 13136 33856
rect 13084 33813 13093 33847
rect 13093 33813 13127 33847
rect 13127 33813 13136 33847
rect 13084 33804 13136 33813
rect 13176 33804 13228 33856
rect 13360 33804 13412 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 4528 33643 4580 33652
rect 4528 33609 4537 33643
rect 4537 33609 4571 33643
rect 4571 33609 4580 33643
rect 4528 33600 4580 33609
rect 3608 33532 3660 33584
rect 4620 33532 4672 33584
rect 2964 33464 3016 33516
rect 4344 33507 4396 33516
rect 4344 33473 4353 33507
rect 4353 33473 4387 33507
rect 4387 33473 4396 33507
rect 4344 33464 4396 33473
rect 4436 33464 4488 33516
rect 6092 33532 6144 33584
rect 4896 33507 4948 33516
rect 4896 33473 4930 33507
rect 4930 33473 4948 33507
rect 4896 33464 4948 33473
rect 6828 33464 6880 33516
rect 9956 33600 10008 33652
rect 10784 33600 10836 33652
rect 11612 33600 11664 33652
rect 11704 33643 11756 33652
rect 11704 33609 11713 33643
rect 11713 33609 11747 33643
rect 11747 33609 11756 33643
rect 11704 33600 11756 33609
rect 10140 33532 10192 33584
rect 12624 33532 12676 33584
rect 8300 33464 8352 33516
rect 8484 33464 8536 33516
rect 8668 33507 8720 33516
rect 8668 33473 8702 33507
rect 8702 33473 8720 33507
rect 8668 33464 8720 33473
rect 7656 33371 7708 33380
rect 7656 33337 7665 33371
rect 7665 33337 7699 33371
rect 7699 33337 7708 33371
rect 7656 33328 7708 33337
rect 3884 33260 3936 33312
rect 4344 33260 4396 33312
rect 4804 33260 4856 33312
rect 5908 33260 5960 33312
rect 8760 33260 8812 33312
rect 9496 33260 9548 33312
rect 9956 33464 10008 33516
rect 10784 33507 10836 33516
rect 10784 33473 10793 33507
rect 10793 33473 10827 33507
rect 10827 33473 10836 33507
rect 10784 33464 10836 33473
rect 11980 33464 12032 33516
rect 12256 33464 12308 33516
rect 11244 33396 11296 33448
rect 12164 33439 12216 33448
rect 12164 33405 12173 33439
rect 12173 33405 12207 33439
rect 12207 33405 12216 33439
rect 12164 33396 12216 33405
rect 10416 33328 10468 33380
rect 12808 33464 12860 33516
rect 13912 33464 13964 33516
rect 10508 33260 10560 33312
rect 10600 33303 10652 33312
rect 10600 33269 10609 33303
rect 10609 33269 10643 33303
rect 10643 33269 10652 33303
rect 10600 33260 10652 33269
rect 10784 33260 10836 33312
rect 12716 33260 12768 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 2964 33099 3016 33108
rect 2964 33065 2973 33099
rect 2973 33065 3007 33099
rect 3007 33065 3016 33099
rect 2964 33056 3016 33065
rect 4068 32988 4120 33040
rect 4804 32920 4856 32972
rect 3884 32852 3936 32904
rect 4252 32895 4304 32904
rect 4252 32861 4261 32895
rect 4261 32861 4295 32895
rect 4295 32861 4304 32895
rect 4252 32852 4304 32861
rect 4620 32895 4672 32904
rect 4620 32861 4629 32895
rect 4629 32861 4663 32895
rect 4663 32861 4672 32895
rect 4620 32852 4672 32861
rect 5540 32895 5592 32904
rect 5540 32861 5549 32895
rect 5549 32861 5583 32895
rect 5583 32861 5592 32895
rect 5540 32852 5592 32861
rect 6828 33056 6880 33108
rect 8024 33099 8076 33108
rect 8024 33065 8033 33099
rect 8033 33065 8067 33099
rect 8067 33065 8076 33099
rect 8024 33056 8076 33065
rect 8668 33056 8720 33108
rect 9312 33099 9364 33108
rect 9312 33065 9321 33099
rect 9321 33065 9355 33099
rect 9355 33065 9364 33099
rect 9312 33056 9364 33065
rect 9864 33056 9916 33108
rect 12808 33099 12860 33108
rect 12808 33065 12817 33099
rect 12817 33065 12851 33099
rect 12851 33065 12860 33099
rect 12808 33056 12860 33065
rect 8300 32988 8352 33040
rect 9404 32988 9456 33040
rect 6092 32852 6144 32904
rect 6460 32852 6512 32904
rect 6920 32895 6972 32904
rect 6920 32861 6954 32895
rect 6954 32861 6972 32895
rect 6920 32852 6972 32861
rect 7380 32852 7432 32904
rect 8300 32895 8352 32904
rect 8300 32861 8309 32895
rect 8309 32861 8343 32895
rect 8343 32861 8352 32895
rect 8300 32852 8352 32861
rect 4344 32784 4396 32836
rect 7012 32784 7064 32836
rect 7472 32784 7524 32836
rect 8760 32852 8812 32904
rect 8576 32784 8628 32836
rect 9036 32852 9088 32904
rect 9956 32963 10008 32972
rect 9956 32929 9965 32963
rect 9965 32929 9999 32963
rect 9999 32929 10008 32963
rect 9956 32920 10008 32929
rect 10140 32920 10192 32972
rect 10876 32920 10928 32972
rect 11152 32963 11204 32972
rect 11152 32929 11161 32963
rect 11161 32929 11195 32963
rect 11195 32929 11204 32963
rect 11152 32920 11204 32929
rect 12164 32920 12216 32972
rect 13084 33056 13136 33108
rect 10048 32895 10100 32904
rect 10048 32861 10057 32895
rect 10057 32861 10091 32895
rect 10091 32861 10100 32895
rect 10048 32852 10100 32861
rect 10600 32852 10652 32904
rect 3516 32716 3568 32768
rect 3976 32716 4028 32768
rect 4068 32716 4120 32768
rect 5816 32716 5868 32768
rect 6276 32716 6328 32768
rect 10232 32784 10284 32836
rect 9128 32759 9180 32768
rect 9128 32725 9137 32759
rect 9137 32725 9171 32759
rect 9171 32725 9180 32759
rect 9128 32716 9180 32725
rect 9220 32716 9272 32768
rect 13912 32852 13964 32904
rect 12900 32784 12952 32836
rect 13176 32827 13228 32836
rect 13176 32793 13185 32827
rect 13185 32793 13219 32827
rect 13219 32793 13228 32827
rect 13176 32784 13228 32793
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 4252 32512 4304 32564
rect 5172 32512 5224 32564
rect 7656 32512 7708 32564
rect 10508 32512 10560 32564
rect 11704 32512 11756 32564
rect 4160 32444 4212 32496
rect 6276 32444 6328 32496
rect 10048 32444 10100 32496
rect 11888 32444 11940 32496
rect 13912 32444 13964 32496
rect 3976 32419 4028 32428
rect 3976 32385 3985 32419
rect 3985 32385 4019 32419
rect 4019 32385 4028 32419
rect 3976 32376 4028 32385
rect 4344 32376 4396 32428
rect 4620 32308 4672 32360
rect 5264 32419 5316 32428
rect 5264 32385 5273 32419
rect 5273 32385 5307 32419
rect 5307 32385 5316 32419
rect 5264 32376 5316 32385
rect 5448 32308 5500 32360
rect 5908 32376 5960 32428
rect 10140 32419 10192 32428
rect 10140 32385 10149 32419
rect 10149 32385 10183 32419
rect 10183 32385 10192 32419
rect 10140 32376 10192 32385
rect 10232 32376 10284 32428
rect 11152 32419 11204 32428
rect 11152 32385 11165 32419
rect 11165 32385 11204 32419
rect 11152 32376 11204 32385
rect 11244 32376 11296 32428
rect 6000 32308 6052 32360
rect 4804 32240 4856 32292
rect 3608 32215 3660 32224
rect 3608 32181 3617 32215
rect 3617 32181 3651 32215
rect 3651 32181 3660 32215
rect 3608 32172 3660 32181
rect 3700 32215 3752 32224
rect 3700 32181 3709 32215
rect 3709 32181 3743 32215
rect 3743 32181 3752 32215
rect 3700 32172 3752 32181
rect 4988 32172 5040 32224
rect 11428 32172 11480 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 3608 31968 3660 32020
rect 4712 31968 4764 32020
rect 3700 31900 3752 31952
rect 5908 31968 5960 32020
rect 7012 31968 7064 32020
rect 5172 31900 5224 31952
rect 2964 31764 3016 31816
rect 4896 31764 4948 31816
rect 4988 31807 5040 31816
rect 4988 31773 4997 31807
rect 4997 31773 5031 31807
rect 5031 31773 5040 31807
rect 4988 31764 5040 31773
rect 5448 31900 5500 31952
rect 6184 31900 6236 31952
rect 5356 31875 5408 31884
rect 5356 31841 5365 31875
rect 5365 31841 5399 31875
rect 5399 31841 5408 31875
rect 5356 31832 5408 31841
rect 5908 31832 5960 31884
rect 4804 31696 4856 31748
rect 6000 31807 6052 31816
rect 6000 31773 6009 31807
rect 6009 31773 6043 31807
rect 6043 31773 6052 31807
rect 6000 31764 6052 31773
rect 7012 31875 7064 31884
rect 7012 31841 7021 31875
rect 7021 31841 7055 31875
rect 7055 31841 7064 31875
rect 7012 31832 7064 31841
rect 6276 31807 6328 31816
rect 6276 31773 6285 31807
rect 6285 31773 6319 31807
rect 6319 31773 6328 31807
rect 6276 31764 6328 31773
rect 6920 31807 6972 31816
rect 6920 31773 6929 31807
rect 6929 31773 6963 31807
rect 6963 31773 6972 31807
rect 6920 31764 6972 31773
rect 5356 31696 5408 31748
rect 6828 31696 6880 31748
rect 8484 31807 8536 31816
rect 8484 31773 8493 31807
rect 8493 31773 8527 31807
rect 8527 31773 8536 31807
rect 8484 31764 8536 31773
rect 9312 31764 9364 31816
rect 10232 31807 10284 31816
rect 10232 31773 10241 31807
rect 10241 31773 10275 31807
rect 10275 31773 10284 31807
rect 10232 31764 10284 31773
rect 11428 31807 11480 31816
rect 4344 31671 4396 31680
rect 4344 31637 4353 31671
rect 4353 31637 4387 31671
rect 4387 31637 4396 31671
rect 4344 31628 4396 31637
rect 6552 31671 6604 31680
rect 6552 31637 6561 31671
rect 6561 31637 6595 31671
rect 6595 31637 6604 31671
rect 6552 31628 6604 31637
rect 7932 31671 7984 31680
rect 7932 31637 7941 31671
rect 7941 31637 7975 31671
rect 7975 31637 7984 31671
rect 7932 31628 7984 31637
rect 8116 31628 8168 31680
rect 9128 31628 9180 31680
rect 9404 31628 9456 31680
rect 9496 31628 9548 31680
rect 11428 31773 11436 31807
rect 11436 31773 11470 31807
rect 11470 31773 11480 31807
rect 11428 31764 11480 31773
rect 11520 31807 11572 31816
rect 11520 31773 11529 31807
rect 11529 31773 11563 31807
rect 11563 31773 11572 31807
rect 11520 31764 11572 31773
rect 12440 31764 12492 31816
rect 12624 31807 12676 31816
rect 12624 31773 12633 31807
rect 12633 31773 12667 31807
rect 12667 31773 12676 31807
rect 12624 31764 12676 31773
rect 12900 31807 12952 31816
rect 12900 31773 12909 31807
rect 12909 31773 12943 31807
rect 12943 31773 12952 31807
rect 12900 31764 12952 31773
rect 12992 31807 13044 31816
rect 12992 31773 13001 31807
rect 13001 31773 13035 31807
rect 13035 31773 13044 31807
rect 12992 31764 13044 31773
rect 11060 31671 11112 31680
rect 11060 31637 11069 31671
rect 11069 31637 11103 31671
rect 11103 31637 11112 31671
rect 11060 31628 11112 31637
rect 13360 31628 13412 31680
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 4712 31424 4764 31476
rect 4804 31424 4856 31476
rect 7012 31424 7064 31476
rect 4344 31356 4396 31408
rect 5172 31331 5224 31340
rect 5172 31297 5181 31331
rect 5181 31297 5215 31331
rect 5215 31297 5224 31331
rect 5172 31288 5224 31297
rect 6828 31356 6880 31408
rect 6920 31356 6972 31408
rect 8484 31424 8536 31476
rect 9312 31467 9364 31476
rect 9312 31433 9321 31467
rect 9321 31433 9355 31467
rect 9355 31433 9364 31467
rect 9312 31424 9364 31433
rect 6184 31331 6236 31340
rect 6184 31297 6193 31331
rect 6193 31297 6227 31331
rect 6227 31297 6236 31331
rect 6184 31288 6236 31297
rect 6368 31288 6420 31340
rect 6460 31331 6512 31340
rect 6460 31297 6469 31331
rect 6469 31297 6503 31331
rect 6503 31297 6512 31331
rect 6460 31288 6512 31297
rect 6736 31331 6788 31340
rect 6736 31297 6770 31331
rect 6770 31297 6788 31331
rect 6736 31288 6788 31297
rect 10876 31356 10928 31408
rect 8208 31331 8260 31340
rect 8208 31297 8242 31331
rect 8242 31297 8260 31331
rect 8208 31288 8260 31297
rect 9128 31288 9180 31340
rect 9956 31288 10008 31340
rect 11520 31288 11572 31340
rect 13176 31356 13228 31408
rect 13360 31399 13412 31408
rect 13360 31365 13394 31399
rect 13394 31365 13412 31399
rect 13360 31356 13412 31365
rect 13544 31356 13596 31408
rect 4712 31263 4764 31272
rect 4712 31229 4721 31263
rect 4721 31229 4755 31263
rect 4755 31229 4764 31263
rect 4712 31220 4764 31229
rect 5632 31220 5684 31272
rect 9404 31220 9456 31272
rect 12992 31220 13044 31272
rect 8944 31152 8996 31204
rect 12624 31152 12676 31204
rect 12808 31152 12860 31204
rect 5540 31084 5592 31136
rect 10692 31084 10744 31136
rect 10784 31084 10836 31136
rect 12992 31084 13044 31136
rect 14096 31084 14148 31136
rect 14464 31127 14516 31136
rect 14464 31093 14473 31127
rect 14473 31093 14507 31127
rect 14507 31093 14516 31127
rect 14464 31084 14516 31093
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 6736 30880 6788 30932
rect 8208 30923 8260 30932
rect 8208 30889 8217 30923
rect 8217 30889 8251 30923
rect 8251 30889 8260 30923
rect 8208 30880 8260 30889
rect 9404 30880 9456 30932
rect 11060 30880 11112 30932
rect 12808 30880 12860 30932
rect 13268 30880 13320 30932
rect 3700 30744 3752 30796
rect 3884 30676 3936 30728
rect 5172 30744 5224 30796
rect 6552 30744 6604 30796
rect 8944 30812 8996 30864
rect 10784 30812 10836 30864
rect 5356 30676 5408 30728
rect 8024 30719 8076 30728
rect 8024 30685 8058 30719
rect 8058 30685 8076 30719
rect 8024 30676 8076 30685
rect 8392 30608 8444 30660
rect 3148 30540 3200 30592
rect 4804 30540 4856 30592
rect 7012 30540 7064 30592
rect 7932 30583 7984 30592
rect 7932 30549 7941 30583
rect 7941 30549 7975 30583
rect 7975 30549 7984 30583
rect 11152 30744 11204 30796
rect 12992 30812 13044 30864
rect 13452 30812 13504 30864
rect 11704 30787 11756 30796
rect 11704 30753 11713 30787
rect 11713 30753 11747 30787
rect 11747 30753 11756 30787
rect 11704 30744 11756 30753
rect 12164 30744 12216 30796
rect 9312 30676 9364 30728
rect 9956 30719 10008 30728
rect 9956 30685 9965 30719
rect 9965 30685 9999 30719
rect 9999 30685 10008 30719
rect 9956 30676 10008 30685
rect 10232 30719 10284 30728
rect 10232 30685 10241 30719
rect 10241 30685 10275 30719
rect 10275 30685 10284 30719
rect 10232 30676 10284 30685
rect 10692 30719 10744 30728
rect 10692 30685 10701 30719
rect 10701 30685 10735 30719
rect 10735 30685 10744 30719
rect 10692 30676 10744 30685
rect 10968 30719 11020 30728
rect 10968 30685 10977 30719
rect 10977 30685 11011 30719
rect 11011 30685 11020 30719
rect 10968 30676 11020 30685
rect 7932 30540 7984 30549
rect 9312 30540 9364 30592
rect 9496 30583 9548 30592
rect 9496 30549 9505 30583
rect 9505 30549 9539 30583
rect 9539 30549 9548 30583
rect 9496 30540 9548 30549
rect 10784 30583 10836 30592
rect 10784 30549 10793 30583
rect 10793 30549 10827 30583
rect 10827 30549 10836 30583
rect 10784 30540 10836 30549
rect 11336 30719 11388 30728
rect 11336 30685 11345 30719
rect 11345 30685 11379 30719
rect 11379 30685 11388 30719
rect 11336 30676 11388 30685
rect 11796 30719 11848 30728
rect 11796 30685 11805 30719
rect 11805 30685 11839 30719
rect 11839 30685 11848 30719
rect 11796 30676 11848 30685
rect 12440 30719 12492 30728
rect 12440 30685 12449 30719
rect 12449 30685 12483 30719
rect 12483 30685 12492 30719
rect 12440 30676 12492 30685
rect 12808 30719 12860 30728
rect 12808 30685 12817 30719
rect 12817 30685 12851 30719
rect 12851 30685 12860 30719
rect 12808 30676 12860 30685
rect 14004 30744 14056 30796
rect 14096 30787 14148 30796
rect 14096 30753 14105 30787
rect 14105 30753 14139 30787
rect 14139 30753 14148 30787
rect 14096 30744 14148 30753
rect 13268 30676 13320 30728
rect 13452 30719 13504 30728
rect 13452 30685 13461 30719
rect 13461 30685 13495 30719
rect 13495 30685 13504 30719
rect 13452 30676 13504 30685
rect 11244 30540 11296 30592
rect 13084 30540 13136 30592
rect 14096 30540 14148 30592
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 2964 30311 3016 30320
rect 2964 30277 2973 30311
rect 2973 30277 3007 30311
rect 3007 30277 3016 30311
rect 2964 30268 3016 30277
rect 3884 30336 3936 30388
rect 5356 30336 5408 30388
rect 5540 30336 5592 30388
rect 8484 30336 8536 30388
rect 3700 30268 3752 30320
rect 4712 30268 4764 30320
rect 6368 30268 6420 30320
rect 8300 30200 8352 30252
rect 9956 30336 10008 30388
rect 12624 30311 12676 30320
rect 12624 30277 12633 30311
rect 12633 30277 12667 30311
rect 12667 30277 12676 30311
rect 12624 30268 12676 30277
rect 12808 30336 12860 30388
rect 13360 30379 13412 30388
rect 13360 30345 13369 30379
rect 13369 30345 13403 30379
rect 13403 30345 13412 30379
rect 13360 30336 13412 30345
rect 13176 30268 13228 30320
rect 14096 30311 14148 30320
rect 9128 30200 9180 30252
rect 9404 30243 9456 30252
rect 9404 30209 9413 30243
rect 9413 30209 9447 30243
rect 9447 30209 9456 30243
rect 9404 30200 9456 30209
rect 9864 30200 9916 30252
rect 11060 30243 11112 30252
rect 11060 30209 11069 30243
rect 11069 30209 11103 30243
rect 11103 30209 11112 30243
rect 11060 30200 11112 30209
rect 11336 30200 11388 30252
rect 11796 30200 11848 30252
rect 5632 30064 5684 30116
rect 6276 30064 6328 30116
rect 12164 30200 12216 30252
rect 12440 30200 12492 30252
rect 14096 30277 14105 30311
rect 14105 30277 14139 30311
rect 14139 30277 14148 30311
rect 14096 30268 14148 30277
rect 3148 30039 3200 30048
rect 3148 30005 3157 30039
rect 3157 30005 3191 30039
rect 3191 30005 3200 30039
rect 3148 29996 3200 30005
rect 8484 30039 8536 30048
rect 8484 30005 8493 30039
rect 8493 30005 8527 30039
rect 8527 30005 8536 30039
rect 8484 29996 8536 30005
rect 8760 30039 8812 30048
rect 8760 30005 8769 30039
rect 8769 30005 8803 30039
rect 8803 30005 8812 30039
rect 8760 29996 8812 30005
rect 9312 30064 9364 30116
rect 9588 30064 9640 30116
rect 9496 29996 9548 30048
rect 11244 30039 11296 30048
rect 11244 30005 11253 30039
rect 11253 30005 11287 30039
rect 11287 30005 11296 30039
rect 11244 29996 11296 30005
rect 11428 29996 11480 30048
rect 12440 30064 12492 30116
rect 13176 30132 13228 30184
rect 13728 30132 13780 30184
rect 13636 30064 13688 30116
rect 12348 30039 12400 30048
rect 12348 30005 12357 30039
rect 12357 30005 12391 30039
rect 12391 30005 12400 30039
rect 12348 29996 12400 30005
rect 12624 29996 12676 30048
rect 14464 30200 14516 30252
rect 14004 30064 14056 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 8484 29835 8536 29844
rect 8484 29801 8493 29835
rect 8493 29801 8527 29835
rect 8527 29801 8536 29835
rect 8484 29792 8536 29801
rect 10416 29792 10468 29844
rect 3700 29656 3752 29708
rect 2228 29631 2280 29640
rect 2228 29597 2237 29631
rect 2237 29597 2271 29631
rect 2271 29597 2280 29631
rect 2228 29588 2280 29597
rect 4712 29656 4764 29708
rect 5816 29656 5868 29708
rect 2504 29563 2556 29572
rect 2504 29529 2538 29563
rect 2538 29529 2556 29563
rect 2504 29520 2556 29529
rect 6184 29631 6236 29640
rect 6184 29597 6192 29631
rect 6192 29597 6226 29631
rect 6226 29597 6236 29631
rect 6184 29588 6236 29597
rect 6276 29631 6328 29640
rect 6276 29597 6285 29631
rect 6285 29597 6319 29631
rect 6319 29597 6328 29631
rect 6276 29588 6328 29597
rect 6368 29588 6420 29640
rect 7012 29699 7064 29708
rect 7012 29665 7021 29699
rect 7021 29665 7055 29699
rect 7055 29665 7064 29699
rect 7012 29656 7064 29665
rect 9404 29724 9456 29776
rect 11244 29792 11296 29844
rect 8760 29656 8812 29708
rect 6828 29588 6880 29640
rect 7380 29588 7432 29640
rect 8576 29631 8628 29640
rect 8576 29597 8585 29631
rect 8585 29597 8619 29631
rect 8619 29597 8628 29631
rect 8576 29588 8628 29597
rect 9496 29631 9548 29640
rect 9496 29597 9505 29631
rect 9505 29597 9539 29631
rect 9539 29597 9548 29631
rect 9496 29588 9548 29597
rect 10416 29699 10468 29708
rect 10416 29665 10425 29699
rect 10425 29665 10459 29699
rect 10459 29665 10468 29699
rect 10416 29656 10468 29665
rect 10692 29631 10744 29640
rect 10692 29597 10699 29631
rect 10699 29597 10744 29631
rect 3608 29495 3660 29504
rect 3608 29461 3617 29495
rect 3617 29461 3651 29495
rect 3651 29461 3660 29495
rect 3608 29452 3660 29461
rect 3792 29495 3844 29504
rect 3792 29461 3801 29495
rect 3801 29461 3835 29495
rect 3835 29461 3844 29495
rect 3792 29452 3844 29461
rect 3884 29452 3936 29504
rect 5356 29452 5408 29504
rect 5540 29495 5592 29504
rect 5540 29461 5549 29495
rect 5549 29461 5583 29495
rect 5583 29461 5592 29495
rect 5540 29452 5592 29461
rect 8668 29520 8720 29572
rect 10232 29520 10284 29572
rect 10692 29588 10744 29597
rect 10784 29631 10836 29640
rect 10784 29597 10793 29631
rect 10793 29597 10827 29631
rect 10827 29597 10836 29631
rect 10784 29588 10836 29597
rect 12900 29724 12952 29776
rect 13176 29724 13228 29776
rect 10876 29563 10928 29572
rect 10876 29529 10885 29563
rect 10885 29529 10919 29563
rect 10919 29529 10928 29563
rect 10876 29520 10928 29529
rect 10600 29452 10652 29504
rect 11980 29588 12032 29640
rect 12348 29588 12400 29640
rect 13452 29631 13504 29640
rect 13452 29597 13461 29631
rect 13461 29597 13495 29631
rect 13495 29597 13504 29631
rect 13452 29588 13504 29597
rect 13636 29631 13688 29640
rect 13636 29597 13645 29631
rect 13645 29597 13679 29631
rect 13679 29597 13688 29631
rect 13636 29588 13688 29597
rect 14832 29588 14884 29640
rect 11612 29520 11664 29572
rect 12164 29520 12216 29572
rect 12900 29452 12952 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 2504 29291 2556 29300
rect 2504 29257 2513 29291
rect 2513 29257 2547 29291
rect 2547 29257 2556 29291
rect 2504 29248 2556 29257
rect 2964 29248 3016 29300
rect 3700 29248 3752 29300
rect 4712 29248 4764 29300
rect 3608 29223 3660 29232
rect 3608 29189 3617 29223
rect 3617 29189 3651 29223
rect 3651 29189 3660 29223
rect 3608 29180 3660 29189
rect 4804 29155 4856 29164
rect 4804 29121 4813 29155
rect 4813 29121 4847 29155
rect 4847 29121 4856 29155
rect 4804 29112 4856 29121
rect 4896 29112 4948 29164
rect 5540 29180 5592 29232
rect 6368 29291 6420 29300
rect 6368 29257 6377 29291
rect 6377 29257 6411 29291
rect 6411 29257 6420 29291
rect 6368 29248 6420 29257
rect 9404 29248 9456 29300
rect 10600 29291 10652 29300
rect 10600 29257 10609 29291
rect 10609 29257 10643 29291
rect 10643 29257 10652 29291
rect 10600 29248 10652 29257
rect 10692 29291 10744 29300
rect 10692 29257 10701 29291
rect 10701 29257 10735 29291
rect 10735 29257 10744 29291
rect 10692 29248 10744 29257
rect 12992 29248 13044 29300
rect 5356 29155 5408 29164
rect 5356 29121 5365 29155
rect 5365 29121 5399 29155
rect 5399 29121 5408 29155
rect 5356 29112 5408 29121
rect 7196 29112 7248 29164
rect 8300 29155 8352 29164
rect 8300 29121 8309 29155
rect 8309 29121 8343 29155
rect 8343 29121 8352 29155
rect 8300 29112 8352 29121
rect 8484 29112 8536 29164
rect 10232 29155 10284 29164
rect 10232 29121 10241 29155
rect 10241 29121 10275 29155
rect 10275 29121 10284 29155
rect 10232 29112 10284 29121
rect 10600 29112 10652 29164
rect 11428 29180 11480 29232
rect 11704 29180 11756 29232
rect 5448 29044 5500 29096
rect 7748 29087 7800 29096
rect 7748 29053 7757 29087
rect 7757 29053 7791 29087
rect 7791 29053 7800 29087
rect 7748 29044 7800 29053
rect 11796 29155 11848 29164
rect 11796 29121 11805 29155
rect 11805 29121 11839 29155
rect 11839 29121 11848 29155
rect 11796 29112 11848 29121
rect 11980 29155 12032 29164
rect 11980 29121 11989 29155
rect 11989 29121 12023 29155
rect 12023 29121 12032 29155
rect 11980 29112 12032 29121
rect 12164 29155 12216 29164
rect 12164 29121 12173 29155
rect 12173 29121 12207 29155
rect 12207 29121 12216 29155
rect 12164 29112 12216 29121
rect 12716 29180 12768 29232
rect 14832 29291 14884 29300
rect 14832 29257 14841 29291
rect 14841 29257 14875 29291
rect 14875 29257 14884 29291
rect 14832 29248 14884 29257
rect 12072 29044 12124 29096
rect 12808 29112 12860 29164
rect 13084 29112 13136 29164
rect 12716 29087 12768 29096
rect 12716 29053 12725 29087
rect 12725 29053 12759 29087
rect 12759 29053 12768 29087
rect 12716 29044 12768 29053
rect 12900 29044 12952 29096
rect 13452 29087 13504 29096
rect 13452 29053 13461 29087
rect 13461 29053 13495 29087
rect 13495 29053 13504 29087
rect 13452 29044 13504 29053
rect 3240 29019 3292 29028
rect 3240 28985 3249 29019
rect 3249 28985 3283 29019
rect 3283 28985 3292 29019
rect 3240 28976 3292 28985
rect 3792 28976 3844 29028
rect 6736 28976 6788 29028
rect 3884 28908 3936 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 4804 28704 4856 28756
rect 5816 28704 5868 28756
rect 7196 28747 7248 28756
rect 7196 28713 7205 28747
rect 7205 28713 7239 28747
rect 7239 28713 7248 28747
rect 7196 28704 7248 28713
rect 10232 28704 10284 28756
rect 11060 28704 11112 28756
rect 4252 28636 4304 28688
rect 5356 28636 5408 28688
rect 7840 28636 7892 28688
rect 13360 28636 13412 28688
rect 3976 28568 4028 28620
rect 4068 28543 4120 28552
rect 4068 28509 4077 28543
rect 4077 28509 4111 28543
rect 4111 28509 4120 28543
rect 4068 28500 4120 28509
rect 4252 28543 4304 28552
rect 4252 28509 4261 28543
rect 4261 28509 4295 28543
rect 4295 28509 4304 28543
rect 4252 28500 4304 28509
rect 4344 28500 4396 28552
rect 4712 28543 4764 28552
rect 4712 28509 4721 28543
rect 4721 28509 4755 28543
rect 4755 28509 4764 28543
rect 4712 28500 4764 28509
rect 6920 28611 6972 28620
rect 6920 28577 6929 28611
rect 6929 28577 6963 28611
rect 6963 28577 6972 28611
rect 6920 28568 6972 28577
rect 7012 28611 7064 28620
rect 7012 28577 7046 28611
rect 7046 28577 7064 28611
rect 7012 28568 7064 28577
rect 8208 28500 8260 28552
rect 3700 28364 3752 28416
rect 4804 28364 4856 28416
rect 7932 28432 7984 28484
rect 8392 28432 8444 28484
rect 10508 28500 10560 28552
rect 10600 28543 10652 28552
rect 10600 28509 10609 28543
rect 10609 28509 10643 28543
rect 10643 28509 10652 28543
rect 10600 28500 10652 28509
rect 11520 28500 11572 28552
rect 13452 28568 13504 28620
rect 10692 28432 10744 28484
rect 11428 28432 11480 28484
rect 11888 28475 11940 28484
rect 11888 28441 11897 28475
rect 11897 28441 11931 28475
rect 11931 28441 11940 28475
rect 11888 28432 11940 28441
rect 12348 28432 12400 28484
rect 13176 28543 13228 28552
rect 13176 28509 13185 28543
rect 13185 28509 13219 28543
rect 13219 28509 13228 28543
rect 13176 28500 13228 28509
rect 13820 28500 13872 28552
rect 12624 28432 12676 28484
rect 13544 28432 13596 28484
rect 13728 28432 13780 28484
rect 6276 28364 6328 28416
rect 12900 28407 12952 28416
rect 12900 28373 12909 28407
rect 12909 28373 12943 28407
rect 12943 28373 12952 28407
rect 12900 28364 12952 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 3608 28160 3660 28212
rect 4068 28160 4120 28212
rect 8668 28160 8720 28212
rect 10600 28160 10652 28212
rect 11520 28203 11572 28212
rect 11520 28169 11529 28203
rect 11529 28169 11563 28203
rect 11563 28169 11572 28203
rect 11520 28160 11572 28169
rect 13728 28160 13780 28212
rect 3240 28067 3292 28076
rect 3240 28033 3249 28067
rect 3249 28033 3283 28067
rect 3283 28033 3292 28067
rect 3240 28024 3292 28033
rect 3884 28024 3936 28076
rect 4252 28092 4304 28144
rect 5264 28092 5316 28144
rect 3792 27956 3844 28008
rect 4344 28067 4396 28076
rect 4344 28033 4353 28067
rect 4353 28033 4387 28067
rect 4387 28033 4396 28067
rect 4344 28024 4396 28033
rect 6276 28092 6328 28144
rect 7748 28092 7800 28144
rect 4620 27956 4672 28008
rect 5724 27999 5776 28008
rect 5724 27965 5733 27999
rect 5733 27965 5767 27999
rect 5767 27965 5776 27999
rect 5724 27956 5776 27965
rect 3700 27888 3752 27940
rect 6368 28067 6420 28076
rect 6368 28033 6377 28067
rect 6377 28033 6411 28067
rect 6411 28033 6420 28067
rect 6368 28024 6420 28033
rect 6736 28024 6788 28076
rect 7380 28067 7432 28076
rect 7380 28033 7389 28067
rect 7389 28033 7423 28067
rect 7423 28033 7432 28067
rect 8484 28092 8536 28144
rect 7380 28024 7432 28033
rect 8300 28067 8352 28076
rect 8300 28033 8309 28067
rect 8309 28033 8343 28067
rect 8343 28033 8352 28067
rect 8300 28024 8352 28033
rect 9864 28067 9916 28076
rect 9864 28033 9882 28067
rect 9882 28033 9916 28067
rect 9864 28024 9916 28033
rect 10324 28092 10376 28144
rect 10416 28024 10468 28076
rect 10508 28024 10560 28076
rect 10692 28067 10744 28076
rect 10692 28033 10701 28067
rect 10701 28033 10735 28067
rect 10735 28033 10744 28067
rect 10692 28024 10744 28033
rect 11704 28067 11756 28076
rect 11704 28033 11713 28067
rect 11713 28033 11747 28067
rect 11747 28033 11756 28067
rect 11704 28024 11756 28033
rect 10140 27999 10192 28008
rect 10140 27965 10149 27999
rect 10149 27965 10183 27999
rect 10183 27965 10192 27999
rect 10140 27956 10192 27965
rect 12900 28092 12952 28144
rect 12072 28024 12124 28076
rect 12348 27956 12400 28008
rect 8392 27888 8444 27940
rect 3884 27863 3936 27872
rect 3884 27829 3893 27863
rect 3893 27829 3927 27863
rect 3927 27829 3936 27863
rect 3884 27820 3936 27829
rect 3976 27820 4028 27872
rect 4712 27820 4764 27872
rect 6276 27820 6328 27872
rect 6920 27863 6972 27872
rect 6920 27829 6929 27863
rect 6929 27829 6963 27863
rect 6963 27829 6972 27863
rect 6920 27820 6972 27829
rect 7564 27863 7616 27872
rect 7564 27829 7573 27863
rect 7573 27829 7607 27863
rect 7607 27829 7616 27863
rect 7564 27820 7616 27829
rect 7932 27820 7984 27872
rect 9128 27820 9180 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 3976 27616 4028 27668
rect 5724 27616 5776 27668
rect 8484 27616 8536 27668
rect 9496 27616 9548 27668
rect 4068 27548 4120 27600
rect 8300 27548 8352 27600
rect 8944 27548 8996 27600
rect 9864 27616 9916 27668
rect 2228 27523 2280 27532
rect 2228 27489 2237 27523
rect 2237 27489 2271 27523
rect 2271 27489 2280 27523
rect 2228 27480 2280 27489
rect 6368 27480 6420 27532
rect 3056 27412 3108 27464
rect 4620 27412 4672 27464
rect 5816 27412 5868 27464
rect 6276 27455 6328 27464
rect 6276 27421 6285 27455
rect 6285 27421 6319 27455
rect 6319 27421 6328 27455
rect 6276 27412 6328 27421
rect 2688 27344 2740 27396
rect 3516 27344 3568 27396
rect 7472 27344 7524 27396
rect 8668 27480 8720 27532
rect 9680 27591 9732 27600
rect 9680 27557 9689 27591
rect 9689 27557 9723 27591
rect 9723 27557 9732 27591
rect 9680 27548 9732 27557
rect 8576 27387 8628 27396
rect 8576 27353 8617 27387
rect 8617 27353 8628 27387
rect 8576 27344 8628 27353
rect 2964 27276 3016 27328
rect 4068 27319 4120 27328
rect 4068 27285 4077 27319
rect 4077 27285 4111 27319
rect 4111 27285 4120 27319
rect 4068 27276 4120 27285
rect 4804 27276 4856 27328
rect 8208 27276 8260 27328
rect 9128 27412 9180 27464
rect 9312 27412 9364 27464
rect 10140 27523 10192 27532
rect 10140 27489 10149 27523
rect 10149 27489 10183 27523
rect 10183 27489 10192 27523
rect 10140 27480 10192 27489
rect 10784 27480 10836 27532
rect 11152 27412 11204 27464
rect 11704 27412 11756 27464
rect 9036 27344 9088 27396
rect 9588 27344 9640 27396
rect 10232 27344 10284 27396
rect 11428 27344 11480 27396
rect 11796 27344 11848 27396
rect 12256 27344 12308 27396
rect 9312 27319 9364 27328
rect 9312 27285 9321 27319
rect 9321 27285 9355 27319
rect 9355 27285 9364 27319
rect 9312 27276 9364 27285
rect 9772 27276 9824 27328
rect 10600 27276 10652 27328
rect 11612 27319 11664 27328
rect 11612 27285 11621 27319
rect 11621 27285 11655 27319
rect 11655 27285 11664 27319
rect 11612 27276 11664 27285
rect 12072 27276 12124 27328
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 2688 27115 2740 27124
rect 2688 27081 2697 27115
rect 2697 27081 2731 27115
rect 2731 27081 2740 27115
rect 2688 27072 2740 27081
rect 2964 27072 3016 27124
rect 3608 27047 3660 27056
rect 3608 27013 3617 27047
rect 3617 27013 3651 27047
rect 3651 27013 3660 27047
rect 3608 27004 3660 27013
rect 4068 27047 4120 27056
rect 4068 27013 4077 27047
rect 4077 27013 4111 27047
rect 4111 27013 4120 27047
rect 4068 27004 4120 27013
rect 7472 27072 7524 27124
rect 7840 27115 7892 27124
rect 7840 27081 7849 27115
rect 7849 27081 7883 27115
rect 7883 27081 7892 27115
rect 7840 27072 7892 27081
rect 7932 27115 7984 27124
rect 7932 27081 7941 27115
rect 7941 27081 7975 27115
rect 7975 27081 7984 27115
rect 7932 27072 7984 27081
rect 8392 27072 8444 27124
rect 8484 27072 8536 27124
rect 9036 27115 9088 27124
rect 9036 27081 9045 27115
rect 9045 27081 9079 27115
rect 9079 27081 9088 27115
rect 9036 27072 9088 27081
rect 10416 27072 10468 27124
rect 12624 27072 12676 27124
rect 5540 27004 5592 27056
rect 10232 27004 10284 27056
rect 10692 27004 10744 27056
rect 12440 27004 12492 27056
rect 12716 27004 12768 27056
rect 3792 26979 3844 26988
rect 3792 26945 3801 26979
rect 3801 26945 3835 26979
rect 3835 26945 3844 26979
rect 3792 26936 3844 26945
rect 4068 26868 4120 26920
rect 3700 26800 3752 26852
rect 848 26732 900 26784
rect 3884 26732 3936 26784
rect 4620 26936 4672 26988
rect 7564 26936 7616 26988
rect 8484 26979 8536 26988
rect 8484 26945 8493 26979
rect 8493 26945 8527 26979
rect 8527 26945 8536 26979
rect 8484 26936 8536 26945
rect 5816 26868 5868 26920
rect 8208 26911 8260 26920
rect 8208 26877 8217 26911
rect 8217 26877 8251 26911
rect 8251 26877 8260 26911
rect 8208 26868 8260 26877
rect 8668 26936 8720 26988
rect 8944 26979 8996 26988
rect 8944 26945 8953 26979
rect 8953 26945 8987 26979
rect 8987 26945 8996 26979
rect 8944 26936 8996 26945
rect 9680 26936 9732 26988
rect 10140 26979 10192 26988
rect 10140 26945 10149 26979
rect 10149 26945 10183 26979
rect 10183 26945 10192 26979
rect 10140 26936 10192 26945
rect 11612 26936 11664 26988
rect 12072 26979 12124 26988
rect 12072 26945 12081 26979
rect 12081 26945 12115 26979
rect 12115 26945 12124 26979
rect 12072 26936 12124 26945
rect 8392 26732 8444 26784
rect 9588 26868 9640 26920
rect 13820 26936 13872 26988
rect 13912 26936 13964 26988
rect 9128 26800 9180 26852
rect 12440 26911 12492 26920
rect 12440 26877 12449 26911
rect 12449 26877 12483 26911
rect 12483 26877 12492 26911
rect 12440 26868 12492 26877
rect 12716 26911 12768 26920
rect 12716 26877 12725 26911
rect 12725 26877 12759 26911
rect 12759 26877 12768 26911
rect 12716 26868 12768 26877
rect 13084 26868 13136 26920
rect 11704 26800 11756 26852
rect 9772 26732 9824 26784
rect 12164 26732 12216 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 7012 26528 7064 26580
rect 7840 26528 7892 26580
rect 9312 26528 9364 26580
rect 11612 26571 11664 26580
rect 11612 26537 11621 26571
rect 11621 26537 11655 26571
rect 11655 26537 11664 26571
rect 11612 26528 11664 26537
rect 11704 26528 11756 26580
rect 5264 26503 5316 26512
rect 5264 26469 5273 26503
rect 5273 26469 5307 26503
rect 5307 26469 5316 26503
rect 5264 26460 5316 26469
rect 11428 26460 11480 26512
rect 8208 26392 8260 26444
rect 4620 26324 4672 26376
rect 4804 26324 4856 26376
rect 5816 26324 5868 26376
rect 5356 26256 5408 26308
rect 6920 26324 6972 26376
rect 9128 26367 9180 26376
rect 9128 26333 9137 26367
rect 9137 26333 9171 26367
rect 9171 26333 9180 26367
rect 9128 26324 9180 26333
rect 10324 26435 10376 26444
rect 10324 26401 10333 26435
rect 10333 26401 10367 26435
rect 10367 26401 10376 26435
rect 10324 26392 10376 26401
rect 10416 26435 10468 26444
rect 10416 26401 10425 26435
rect 10425 26401 10459 26435
rect 10459 26401 10468 26435
rect 10416 26392 10468 26401
rect 10692 26324 10744 26376
rect 10784 26367 10836 26376
rect 10784 26333 10793 26367
rect 10793 26333 10827 26367
rect 10827 26333 10836 26367
rect 10784 26324 10836 26333
rect 6368 26299 6420 26308
rect 6368 26265 6402 26299
rect 6402 26265 6420 26299
rect 4252 26188 4304 26240
rect 6368 26256 6420 26265
rect 11152 26367 11204 26376
rect 11152 26333 11161 26367
rect 11161 26333 11195 26367
rect 11195 26333 11204 26367
rect 11152 26324 11204 26333
rect 12072 26571 12124 26580
rect 12072 26537 12081 26571
rect 12081 26537 12115 26571
rect 12115 26537 12124 26571
rect 12072 26528 12124 26537
rect 12256 26528 12308 26580
rect 13084 26528 13136 26580
rect 11796 26299 11848 26308
rect 11796 26265 11823 26299
rect 11823 26265 11848 26299
rect 11796 26256 11848 26265
rect 11980 26299 12032 26308
rect 11980 26265 11989 26299
rect 11989 26265 12023 26299
rect 12023 26265 12032 26299
rect 11980 26256 12032 26265
rect 7932 26188 7984 26240
rect 10692 26231 10744 26240
rect 10692 26197 10701 26231
rect 10701 26197 10735 26231
rect 10735 26197 10744 26231
rect 10692 26188 10744 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 3516 25984 3568 26036
rect 4712 25984 4764 26036
rect 8208 25916 8260 25968
rect 9312 25984 9364 26036
rect 11152 25984 11204 26036
rect 11980 25984 12032 26036
rect 9036 25916 9088 25968
rect 10692 25916 10744 25968
rect 7012 25848 7064 25900
rect 7840 25848 7892 25900
rect 7932 25891 7984 25900
rect 7932 25857 7941 25891
rect 7941 25857 7975 25891
rect 7975 25857 7984 25891
rect 7932 25848 7984 25857
rect 8392 25891 8444 25900
rect 8392 25857 8401 25891
rect 8401 25857 8435 25891
rect 8435 25857 8444 25891
rect 8392 25848 8444 25857
rect 4620 25823 4672 25832
rect 4620 25789 4629 25823
rect 4629 25789 4663 25823
rect 4663 25789 4672 25823
rect 4620 25780 4672 25789
rect 5632 25823 5684 25832
rect 5632 25789 5641 25823
rect 5641 25789 5675 25823
rect 5675 25789 5684 25823
rect 5632 25780 5684 25789
rect 8484 25823 8536 25832
rect 8484 25789 8493 25823
rect 8493 25789 8527 25823
rect 8527 25789 8536 25823
rect 8484 25780 8536 25789
rect 10048 25848 10100 25900
rect 12348 25916 12400 25968
rect 13268 25916 13320 25968
rect 13728 25916 13780 25968
rect 11980 25891 12032 25900
rect 11980 25857 12014 25891
rect 12014 25857 12032 25891
rect 11980 25848 12032 25857
rect 6368 25755 6420 25764
rect 6368 25721 6377 25755
rect 6377 25721 6411 25755
rect 6411 25721 6420 25755
rect 6368 25712 6420 25721
rect 8208 25712 8260 25764
rect 4252 25644 4304 25696
rect 4712 25644 4764 25696
rect 5356 25644 5408 25696
rect 6000 25644 6052 25696
rect 7012 25687 7064 25696
rect 7012 25653 7021 25687
rect 7021 25653 7055 25687
rect 7055 25653 7064 25687
rect 7012 25644 7064 25653
rect 7564 25644 7616 25696
rect 9496 25687 9548 25696
rect 9496 25653 9505 25687
rect 9505 25653 9539 25687
rect 9539 25653 9548 25687
rect 9496 25644 9548 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 10600 25483 10652 25492
rect 10600 25449 10609 25483
rect 10609 25449 10643 25483
rect 10643 25449 10652 25483
rect 10600 25440 10652 25449
rect 11980 25440 12032 25492
rect 6920 25372 6972 25424
rect 5264 25304 5316 25356
rect 5816 25236 5868 25288
rect 6000 25279 6052 25288
rect 6000 25245 6034 25279
rect 6034 25245 6052 25279
rect 6000 25236 6052 25245
rect 4160 25168 4212 25220
rect 6552 25236 6604 25288
rect 7104 25236 7156 25288
rect 3792 25143 3844 25152
rect 3792 25109 3801 25143
rect 3801 25109 3835 25143
rect 3835 25109 3844 25143
rect 3792 25100 3844 25109
rect 6552 25100 6604 25152
rect 7564 25279 7616 25288
rect 7564 25245 7573 25279
rect 7573 25245 7607 25279
rect 7607 25245 7616 25279
rect 7564 25236 7616 25245
rect 7932 25304 7984 25356
rect 12440 25372 12492 25424
rect 8300 25236 8352 25288
rect 12164 25304 12216 25356
rect 10048 25236 10100 25288
rect 11428 25236 11480 25288
rect 7472 25168 7524 25220
rect 9496 25211 9548 25220
rect 9496 25177 9530 25211
rect 9530 25177 9548 25211
rect 9496 25168 9548 25177
rect 7656 25100 7708 25152
rect 8392 25100 8444 25152
rect 9312 25100 9364 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 4160 24939 4212 24948
rect 4160 24905 4169 24939
rect 4169 24905 4203 24939
rect 4203 24905 4212 24939
rect 4160 24896 4212 24905
rect 5632 24939 5684 24948
rect 5632 24905 5641 24939
rect 5641 24905 5675 24939
rect 5675 24905 5684 24939
rect 5632 24896 5684 24905
rect 5448 24760 5500 24812
rect 7564 24828 7616 24880
rect 7472 24760 7524 24812
rect 7656 24803 7708 24812
rect 7656 24769 7665 24803
rect 7665 24769 7699 24803
rect 7699 24769 7708 24803
rect 7656 24760 7708 24769
rect 5908 24735 5960 24744
rect 5908 24701 5917 24735
rect 5917 24701 5951 24735
rect 5951 24701 5960 24735
rect 5908 24692 5960 24701
rect 6460 24692 6512 24744
rect 6828 24692 6880 24744
rect 7288 24735 7340 24744
rect 7288 24701 7297 24735
rect 7297 24701 7331 24735
rect 7331 24701 7340 24735
rect 7288 24692 7340 24701
rect 7564 24692 7616 24744
rect 7748 24735 7800 24744
rect 7748 24701 7757 24735
rect 7757 24701 7791 24735
rect 7791 24701 7800 24735
rect 7748 24692 7800 24701
rect 5816 24624 5868 24676
rect 9128 24624 9180 24676
rect 6368 24556 6420 24608
rect 6828 24556 6880 24608
rect 7196 24599 7248 24608
rect 7196 24565 7205 24599
rect 7205 24565 7239 24599
rect 7239 24565 7248 24599
rect 7196 24556 7248 24565
rect 7380 24556 7432 24608
rect 7564 24556 7616 24608
rect 8208 24556 8260 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 5448 24395 5500 24404
rect 5448 24361 5457 24395
rect 5457 24361 5491 24395
rect 5491 24361 5500 24395
rect 5448 24352 5500 24361
rect 6460 24395 6512 24404
rect 6460 24361 6469 24395
rect 6469 24361 6503 24395
rect 6503 24361 6512 24395
rect 6460 24352 6512 24361
rect 7012 24352 7064 24404
rect 7472 24352 7524 24404
rect 5908 24284 5960 24336
rect 6736 24284 6788 24336
rect 7840 24352 7892 24404
rect 8116 24395 8168 24404
rect 8116 24361 8125 24395
rect 8125 24361 8159 24395
rect 8159 24361 8168 24395
rect 8116 24352 8168 24361
rect 3792 24216 3844 24268
rect 5816 24259 5868 24268
rect 5816 24225 5825 24259
rect 5825 24225 5859 24259
rect 5859 24225 5868 24259
rect 5816 24216 5868 24225
rect 6000 24148 6052 24200
rect 8300 24259 8352 24268
rect 8300 24225 8309 24259
rect 8309 24225 8343 24259
rect 8343 24225 8352 24259
rect 8300 24216 8352 24225
rect 6276 24191 6328 24200
rect 6276 24157 6285 24191
rect 6285 24157 6319 24191
rect 6319 24157 6328 24191
rect 6276 24148 6328 24157
rect 6368 24191 6420 24200
rect 6368 24157 6377 24191
rect 6377 24157 6411 24191
rect 6411 24157 6420 24191
rect 6368 24148 6420 24157
rect 6552 24080 6604 24132
rect 4804 24012 4856 24064
rect 7380 24148 7432 24200
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 10416 24191 10468 24200
rect 10416 24157 10425 24191
rect 10425 24157 10459 24191
rect 10459 24157 10468 24191
rect 10416 24148 10468 24157
rect 11980 24191 12032 24200
rect 11980 24157 11989 24191
rect 11989 24157 12023 24191
rect 12023 24157 12032 24191
rect 11980 24148 12032 24157
rect 12072 24191 12124 24200
rect 12072 24157 12081 24191
rect 12081 24157 12115 24191
rect 12115 24157 12124 24191
rect 12072 24148 12124 24157
rect 7196 24080 7248 24132
rect 7748 24012 7800 24064
rect 8668 24012 8720 24064
rect 11612 24080 11664 24132
rect 12256 24148 12308 24200
rect 9772 24012 9824 24064
rect 10784 24012 10836 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 4620 23808 4672 23860
rect 7748 23808 7800 23860
rect 8208 23808 8260 23860
rect 3056 23715 3108 23724
rect 3056 23681 3065 23715
rect 3065 23681 3099 23715
rect 3099 23681 3108 23715
rect 3056 23672 3108 23681
rect 3148 23672 3200 23724
rect 8116 23715 8168 23724
rect 8116 23681 8125 23715
rect 8125 23681 8159 23715
rect 8159 23681 8168 23715
rect 8116 23672 8168 23681
rect 8392 23715 8444 23724
rect 8392 23681 8401 23715
rect 8401 23681 8435 23715
rect 8435 23681 8444 23715
rect 8392 23672 8444 23681
rect 10048 23740 10100 23792
rect 9772 23715 9824 23724
rect 9772 23681 9806 23715
rect 9806 23681 9824 23715
rect 9772 23672 9824 23681
rect 6644 23536 6696 23588
rect 11888 23672 11940 23724
rect 13176 23672 13228 23724
rect 13268 23715 13320 23724
rect 13268 23681 13277 23715
rect 13277 23681 13311 23715
rect 13311 23681 13320 23715
rect 13268 23672 13320 23681
rect 13820 23672 13872 23724
rect 7472 23511 7524 23520
rect 7472 23477 7481 23511
rect 7481 23477 7515 23511
rect 7515 23477 7524 23511
rect 7472 23468 7524 23477
rect 12164 23468 12216 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 3148 23307 3200 23316
rect 3148 23273 3157 23307
rect 3157 23273 3191 23307
rect 3191 23273 3200 23307
rect 3148 23264 3200 23273
rect 3332 23264 3384 23316
rect 4712 23264 4764 23316
rect 11888 23307 11940 23316
rect 11888 23273 11897 23307
rect 11897 23273 11931 23307
rect 11931 23273 11940 23307
rect 11888 23264 11940 23273
rect 11980 23307 12032 23316
rect 11980 23273 11989 23307
rect 11989 23273 12023 23307
rect 12023 23273 12032 23307
rect 11980 23264 12032 23273
rect 13176 23264 13228 23316
rect 3056 23171 3108 23180
rect 3056 23137 3065 23171
rect 3065 23137 3099 23171
rect 3099 23137 3108 23171
rect 3056 23128 3108 23137
rect 3332 23103 3384 23112
rect 3332 23069 3341 23103
rect 3341 23069 3375 23103
rect 3375 23069 3384 23103
rect 3332 23060 3384 23069
rect 3424 23060 3476 23112
rect 3240 22992 3292 23044
rect 2044 22924 2096 22976
rect 3332 22924 3384 22976
rect 3700 22992 3752 23044
rect 4620 22924 4672 22976
rect 6644 23103 6696 23112
rect 6644 23069 6653 23103
rect 6653 23069 6687 23103
rect 6687 23069 6696 23103
rect 6644 23060 6696 23069
rect 8484 23060 8536 23112
rect 10048 23060 10100 23112
rect 10784 23103 10836 23112
rect 10784 23069 10818 23103
rect 10818 23069 10836 23103
rect 10784 23060 10836 23069
rect 12164 23060 12216 23112
rect 12808 23060 12860 23112
rect 13084 23103 13136 23112
rect 13084 23069 13093 23103
rect 13093 23069 13127 23103
rect 13127 23069 13136 23103
rect 13084 23060 13136 23069
rect 9220 23035 9272 23044
rect 9220 23001 9254 23035
rect 9254 23001 9272 23035
rect 9220 22992 9272 23001
rect 11704 22992 11756 23044
rect 12992 23035 13044 23044
rect 12992 23001 13001 23035
rect 13001 23001 13035 23035
rect 13035 23001 13044 23035
rect 12992 22992 13044 23001
rect 5264 22967 5316 22976
rect 5264 22933 5273 22967
rect 5273 22933 5307 22967
rect 5307 22933 5316 22967
rect 5264 22924 5316 22933
rect 6000 22924 6052 22976
rect 9864 22924 9916 22976
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 3240 22695 3292 22704
rect 3240 22661 3249 22695
rect 3249 22661 3283 22695
rect 3283 22661 3292 22695
rect 6276 22720 6328 22772
rect 10416 22720 10468 22772
rect 11704 22763 11756 22772
rect 11704 22729 11713 22763
rect 11713 22729 11747 22763
rect 11747 22729 11756 22763
rect 11704 22720 11756 22729
rect 12072 22720 12124 22772
rect 3240 22652 3292 22661
rect 3884 22652 3936 22704
rect 5264 22652 5316 22704
rect 848 22584 900 22636
rect 3424 22627 3476 22636
rect 3424 22593 3433 22627
rect 3433 22593 3467 22627
rect 3467 22593 3476 22627
rect 3424 22584 3476 22593
rect 4804 22627 4856 22636
rect 4804 22593 4813 22627
rect 4813 22593 4847 22627
rect 4847 22593 4856 22627
rect 4804 22584 4856 22593
rect 3884 22516 3936 22568
rect 1768 22448 1820 22500
rect 3700 22448 3752 22500
rect 4620 22448 4672 22500
rect 5816 22559 5868 22568
rect 5816 22525 5825 22559
rect 5825 22525 5859 22559
rect 5859 22525 5868 22559
rect 5816 22516 5868 22525
rect 6000 22627 6052 22636
rect 6000 22593 6009 22627
rect 6009 22593 6043 22627
rect 6043 22593 6052 22627
rect 6000 22584 6052 22593
rect 6552 22584 6604 22636
rect 6828 22584 6880 22636
rect 7288 22584 7340 22636
rect 7472 22627 7524 22636
rect 7472 22593 7481 22627
rect 7481 22593 7515 22627
rect 7515 22593 7524 22627
rect 7472 22584 7524 22593
rect 6736 22559 6788 22568
rect 6736 22525 6745 22559
rect 6745 22525 6779 22559
rect 6779 22525 6788 22559
rect 6736 22516 6788 22525
rect 7012 22448 7064 22500
rect 7472 22448 7524 22500
rect 8484 22627 8536 22636
rect 8484 22593 8493 22627
rect 8493 22593 8527 22627
rect 8527 22593 8536 22627
rect 8484 22584 8536 22593
rect 8760 22627 8812 22636
rect 8760 22593 8794 22627
rect 8794 22593 8812 22627
rect 8760 22584 8812 22593
rect 11612 22627 11664 22636
rect 11612 22593 11621 22627
rect 11621 22593 11655 22627
rect 11655 22593 11664 22627
rect 11612 22584 11664 22593
rect 8392 22559 8444 22568
rect 8392 22525 8401 22559
rect 8401 22525 8435 22559
rect 8435 22525 8444 22559
rect 8392 22516 8444 22525
rect 12164 22627 12216 22636
rect 12164 22593 12173 22627
rect 12173 22593 12207 22627
rect 12207 22593 12216 22627
rect 12164 22584 12216 22593
rect 12440 22584 12492 22636
rect 16120 22584 16172 22636
rect 12808 22516 12860 22568
rect 16396 22491 16448 22500
rect 16396 22457 16405 22491
rect 16405 22457 16439 22491
rect 16439 22457 16448 22491
rect 16396 22448 16448 22457
rect 4804 22380 4856 22432
rect 5632 22423 5684 22432
rect 5632 22389 5641 22423
rect 5641 22389 5675 22423
rect 5675 22389 5684 22423
rect 5632 22380 5684 22389
rect 5908 22380 5960 22432
rect 7196 22380 7248 22432
rect 7564 22423 7616 22432
rect 7564 22389 7573 22423
rect 7573 22389 7607 22423
rect 7607 22389 7616 22423
rect 7564 22380 7616 22389
rect 14280 22380 14332 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 9956 22176 10008 22228
rect 16120 22219 16172 22228
rect 16120 22185 16129 22219
rect 16129 22185 16163 22219
rect 16163 22185 16172 22219
rect 16120 22176 16172 22185
rect 8392 22108 8444 22160
rect 12440 22151 12492 22160
rect 12440 22117 12449 22151
rect 12449 22117 12483 22151
rect 12483 22117 12492 22151
rect 12440 22108 12492 22117
rect 7380 22083 7432 22092
rect 7380 22049 7389 22083
rect 7389 22049 7423 22083
rect 7423 22049 7432 22083
rect 7380 22040 7432 22049
rect 848 21972 900 22024
rect 1860 21972 1912 22024
rect 112 21904 164 21956
rect 2780 21972 2832 22024
rect 3056 21972 3108 22024
rect 4712 21972 4764 22024
rect 2320 21879 2372 21888
rect 2320 21845 2329 21879
rect 2329 21845 2363 21879
rect 2363 21845 2372 21879
rect 2320 21836 2372 21845
rect 3792 21904 3844 21956
rect 5816 21836 5868 21888
rect 6552 21836 6604 21888
rect 6736 21879 6788 21888
rect 6736 21845 6745 21879
rect 6745 21845 6779 21879
rect 6779 21845 6788 21879
rect 6736 21836 6788 21845
rect 7012 22015 7064 22024
rect 7012 21981 7021 22015
rect 7021 21981 7055 22015
rect 7055 21981 7064 22015
rect 7012 21972 7064 21981
rect 7196 22015 7248 22024
rect 7196 21981 7205 22015
rect 7205 21981 7239 22015
rect 7239 21981 7248 22015
rect 7196 21972 7248 21981
rect 7288 22015 7340 22024
rect 7288 21981 7294 22015
rect 7294 21981 7328 22015
rect 7328 21981 7340 22015
rect 10048 22040 10100 22092
rect 7288 21972 7340 21981
rect 7380 21904 7432 21956
rect 7656 21947 7708 21956
rect 7656 21913 7690 21947
rect 7690 21913 7708 21947
rect 7656 21904 7708 21913
rect 11336 21972 11388 22024
rect 9864 21947 9916 21956
rect 9864 21913 9873 21947
rect 9873 21913 9907 21947
rect 9907 21913 9916 21947
rect 9864 21904 9916 21913
rect 12532 21972 12584 22024
rect 12992 21972 13044 22024
rect 13820 22015 13872 22024
rect 13820 21981 13829 22015
rect 13829 21981 13863 22015
rect 13863 21981 13872 22015
rect 13820 21972 13872 21981
rect 14372 21972 14424 22024
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 16120 21972 16172 22024
rect 12624 21904 12676 21956
rect 13360 21904 13412 21956
rect 9680 21836 9732 21888
rect 11428 21836 11480 21888
rect 11796 21836 11848 21888
rect 12164 21836 12216 21888
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 13268 21836 13320 21888
rect 16396 21879 16448 21888
rect 16396 21845 16405 21879
rect 16405 21845 16439 21879
rect 16439 21845 16448 21879
rect 16396 21836 16448 21845
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 2872 21632 2924 21684
rect 3056 21632 3108 21684
rect 5632 21564 5684 21616
rect 1768 21496 1820 21548
rect 2044 21539 2096 21548
rect 2044 21505 2053 21539
rect 2053 21505 2087 21539
rect 2087 21505 2096 21539
rect 2044 21496 2096 21505
rect 2780 21539 2832 21548
rect 2780 21505 2789 21539
rect 2789 21505 2823 21539
rect 2823 21505 2832 21539
rect 2780 21496 2832 21505
rect 3056 21539 3108 21548
rect 3056 21505 3090 21539
rect 3090 21505 3108 21539
rect 3056 21496 3108 21505
rect 3884 21496 3936 21548
rect 4620 21496 4672 21548
rect 4712 21539 4764 21548
rect 4712 21505 4721 21539
rect 4721 21505 4755 21539
rect 4755 21505 4764 21539
rect 4712 21496 4764 21505
rect 5724 21496 5776 21548
rect 7012 21632 7064 21684
rect 6736 21564 6788 21616
rect 7656 21675 7708 21684
rect 7656 21641 7665 21675
rect 7665 21641 7699 21675
rect 7699 21641 7708 21675
rect 7656 21632 7708 21641
rect 11336 21675 11388 21684
rect 11336 21641 11345 21675
rect 11345 21641 11379 21675
rect 11379 21641 11388 21675
rect 11336 21632 11388 21641
rect 11428 21632 11480 21684
rect 6644 21496 6696 21548
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 7288 21496 7340 21548
rect 7472 21496 7524 21548
rect 1952 21471 2004 21480
rect 1952 21437 1961 21471
rect 1961 21437 1995 21471
rect 1995 21437 2004 21471
rect 1952 21428 2004 21437
rect 7564 21428 7616 21480
rect 2136 21292 2188 21344
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 9864 21539 9916 21548
rect 9864 21505 9873 21539
rect 9873 21505 9907 21539
rect 9907 21505 9916 21539
rect 9864 21496 9916 21505
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 11152 21539 11204 21548
rect 11152 21505 11161 21539
rect 11161 21505 11195 21539
rect 11195 21505 11204 21539
rect 11152 21496 11204 21505
rect 12532 21632 12584 21684
rect 12624 21564 12676 21616
rect 13084 21564 13136 21616
rect 12348 21496 12400 21548
rect 13452 21496 13504 21548
rect 14372 21539 14424 21548
rect 14372 21505 14381 21539
rect 14381 21505 14415 21539
rect 14415 21505 14424 21539
rect 14372 21496 14424 21505
rect 14648 21539 14700 21548
rect 14648 21505 14682 21539
rect 14682 21505 14700 21539
rect 14648 21496 14700 21505
rect 9772 21428 9824 21480
rect 11244 21360 11296 21412
rect 11796 21471 11848 21480
rect 11796 21437 11805 21471
rect 11805 21437 11839 21471
rect 11839 21437 11848 21471
rect 11796 21428 11848 21437
rect 11980 21471 12032 21480
rect 11980 21437 12014 21471
rect 12014 21437 12032 21471
rect 11980 21428 12032 21437
rect 12164 21360 12216 21412
rect 12532 21360 12584 21412
rect 12900 21360 12952 21412
rect 13268 21428 13320 21480
rect 3976 21292 4028 21344
rect 4068 21292 4120 21344
rect 6460 21292 6512 21344
rect 6552 21335 6604 21344
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 7380 21292 7432 21344
rect 11612 21292 11664 21344
rect 14188 21360 14240 21412
rect 15936 21428 15988 21480
rect 13360 21335 13412 21344
rect 13360 21301 13369 21335
rect 13369 21301 13403 21335
rect 13403 21301 13412 21335
rect 13360 21292 13412 21301
rect 15844 21335 15896 21344
rect 15844 21301 15853 21335
rect 15853 21301 15887 21335
rect 15887 21301 15896 21335
rect 15844 21292 15896 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 2688 21088 2740 21140
rect 3056 21131 3108 21140
rect 3056 21097 3065 21131
rect 3065 21097 3099 21131
rect 3099 21097 3108 21131
rect 3056 21088 3108 21097
rect 3884 21088 3936 21140
rect 3976 21131 4028 21140
rect 3976 21097 3985 21131
rect 3985 21097 4019 21131
rect 4019 21097 4028 21131
rect 3976 21088 4028 21097
rect 3148 20995 3200 21004
rect 3148 20961 3157 20995
rect 3157 20961 3191 20995
rect 3191 20961 3200 20995
rect 3148 20952 3200 20961
rect 2780 20884 2832 20936
rect 2964 20884 3016 20936
rect 3332 20884 3384 20936
rect 3700 21020 3752 21072
rect 4068 21020 4120 21072
rect 5724 21088 5776 21140
rect 6920 21088 6972 21140
rect 6368 21020 6420 21072
rect 6552 21020 6604 21072
rect 10232 21131 10284 21140
rect 10232 21097 10241 21131
rect 10241 21097 10275 21131
rect 10275 21097 10284 21131
rect 10232 21088 10284 21097
rect 11152 21088 11204 21140
rect 11520 21088 11572 21140
rect 9864 21020 9916 21072
rect 3608 20927 3660 20936
rect 3608 20893 3617 20927
rect 3617 20893 3651 20927
rect 3651 20893 3660 20927
rect 3608 20884 3660 20893
rect 1492 20816 1544 20868
rect 1768 20816 1820 20868
rect 3792 20816 3844 20868
rect 4620 20884 4672 20936
rect 5816 20952 5868 21004
rect 12256 21088 12308 21140
rect 12900 21131 12952 21140
rect 12900 21097 12909 21131
rect 12909 21097 12943 21131
rect 12943 21097 12952 21131
rect 12900 21088 12952 21097
rect 13084 21088 13136 21140
rect 13452 21131 13504 21140
rect 13452 21097 13461 21131
rect 13461 21097 13495 21131
rect 13495 21097 13504 21131
rect 13452 21088 13504 21097
rect 14648 21088 14700 21140
rect 16120 21131 16172 21140
rect 16120 21097 16129 21131
rect 16129 21097 16163 21131
rect 16163 21097 16172 21131
rect 16120 21088 16172 21097
rect 12164 21020 12216 21072
rect 12808 21063 12860 21072
rect 12808 21029 12817 21063
rect 12817 21029 12851 21063
rect 12851 21029 12860 21063
rect 12808 21020 12860 21029
rect 13544 21020 13596 21072
rect 5908 20884 5960 20936
rect 4712 20816 4764 20868
rect 6828 20884 6880 20936
rect 5724 20791 5776 20800
rect 5724 20757 5733 20791
rect 5733 20757 5767 20791
rect 5767 20757 5776 20791
rect 5724 20748 5776 20757
rect 6184 20816 6236 20868
rect 7288 20927 7340 20936
rect 7288 20893 7297 20927
rect 7297 20893 7331 20927
rect 7331 20893 7340 20927
rect 7288 20884 7340 20893
rect 7472 20884 7524 20936
rect 7564 20927 7616 20936
rect 7564 20893 7573 20927
rect 7573 20893 7607 20927
rect 7607 20893 7616 20927
rect 7564 20884 7616 20893
rect 11796 20884 11848 20936
rect 12164 20884 12216 20936
rect 7840 20816 7892 20868
rect 8392 20859 8444 20868
rect 8392 20825 8401 20859
rect 8401 20825 8435 20859
rect 8435 20825 8444 20859
rect 8392 20816 8444 20825
rect 9772 20816 9824 20868
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 8576 20791 8628 20800
rect 8576 20757 8601 20791
rect 8601 20757 8628 20791
rect 8576 20748 8628 20757
rect 8760 20791 8812 20800
rect 8760 20757 8769 20791
rect 8769 20757 8803 20791
rect 8803 20757 8812 20791
rect 8760 20748 8812 20757
rect 12256 20791 12308 20800
rect 12256 20757 12265 20791
rect 12265 20757 12299 20791
rect 12299 20757 12308 20791
rect 12256 20748 12308 20757
rect 12440 20791 12492 20800
rect 12440 20757 12449 20791
rect 12449 20757 12483 20791
rect 12483 20757 12492 20791
rect 12440 20748 12492 20757
rect 14188 20927 14240 20936
rect 14188 20893 14198 20927
rect 14198 20893 14232 20927
rect 14232 20893 14240 20927
rect 14188 20884 14240 20893
rect 15844 20884 15896 20936
rect 15936 20927 15988 20936
rect 15936 20893 15945 20927
rect 15945 20893 15979 20927
rect 15979 20893 15988 20927
rect 15936 20884 15988 20893
rect 13820 20748 13872 20800
rect 15016 20748 15068 20800
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 1492 20587 1544 20596
rect 1492 20553 1501 20587
rect 1501 20553 1535 20587
rect 1535 20553 1544 20587
rect 1492 20544 1544 20553
rect 3148 20544 3200 20596
rect 6184 20587 6236 20596
rect 6184 20553 6193 20587
rect 6193 20553 6227 20587
rect 6227 20553 6236 20587
rect 6184 20544 6236 20553
rect 6368 20544 6420 20596
rect 6828 20544 6880 20596
rect 1768 20519 1820 20528
rect 1768 20485 1777 20519
rect 1777 20485 1811 20519
rect 1811 20485 1820 20519
rect 1768 20476 1820 20485
rect 1860 20519 1912 20528
rect 1860 20485 1869 20519
rect 1869 20485 1903 20519
rect 1903 20485 1912 20519
rect 1860 20476 1912 20485
rect 2320 20476 2372 20528
rect 2136 20451 2188 20460
rect 2136 20417 2145 20451
rect 2145 20417 2179 20451
rect 2179 20417 2188 20451
rect 2136 20408 2188 20417
rect 2688 20408 2740 20460
rect 2872 20476 2924 20528
rect 3516 20476 3568 20528
rect 5724 20476 5776 20528
rect 3056 20451 3108 20460
rect 3056 20417 3065 20451
rect 3065 20417 3099 20451
rect 3099 20417 3108 20451
rect 3056 20408 3108 20417
rect 3700 20451 3752 20460
rect 3700 20417 3709 20451
rect 3709 20417 3743 20451
rect 3743 20417 3752 20451
rect 3700 20408 3752 20417
rect 3792 20408 3844 20460
rect 1952 20340 2004 20392
rect 1308 20272 1360 20324
rect 3148 20340 3200 20392
rect 3608 20340 3660 20392
rect 6368 20451 6420 20460
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 7012 20408 7064 20460
rect 7472 20544 7524 20596
rect 9864 20587 9916 20596
rect 9864 20553 9889 20587
rect 9889 20553 9916 20587
rect 9864 20544 9916 20553
rect 11244 20544 11296 20596
rect 11888 20544 11940 20596
rect 13636 20544 13688 20596
rect 9680 20519 9732 20528
rect 9680 20485 9689 20519
rect 9689 20485 9723 20519
rect 9723 20485 9732 20519
rect 9680 20476 9732 20485
rect 11796 20476 11848 20528
rect 11980 20476 12032 20528
rect 7748 20408 7800 20460
rect 11520 20451 11572 20460
rect 11520 20417 11529 20451
rect 11529 20417 11563 20451
rect 11563 20417 11572 20451
rect 11520 20408 11572 20417
rect 12256 20408 12308 20460
rect 13452 20408 13504 20460
rect 7196 20383 7248 20392
rect 7196 20349 7205 20383
rect 7205 20349 7239 20383
rect 7239 20349 7248 20383
rect 7196 20340 7248 20349
rect 9220 20340 9272 20392
rect 9496 20340 9548 20392
rect 13176 20340 13228 20392
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 15384 20544 15436 20596
rect 3332 20272 3384 20324
rect 3608 20247 3660 20256
rect 3608 20213 3617 20247
rect 3617 20213 3651 20247
rect 3651 20213 3660 20247
rect 3608 20204 3660 20213
rect 3700 20204 3752 20256
rect 14464 20272 14516 20324
rect 15936 20340 15988 20392
rect 8392 20204 8444 20256
rect 8852 20247 8904 20256
rect 8852 20213 8861 20247
rect 8861 20213 8895 20247
rect 8895 20213 8904 20247
rect 8852 20204 8904 20213
rect 9772 20204 9824 20256
rect 10784 20247 10836 20256
rect 10784 20213 10793 20247
rect 10793 20213 10827 20247
rect 10827 20213 10836 20247
rect 10784 20204 10836 20213
rect 11520 20204 11572 20256
rect 11980 20204 12032 20256
rect 13176 20204 13228 20256
rect 13452 20204 13504 20256
rect 13820 20204 13872 20256
rect 15292 20204 15344 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 2780 20000 2832 20052
rect 2964 20000 3016 20052
rect 6368 20000 6420 20052
rect 7104 20000 7156 20052
rect 7748 20043 7800 20052
rect 7748 20009 7757 20043
rect 7757 20009 7791 20043
rect 7791 20009 7800 20043
rect 7748 20000 7800 20009
rect 8576 20000 8628 20052
rect 9496 20000 9548 20052
rect 15936 20043 15988 20052
rect 15936 20009 15945 20043
rect 15945 20009 15979 20043
rect 15979 20009 15988 20043
rect 15936 20000 15988 20009
rect 848 19796 900 19848
rect 2044 19796 2096 19848
rect 3240 19932 3292 19984
rect 3148 19907 3200 19916
rect 3148 19873 3157 19907
rect 3157 19873 3191 19907
rect 3191 19873 3200 19907
rect 3148 19864 3200 19873
rect 3792 19907 3844 19916
rect 3792 19873 3801 19907
rect 3801 19873 3835 19907
rect 3835 19873 3844 19907
rect 3792 19864 3844 19873
rect 12072 19932 12124 19984
rect 7380 19907 7432 19916
rect 2320 19839 2372 19848
rect 2320 19805 2329 19839
rect 2329 19805 2363 19839
rect 2363 19805 2372 19839
rect 2320 19796 2372 19805
rect 3700 19796 3752 19848
rect 3148 19728 3200 19780
rect 2136 19703 2188 19712
rect 2136 19669 2145 19703
rect 2145 19669 2179 19703
rect 2179 19669 2188 19703
rect 2136 19660 2188 19669
rect 2872 19703 2924 19712
rect 2872 19669 2881 19703
rect 2881 19669 2915 19703
rect 2915 19669 2924 19703
rect 2872 19660 2924 19669
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 6828 19796 6880 19848
rect 7380 19873 7389 19907
rect 7389 19873 7423 19907
rect 7423 19873 7432 19907
rect 7380 19864 7432 19873
rect 10784 19864 10836 19916
rect 7012 19839 7064 19848
rect 7012 19805 7021 19839
rect 7021 19805 7055 19839
rect 7055 19805 7064 19839
rect 7012 19796 7064 19805
rect 7472 19796 7524 19848
rect 7564 19839 7616 19848
rect 7564 19805 7573 19839
rect 7573 19805 7607 19839
rect 7607 19805 7616 19839
rect 7564 19796 7616 19805
rect 9864 19796 9916 19848
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 11796 19839 11848 19848
rect 11796 19805 11805 19839
rect 11805 19805 11839 19839
rect 11839 19805 11848 19839
rect 11796 19796 11848 19805
rect 11888 19796 11940 19848
rect 13912 19932 13964 19984
rect 13452 19864 13504 19916
rect 13820 19864 13872 19916
rect 9588 19728 9640 19780
rect 6736 19660 6788 19712
rect 11704 19660 11756 19712
rect 13360 19728 13412 19780
rect 14556 19839 14608 19848
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 14924 19728 14976 19780
rect 13452 19660 13504 19712
rect 15476 19660 15528 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 3148 19499 3200 19508
rect 3148 19465 3157 19499
rect 3157 19465 3191 19499
rect 3191 19465 3200 19499
rect 3148 19456 3200 19465
rect 3240 19499 3292 19508
rect 3240 19465 3249 19499
rect 3249 19465 3283 19499
rect 3283 19465 3292 19499
rect 3240 19456 3292 19465
rect 6644 19456 6696 19508
rect 9220 19499 9272 19508
rect 9220 19465 9229 19499
rect 9229 19465 9263 19499
rect 9263 19465 9272 19499
rect 9220 19456 9272 19465
rect 11428 19456 11480 19508
rect 7196 19388 7248 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 2872 19320 2924 19372
rect 3516 19295 3568 19304
rect 3516 19261 3525 19295
rect 3525 19261 3559 19295
rect 3559 19261 3568 19295
rect 3516 19252 3568 19261
rect 3700 19252 3752 19304
rect 7656 19320 7708 19372
rect 8208 19388 8260 19440
rect 9772 19388 9824 19440
rect 11612 19456 11664 19508
rect 11980 19499 12032 19508
rect 11980 19465 11989 19499
rect 11989 19465 12023 19499
rect 12023 19465 12032 19499
rect 11980 19456 12032 19465
rect 13360 19499 13412 19508
rect 13360 19465 13369 19499
rect 13369 19465 13403 19499
rect 13403 19465 13412 19499
rect 13360 19456 13412 19465
rect 13728 19456 13780 19508
rect 14924 19499 14976 19508
rect 14924 19465 14933 19499
rect 14933 19465 14967 19499
rect 14967 19465 14976 19499
rect 14924 19456 14976 19465
rect 15292 19499 15344 19508
rect 15292 19465 15301 19499
rect 15301 19465 15335 19499
rect 15335 19465 15344 19499
rect 15292 19456 15344 19465
rect 8116 19363 8168 19372
rect 8116 19329 8150 19363
rect 8150 19329 8168 19363
rect 8116 19320 8168 19329
rect 9680 19363 9732 19372
rect 9680 19329 9689 19363
rect 9689 19329 9723 19363
rect 9723 19329 9732 19363
rect 9680 19320 9732 19329
rect 11704 19320 11756 19372
rect 12256 19320 12308 19372
rect 13268 19320 13320 19372
rect 13544 19363 13596 19372
rect 13544 19329 13553 19363
rect 13553 19329 13587 19363
rect 13587 19329 13596 19363
rect 13544 19320 13596 19329
rect 13636 19320 13688 19372
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 12072 19252 12124 19261
rect 12532 19252 12584 19304
rect 13360 19252 13412 19304
rect 7840 19184 7892 19236
rect 2780 19159 2832 19168
rect 2780 19125 2789 19159
rect 2789 19125 2823 19159
rect 2823 19125 2832 19159
rect 2780 19116 2832 19125
rect 2872 19159 2924 19168
rect 2872 19125 2881 19159
rect 2881 19125 2915 19159
rect 2915 19125 2924 19159
rect 2872 19116 2924 19125
rect 5264 19116 5316 19168
rect 9588 19159 9640 19168
rect 9588 19125 9597 19159
rect 9597 19125 9631 19159
rect 9631 19125 9640 19159
rect 9588 19116 9640 19125
rect 9864 19184 9916 19236
rect 12992 19227 13044 19236
rect 12992 19193 13001 19227
rect 13001 19193 13035 19227
rect 13035 19193 13044 19227
rect 12992 19184 13044 19193
rect 13544 19227 13596 19236
rect 13544 19193 13553 19227
rect 13553 19193 13587 19227
rect 13587 19193 13596 19227
rect 13544 19184 13596 19193
rect 13728 19184 13780 19236
rect 14372 19363 14424 19372
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 14372 19320 14424 19329
rect 14096 19252 14148 19304
rect 15384 19295 15436 19304
rect 15384 19261 15393 19295
rect 15393 19261 15427 19295
rect 15427 19261 15436 19295
rect 15384 19252 15436 19261
rect 15476 19295 15528 19304
rect 15476 19261 15485 19295
rect 15485 19261 15519 19295
rect 15519 19261 15528 19295
rect 15476 19252 15528 19261
rect 13912 19184 13964 19236
rect 14740 19227 14792 19236
rect 14740 19193 14749 19227
rect 14749 19193 14783 19227
rect 14783 19193 14792 19227
rect 14740 19184 14792 19193
rect 14004 19116 14056 19168
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 2136 18912 2188 18964
rect 2320 18955 2372 18964
rect 2320 18921 2329 18955
rect 2329 18921 2363 18955
rect 2363 18921 2372 18955
rect 2320 18912 2372 18921
rect 6000 18912 6052 18964
rect 8116 18912 8168 18964
rect 12256 18912 12308 18964
rect 13360 18955 13412 18964
rect 13360 18921 13369 18955
rect 13369 18921 13403 18955
rect 13403 18921 13412 18955
rect 13360 18912 13412 18921
rect 13452 18912 13504 18964
rect 3792 18776 3844 18828
rect 8576 18844 8628 18896
rect 7472 18776 7524 18828
rect 8668 18819 8720 18828
rect 8668 18785 8677 18819
rect 8677 18785 8711 18819
rect 8711 18785 8720 18819
rect 8668 18776 8720 18785
rect 2780 18708 2832 18760
rect 8852 18708 8904 18760
rect 13268 18844 13320 18896
rect 14096 18912 14148 18964
rect 15384 18912 15436 18964
rect 14004 18844 14056 18896
rect 9588 18819 9640 18828
rect 9588 18785 9597 18819
rect 9597 18785 9631 18819
rect 9631 18785 9640 18819
rect 9588 18776 9640 18785
rect 10140 18776 10192 18828
rect 11520 18776 11572 18828
rect 14464 18819 14516 18828
rect 14464 18785 14473 18819
rect 14473 18785 14507 18819
rect 14507 18785 14516 18819
rect 14464 18776 14516 18785
rect 10784 18751 10836 18760
rect 10784 18717 10793 18751
rect 10793 18717 10827 18751
rect 10827 18717 10836 18751
rect 10784 18708 10836 18717
rect 12072 18708 12124 18760
rect 12348 18751 12400 18760
rect 12348 18717 12357 18751
rect 12357 18717 12391 18751
rect 12391 18717 12400 18751
rect 12348 18708 12400 18717
rect 12532 18751 12584 18760
rect 12532 18717 12541 18751
rect 12541 18717 12575 18751
rect 12575 18717 12584 18751
rect 12532 18708 12584 18717
rect 12992 18708 13044 18760
rect 13360 18751 13412 18760
rect 13360 18717 13369 18751
rect 13369 18717 13403 18751
rect 13403 18717 13412 18751
rect 13360 18708 13412 18717
rect 2964 18640 3016 18692
rect 3516 18640 3568 18692
rect 5540 18683 5592 18692
rect 5540 18649 5574 18683
rect 5574 18649 5592 18683
rect 5540 18640 5592 18649
rect 9496 18640 9548 18692
rect 12164 18640 12216 18692
rect 11888 18615 11940 18624
rect 11888 18581 11897 18615
rect 11897 18581 11931 18615
rect 11931 18581 11940 18615
rect 11888 18572 11940 18581
rect 12900 18640 12952 18692
rect 12440 18615 12492 18624
rect 12440 18581 12449 18615
rect 12449 18581 12483 18615
rect 12483 18581 12492 18615
rect 12440 18572 12492 18581
rect 13728 18572 13780 18624
rect 14648 18615 14700 18624
rect 14648 18581 14657 18615
rect 14657 18581 14691 18615
rect 14691 18581 14700 18615
rect 14648 18572 14700 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 3056 18368 3108 18420
rect 3700 18368 3752 18420
rect 5264 18368 5316 18420
rect 5540 18368 5592 18420
rect 7472 18411 7524 18420
rect 7472 18377 7497 18411
rect 7497 18377 7524 18411
rect 7472 18368 7524 18377
rect 2136 18300 2188 18352
rect 6000 18300 6052 18352
rect 7288 18343 7340 18352
rect 7288 18309 7297 18343
rect 7297 18309 7331 18343
rect 7331 18309 7340 18343
rect 7288 18300 7340 18309
rect 2228 18207 2280 18216
rect 2228 18173 2237 18207
rect 2237 18173 2271 18207
rect 2271 18173 2280 18207
rect 2228 18164 2280 18173
rect 2964 18232 3016 18284
rect 3792 18232 3844 18284
rect 3976 18275 4028 18284
rect 3976 18241 4010 18275
rect 4010 18241 4028 18275
rect 3976 18232 4028 18241
rect 6828 18275 6880 18284
rect 6828 18241 6837 18275
rect 6837 18241 6871 18275
rect 6871 18241 6880 18275
rect 6828 18232 6880 18241
rect 10784 18368 10836 18420
rect 14648 18368 14700 18420
rect 15016 18368 15068 18420
rect 11796 18343 11848 18352
rect 11796 18309 11805 18343
rect 11805 18309 11839 18343
rect 11839 18309 11848 18343
rect 11796 18300 11848 18309
rect 2688 18164 2740 18216
rect 3516 18164 3568 18216
rect 6092 18207 6144 18216
rect 6092 18173 6101 18207
rect 6101 18173 6135 18207
rect 6135 18173 6144 18207
rect 6092 18164 6144 18173
rect 9588 18164 9640 18216
rect 2964 18096 3016 18148
rect 3424 18096 3476 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 2780 18071 2832 18080
rect 2780 18037 2789 18071
rect 2789 18037 2823 18071
rect 2823 18037 2832 18071
rect 2780 18028 2832 18037
rect 7472 18071 7524 18080
rect 7472 18037 7481 18071
rect 7481 18037 7515 18071
rect 7515 18037 7524 18071
rect 7472 18028 7524 18037
rect 8116 18028 8168 18080
rect 9864 18028 9916 18080
rect 12072 18275 12124 18284
rect 12072 18241 12081 18275
rect 12081 18241 12115 18275
rect 12115 18241 12124 18275
rect 12072 18232 12124 18241
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 12256 18164 12308 18216
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 12992 18232 13044 18284
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 14004 18232 14056 18284
rect 14464 18232 14516 18284
rect 13084 18164 13136 18216
rect 13820 18164 13872 18216
rect 14280 18164 14332 18216
rect 14004 18096 14056 18148
rect 11888 18028 11940 18080
rect 12348 18028 12400 18080
rect 12808 18028 12860 18080
rect 14188 18028 14240 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 2964 17824 3016 17876
rect 3332 17867 3384 17876
rect 3332 17833 3341 17867
rect 3341 17833 3375 17867
rect 3375 17833 3384 17867
rect 3332 17824 3384 17833
rect 3608 17824 3660 17876
rect 3976 17824 4028 17876
rect 8300 17824 8352 17876
rect 1400 17731 1452 17740
rect 1400 17697 1409 17731
rect 1409 17697 1443 17731
rect 1443 17697 1452 17731
rect 1400 17688 1452 17697
rect 2780 17620 2832 17672
rect 1676 17595 1728 17604
rect 1676 17561 1710 17595
rect 1710 17561 1728 17595
rect 1676 17552 1728 17561
rect 2228 17552 2280 17604
rect 3056 17688 3108 17740
rect 6184 17688 6236 17740
rect 6828 17688 6880 17740
rect 3516 17620 3568 17672
rect 3976 17620 4028 17672
rect 3056 17552 3108 17604
rect 5264 17552 5316 17604
rect 7840 17552 7892 17604
rect 8116 17620 8168 17672
rect 12164 17688 12216 17740
rect 12992 17824 13044 17876
rect 14464 17731 14516 17740
rect 14464 17697 14473 17731
rect 14473 17697 14507 17731
rect 14507 17697 14516 17731
rect 14464 17688 14516 17697
rect 8944 17552 8996 17604
rect 11888 17595 11940 17604
rect 11888 17561 11897 17595
rect 11897 17561 11931 17595
rect 11931 17561 11940 17595
rect 11888 17552 11940 17561
rect 12532 17552 12584 17604
rect 12992 17620 13044 17672
rect 14188 17663 14240 17672
rect 14188 17629 14197 17663
rect 14197 17629 14231 17663
rect 14231 17629 14240 17663
rect 14188 17620 14240 17629
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 14280 17620 14332 17629
rect 14832 17620 14884 17672
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 2872 17484 2924 17536
rect 6736 17484 6788 17536
rect 8392 17527 8444 17536
rect 8392 17493 8401 17527
rect 8401 17493 8435 17527
rect 8435 17493 8444 17527
rect 8392 17484 8444 17493
rect 12440 17484 12492 17536
rect 14004 17484 14056 17536
rect 15844 17527 15896 17536
rect 15844 17493 15853 17527
rect 15853 17493 15887 17527
rect 15887 17493 15896 17527
rect 15844 17484 15896 17493
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 2136 17280 2188 17332
rect 3332 17280 3384 17332
rect 3700 17280 3752 17332
rect 2228 17187 2280 17196
rect 2228 17153 2237 17187
rect 2237 17153 2271 17187
rect 2271 17153 2280 17187
rect 2228 17144 2280 17153
rect 2780 17212 2832 17264
rect 6184 17323 6236 17332
rect 6184 17289 6193 17323
rect 6193 17289 6227 17323
rect 6227 17289 6236 17323
rect 6184 17280 6236 17289
rect 2872 17144 2924 17196
rect 3884 17212 3936 17264
rect 6736 17323 6788 17332
rect 6736 17289 6745 17323
rect 6745 17289 6779 17323
rect 6779 17289 6788 17323
rect 6736 17280 6788 17289
rect 7012 17280 7064 17332
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 8852 17280 8904 17332
rect 8944 17323 8996 17332
rect 8944 17289 8953 17323
rect 8953 17289 8987 17323
rect 8987 17289 8996 17323
rect 8944 17280 8996 17289
rect 12164 17280 12216 17332
rect 12900 17323 12952 17332
rect 12900 17289 12909 17323
rect 12909 17289 12943 17323
rect 12943 17289 12952 17323
rect 12900 17280 12952 17289
rect 13360 17280 13412 17332
rect 15936 17280 15988 17332
rect 16396 17280 16448 17332
rect 7288 17144 7340 17196
rect 9772 17212 9824 17264
rect 12348 17212 12400 17264
rect 3792 17076 3844 17128
rect 5816 17076 5868 17128
rect 8024 17187 8076 17196
rect 8024 17153 8033 17187
rect 8033 17153 8067 17187
rect 8067 17153 8076 17187
rect 8024 17144 8076 17153
rect 8392 17144 8444 17196
rect 8852 17187 8904 17196
rect 8852 17153 8861 17187
rect 8861 17153 8895 17187
rect 8895 17153 8904 17187
rect 8852 17144 8904 17153
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 11796 17187 11848 17196
rect 11796 17153 11805 17187
rect 11805 17153 11839 17187
rect 11839 17153 11848 17187
rect 11796 17144 11848 17153
rect 3332 17008 3384 17060
rect 3056 16940 3108 16992
rect 3700 16983 3752 16992
rect 3700 16949 3709 16983
rect 3709 16949 3743 16983
rect 3743 16949 3752 16983
rect 3700 16940 3752 16949
rect 8300 17008 8352 17060
rect 9864 17119 9916 17128
rect 9864 17085 9873 17119
rect 9873 17085 9907 17119
rect 9907 17085 9916 17119
rect 9864 17076 9916 17085
rect 11612 17076 11664 17128
rect 12164 17187 12216 17196
rect 12164 17153 12173 17187
rect 12173 17153 12207 17187
rect 12207 17153 12216 17187
rect 12164 17144 12216 17153
rect 12532 17144 12584 17196
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 14188 17255 14240 17264
rect 14188 17221 14197 17255
rect 14197 17221 14231 17255
rect 14231 17221 14240 17255
rect 14188 17212 14240 17221
rect 14464 17212 14516 17264
rect 14280 17187 14332 17196
rect 14280 17153 14289 17187
rect 14289 17153 14323 17187
rect 14323 17153 14332 17187
rect 14280 17144 14332 17153
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 14556 17144 14608 17196
rect 15016 17187 15068 17196
rect 15016 17153 15050 17187
rect 15050 17153 15068 17187
rect 15016 17144 15068 17153
rect 16212 17187 16264 17196
rect 16212 17153 16221 17187
rect 16221 17153 16255 17187
rect 16255 17153 16264 17187
rect 16212 17144 16264 17153
rect 9128 17051 9180 17060
rect 9128 17017 9137 17051
rect 9137 17017 9171 17051
rect 9171 17017 9180 17051
rect 9128 17008 9180 17017
rect 13268 17119 13320 17128
rect 13268 17085 13277 17119
rect 13277 17085 13311 17119
rect 13311 17085 13320 17119
rect 13268 17076 13320 17085
rect 13452 17076 13504 17128
rect 16396 17051 16448 17060
rect 16396 17017 16405 17051
rect 16405 17017 16439 17051
rect 16439 17017 16448 17051
rect 16396 17008 16448 17017
rect 4620 16940 4672 16992
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 11428 16940 11480 16992
rect 12164 16940 12216 16992
rect 13268 16940 13320 16992
rect 13544 16940 13596 16992
rect 15384 16940 15436 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 2872 16779 2924 16788
rect 2872 16745 2881 16779
rect 2881 16745 2915 16779
rect 2915 16745 2924 16779
rect 2872 16736 2924 16745
rect 3884 16736 3936 16788
rect 7472 16736 7524 16788
rect 8484 16736 8536 16788
rect 12072 16736 12124 16788
rect 12348 16736 12400 16788
rect 3148 16668 3200 16720
rect 7288 16668 7340 16720
rect 8116 16711 8168 16720
rect 8116 16677 8125 16711
rect 8125 16677 8159 16711
rect 8159 16677 8168 16711
rect 8116 16668 8168 16677
rect 8300 16668 8352 16720
rect 8668 16668 8720 16720
rect 13544 16736 13596 16788
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 3516 16600 3568 16652
rect 3792 16600 3844 16652
rect 9588 16643 9640 16652
rect 9588 16609 9597 16643
rect 9597 16609 9631 16643
rect 9631 16609 9640 16643
rect 9588 16600 9640 16609
rect 9864 16643 9916 16652
rect 9864 16609 9873 16643
rect 9873 16609 9907 16643
rect 9907 16609 9916 16643
rect 9864 16600 9916 16609
rect 2872 16464 2924 16516
rect 4068 16464 4120 16516
rect 11520 16575 11572 16584
rect 11520 16541 11529 16575
rect 11529 16541 11563 16575
rect 11563 16541 11572 16575
rect 11520 16532 11572 16541
rect 11704 16532 11756 16584
rect 7564 16507 7616 16516
rect 7564 16473 7573 16507
rect 7573 16473 7607 16507
rect 7607 16473 7616 16507
rect 7564 16464 7616 16473
rect 8484 16507 8536 16516
rect 8484 16473 8493 16507
rect 8493 16473 8527 16507
rect 8527 16473 8536 16507
rect 8484 16464 8536 16473
rect 9036 16464 9088 16516
rect 2504 16396 2556 16448
rect 2964 16396 3016 16448
rect 5356 16439 5408 16448
rect 5356 16405 5365 16439
rect 5365 16405 5399 16439
rect 5399 16405 5408 16439
rect 5356 16396 5408 16405
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 7748 16439 7800 16448
rect 7748 16405 7757 16439
rect 7757 16405 7791 16439
rect 7791 16405 7800 16439
rect 7748 16396 7800 16405
rect 8300 16396 8352 16448
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 9956 16396 10008 16448
rect 11612 16396 11664 16448
rect 11980 16532 12032 16584
rect 12164 16575 12216 16584
rect 12164 16541 12173 16575
rect 12173 16541 12207 16575
rect 12207 16541 12216 16575
rect 12164 16532 12216 16541
rect 13084 16600 13136 16652
rect 14004 16668 14056 16720
rect 13820 16600 13872 16652
rect 12532 16532 12584 16584
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 13360 16532 13412 16584
rect 15016 16736 15068 16788
rect 16212 16736 16264 16788
rect 13728 16507 13780 16516
rect 13728 16473 13737 16507
rect 13737 16473 13771 16507
rect 13771 16473 13780 16507
rect 13728 16464 13780 16473
rect 13912 16464 13964 16516
rect 12532 16439 12584 16448
rect 12532 16405 12541 16439
rect 12541 16405 12575 16439
rect 12575 16405 12584 16439
rect 12532 16396 12584 16405
rect 13636 16396 13688 16448
rect 14740 16532 14792 16584
rect 15844 16532 15896 16584
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 15384 16464 15436 16516
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 4068 16235 4120 16244
rect 4068 16201 4077 16235
rect 4077 16201 4111 16235
rect 4111 16201 4120 16235
rect 4068 16192 4120 16201
rect 7564 16192 7616 16244
rect 8024 16192 8076 16244
rect 9772 16192 9824 16244
rect 3976 16124 4028 16176
rect 4712 16056 4764 16108
rect 5356 16056 5408 16108
rect 6920 16124 6972 16176
rect 8208 16124 8260 16176
rect 8300 16167 8352 16176
rect 8300 16133 8309 16167
rect 8309 16133 8343 16167
rect 8343 16133 8352 16167
rect 8300 16124 8352 16133
rect 8944 16124 8996 16176
rect 6644 16099 6696 16108
rect 6644 16065 6678 16099
rect 6678 16065 6696 16099
rect 6644 16056 6696 16065
rect 7840 16056 7892 16108
rect 9956 16235 10008 16244
rect 9956 16201 9965 16235
rect 9965 16201 9999 16235
rect 9999 16201 10008 16235
rect 9956 16192 10008 16201
rect 11796 16192 11848 16244
rect 12256 16192 12308 16244
rect 12532 16192 12584 16244
rect 12716 16192 12768 16244
rect 13268 16192 13320 16244
rect 12992 16124 13044 16176
rect 13820 16167 13872 16176
rect 13820 16133 13829 16167
rect 13829 16133 13863 16167
rect 13863 16133 13872 16167
rect 13820 16124 13872 16133
rect 11704 16099 11756 16108
rect 11704 16065 11713 16099
rect 11713 16065 11747 16099
rect 11747 16065 11756 16099
rect 11704 16056 11756 16065
rect 4620 16031 4672 16040
rect 4620 15997 4629 16031
rect 4629 15997 4663 16031
rect 4663 15997 4672 16031
rect 4620 15988 4672 15997
rect 7748 15988 7800 16040
rect 8208 15988 8260 16040
rect 5356 15852 5408 15904
rect 8300 15895 8352 15904
rect 8300 15861 8309 15895
rect 8309 15861 8343 15895
rect 8343 15861 8352 15895
rect 8300 15852 8352 15861
rect 14280 16056 14332 16108
rect 16120 16056 16172 16108
rect 12900 15988 12952 16040
rect 12440 15963 12492 15972
rect 12440 15929 12449 15963
rect 12449 15929 12483 15963
rect 12483 15929 12492 15963
rect 12440 15920 12492 15929
rect 12072 15895 12124 15904
rect 12072 15861 12081 15895
rect 12081 15861 12115 15895
rect 12115 15861 12124 15895
rect 12072 15852 12124 15861
rect 13360 15920 13412 15972
rect 12992 15852 13044 15904
rect 13636 15895 13688 15904
rect 13636 15861 13645 15895
rect 13645 15861 13679 15895
rect 13679 15861 13688 15895
rect 13636 15852 13688 15861
rect 15752 15895 15804 15904
rect 15752 15861 15761 15895
rect 15761 15861 15795 15895
rect 15795 15861 15804 15895
rect 15752 15852 15804 15861
rect 15844 15895 15896 15904
rect 15844 15861 15853 15895
rect 15853 15861 15887 15895
rect 15887 15861 15896 15895
rect 15844 15852 15896 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 2964 15648 3016 15700
rect 3332 15648 3384 15700
rect 6644 15648 6696 15700
rect 8300 15648 8352 15700
rect 9036 15648 9088 15700
rect 9312 15648 9364 15700
rect 12072 15648 12124 15700
rect 15660 15648 15712 15700
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 16396 15691 16448 15700
rect 16396 15657 16405 15691
rect 16405 15657 16439 15691
rect 16439 15657 16448 15691
rect 16396 15648 16448 15657
rect 2872 15580 2924 15632
rect 2504 15487 2556 15496
rect 2504 15453 2513 15487
rect 2513 15453 2547 15487
rect 2547 15453 2556 15487
rect 2504 15444 2556 15453
rect 3148 15512 3200 15564
rect 2964 15444 3016 15496
rect 5540 15580 5592 15632
rect 6092 15512 6144 15564
rect 2688 15419 2740 15428
rect 2688 15385 2697 15419
rect 2697 15385 2731 15419
rect 2731 15385 2740 15419
rect 2688 15376 2740 15385
rect 2136 15308 2188 15360
rect 2596 15308 2648 15360
rect 3148 15376 3200 15428
rect 3976 15444 4028 15496
rect 6460 15555 6512 15564
rect 6460 15521 6469 15555
rect 6469 15521 6503 15555
rect 6503 15521 6512 15555
rect 6460 15512 6512 15521
rect 7656 15512 7708 15564
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 10140 15512 10192 15564
rect 13176 15580 13228 15632
rect 13820 15580 13872 15632
rect 6828 15444 6880 15496
rect 10048 15444 10100 15496
rect 12624 15444 12676 15496
rect 13176 15487 13228 15496
rect 13176 15453 13185 15487
rect 13185 15453 13219 15487
rect 13219 15453 13228 15487
rect 13176 15444 13228 15453
rect 8852 15376 8904 15428
rect 11704 15376 11756 15428
rect 12256 15419 12308 15428
rect 12256 15385 12281 15419
rect 12281 15385 12308 15419
rect 12256 15376 12308 15385
rect 4252 15308 4304 15360
rect 5540 15308 5592 15360
rect 7012 15308 7064 15360
rect 7380 15351 7432 15360
rect 7380 15317 7389 15351
rect 7389 15317 7423 15351
rect 7423 15317 7432 15351
rect 7380 15308 7432 15317
rect 8760 15351 8812 15360
rect 8760 15317 8769 15351
rect 8769 15317 8803 15351
rect 8803 15317 8812 15351
rect 8760 15308 8812 15317
rect 9496 15308 9548 15360
rect 10324 15308 10376 15360
rect 12440 15351 12492 15360
rect 12440 15317 12449 15351
rect 12449 15317 12483 15351
rect 12483 15317 12492 15351
rect 13544 15487 13596 15496
rect 13544 15453 13553 15487
rect 13553 15453 13587 15487
rect 13587 15453 13596 15487
rect 13544 15444 13596 15453
rect 13636 15444 13688 15496
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 14188 15444 14240 15496
rect 14556 15512 14608 15564
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 15752 15444 15804 15496
rect 14740 15376 14792 15428
rect 15108 15376 15160 15428
rect 12440 15308 12492 15317
rect 14280 15308 14332 15360
rect 15568 15308 15620 15360
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 2964 15147 3016 15156
rect 2964 15113 2973 15147
rect 2973 15113 3007 15147
rect 3007 15113 3016 15147
rect 2964 15104 3016 15113
rect 5540 15147 5592 15156
rect 5540 15113 5549 15147
rect 5549 15113 5583 15147
rect 5583 15113 5592 15147
rect 5540 15104 5592 15113
rect 7656 15104 7708 15156
rect 8116 15104 8168 15156
rect 10048 15104 10100 15156
rect 2780 15036 2832 15088
rect 1860 15011 1912 15020
rect 1860 14977 1894 15011
rect 1894 14977 1912 15011
rect 1860 14968 1912 14977
rect 3148 14968 3200 15020
rect 4252 14968 4304 15020
rect 6920 15036 6972 15088
rect 8852 15036 8904 15088
rect 9588 15036 9640 15088
rect 6644 15011 6696 15020
rect 6644 14977 6678 15011
rect 6678 14977 6696 15011
rect 6644 14968 6696 14977
rect 9036 15011 9088 15020
rect 9036 14977 9054 15011
rect 9054 14977 9088 15011
rect 9036 14968 9088 14977
rect 11244 14968 11296 15020
rect 12532 15104 12584 15156
rect 13084 15147 13136 15156
rect 13084 15113 13093 15147
rect 13093 15113 13127 15147
rect 13127 15113 13136 15147
rect 13084 15104 13136 15113
rect 11888 14968 11940 15020
rect 12440 15036 12492 15088
rect 13176 15036 13228 15088
rect 14096 15104 14148 15156
rect 15108 15147 15160 15156
rect 15108 15113 15117 15147
rect 15117 15113 15151 15147
rect 15151 15113 15160 15147
rect 15108 15104 15160 15113
rect 15844 15104 15896 15156
rect 15568 15079 15620 15088
rect 15568 15045 15577 15079
rect 15577 15045 15611 15079
rect 15611 15045 15620 15079
rect 15568 15036 15620 15045
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 12808 14968 12860 15020
rect 3424 14832 3476 14884
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 8944 14764 8996 14816
rect 12532 14943 12584 14952
rect 12532 14909 12541 14943
rect 12541 14909 12575 14943
rect 12575 14909 12584 14943
rect 12532 14900 12584 14909
rect 12716 14900 12768 14952
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 14096 14968 14148 15020
rect 16120 14968 16172 15020
rect 14372 14900 14424 14952
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 11888 14875 11940 14884
rect 11888 14841 11897 14875
rect 11897 14841 11931 14875
rect 11931 14841 11940 14875
rect 11888 14832 11940 14841
rect 13268 14832 13320 14884
rect 13544 14832 13596 14884
rect 16212 14764 16264 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 1860 14560 1912 14612
rect 2964 14560 3016 14612
rect 3148 14603 3200 14612
rect 3148 14569 3157 14603
rect 3157 14569 3191 14603
rect 3191 14569 3200 14603
rect 3148 14560 3200 14569
rect 6644 14560 6696 14612
rect 6828 14492 6880 14544
rect 8852 14560 8904 14612
rect 9036 14560 9088 14612
rect 2044 14424 2096 14476
rect 2688 14424 2740 14476
rect 7380 14467 7432 14476
rect 7380 14433 7389 14467
rect 7389 14433 7423 14467
rect 7423 14433 7432 14467
rect 7380 14424 7432 14433
rect 2136 14399 2188 14408
rect 2136 14365 2145 14399
rect 2145 14365 2179 14399
rect 2179 14365 2188 14399
rect 2136 14356 2188 14365
rect 2964 14356 3016 14408
rect 3516 14356 3568 14408
rect 6920 14356 6972 14408
rect 7932 14356 7984 14408
rect 8760 14424 8812 14476
rect 9588 14467 9640 14476
rect 9588 14433 9597 14467
rect 9597 14433 9631 14467
rect 9631 14433 9640 14467
rect 9588 14424 9640 14433
rect 12992 14560 13044 14612
rect 13728 14560 13780 14612
rect 16120 14603 16172 14612
rect 16120 14569 16129 14603
rect 16129 14569 16163 14603
rect 16163 14569 16172 14603
rect 16120 14560 16172 14569
rect 11888 14492 11940 14544
rect 8944 14356 8996 14408
rect 9864 14356 9916 14408
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 11612 14356 11664 14408
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 12532 14467 12584 14476
rect 12532 14433 12541 14467
rect 12541 14433 12575 14467
rect 12575 14433 12584 14467
rect 12532 14424 12584 14433
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 13084 14424 13136 14476
rect 13820 14424 13872 14476
rect 14188 14424 14240 14476
rect 14556 14424 14608 14476
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 13360 14399 13412 14408
rect 13360 14365 13369 14399
rect 13369 14365 13403 14399
rect 13403 14365 13412 14399
rect 13360 14356 13412 14365
rect 13452 14356 13504 14408
rect 16028 14356 16080 14408
rect 16212 14399 16264 14408
rect 16212 14365 16221 14399
rect 16221 14365 16255 14399
rect 16255 14365 16264 14399
rect 16212 14356 16264 14365
rect 2596 14288 2648 14340
rect 4068 14288 4120 14340
rect 2872 14263 2924 14272
rect 2872 14229 2881 14263
rect 2881 14229 2915 14263
rect 2915 14229 2924 14263
rect 2872 14220 2924 14229
rect 3608 14263 3660 14272
rect 3608 14229 3617 14263
rect 3617 14229 3651 14263
rect 3651 14229 3660 14263
rect 3608 14220 3660 14229
rect 6000 14288 6052 14340
rect 8116 14263 8168 14272
rect 8116 14229 8125 14263
rect 8125 14229 8159 14263
rect 8159 14229 8168 14263
rect 8116 14220 8168 14229
rect 9312 14263 9364 14272
rect 9312 14229 9321 14263
rect 9321 14229 9355 14263
rect 9355 14229 9364 14263
rect 9312 14220 9364 14229
rect 12532 14288 12584 14340
rect 13084 14288 13136 14340
rect 14648 14288 14700 14340
rect 15016 14331 15068 14340
rect 15016 14297 15050 14331
rect 15050 14297 15068 14331
rect 15016 14288 15068 14297
rect 13176 14220 13228 14272
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 13544 14220 13596 14272
rect 14832 14220 14884 14272
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 2964 14016 3016 14068
rect 3976 14016 4028 14068
rect 4068 14059 4120 14068
rect 4068 14025 4077 14059
rect 4077 14025 4111 14059
rect 4111 14025 4120 14059
rect 4068 14016 4120 14025
rect 2780 13948 2832 14000
rect 3792 13948 3844 14000
rect 6368 13948 6420 14000
rect 10232 14016 10284 14068
rect 11888 14016 11940 14068
rect 12440 14016 12492 14068
rect 12532 14059 12584 14068
rect 12532 14025 12541 14059
rect 12541 14025 12575 14059
rect 12575 14025 12584 14059
rect 12532 14016 12584 14025
rect 12624 14016 12676 14068
rect 13176 14016 13228 14068
rect 6644 13948 6696 14000
rect 6920 13948 6972 14000
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 2044 13855 2096 13864
rect 2044 13821 2053 13855
rect 2053 13821 2087 13855
rect 2087 13821 2096 13855
rect 2044 13812 2096 13821
rect 2964 13880 3016 13932
rect 9128 13948 9180 14000
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 6000 13812 6052 13864
rect 9128 13812 9180 13864
rect 2596 13744 2648 13796
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 11704 13948 11756 14000
rect 11244 13880 11296 13932
rect 12164 13923 12216 13932
rect 12164 13889 12173 13923
rect 12173 13889 12207 13923
rect 12207 13889 12216 13923
rect 12164 13880 12216 13889
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2228 13676 2280 13728
rect 9680 13744 9732 13796
rect 12532 13744 12584 13796
rect 13176 13923 13228 13932
rect 13176 13889 13185 13923
rect 13185 13889 13219 13923
rect 13219 13889 13228 13923
rect 13176 13880 13228 13889
rect 13636 13948 13688 14000
rect 13820 14016 13872 14068
rect 14464 14016 14516 14068
rect 15016 14059 15068 14068
rect 15016 14025 15025 14059
rect 15025 14025 15059 14059
rect 15059 14025 15068 14059
rect 15016 14016 15068 14025
rect 13268 13812 13320 13864
rect 13912 13880 13964 13932
rect 14004 13923 14056 13932
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 13636 13812 13688 13864
rect 14280 13880 14332 13932
rect 16120 13880 16172 13932
rect 14372 13812 14424 13864
rect 11796 13676 11848 13728
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 13544 13676 13596 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 2320 13472 2372 13524
rect 2596 13472 2648 13524
rect 13176 13515 13228 13524
rect 13176 13481 13185 13515
rect 13185 13481 13219 13515
rect 13219 13481 13228 13515
rect 13176 13472 13228 13481
rect 13544 13515 13596 13524
rect 13544 13481 13553 13515
rect 13553 13481 13587 13515
rect 13587 13481 13596 13515
rect 13544 13472 13596 13481
rect 14004 13472 14056 13524
rect 2688 13404 2740 13456
rect 3424 13404 3476 13456
rect 12900 13404 12952 13456
rect 13268 13404 13320 13456
rect 13820 13404 13872 13456
rect 14280 13404 14332 13456
rect 3792 13379 3844 13388
rect 3792 13345 3801 13379
rect 3801 13345 3835 13379
rect 3835 13345 3844 13379
rect 3792 13336 3844 13345
rect 2780 13268 2832 13320
rect 1492 13200 1544 13252
rect 4252 13200 4304 13252
rect 8852 13336 8904 13388
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 11244 13336 11296 13388
rect 12072 13336 12124 13388
rect 6644 13268 6696 13320
rect 8208 13268 8260 13320
rect 10232 13268 10284 13320
rect 11520 13268 11572 13320
rect 5264 13132 5316 13184
rect 5724 13175 5776 13184
rect 5724 13141 5733 13175
rect 5733 13141 5767 13175
rect 5767 13141 5776 13175
rect 5724 13132 5776 13141
rect 6092 13175 6144 13184
rect 6092 13141 6101 13175
rect 6101 13141 6135 13175
rect 6135 13141 6144 13175
rect 6092 13132 6144 13141
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 9864 13200 9916 13252
rect 12532 13311 12584 13320
rect 12532 13277 12541 13311
rect 12541 13277 12575 13311
rect 12575 13277 12584 13311
rect 12532 13268 12584 13277
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 11796 13200 11848 13252
rect 8392 13175 8444 13184
rect 8392 13141 8401 13175
rect 8401 13141 8435 13175
rect 8435 13141 8444 13175
rect 8392 13132 8444 13141
rect 11888 13132 11940 13184
rect 12716 13200 12768 13252
rect 13084 13311 13136 13320
rect 13084 13277 13093 13311
rect 13093 13277 13127 13311
rect 13127 13277 13136 13311
rect 13084 13268 13136 13277
rect 13452 13379 13504 13388
rect 13452 13345 13461 13379
rect 13461 13345 13495 13379
rect 13495 13345 13504 13379
rect 13452 13336 13504 13345
rect 14464 13336 14516 13388
rect 13176 13200 13228 13252
rect 14280 13311 14332 13320
rect 14280 13277 14289 13311
rect 14289 13277 14323 13311
rect 14323 13277 14332 13311
rect 14280 13268 14332 13277
rect 15936 13268 15988 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 14188 13200 14240 13252
rect 14372 13200 14424 13252
rect 15016 13200 15068 13252
rect 15384 13132 15436 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 15844 13175 15896 13184
rect 15844 13141 15853 13175
rect 15853 13141 15887 13175
rect 15887 13141 15896 13175
rect 15844 13132 15896 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 1308 12928 1360 12980
rect 2780 12860 2832 12912
rect 2228 12835 2280 12844
rect 2228 12801 2262 12835
rect 2262 12801 2280 12835
rect 2228 12792 2280 12801
rect 3976 12928 4028 12980
rect 4252 12971 4304 12980
rect 4252 12937 4261 12971
rect 4261 12937 4295 12971
rect 4295 12937 4304 12971
rect 4252 12928 4304 12937
rect 6092 12928 6144 12980
rect 7104 12928 7156 12980
rect 8116 12928 8168 12980
rect 9312 12928 9364 12980
rect 9864 12971 9916 12980
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 3424 12860 3476 12912
rect 3608 12767 3660 12776
rect 3608 12733 3617 12767
rect 3617 12733 3651 12767
rect 3651 12733 3660 12767
rect 3608 12724 3660 12733
rect 4068 12724 4120 12776
rect 7104 12835 7156 12844
rect 7104 12801 7113 12835
rect 7113 12801 7147 12835
rect 7147 12801 7156 12835
rect 7104 12792 7156 12801
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7380 12792 7432 12844
rect 4712 12724 4764 12776
rect 8300 12792 8352 12844
rect 10232 12792 10284 12844
rect 11888 12971 11940 12980
rect 11888 12937 11897 12971
rect 11897 12937 11931 12971
rect 11931 12937 11940 12971
rect 11888 12928 11940 12937
rect 12164 12792 12216 12844
rect 12624 12792 12676 12844
rect 12900 12792 12952 12844
rect 13176 12835 13228 12844
rect 13176 12801 13185 12835
rect 13185 12801 13219 12835
rect 13219 12801 13228 12835
rect 13176 12792 13228 12801
rect 8116 12767 8168 12776
rect 8116 12733 8125 12767
rect 8125 12733 8159 12767
rect 8159 12733 8168 12767
rect 8116 12724 8168 12733
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 9036 12656 9088 12708
rect 2320 12588 2372 12640
rect 2688 12588 2740 12640
rect 7932 12588 7984 12640
rect 11336 12724 11388 12776
rect 12348 12724 12400 12776
rect 15752 12928 15804 12980
rect 16120 12928 16172 12980
rect 16396 12928 16448 12980
rect 13912 12860 13964 12912
rect 14372 12903 14424 12912
rect 14372 12869 14381 12903
rect 14381 12869 14415 12903
rect 14415 12869 14424 12903
rect 14372 12860 14424 12869
rect 15200 12860 15252 12912
rect 13728 12835 13780 12844
rect 13728 12801 13737 12835
rect 13737 12801 13771 12835
rect 13771 12801 13780 12835
rect 13728 12792 13780 12801
rect 13820 12835 13872 12844
rect 13820 12801 13829 12835
rect 13829 12801 13863 12835
rect 13863 12801 13872 12835
rect 13820 12792 13872 12801
rect 14188 12835 14240 12844
rect 14188 12801 14197 12835
rect 14197 12801 14231 12835
rect 14231 12801 14240 12835
rect 14188 12792 14240 12801
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 14740 12792 14792 12844
rect 14924 12792 14976 12844
rect 16488 12835 16540 12844
rect 16488 12801 16497 12835
rect 16497 12801 16531 12835
rect 16531 12801 16540 12835
rect 16488 12792 16540 12801
rect 12808 12656 12860 12708
rect 13728 12656 13780 12708
rect 13912 12656 13964 12708
rect 14556 12656 14608 12708
rect 16028 12656 16080 12708
rect 10140 12588 10192 12640
rect 10508 12588 10560 12640
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 15568 12588 15620 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 4068 12384 4120 12436
rect 5264 12384 5316 12436
rect 6552 12384 6604 12436
rect 7104 12384 7156 12436
rect 8300 12384 8352 12436
rect 8484 12384 8536 12436
rect 10324 12427 10376 12436
rect 10324 12393 10333 12427
rect 10333 12393 10367 12427
rect 10367 12393 10376 12427
rect 10324 12384 10376 12393
rect 14188 12384 14240 12436
rect 15200 12427 15252 12436
rect 15200 12393 15209 12427
rect 15209 12393 15243 12427
rect 15243 12393 15252 12427
rect 15200 12384 15252 12393
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 5356 12316 5408 12368
rect 3884 12248 3936 12300
rect 2964 12180 3016 12232
rect 8208 12248 8260 12300
rect 8944 12291 8996 12300
rect 8944 12257 8953 12291
rect 8953 12257 8987 12291
rect 8987 12257 8996 12291
rect 8944 12248 8996 12257
rect 16396 12359 16448 12368
rect 16396 12325 16405 12359
rect 16405 12325 16439 12359
rect 16439 12325 16448 12359
rect 16396 12316 16448 12325
rect 11980 12248 12032 12300
rect 3884 12112 3936 12164
rect 848 12044 900 12096
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 3056 12044 3108 12096
rect 3608 12044 3660 12096
rect 4068 12044 4120 12096
rect 4436 12223 4488 12232
rect 4436 12189 4445 12223
rect 4445 12189 4479 12223
rect 4479 12189 4488 12223
rect 4436 12180 4488 12189
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 6644 12180 6696 12232
rect 8116 12180 8168 12232
rect 8760 12180 8812 12232
rect 10048 12180 10100 12232
rect 11612 12180 11664 12232
rect 12072 12223 12124 12232
rect 12072 12189 12081 12223
rect 12081 12189 12115 12223
rect 12115 12189 12124 12223
rect 12072 12180 12124 12189
rect 12532 12248 12584 12300
rect 13176 12248 13228 12300
rect 13820 12248 13872 12300
rect 14740 12248 14792 12300
rect 15568 12248 15620 12300
rect 15752 12291 15804 12300
rect 15752 12257 15761 12291
rect 15761 12257 15795 12291
rect 15795 12257 15804 12291
rect 15752 12248 15804 12257
rect 12992 12180 13044 12232
rect 14004 12180 14056 12232
rect 14372 12180 14424 12232
rect 16028 12180 16080 12232
rect 16304 12180 16356 12232
rect 4344 12044 4396 12096
rect 5724 12112 5776 12164
rect 9496 12112 9548 12164
rect 11520 12112 11572 12164
rect 11980 12112 12032 12164
rect 15844 12112 15896 12164
rect 4804 12044 4856 12096
rect 7380 12087 7432 12096
rect 7380 12053 7389 12087
rect 7389 12053 7423 12087
rect 7423 12053 7432 12087
rect 7380 12044 7432 12053
rect 7840 12087 7892 12096
rect 7840 12053 7849 12087
rect 7849 12053 7883 12087
rect 7883 12053 7892 12087
rect 7840 12044 7892 12053
rect 8300 12044 8352 12096
rect 8944 12044 8996 12096
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 11796 12087 11848 12096
rect 11796 12053 11805 12087
rect 11805 12053 11839 12087
rect 11839 12053 11848 12087
rect 11796 12044 11848 12053
rect 11888 12087 11940 12096
rect 11888 12053 11897 12087
rect 11897 12053 11931 12087
rect 11931 12053 11940 12087
rect 11888 12044 11940 12053
rect 15476 12044 15528 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 3792 11840 3844 11892
rect 4344 11840 4396 11892
rect 4712 11840 4764 11892
rect 8668 11840 8720 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 10048 11840 10100 11892
rect 2872 11772 2924 11824
rect 2780 11704 2832 11756
rect 3608 11747 3660 11756
rect 3608 11713 3642 11747
rect 3642 11713 3660 11747
rect 3608 11704 3660 11713
rect 4896 11772 4948 11824
rect 5540 11772 5592 11824
rect 7380 11772 7432 11824
rect 10416 11772 10468 11824
rect 11796 11840 11848 11892
rect 11888 11815 11940 11824
rect 11888 11781 11897 11815
rect 11897 11781 11931 11815
rect 11931 11781 11940 11815
rect 11888 11772 11940 11781
rect 5080 11747 5132 11756
rect 5080 11713 5114 11747
rect 5114 11713 5132 11747
rect 5080 11704 5132 11713
rect 6644 11704 6696 11756
rect 11336 11747 11388 11756
rect 11336 11713 11345 11747
rect 11345 11713 11379 11747
rect 11379 11713 11388 11747
rect 11336 11704 11388 11713
rect 11612 11704 11664 11756
rect 11796 11747 11848 11756
rect 11796 11713 11805 11747
rect 11805 11713 11839 11747
rect 11839 11713 11848 11747
rect 11796 11704 11848 11713
rect 12624 11840 12676 11892
rect 14280 11840 14332 11892
rect 15476 11883 15528 11892
rect 15476 11849 15485 11883
rect 15485 11849 15519 11883
rect 15519 11849 15528 11883
rect 15476 11840 15528 11849
rect 15936 11883 15988 11892
rect 15936 11849 15945 11883
rect 15945 11849 15979 11883
rect 15979 11849 15988 11883
rect 15936 11840 15988 11849
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 12164 11704 12216 11713
rect 13360 11772 13412 11824
rect 2964 11679 3016 11688
rect 2964 11645 2973 11679
rect 2973 11645 3007 11679
rect 3007 11645 3016 11679
rect 2964 11636 3016 11645
rect 3240 11679 3292 11688
rect 3240 11645 3249 11679
rect 3249 11645 3283 11679
rect 3283 11645 3292 11679
rect 3240 11636 3292 11645
rect 8944 11679 8996 11688
rect 8944 11645 8953 11679
rect 8953 11645 8987 11679
rect 8987 11645 8996 11679
rect 8944 11636 8996 11645
rect 9588 11636 9640 11688
rect 13820 11704 13872 11756
rect 14004 11704 14056 11756
rect 14648 11747 14700 11756
rect 14648 11713 14657 11747
rect 14657 11713 14691 11747
rect 14691 11713 14700 11747
rect 14648 11704 14700 11713
rect 13176 11636 13228 11688
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 16212 11747 16264 11756
rect 16212 11713 16221 11747
rect 16221 11713 16255 11747
rect 16255 11713 16264 11747
rect 16212 11704 16264 11713
rect 15568 11679 15620 11688
rect 15568 11645 15577 11679
rect 15577 11645 15611 11679
rect 15611 11645 15620 11679
rect 15568 11636 15620 11645
rect 1676 11568 1728 11620
rect 2136 11500 2188 11552
rect 13912 11568 13964 11620
rect 16396 11611 16448 11620
rect 16396 11577 16405 11611
rect 16405 11577 16439 11611
rect 16439 11577 16448 11611
rect 16396 11568 16448 11577
rect 3976 11500 4028 11552
rect 5540 11500 5592 11552
rect 12440 11500 12492 11552
rect 13176 11500 13228 11552
rect 14556 11500 14608 11552
rect 15108 11543 15160 11552
rect 15108 11509 15117 11543
rect 15117 11509 15151 11543
rect 15151 11509 15160 11543
rect 15108 11500 15160 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 1124 11296 1176 11348
rect 2964 11296 3016 11348
rect 3700 11296 3752 11348
rect 4068 11296 4120 11348
rect 5080 11296 5132 11348
rect 7012 11296 7064 11348
rect 8392 11296 8444 11348
rect 9956 11296 10008 11348
rect 11796 11296 11848 11348
rect 12900 11296 12952 11348
rect 12992 11296 13044 11348
rect 13820 11296 13872 11348
rect 13912 11339 13964 11348
rect 13912 11305 13921 11339
rect 13921 11305 13955 11339
rect 13955 11305 13964 11339
rect 13912 11296 13964 11305
rect 15568 11296 15620 11348
rect 16028 11296 16080 11348
rect 2872 11228 2924 11280
rect 3424 11228 3476 11280
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 2872 11092 2924 11144
rect 3792 11135 3844 11144
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 3976 11135 4028 11144
rect 3976 11101 3985 11135
rect 3985 11101 4019 11135
rect 4019 11101 4028 11135
rect 3976 11092 4028 11101
rect 2044 11067 2096 11076
rect 2044 11033 2078 11067
rect 2078 11033 2096 11067
rect 2044 11024 2096 11033
rect 2228 11024 2280 11076
rect 3056 11024 3108 11076
rect 4620 11228 4672 11280
rect 6552 11228 6604 11280
rect 11520 11228 11572 11280
rect 4804 11160 4856 11212
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 4252 11024 4304 11076
rect 4896 11092 4948 11144
rect 6644 11092 6696 11144
rect 8668 11092 8720 11144
rect 10048 11160 10100 11212
rect 10508 11160 10560 11212
rect 11336 11092 11388 11144
rect 11796 11135 11848 11144
rect 11796 11101 11805 11135
rect 11805 11101 11839 11135
rect 11839 11101 11848 11135
rect 11796 11092 11848 11101
rect 11980 11160 12032 11212
rect 13084 11228 13136 11280
rect 13268 11160 13320 11212
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13544 11160 13596 11169
rect 12164 11135 12216 11144
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 12256 11135 12308 11144
rect 12256 11101 12265 11135
rect 12265 11101 12299 11135
rect 12299 11101 12308 11135
rect 12256 11092 12308 11101
rect 6276 11024 6328 11076
rect 9496 11024 9548 11076
rect 11980 11067 12032 11076
rect 11980 11033 11989 11067
rect 11989 11033 12023 11067
rect 12023 11033 12032 11067
rect 11980 11024 12032 11033
rect 2320 10956 2372 11008
rect 2688 10956 2740 11008
rect 4160 10956 4212 11008
rect 4712 10956 4764 11008
rect 7288 10999 7340 11008
rect 7288 10965 7297 10999
rect 7297 10965 7331 10999
rect 7331 10965 7340 10999
rect 7288 10956 7340 10965
rect 10508 10956 10560 11008
rect 11704 10956 11756 11008
rect 12256 10956 12308 11008
rect 12532 11092 12584 11144
rect 12624 11092 12676 11144
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 12900 11135 12952 11144
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 12992 11135 13044 11144
rect 12992 11101 13001 11135
rect 13001 11101 13035 11135
rect 13035 11101 13044 11135
rect 12992 11092 13044 11101
rect 13176 11135 13228 11144
rect 13176 11101 13185 11135
rect 13185 11101 13219 11135
rect 13219 11101 13228 11135
rect 13176 11092 13228 11101
rect 13636 11092 13688 11144
rect 13728 11135 13780 11144
rect 13728 11101 13737 11135
rect 13737 11101 13771 11135
rect 13771 11101 13780 11135
rect 13728 11092 13780 11101
rect 14740 11160 14792 11212
rect 14188 11092 14240 11144
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 15108 11135 15160 11144
rect 15108 11101 15142 11135
rect 15142 11101 15160 11135
rect 15108 11092 15160 11101
rect 16304 11339 16356 11348
rect 16304 11305 16313 11339
rect 16313 11305 16347 11339
rect 16347 11305 16356 11339
rect 16304 11296 16356 11305
rect 13084 11024 13136 11076
rect 12624 10956 12676 11008
rect 12716 10956 12768 11008
rect 13636 10956 13688 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 2044 10752 2096 10804
rect 2780 10752 2832 10804
rect 2596 10684 2648 10736
rect 5816 10752 5868 10804
rect 6276 10752 6328 10804
rect 7840 10752 7892 10804
rect 12164 10795 12216 10804
rect 12164 10761 12173 10795
rect 12173 10761 12207 10795
rect 12207 10761 12216 10795
rect 12164 10752 12216 10761
rect 3884 10684 3936 10736
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 2228 10616 2280 10668
rect 2412 10616 2464 10668
rect 2777 10659 2829 10668
rect 2777 10625 2786 10659
rect 2786 10625 2820 10659
rect 2820 10625 2829 10659
rect 2777 10616 2829 10625
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 2964 10480 3016 10532
rect 3332 10616 3384 10668
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 3700 10616 3752 10668
rect 4252 10684 4304 10736
rect 5540 10684 5592 10736
rect 3424 10480 3476 10532
rect 2412 10455 2464 10464
rect 2412 10421 2421 10455
rect 2421 10421 2455 10455
rect 2455 10421 2464 10455
rect 2412 10412 2464 10421
rect 2504 10412 2556 10464
rect 3240 10412 3292 10464
rect 4160 10659 4212 10668
rect 4160 10625 4169 10659
rect 4169 10625 4203 10659
rect 4203 10625 4212 10659
rect 4160 10616 4212 10625
rect 4620 10616 4672 10668
rect 7288 10616 7340 10668
rect 8116 10659 8168 10668
rect 8116 10625 8125 10659
rect 8125 10625 8159 10659
rect 8159 10625 8168 10659
rect 8116 10616 8168 10625
rect 9496 10684 9548 10736
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 8300 10548 8352 10600
rect 8484 10659 8536 10668
rect 8484 10625 8493 10659
rect 8493 10625 8527 10659
rect 8527 10625 8536 10659
rect 8484 10616 8536 10625
rect 12256 10659 12308 10668
rect 12256 10625 12265 10659
rect 12265 10625 12299 10659
rect 12299 10625 12308 10659
rect 12256 10616 12308 10625
rect 12900 10752 12952 10804
rect 14004 10795 14056 10804
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 12716 10684 12768 10736
rect 12808 10616 12860 10668
rect 13268 10684 13320 10736
rect 12992 10616 13044 10668
rect 9128 10548 9180 10600
rect 9404 10591 9456 10600
rect 9404 10557 9413 10591
rect 9413 10557 9447 10591
rect 9447 10557 9456 10591
rect 9404 10548 9456 10557
rect 9588 10591 9640 10600
rect 9588 10557 9597 10591
rect 9597 10557 9631 10591
rect 9631 10557 9640 10591
rect 9588 10548 9640 10557
rect 10232 10548 10284 10600
rect 10508 10548 10560 10600
rect 11612 10548 11664 10600
rect 11980 10480 12032 10532
rect 12624 10591 12676 10600
rect 12624 10557 12633 10591
rect 12633 10557 12667 10591
rect 12667 10557 12676 10591
rect 12624 10548 12676 10557
rect 13820 10684 13872 10736
rect 14372 10684 14424 10736
rect 13728 10616 13780 10668
rect 14648 10616 14700 10668
rect 14832 10659 14884 10668
rect 14832 10625 14866 10659
rect 14866 10625 14884 10659
rect 14832 10616 14884 10625
rect 15200 10616 15252 10668
rect 14464 10548 14516 10600
rect 4712 10412 4764 10464
rect 5448 10412 5500 10464
rect 8944 10455 8996 10464
rect 8944 10421 8953 10455
rect 8953 10421 8987 10455
rect 8987 10421 8996 10455
rect 8944 10412 8996 10421
rect 10600 10455 10652 10464
rect 10600 10421 10609 10455
rect 10609 10421 10643 10455
rect 10643 10421 10652 10455
rect 10600 10412 10652 10421
rect 12440 10412 12492 10464
rect 13544 10412 13596 10464
rect 15476 10412 15528 10464
rect 15936 10455 15988 10464
rect 15936 10421 15945 10455
rect 15945 10421 15979 10455
rect 15979 10421 15988 10455
rect 15936 10412 15988 10421
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 2964 10208 3016 10260
rect 1768 10072 1820 10124
rect 1400 9979 1452 9988
rect 1400 9945 1409 9979
rect 1409 9945 1443 9979
rect 1443 9945 1452 9979
rect 1400 9936 1452 9945
rect 2412 9936 2464 9988
rect 3516 10004 3568 10056
rect 6828 10208 6880 10260
rect 9404 10208 9456 10260
rect 9496 10208 9548 10260
rect 10508 10251 10560 10260
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 11336 10208 11388 10260
rect 13636 10183 13688 10192
rect 13636 10149 13645 10183
rect 13645 10149 13679 10183
rect 13679 10149 13688 10183
rect 13636 10140 13688 10149
rect 14648 10140 14700 10192
rect 4160 9936 4212 9988
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 1676 9868 1728 9920
rect 8116 10004 8168 10056
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 5356 9936 5408 9988
rect 8760 10047 8812 10056
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 14832 10208 14884 10260
rect 10692 10004 10744 10056
rect 11704 10047 11756 10056
rect 11704 10013 11722 10047
rect 11722 10013 11756 10047
rect 11704 10004 11756 10013
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 15476 10115 15528 10124
rect 15476 10081 15485 10115
rect 15485 10081 15519 10115
rect 15519 10081 15528 10115
rect 15476 10072 15528 10081
rect 15936 10072 15988 10124
rect 16488 10072 16540 10124
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 13820 10004 13872 10056
rect 9220 9936 9272 9988
rect 10140 9936 10192 9988
rect 12716 9936 12768 9988
rect 10876 9868 10928 9920
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 4068 9664 4120 9716
rect 5080 9664 5132 9716
rect 5172 9664 5224 9716
rect 5632 9664 5684 9716
rect 10140 9707 10192 9716
rect 10140 9673 10149 9707
rect 10149 9673 10183 9707
rect 10183 9673 10192 9707
rect 10140 9664 10192 9673
rect 10600 9664 10652 9716
rect 10692 9664 10744 9716
rect 14004 9664 14056 9716
rect 3792 9596 3844 9648
rect 6368 9596 6420 9648
rect 8944 9639 8996 9648
rect 8944 9605 8978 9639
rect 8978 9605 8996 9639
rect 8944 9596 8996 9605
rect 13912 9596 13964 9648
rect 1676 9571 1728 9580
rect 1676 9537 1685 9571
rect 1685 9537 1719 9571
rect 1719 9537 1728 9571
rect 1676 9528 1728 9537
rect 2504 9528 2556 9580
rect 1032 9392 1084 9444
rect 5356 9528 5408 9580
rect 4160 9460 4212 9512
rect 4620 9460 4672 9512
rect 4712 9460 4764 9512
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 6920 9571 6972 9580
rect 6920 9537 6929 9571
rect 6929 9537 6963 9571
rect 6963 9537 6972 9571
rect 6920 9528 6972 9537
rect 7288 9528 7340 9580
rect 7472 9571 7524 9580
rect 7472 9537 7506 9571
rect 7506 9537 7524 9571
rect 7472 9528 7524 9537
rect 9220 9528 9272 9580
rect 14096 9571 14148 9580
rect 14096 9537 14105 9571
rect 14105 9537 14139 9571
rect 14139 9537 14148 9571
rect 14096 9528 14148 9537
rect 16488 9571 16540 9580
rect 16488 9537 16497 9571
rect 16497 9537 16531 9571
rect 16531 9537 16540 9571
rect 16488 9528 16540 9537
rect 1308 9324 1360 9376
rect 1676 9324 1728 9376
rect 6736 9392 6788 9444
rect 6920 9392 6972 9444
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 8576 9435 8628 9444
rect 8576 9401 8585 9435
rect 8585 9401 8619 9435
rect 8619 9401 8628 9435
rect 8576 9392 8628 9401
rect 10232 9392 10284 9444
rect 4068 9324 4120 9376
rect 7932 9324 7984 9376
rect 8300 9324 8352 9376
rect 9588 9324 9640 9376
rect 16212 9392 16264 9444
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 4436 9120 4488 9172
rect 5908 9120 5960 9172
rect 6736 9120 6788 9172
rect 7472 9120 7524 9172
rect 9036 9120 9088 9172
rect 10876 9163 10928 9172
rect 10876 9129 10885 9163
rect 10885 9129 10919 9163
rect 10919 9129 10928 9163
rect 10876 9120 10928 9129
rect 11060 9120 11112 9172
rect 12808 9120 12860 9172
rect 848 9052 900 9104
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 2780 9052 2832 9104
rect 3516 9052 3568 9104
rect 7288 9052 7340 9104
rect 2044 8916 2096 8968
rect 2596 8984 2648 9036
rect 2320 8959 2372 8968
rect 2320 8925 2329 8959
rect 2329 8925 2363 8959
rect 2363 8925 2372 8959
rect 2320 8916 2372 8925
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 3700 8916 3752 8968
rect 2596 8823 2648 8832
rect 2596 8789 2605 8823
rect 2605 8789 2639 8823
rect 2639 8789 2648 8823
rect 2596 8780 2648 8789
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 2780 8780 2832 8789
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4068 8916 4120 8925
rect 4344 8984 4396 9036
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 7932 8984 7984 9036
rect 8300 8984 8352 9036
rect 8576 8984 8628 9036
rect 9588 8984 9640 9036
rect 4712 8916 4764 8968
rect 5448 8916 5500 8968
rect 6920 8916 6972 8968
rect 5080 8848 5132 8900
rect 5356 8848 5408 8900
rect 6460 8848 6512 8900
rect 9680 8891 9732 8900
rect 9680 8857 9689 8891
rect 9689 8857 9723 8891
rect 9723 8857 9732 8891
rect 9680 8848 9732 8857
rect 6644 8780 6696 8832
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 7472 8780 7524 8789
rect 9864 8823 9916 8832
rect 9864 8789 9873 8823
rect 9873 8789 9907 8823
rect 9907 8789 9916 8823
rect 9864 8780 9916 8789
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 13268 8984 13320 9036
rect 11428 8959 11480 8968
rect 11428 8925 11437 8959
rect 11437 8925 11471 8959
rect 11471 8925 11480 8959
rect 11428 8916 11480 8925
rect 10968 8848 11020 8900
rect 12164 8916 12216 8968
rect 12532 8916 12584 8968
rect 12808 8959 12860 8968
rect 12808 8925 12817 8959
rect 12817 8925 12851 8959
rect 12851 8925 12860 8959
rect 12808 8916 12860 8925
rect 11704 8848 11756 8900
rect 12900 8848 12952 8900
rect 12164 8780 12216 8832
rect 13268 8891 13320 8900
rect 13268 8857 13277 8891
rect 13277 8857 13311 8891
rect 13311 8857 13320 8891
rect 13268 8848 13320 8857
rect 13452 8891 13504 8900
rect 13452 8857 13461 8891
rect 13461 8857 13495 8891
rect 13495 8857 13504 8891
rect 13452 8848 13504 8857
rect 14280 8959 14332 8968
rect 14280 8925 14289 8959
rect 14289 8925 14323 8959
rect 14323 8925 14332 8959
rect 14280 8916 14332 8925
rect 14372 8959 14424 8968
rect 14372 8925 14381 8959
rect 14381 8925 14415 8959
rect 14415 8925 14424 8959
rect 14372 8916 14424 8925
rect 14464 8959 14516 8968
rect 14464 8925 14473 8959
rect 14473 8925 14507 8959
rect 14507 8925 14516 8959
rect 14464 8916 14516 8925
rect 15384 8848 15436 8900
rect 13084 8823 13136 8832
rect 13084 8789 13093 8823
rect 13093 8789 13127 8823
rect 13127 8789 13136 8823
rect 13084 8780 13136 8789
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 1400 8508 1452 8560
rect 3148 8576 3200 8628
rect 2596 8508 2648 8560
rect 2964 8508 3016 8560
rect 6184 8576 6236 8628
rect 13268 8576 13320 8628
rect 15200 8576 15252 8628
rect 3884 8440 3936 8492
rect 1768 8372 1820 8424
rect 3516 8372 3568 8424
rect 3792 8372 3844 8424
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 4620 8372 4672 8424
rect 6368 8551 6420 8560
rect 6368 8517 6377 8551
rect 6377 8517 6411 8551
rect 6411 8517 6420 8551
rect 6368 8508 6420 8517
rect 6736 8508 6788 8560
rect 6920 8440 6972 8492
rect 7472 8440 7524 8492
rect 7380 8372 7432 8424
rect 6184 8347 6236 8356
rect 6184 8313 6193 8347
rect 6193 8313 6227 8347
rect 6227 8313 6236 8347
rect 6184 8304 6236 8313
rect 3056 8236 3108 8288
rect 9588 8508 9640 8560
rect 11888 8508 11940 8560
rect 8392 8440 8444 8492
rect 8852 8440 8904 8492
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9220 8440 9272 8492
rect 9772 8483 9824 8492
rect 9772 8449 9781 8483
rect 9781 8449 9815 8483
rect 9815 8449 9824 8483
rect 9772 8440 9824 8449
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 10968 8440 11020 8492
rect 11704 8440 11756 8492
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 11888 8372 11940 8424
rect 12256 8483 12308 8492
rect 12256 8449 12265 8483
rect 12265 8449 12299 8483
rect 12299 8449 12308 8483
rect 12256 8440 12308 8449
rect 14096 8508 14148 8560
rect 13176 8440 13228 8492
rect 16212 8483 16264 8492
rect 16212 8449 16221 8483
rect 16221 8449 16255 8483
rect 16255 8449 16264 8483
rect 16212 8440 16264 8449
rect 9864 8304 9916 8356
rect 16580 8304 16632 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 1768 8032 1820 8084
rect 2504 8032 2556 8084
rect 4620 8032 4672 8084
rect 6460 8032 6512 8084
rect 3608 7964 3660 8016
rect 6092 7964 6144 8016
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 3424 7828 3476 7880
rect 3976 7828 4028 7880
rect 4528 7896 4580 7948
rect 5356 7896 5408 7948
rect 9036 8032 9088 8084
rect 10692 8032 10744 8084
rect 12900 8032 12952 8084
rect 13176 8075 13228 8084
rect 13176 8041 13185 8075
rect 13185 8041 13219 8075
rect 13219 8041 13228 8075
rect 13176 8032 13228 8041
rect 14280 8032 14332 8084
rect 4252 7828 4304 7880
rect 5264 7828 5316 7880
rect 6000 7828 6052 7880
rect 6736 7871 6788 7880
rect 6736 7837 6745 7871
rect 6745 7837 6779 7871
rect 6779 7837 6788 7871
rect 6736 7828 6788 7837
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 8852 7828 8904 7880
rect 9772 7828 9824 7880
rect 11888 7828 11940 7880
rect 12164 7828 12216 7880
rect 13084 7896 13136 7948
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 1676 7803 1728 7812
rect 1676 7769 1710 7803
rect 1710 7769 1728 7803
rect 1676 7760 1728 7769
rect 4620 7803 4672 7812
rect 4620 7769 4629 7803
rect 4629 7769 4663 7803
rect 4663 7769 4672 7803
rect 4620 7760 4672 7769
rect 2964 7735 3016 7744
rect 2964 7701 2973 7735
rect 2973 7701 3007 7735
rect 3007 7701 3016 7735
rect 2964 7692 3016 7701
rect 8024 7760 8076 7812
rect 8300 7760 8352 7812
rect 8668 7760 8720 7812
rect 9496 7803 9548 7812
rect 9496 7769 9530 7803
rect 9530 7769 9548 7803
rect 9496 7760 9548 7769
rect 10140 7760 10192 7812
rect 11520 7760 11572 7812
rect 12440 7760 12492 7812
rect 12992 7828 13044 7880
rect 9312 7692 9364 7744
rect 9680 7692 9732 7744
rect 10876 7692 10928 7744
rect 12624 7692 12676 7744
rect 12808 7692 12860 7744
rect 13084 7692 13136 7744
rect 13360 7692 13412 7744
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 15108 7828 15160 7880
rect 14740 7760 14792 7812
rect 16212 7692 16264 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1676 7488 1728 7540
rect 4804 7488 4856 7540
rect 8024 7531 8076 7540
rect 8024 7497 8033 7531
rect 8033 7497 8067 7531
rect 8067 7497 8076 7531
rect 8024 7488 8076 7497
rect 9036 7488 9088 7540
rect 9404 7488 9456 7540
rect 1952 7395 2004 7404
rect 1952 7361 1961 7395
rect 1961 7361 1995 7395
rect 1995 7361 2004 7395
rect 1952 7352 2004 7361
rect 2504 7463 2556 7472
rect 2504 7429 2513 7463
rect 2513 7429 2547 7463
rect 2547 7429 2556 7463
rect 2504 7420 2556 7429
rect 2596 7352 2648 7404
rect 2872 7420 2924 7472
rect 2964 7395 3016 7404
rect 2964 7361 2973 7395
rect 2973 7361 3007 7395
rect 3007 7361 3016 7395
rect 2964 7352 3016 7361
rect 4160 7420 4212 7472
rect 4528 7420 4580 7472
rect 3700 7284 3752 7336
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 4620 7352 4672 7404
rect 5356 7352 5408 7404
rect 6184 7420 6236 7472
rect 9312 7463 9364 7472
rect 9312 7429 9321 7463
rect 9321 7429 9355 7463
rect 9355 7429 9364 7463
rect 9312 7420 9364 7429
rect 11336 7488 11388 7540
rect 11520 7531 11572 7540
rect 11520 7497 11529 7531
rect 11529 7497 11563 7531
rect 11563 7497 11572 7531
rect 11520 7488 11572 7497
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 12256 7420 12308 7472
rect 12716 7420 12768 7472
rect 9864 7352 9916 7404
rect 10876 7352 10928 7404
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11796 7395 11848 7404
rect 11796 7361 11805 7395
rect 11805 7361 11839 7395
rect 11839 7361 11848 7395
rect 11796 7352 11848 7361
rect 5448 7284 5500 7336
rect 8392 7284 8444 7336
rect 8668 7327 8720 7336
rect 8668 7293 8677 7327
rect 8677 7293 8711 7327
rect 8711 7293 8720 7327
rect 8668 7284 8720 7293
rect 10140 7284 10192 7336
rect 10692 7284 10744 7336
rect 12164 7395 12216 7404
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 12348 7352 12400 7361
rect 12624 7352 12676 7404
rect 12900 7352 12952 7404
rect 13544 7352 13596 7404
rect 14280 7352 14332 7404
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 2688 7148 2740 7200
rect 2964 7148 3016 7200
rect 4620 7148 4672 7200
rect 10600 7216 10652 7268
rect 8576 7148 8628 7200
rect 8944 7191 8996 7200
rect 8944 7157 8953 7191
rect 8953 7157 8987 7191
rect 8987 7157 8996 7191
rect 8944 7148 8996 7157
rect 9036 7148 9088 7200
rect 10508 7148 10560 7200
rect 13084 7284 13136 7336
rect 14372 7284 14424 7336
rect 14924 7352 14976 7404
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 11060 7148 11112 7200
rect 12348 7216 12400 7268
rect 11796 7148 11848 7200
rect 14464 7216 14516 7268
rect 15384 7216 15436 7268
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13452 7148 13504 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 2780 6944 2832 6996
rect 3056 6944 3108 6996
rect 1768 6808 1820 6860
rect 2044 6851 2096 6860
rect 2044 6817 2053 6851
rect 2053 6817 2087 6851
rect 2087 6817 2096 6851
rect 2044 6808 2096 6817
rect 3792 6740 3844 6792
rect 4436 6783 4488 6792
rect 4436 6749 4445 6783
rect 4445 6749 4479 6783
rect 4479 6749 4488 6783
rect 4436 6740 4488 6749
rect 4528 6740 4580 6792
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 14648 6944 14700 6996
rect 8392 6876 8444 6928
rect 13360 6876 13412 6928
rect 8668 6808 8720 6860
rect 10876 6851 10928 6860
rect 10876 6817 10885 6851
rect 10885 6817 10919 6851
rect 10919 6817 10928 6851
rect 10876 6808 10928 6817
rect 4804 6783 4856 6792
rect 4804 6749 4813 6783
rect 4813 6749 4847 6783
rect 4847 6749 4856 6783
rect 4804 6740 4856 6749
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 5356 6740 5408 6792
rect 5448 6740 5500 6792
rect 6552 6740 6604 6792
rect 7380 6783 7432 6792
rect 2688 6672 2740 6724
rect 2872 6604 2924 6656
rect 4160 6715 4212 6724
rect 4160 6681 4169 6715
rect 4169 6681 4203 6715
rect 4203 6681 4212 6715
rect 4160 6672 4212 6681
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 3792 6647 3844 6656
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4620 6604 4672 6656
rect 4712 6604 4764 6656
rect 6000 6647 6052 6656
rect 6000 6613 6009 6647
rect 6009 6613 6043 6647
rect 6043 6613 6052 6647
rect 6000 6604 6052 6613
rect 6920 6672 6972 6724
rect 7840 6783 7892 6792
rect 7840 6749 7849 6783
rect 7849 6749 7883 6783
rect 7883 6749 7892 6783
rect 7840 6740 7892 6749
rect 7932 6783 7984 6792
rect 7932 6749 7941 6783
rect 7941 6749 7975 6783
rect 7975 6749 7984 6783
rect 7932 6740 7984 6749
rect 8024 6740 8076 6792
rect 11796 6740 11848 6792
rect 14280 6783 14332 6792
rect 14280 6749 14289 6783
rect 14289 6749 14323 6783
rect 14323 6749 14332 6783
rect 14280 6740 14332 6749
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 14924 6808 14976 6860
rect 11152 6715 11204 6724
rect 11152 6681 11161 6715
rect 11161 6681 11195 6715
rect 11195 6681 11204 6715
rect 11152 6672 11204 6681
rect 13452 6672 13504 6724
rect 14372 6672 14424 6724
rect 10048 6604 10100 6656
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 13268 6604 13320 6656
rect 15108 6740 15160 6792
rect 15844 6604 15896 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 2688 6443 2740 6452
rect 2688 6409 2697 6443
rect 2697 6409 2731 6443
rect 2731 6409 2740 6443
rect 2688 6400 2740 6409
rect 4528 6443 4580 6452
rect 4528 6409 4537 6443
rect 4537 6409 4571 6443
rect 4571 6409 4580 6443
rect 4528 6400 4580 6409
rect 4620 6400 4672 6452
rect 5264 6400 5316 6452
rect 7012 6400 7064 6452
rect 7932 6400 7984 6452
rect 8668 6400 8720 6452
rect 11152 6400 11204 6452
rect 11888 6400 11940 6452
rect 14464 6400 14516 6452
rect 2964 6307 3016 6316
rect 2964 6273 2973 6307
rect 2973 6273 3007 6307
rect 3007 6273 3016 6307
rect 2964 6264 3016 6273
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3792 6332 3844 6384
rect 4436 6332 4488 6384
rect 4160 6307 4212 6316
rect 4160 6273 4169 6307
rect 4169 6273 4203 6307
rect 4203 6273 4212 6307
rect 4160 6264 4212 6273
rect 5448 6332 5500 6384
rect 6000 6332 6052 6384
rect 9588 6332 9640 6384
rect 12348 6332 12400 6384
rect 13544 6332 13596 6384
rect 3884 6060 3936 6112
rect 4712 6264 4764 6316
rect 4804 6060 4856 6112
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7012 6307 7064 6316
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 8852 6264 8904 6316
rect 9036 6264 9088 6316
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 9864 6264 9916 6316
rect 11244 6264 11296 6316
rect 7104 6196 7156 6248
rect 8944 6128 8996 6180
rect 10140 6060 10192 6112
rect 10232 6060 10284 6112
rect 11428 6060 11480 6112
rect 12808 6239 12860 6248
rect 12808 6205 12817 6239
rect 12817 6205 12851 6239
rect 12851 6205 12860 6239
rect 12808 6196 12860 6205
rect 13268 6239 13320 6248
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 13912 6264 13964 6316
rect 14372 6332 14424 6384
rect 16212 6400 16264 6452
rect 15384 6375 15436 6384
rect 15384 6341 15418 6375
rect 15418 6341 15436 6375
rect 15384 6332 15436 6341
rect 14464 6307 14516 6316
rect 14464 6273 14473 6307
rect 14473 6273 14507 6307
rect 14507 6273 14516 6307
rect 14464 6264 14516 6273
rect 14648 6307 14700 6316
rect 14648 6273 14657 6307
rect 14657 6273 14691 6307
rect 14691 6273 14700 6307
rect 14648 6264 14700 6273
rect 14832 6307 14884 6316
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 15844 6264 15896 6316
rect 15108 6239 15160 6248
rect 15108 6205 15117 6239
rect 15117 6205 15151 6239
rect 15151 6205 15160 6239
rect 15108 6196 15160 6205
rect 13820 6128 13872 6180
rect 14004 6128 14056 6180
rect 14464 6128 14516 6180
rect 14924 6128 14976 6180
rect 14648 6060 14700 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2228 5788 2280 5840
rect 2596 5788 2648 5840
rect 3056 5788 3108 5840
rect 2872 5720 2924 5772
rect 7012 5788 7064 5840
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 1768 5652 1820 5704
rect 2228 5695 2280 5704
rect 2228 5661 2237 5695
rect 2237 5661 2271 5695
rect 2271 5661 2280 5695
rect 2228 5652 2280 5661
rect 2320 5652 2372 5704
rect 5356 5720 5408 5772
rect 3240 5695 3292 5704
rect 3240 5661 3249 5695
rect 3249 5661 3283 5695
rect 3283 5661 3292 5695
rect 3240 5652 3292 5661
rect 3516 5652 3568 5704
rect 3884 5652 3936 5704
rect 2136 5584 2188 5636
rect 8392 5720 8444 5772
rect 7012 5652 7064 5704
rect 7564 5584 7616 5636
rect 8852 5720 8904 5772
rect 8760 5652 8812 5704
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 1584 5516 1636 5568
rect 1952 5516 2004 5568
rect 2780 5559 2832 5568
rect 2780 5525 2789 5559
rect 2789 5525 2823 5559
rect 2823 5525 2832 5559
rect 2780 5516 2832 5525
rect 7656 5559 7708 5568
rect 7656 5525 7665 5559
rect 7665 5525 7699 5559
rect 7699 5525 7708 5559
rect 7656 5516 7708 5525
rect 8668 5584 8720 5636
rect 9588 5695 9640 5704
rect 9588 5661 9597 5695
rect 9597 5661 9631 5695
rect 9631 5661 9640 5695
rect 9588 5652 9640 5661
rect 10140 5720 10192 5772
rect 11060 5652 11112 5704
rect 11244 5652 11296 5704
rect 11980 5652 12032 5704
rect 15200 5788 15252 5840
rect 13084 5652 13136 5704
rect 16212 5695 16264 5704
rect 16212 5661 16221 5695
rect 16221 5661 16255 5695
rect 16255 5661 16264 5695
rect 16212 5652 16264 5661
rect 8944 5516 8996 5568
rect 9956 5584 10008 5636
rect 10232 5584 10284 5636
rect 10416 5584 10468 5636
rect 10508 5516 10560 5568
rect 11060 5516 11112 5568
rect 12440 5516 12492 5568
rect 12992 5584 13044 5636
rect 13452 5584 13504 5636
rect 14372 5627 14424 5636
rect 14372 5593 14381 5627
rect 14381 5593 14415 5627
rect 14415 5593 14424 5627
rect 14372 5584 14424 5593
rect 14556 5559 14608 5568
rect 14556 5525 14565 5559
rect 14565 5525 14599 5559
rect 14599 5525 14608 5559
rect 14556 5516 14608 5525
rect 16580 5516 16632 5568
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 2320 5312 2372 5364
rect 3240 5312 3292 5364
rect 3884 5312 3936 5364
rect 2780 5244 2832 5296
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 1952 5219 2004 5228
rect 1952 5185 1961 5219
rect 1961 5185 1995 5219
rect 1995 5185 2004 5219
rect 1952 5176 2004 5185
rect 3516 5176 3568 5228
rect 2044 5108 2096 5160
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 2964 4972 3016 5024
rect 4068 5219 4120 5228
rect 4068 5185 4077 5219
rect 4077 5185 4111 5219
rect 4111 5185 4120 5219
rect 4068 5176 4120 5185
rect 4712 5219 4764 5228
rect 4712 5185 4721 5219
rect 4721 5185 4755 5219
rect 4755 5185 4764 5219
rect 4712 5176 4764 5185
rect 8024 5312 8076 5364
rect 5172 5176 5224 5228
rect 6828 5244 6880 5296
rect 5356 5219 5408 5228
rect 5356 5185 5365 5219
rect 5365 5185 5399 5219
rect 5399 5185 5408 5219
rect 5356 5176 5408 5185
rect 5540 5176 5592 5228
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 7012 5176 7064 5228
rect 7196 5219 7248 5228
rect 7196 5185 7230 5219
rect 7230 5185 7248 5219
rect 7196 5176 7248 5185
rect 10140 5244 10192 5296
rect 8944 5219 8996 5228
rect 8944 5185 8978 5219
rect 8978 5185 8996 5219
rect 8944 5176 8996 5185
rect 9220 5176 9272 5228
rect 10600 5219 10652 5228
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 10600 5176 10652 5185
rect 11336 5312 11388 5364
rect 12348 5312 12400 5364
rect 12992 5355 13044 5364
rect 12992 5321 13001 5355
rect 13001 5321 13035 5355
rect 13035 5321 13044 5355
rect 12992 5312 13044 5321
rect 14372 5312 14424 5364
rect 11980 5287 12032 5296
rect 11980 5253 11989 5287
rect 11989 5253 12023 5287
rect 12023 5253 12032 5287
rect 11980 5244 12032 5253
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 9680 5108 9732 5160
rect 11060 5176 11112 5228
rect 11244 5176 11296 5228
rect 11888 5219 11940 5228
rect 11888 5185 11897 5219
rect 11897 5185 11931 5219
rect 11931 5185 11940 5219
rect 11888 5176 11940 5185
rect 12072 5219 12124 5228
rect 12072 5185 12081 5219
rect 12081 5185 12115 5219
rect 12115 5185 12124 5219
rect 12072 5176 12124 5185
rect 12440 5176 12492 5228
rect 12808 5244 12860 5296
rect 13084 5244 13136 5296
rect 15108 5244 15160 5296
rect 15660 5244 15712 5296
rect 4620 4972 4672 5024
rect 5540 5040 5592 5092
rect 5908 5040 5960 5092
rect 10416 5040 10468 5092
rect 5724 5015 5776 5024
rect 5724 4981 5733 5015
rect 5733 4981 5767 5015
rect 5767 4981 5776 5015
rect 5724 4972 5776 4981
rect 7564 4972 7616 5024
rect 9588 4972 9640 5024
rect 10968 5040 11020 5092
rect 11888 5040 11940 5092
rect 12348 5040 12400 5092
rect 14096 5176 14148 5228
rect 14188 5176 14240 5228
rect 14924 5176 14976 5228
rect 14648 5108 14700 5160
rect 15568 5219 15620 5228
rect 15568 5185 15577 5219
rect 15577 5185 15611 5219
rect 15611 5185 15620 5219
rect 15568 5176 15620 5185
rect 14740 4972 14792 5024
rect 15016 5015 15068 5024
rect 15016 4981 15025 5015
rect 15025 4981 15059 5015
rect 15059 4981 15068 5015
rect 15016 4972 15068 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2136 4768 2188 4820
rect 2044 4564 2096 4616
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 3976 4768 4028 4820
rect 7012 4768 7064 4820
rect 7196 4811 7248 4820
rect 7196 4777 7205 4811
rect 7205 4777 7239 4811
rect 7239 4777 7248 4811
rect 7196 4768 7248 4777
rect 7840 4700 7892 4752
rect 8944 4743 8996 4752
rect 8944 4709 8953 4743
rect 8953 4709 8987 4743
rect 8987 4709 8996 4743
rect 8944 4700 8996 4709
rect 14096 4811 14148 4820
rect 14096 4777 14105 4811
rect 14105 4777 14139 4811
rect 14139 4777 14148 4811
rect 14096 4768 14148 4777
rect 15016 4700 15068 4752
rect 2964 4564 3016 4616
rect 3516 4564 3568 4616
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4068 4564 4120 4573
rect 4620 4564 4672 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 8208 4632 8260 4684
rect 1492 4496 1544 4548
rect 5724 4496 5776 4548
rect 5908 4496 5960 4548
rect 6828 4496 6880 4548
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 8024 4564 8076 4616
rect 9220 4607 9272 4616
rect 8392 4539 8444 4548
rect 8392 4505 8401 4539
rect 8401 4505 8435 4539
rect 8435 4505 8444 4539
rect 8392 4496 8444 4505
rect 2872 4428 2924 4480
rect 4620 4428 4672 4480
rect 5632 4428 5684 4480
rect 9220 4573 9229 4607
rect 9229 4573 9263 4607
rect 9263 4573 9272 4607
rect 9220 4564 9272 4573
rect 13268 4632 13320 4684
rect 12164 4564 12216 4616
rect 9680 4496 9732 4548
rect 13912 4564 13964 4616
rect 14096 4632 14148 4684
rect 14280 4564 14332 4616
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 14648 4632 14700 4684
rect 15108 4675 15160 4684
rect 15108 4641 15117 4675
rect 15117 4641 15151 4675
rect 15151 4641 15160 4675
rect 15108 4632 15160 4641
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 8852 4428 8904 4480
rect 9496 4428 9548 4480
rect 9588 4428 9640 4480
rect 14556 4428 14608 4480
rect 15108 4496 15160 4548
rect 15568 4428 15620 4480
rect 16488 4471 16540 4480
rect 16488 4437 16497 4471
rect 16497 4437 16531 4471
rect 16531 4437 16540 4471
rect 16488 4428 16540 4437
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 4712 4224 4764 4276
rect 7196 4224 7248 4276
rect 2872 4156 2924 4208
rect 3976 4156 4028 4208
rect 4620 4156 4672 4208
rect 6552 4156 6604 4208
rect 2136 4088 2188 4140
rect 2780 4088 2832 4140
rect 3516 4088 3568 4140
rect 3700 4088 3752 4140
rect 7564 4156 7616 4208
rect 7840 4199 7892 4208
rect 7840 4165 7849 4199
rect 7849 4165 7883 4199
rect 7883 4165 7892 4199
rect 7840 4156 7892 4165
rect 8392 4224 8444 4276
rect 9680 4224 9732 4276
rect 11612 4224 11664 4276
rect 7196 4088 7248 4140
rect 8760 4156 8812 4208
rect 9588 4156 9640 4208
rect 6828 4020 6880 4072
rect 10048 4088 10100 4140
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 8300 4020 8352 4072
rect 9772 4020 9824 4072
rect 11244 4088 11296 4140
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 3148 3952 3200 4004
rect 3332 3952 3384 4004
rect 7288 3995 7340 4004
rect 7288 3961 7297 3995
rect 7297 3961 7331 3995
rect 7331 3961 7340 3995
rect 7288 3952 7340 3961
rect 8484 3952 8536 4004
rect 9680 3952 9732 4004
rect 11612 4020 11664 4072
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 11980 4088 12032 4140
rect 12808 4224 12860 4276
rect 14096 4224 14148 4276
rect 14280 4224 14332 4276
rect 14372 4224 14424 4276
rect 13452 4156 13504 4208
rect 13544 4156 13596 4208
rect 12256 4020 12308 4072
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13820 4088 13872 4140
rect 14188 4131 14240 4140
rect 14188 4097 14197 4131
rect 14197 4097 14231 4131
rect 14231 4097 14240 4131
rect 14188 4088 14240 4097
rect 14280 4088 14332 4140
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 14556 4088 14608 4140
rect 14924 4156 14976 4208
rect 15568 4088 15620 4140
rect 15844 4131 15896 4140
rect 15844 4097 15853 4131
rect 15853 4097 15887 4131
rect 15887 4097 15896 4131
rect 15844 4088 15896 4097
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 15108 4063 15160 4072
rect 15108 4029 15117 4063
rect 15117 4029 15151 4063
rect 15151 4029 15160 4063
rect 15108 4020 15160 4029
rect 11520 3995 11572 4004
rect 11520 3961 11529 3995
rect 11529 3961 11563 3995
rect 11563 3961 11572 3995
rect 11520 3952 11572 3961
rect 12532 3952 12584 4004
rect 17408 4020 17460 4072
rect 16764 3952 16816 4004
rect 1400 3884 1452 3936
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 2320 3884 2372 3936
rect 3424 3884 3476 3936
rect 10232 3927 10284 3936
rect 10232 3893 10241 3927
rect 10241 3893 10275 3927
rect 10275 3893 10284 3927
rect 10232 3884 10284 3893
rect 11888 3884 11940 3936
rect 14096 3884 14148 3936
rect 14464 3884 14516 3936
rect 16120 3884 16172 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 3608 3680 3660 3732
rect 3056 3612 3108 3664
rect 2412 3544 2464 3596
rect 6828 3680 6880 3732
rect 7288 3680 7340 3732
rect 10048 3680 10100 3732
rect 12348 3680 12400 3732
rect 13084 3680 13136 3732
rect 13360 3680 13412 3732
rect 14372 3612 14424 3664
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 1952 3519 2004 3528
rect 1952 3485 1961 3519
rect 1961 3485 1995 3519
rect 1995 3485 2004 3519
rect 1952 3476 2004 3485
rect 2964 3476 3016 3528
rect 3240 3519 3292 3528
rect 3240 3485 3249 3519
rect 3249 3485 3283 3519
rect 3283 3485 3292 3519
rect 3240 3476 3292 3485
rect 3884 3519 3936 3528
rect 3884 3485 3893 3519
rect 3893 3485 3927 3519
rect 3927 3485 3936 3519
rect 3884 3476 3936 3485
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 2504 3383 2556 3392
rect 2504 3349 2513 3383
rect 2513 3349 2547 3383
rect 2547 3349 2556 3383
rect 2504 3340 2556 3349
rect 2596 3340 2648 3392
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 4252 3476 4304 3485
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5448 3476 5500 3528
rect 7288 3519 7340 3528
rect 7288 3485 7297 3519
rect 7297 3485 7331 3519
rect 7331 3485 7340 3519
rect 7288 3476 7340 3485
rect 8208 3544 8260 3596
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 8024 3476 8076 3528
rect 5172 3408 5224 3460
rect 8576 3519 8628 3528
rect 8576 3485 8585 3519
rect 8585 3485 8619 3519
rect 8619 3485 8628 3519
rect 8576 3476 8628 3485
rect 13268 3544 13320 3596
rect 9588 3476 9640 3528
rect 9680 3519 9732 3528
rect 9680 3485 9689 3519
rect 9689 3485 9723 3519
rect 9723 3485 9732 3519
rect 9680 3476 9732 3485
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10232 3476 10284 3528
rect 12440 3476 12492 3528
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 13820 3544 13872 3596
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 14372 3519 14424 3528
rect 14372 3485 14381 3519
rect 14381 3485 14415 3519
rect 14415 3485 14424 3519
rect 14372 3476 14424 3485
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 14556 3519 14608 3528
rect 14556 3485 14565 3519
rect 14565 3485 14599 3519
rect 14599 3485 14608 3519
rect 14556 3476 14608 3485
rect 14740 3476 14792 3528
rect 15476 3612 15528 3664
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 16028 3519 16080 3528
rect 16028 3485 16037 3519
rect 16037 3485 16071 3519
rect 16071 3485 16080 3519
rect 16028 3476 16080 3485
rect 11888 3451 11940 3460
rect 4160 3340 4212 3392
rect 4528 3383 4580 3392
rect 4528 3349 4537 3383
rect 4537 3349 4571 3383
rect 4571 3349 4580 3383
rect 4528 3340 4580 3349
rect 4988 3340 5040 3392
rect 11888 3417 11922 3451
rect 11922 3417 11940 3451
rect 11888 3408 11940 3417
rect 7012 3383 7064 3392
rect 7012 3349 7021 3383
rect 7021 3349 7055 3383
rect 7055 3349 7064 3383
rect 7012 3340 7064 3349
rect 8116 3383 8168 3392
rect 8116 3349 8125 3383
rect 8125 3349 8159 3383
rect 8159 3349 8168 3383
rect 8116 3340 8168 3349
rect 9588 3340 9640 3392
rect 10048 3340 10100 3392
rect 10968 3340 11020 3392
rect 11980 3340 12032 3392
rect 13084 3383 13136 3392
rect 13084 3349 13093 3383
rect 13093 3349 13127 3383
rect 13127 3349 13136 3383
rect 13084 3340 13136 3349
rect 14188 3340 14240 3392
rect 14740 3340 14792 3392
rect 14924 3340 14976 3392
rect 15108 3340 15160 3392
rect 15384 3340 15436 3392
rect 15844 3383 15896 3392
rect 15844 3349 15853 3383
rect 15853 3349 15887 3383
rect 15887 3349 15896 3383
rect 15844 3340 15896 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 1676 3068 1728 3120
rect 2780 3136 2832 3188
rect 4160 3179 4212 3188
rect 4160 3145 4169 3179
rect 4169 3145 4203 3179
rect 4203 3145 4212 3179
rect 4160 3136 4212 3145
rect 4804 3136 4856 3188
rect 8300 3136 8352 3188
rect 9864 3136 9916 3188
rect 4528 3111 4580 3120
rect 2044 3000 2096 3052
rect 4528 3077 4562 3111
rect 4562 3077 4580 3111
rect 4528 3068 4580 3077
rect 5448 3068 5500 3120
rect 6828 3068 6880 3120
rect 7012 3068 7064 3120
rect 2228 3000 2280 3052
rect 2596 3043 2648 3052
rect 2596 3009 2630 3043
rect 2630 3009 2648 3043
rect 2596 3000 2648 3009
rect 3148 3000 3200 3052
rect 3884 3000 3936 3052
rect 4068 3000 4120 3052
rect 3700 2839 3752 2848
rect 3700 2805 3709 2839
rect 3709 2805 3743 2839
rect 3743 2805 3752 2839
rect 3700 2796 3752 2805
rect 5816 2932 5868 2984
rect 8116 3000 8168 3052
rect 10140 3068 10192 3120
rect 11244 3068 11296 3120
rect 12992 3136 13044 3188
rect 13544 3136 13596 3188
rect 14464 3136 14516 3188
rect 16028 3179 16080 3188
rect 16028 3145 16037 3179
rect 16037 3145 16071 3179
rect 16071 3145 16080 3179
rect 16028 3136 16080 3145
rect 11888 3111 11940 3120
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 9588 3000 9640 3052
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 14648 3068 14700 3120
rect 4068 2864 4120 2916
rect 6552 2864 6604 2916
rect 11428 2932 11480 2984
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 13084 3000 13136 3052
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 12440 2932 12492 2941
rect 10968 2864 11020 2916
rect 6184 2796 6236 2848
rect 9128 2796 9180 2848
rect 13912 2864 13964 2916
rect 14280 3000 14332 3052
rect 14924 3043 14976 3052
rect 14924 3009 14958 3043
rect 14958 3009 14976 3043
rect 14924 3000 14976 3009
rect 15200 3000 15252 3052
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 14556 2796 14608 2848
rect 16304 2839 16356 2848
rect 16304 2805 16313 2839
rect 16313 2805 16347 2839
rect 16347 2805 16356 2839
rect 16304 2796 16356 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 2780 2635 2832 2644
rect 2780 2601 2789 2635
rect 2789 2601 2823 2635
rect 2823 2601 2832 2635
rect 2780 2592 2832 2601
rect 3240 2592 3292 2644
rect 2228 2388 2280 2440
rect 3700 2388 3752 2440
rect 4620 2388 4672 2440
rect 4712 2431 4764 2440
rect 4712 2397 4721 2431
rect 4721 2397 4755 2431
rect 4755 2397 4764 2431
rect 4712 2388 4764 2397
rect 6920 2592 6972 2644
rect 7472 2592 7524 2644
rect 8576 2592 8628 2644
rect 14372 2592 14424 2644
rect 15108 2592 15160 2644
rect 5816 2524 5868 2576
rect 8024 2524 8076 2576
rect 5448 2431 5500 2440
rect 5448 2397 5457 2431
rect 5457 2397 5491 2431
rect 5491 2397 5500 2431
rect 5448 2388 5500 2397
rect 6000 2388 6052 2440
rect 6184 2431 6236 2440
rect 6184 2397 6193 2431
rect 6193 2397 6227 2431
rect 6227 2397 6236 2431
rect 6184 2388 6236 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 6644 2388 6696 2440
rect 7288 2388 7340 2440
rect 9496 2456 9548 2508
rect 7564 2388 7616 2440
rect 8300 2388 8352 2440
rect 9956 2388 10008 2440
rect 12256 2456 12308 2508
rect 1492 2320 1544 2372
rect 3792 2320 3844 2372
rect 3884 2252 3936 2304
rect 4528 2295 4580 2304
rect 4528 2261 4537 2295
rect 4537 2261 4571 2295
rect 4571 2261 4580 2295
rect 4528 2252 4580 2261
rect 5172 2252 5224 2304
rect 6460 2320 6512 2372
rect 8392 2363 8444 2372
rect 8392 2329 8401 2363
rect 8401 2329 8435 2363
rect 8435 2329 8444 2363
rect 8392 2320 8444 2329
rect 11428 2388 11480 2440
rect 11980 2431 12032 2440
rect 11980 2397 11989 2431
rect 11989 2397 12023 2431
rect 12023 2397 12032 2431
rect 11980 2388 12032 2397
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 14464 2456 14516 2508
rect 14648 2456 14700 2508
rect 15384 2431 15436 2440
rect 15384 2397 15418 2431
rect 15418 2397 15436 2431
rect 15384 2388 15436 2397
rect 11060 2320 11112 2372
rect 13268 2320 13320 2372
rect 15568 2320 15620 2372
rect 7012 2252 7064 2304
rect 7748 2295 7800 2304
rect 7748 2261 7757 2295
rect 7757 2261 7791 2295
rect 7791 2261 7800 2295
rect 7748 2252 7800 2261
rect 8300 2252 8352 2304
rect 9036 2252 9088 2304
rect 9680 2252 9732 2304
rect 10324 2252 10376 2304
rect 10968 2252 11020 2304
rect 11612 2252 11664 2304
rect 12256 2252 12308 2304
rect 12900 2252 12952 2304
rect 13544 2252 13596 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 20 1300 72 1352
rect 1584 1300 1636 1352
rect 14188 1300 14240 1352
rect 16304 1300 16356 1352
rect 664 1232 716 1284
rect 2320 1232 2372 1284
rect 14832 1096 14884 1148
rect 15844 1096 15896 1148
<< metal2 >>
rect 10966 41200 11022 42000
rect 12898 41200 12954 42000
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 8668 39636 8720 39642
rect 8668 39578 8720 39584
rect 8208 39364 8260 39370
rect 8208 39306 8260 39312
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 110 39128 166 39137
rect 4874 39131 5182 39140
rect 110 39063 166 39072
rect 124 21962 152 39063
rect 7012 39024 7064 39030
rect 7012 38966 7064 38972
rect 7380 39024 7432 39030
rect 7380 38966 7432 38972
rect 6920 38956 6972 38962
rect 6920 38898 6972 38904
rect 6092 38888 6144 38894
rect 6092 38830 6144 38836
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 6104 38418 6132 38830
rect 6092 38412 6144 38418
rect 6092 38354 6144 38360
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 2964 36848 3016 36854
rect 2964 36790 3016 36796
rect 2044 36712 2096 36718
rect 2044 36654 2096 36660
rect 2056 36378 2084 36654
rect 2780 36576 2832 36582
rect 2780 36518 2832 36524
rect 2044 36372 2096 36378
rect 2044 36314 2096 36320
rect 2792 36174 2820 36518
rect 2136 36168 2188 36174
rect 2136 36110 2188 36116
rect 2780 36168 2832 36174
rect 2780 36110 2832 36116
rect 2148 35698 2176 36110
rect 2976 35834 3004 36790
rect 6104 36786 6132 38354
rect 6644 38276 6696 38282
rect 6644 38218 6696 38224
rect 6656 38010 6684 38218
rect 6644 38004 6696 38010
rect 6644 37946 6696 37952
rect 6932 37670 6960 38898
rect 7024 37942 7052 38966
rect 7104 38956 7156 38962
rect 7156 38916 7236 38944
rect 7104 38898 7156 38904
rect 7104 38752 7156 38758
rect 7104 38694 7156 38700
rect 7116 38010 7144 38694
rect 7208 38010 7236 38916
rect 7392 38486 7420 38966
rect 8220 38962 8248 39306
rect 8208 38956 8260 38962
rect 8208 38898 8260 38904
rect 7932 38752 7984 38758
rect 7932 38694 7984 38700
rect 7944 38554 7972 38694
rect 7748 38548 7800 38554
rect 7748 38490 7800 38496
rect 7932 38548 7984 38554
rect 7932 38490 7984 38496
rect 7380 38480 7432 38486
rect 7380 38422 7432 38428
rect 7564 38208 7616 38214
rect 7564 38150 7616 38156
rect 7656 38208 7708 38214
rect 7656 38150 7708 38156
rect 7104 38004 7156 38010
rect 7104 37946 7156 37952
rect 7196 38004 7248 38010
rect 7196 37946 7248 37952
rect 7012 37936 7064 37942
rect 7012 37878 7064 37884
rect 6828 37664 6880 37670
rect 6828 37606 6880 37612
rect 6920 37664 6972 37670
rect 6920 37606 6972 37612
rect 6840 37466 6868 37606
rect 6828 37460 6880 37466
rect 6828 37402 6880 37408
rect 6736 37120 6788 37126
rect 6736 37062 6788 37068
rect 6748 36854 6776 37062
rect 6736 36848 6788 36854
rect 6736 36790 6788 36796
rect 4068 36780 4120 36786
rect 4068 36722 4120 36728
rect 6092 36780 6144 36786
rect 6092 36722 6144 36728
rect 3608 36712 3660 36718
rect 3608 36654 3660 36660
rect 3620 36174 3648 36654
rect 3976 36576 4028 36582
rect 3976 36518 4028 36524
rect 3988 36258 4016 36518
rect 4080 36378 4108 36722
rect 5356 36576 5408 36582
rect 5356 36518 5408 36524
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4068 36372 4120 36378
rect 4068 36314 4120 36320
rect 4160 36372 4212 36378
rect 4160 36314 4212 36320
rect 4172 36258 4200 36314
rect 3988 36230 4200 36258
rect 3608 36168 3660 36174
rect 3608 36110 3660 36116
rect 3240 36032 3292 36038
rect 3240 35974 3292 35980
rect 2964 35828 3016 35834
rect 2964 35770 3016 35776
rect 3252 35766 3280 35974
rect 3240 35760 3292 35766
rect 3240 35702 3292 35708
rect 2136 35692 2188 35698
rect 2136 35634 2188 35640
rect 2148 35290 2176 35634
rect 2136 35284 2188 35290
rect 2136 35226 2188 35232
rect 2148 34678 2176 35226
rect 3620 35086 3648 36110
rect 4172 35578 4200 36230
rect 4712 36236 4764 36242
rect 4712 36178 4764 36184
rect 4816 36230 5028 36258
rect 4528 36168 4580 36174
rect 4528 36110 4580 36116
rect 4540 35766 4568 36110
rect 4620 36032 4672 36038
rect 4620 35974 4672 35980
rect 4528 35760 4580 35766
rect 4528 35702 4580 35708
rect 3988 35550 4200 35578
rect 3608 35080 3660 35086
rect 3608 35022 3660 35028
rect 3988 35034 4016 35550
rect 4160 35488 4212 35494
rect 4080 35448 4160 35476
rect 4080 35222 4108 35448
rect 4160 35430 4212 35436
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4632 35290 4660 35974
rect 4724 35680 4752 36178
rect 4816 36174 4844 36230
rect 4804 36168 4856 36174
rect 4804 36110 4856 36116
rect 4896 36168 4948 36174
rect 4896 36110 4948 36116
rect 4908 36020 4936 36110
rect 5000 36038 5028 36230
rect 5368 36174 5396 36518
rect 5356 36168 5408 36174
rect 5356 36110 5408 36116
rect 5632 36168 5684 36174
rect 5632 36110 5684 36116
rect 5908 36168 5960 36174
rect 5908 36110 5960 36116
rect 5172 36100 5224 36106
rect 5224 36060 5304 36088
rect 5172 36042 5224 36048
rect 4816 35992 4936 36020
rect 4988 36032 5040 36038
rect 4816 35834 4844 35992
rect 4988 35974 5040 35980
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 5276 35834 5304 36060
rect 5356 36032 5408 36038
rect 5356 35974 5408 35980
rect 4804 35828 4856 35834
rect 4804 35770 4856 35776
rect 5264 35828 5316 35834
rect 5264 35770 5316 35776
rect 4804 35692 4856 35698
rect 4724 35652 4804 35680
rect 4804 35634 4856 35640
rect 5368 35630 5396 35974
rect 5540 35828 5592 35834
rect 5540 35770 5592 35776
rect 5552 35698 5580 35770
rect 5644 35698 5672 36110
rect 5540 35692 5592 35698
rect 5540 35634 5592 35640
rect 5632 35692 5684 35698
rect 5632 35634 5684 35640
rect 5724 35692 5776 35698
rect 5724 35634 5776 35640
rect 5356 35624 5408 35630
rect 5356 35566 5408 35572
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 5356 35488 5408 35494
rect 5356 35430 5408 35436
rect 4620 35284 4672 35290
rect 4620 35226 4672 35232
rect 4068 35216 4120 35222
rect 4068 35158 4120 35164
rect 3056 35012 3108 35018
rect 3056 34954 3108 34960
rect 3068 34746 3096 34954
rect 3056 34740 3108 34746
rect 3056 34682 3108 34688
rect 2136 34672 2188 34678
rect 2136 34614 2188 34620
rect 2872 34468 2924 34474
rect 2872 34410 2924 34416
rect 2884 31804 2912 34410
rect 3620 33590 3648 35022
rect 3988 35006 4200 35034
rect 4172 34950 4200 35006
rect 4160 34944 4212 34950
rect 4160 34886 4212 34892
rect 4172 34474 4200 34886
rect 4160 34468 4212 34474
rect 4160 34410 4212 34416
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4528 34196 4580 34202
rect 4528 34138 4580 34144
rect 4160 34128 4212 34134
rect 4160 34070 4212 34076
rect 3976 33924 4028 33930
rect 3976 33866 4028 33872
rect 3608 33584 3660 33590
rect 3608 33526 3660 33532
rect 2964 33516 3016 33522
rect 2964 33458 3016 33464
rect 2976 33114 3004 33458
rect 3884 33312 3936 33318
rect 3884 33254 3936 33260
rect 2964 33108 3016 33114
rect 2964 33050 3016 33056
rect 3896 32910 3924 33254
rect 3884 32904 3936 32910
rect 3884 32846 3936 32852
rect 3988 32774 4016 33866
rect 4172 33300 4200 34070
rect 4436 34060 4488 34066
rect 4436 34002 4488 34008
rect 4344 33992 4396 33998
rect 4344 33934 4396 33940
rect 4356 33522 4384 33934
rect 4448 33522 4476 34002
rect 4540 33658 4568 34138
rect 4724 33998 4752 35430
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4712 33992 4764 33998
rect 4712 33934 4764 33940
rect 4620 33856 4672 33862
rect 4620 33798 4672 33804
rect 4804 33856 4856 33862
rect 4804 33798 4856 33804
rect 4632 33674 4660 33798
rect 4528 33652 4580 33658
rect 4632 33646 4752 33674
rect 4528 33594 4580 33600
rect 4620 33584 4672 33590
rect 4620 33526 4672 33532
rect 4344 33516 4396 33522
rect 4344 33458 4396 33464
rect 4436 33516 4488 33522
rect 4436 33458 4488 33464
rect 4356 33318 4384 33458
rect 4080 33272 4200 33300
rect 4344 33312 4396 33318
rect 4080 33046 4108 33272
rect 4344 33254 4396 33260
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4068 33040 4120 33046
rect 4120 32988 4200 32994
rect 4068 32982 4200 32988
rect 4080 32966 4200 32982
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 3976 32768 4028 32774
rect 3976 32710 4028 32716
rect 4068 32768 4120 32774
rect 4068 32710 4120 32716
rect 2964 31816 3016 31822
rect 2884 31776 2964 31804
rect 2964 31758 3016 31764
rect 2976 30326 3004 31758
rect 3148 30592 3200 30598
rect 3148 30534 3200 30540
rect 2964 30320 3016 30326
rect 2964 30262 3016 30268
rect 2228 29640 2280 29646
rect 2228 29582 2280 29588
rect 2240 27538 2268 29582
rect 2504 29572 2556 29578
rect 2504 29514 2556 29520
rect 2516 29306 2544 29514
rect 2976 29306 3004 30262
rect 3160 30054 3188 30534
rect 3148 30048 3200 30054
rect 3148 29990 3200 29996
rect 2504 29300 2556 29306
rect 2504 29242 2556 29248
rect 2964 29300 3016 29306
rect 2964 29242 3016 29248
rect 2228 27532 2280 27538
rect 2228 27474 2280 27480
rect 2688 27396 2740 27402
rect 2688 27338 2740 27344
rect 2700 27130 2728 27338
rect 2976 27334 3004 29242
rect 3240 29028 3292 29034
rect 3240 28970 3292 28976
rect 3252 28082 3280 28970
rect 3240 28076 3292 28082
rect 3240 28018 3292 28024
rect 3056 27464 3108 27470
rect 3056 27406 3108 27412
rect 2964 27328 3016 27334
rect 2964 27270 3016 27276
rect 2976 27130 3004 27270
rect 2688 27124 2740 27130
rect 2688 27066 2740 27072
rect 2964 27124 3016 27130
rect 2964 27066 3016 27072
rect 848 26784 900 26790
rect 846 26752 848 26761
rect 900 26752 902 26761
rect 846 26687 902 26696
rect 3068 23730 3096 27406
rect 3528 27402 3556 32710
rect 4080 32450 4108 32710
rect 4172 32502 4200 32966
rect 4632 32910 4660 33526
rect 4252 32904 4304 32910
rect 4252 32846 4304 32852
rect 4620 32904 4672 32910
rect 4620 32846 4672 32852
rect 4264 32570 4292 32846
rect 4344 32836 4396 32842
rect 4344 32778 4396 32784
rect 4252 32564 4304 32570
rect 4252 32506 4304 32512
rect 3988 32434 4108 32450
rect 4160 32496 4212 32502
rect 4160 32438 4212 32444
rect 4356 32434 4384 32778
rect 3976 32428 4108 32434
rect 4028 32422 4108 32428
rect 4344 32428 4396 32434
rect 3976 32370 4028 32376
rect 4344 32370 4396 32376
rect 4632 32366 4660 32846
rect 4620 32360 4672 32366
rect 4620 32302 4672 32308
rect 3608 32224 3660 32230
rect 3608 32166 3660 32172
rect 3700 32224 3752 32230
rect 3700 32166 3752 32172
rect 3620 32026 3648 32166
rect 3608 32020 3660 32026
rect 3608 31962 3660 31968
rect 3712 31958 3740 32166
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 3700 31952 3752 31958
rect 3700 31894 3752 31900
rect 3712 30802 3740 31894
rect 4344 31680 4396 31686
rect 4344 31622 4396 31628
rect 4356 31414 4384 31622
rect 4344 31408 4396 31414
rect 4344 31350 4396 31356
rect 4632 31362 4660 32302
rect 4724 32026 4752 33646
rect 4816 33504 4844 33798
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4896 33516 4948 33522
rect 4816 33476 4896 33504
rect 4896 33458 4948 33464
rect 4804 33312 4856 33318
rect 4804 33254 4856 33260
rect 4816 32978 4844 33254
rect 4804 32972 4856 32978
rect 4804 32914 4856 32920
rect 4816 32450 4844 32914
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 4816 32422 4936 32450
rect 4804 32292 4856 32298
rect 4804 32234 4856 32240
rect 4712 32020 4764 32026
rect 4712 31962 4764 31968
rect 4816 31906 4844 32234
rect 4724 31878 4844 31906
rect 4724 31482 4752 31878
rect 4908 31822 4936 32422
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 5000 31822 5028 32166
rect 5184 31958 5212 32506
rect 5264 32428 5316 32434
rect 5264 32370 5316 32376
rect 5172 31952 5224 31958
rect 5172 31894 5224 31900
rect 4896 31816 4948 31822
rect 4896 31758 4948 31764
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 4804 31748 4856 31754
rect 4804 31690 4856 31696
rect 4816 31482 4844 31690
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4712 31476 4764 31482
rect 4712 31418 4764 31424
rect 4804 31476 4856 31482
rect 4804 31418 4856 31424
rect 4632 31334 4752 31362
rect 4724 31278 4752 31334
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 4712 31272 4764 31278
rect 4712 31214 4764 31220
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3700 30796 3752 30802
rect 3700 30738 3752 30744
rect 3712 30326 3740 30738
rect 3884 30728 3936 30734
rect 3884 30670 3936 30676
rect 3896 30394 3924 30670
rect 3884 30388 3936 30394
rect 3884 30330 3936 30336
rect 3700 30320 3752 30326
rect 3700 30262 3752 30268
rect 3712 29714 3740 30262
rect 3700 29708 3752 29714
rect 3700 29650 3752 29656
rect 3608 29504 3660 29510
rect 3608 29446 3660 29452
rect 3620 29238 3648 29446
rect 3712 29306 3740 29650
rect 3896 29510 3924 30330
rect 4724 30326 4752 31214
rect 5184 30802 5212 31282
rect 5172 30796 5224 30802
rect 5172 30738 5224 30744
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4712 30320 4764 30326
rect 4712 30262 4764 30268
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4712 29708 4764 29714
rect 4712 29650 4764 29656
rect 3792 29504 3844 29510
rect 3792 29446 3844 29452
rect 3884 29504 3936 29510
rect 3884 29446 3936 29452
rect 3700 29300 3752 29306
rect 3700 29242 3752 29248
rect 3608 29232 3660 29238
rect 3608 29174 3660 29180
rect 3804 29034 3832 29446
rect 3792 29028 3844 29034
rect 3792 28970 3844 28976
rect 3896 28966 3924 29446
rect 4724 29306 4752 29650
rect 4712 29300 4764 29306
rect 4816 29288 4844 30534
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4816 29260 4936 29288
rect 4712 29242 4764 29248
rect 3884 28960 3936 28966
rect 3884 28902 3936 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4252 28688 4304 28694
rect 4252 28630 4304 28636
rect 3976 28620 4028 28626
rect 3976 28562 4028 28568
rect 3700 28416 3752 28422
rect 3700 28358 3752 28364
rect 3608 28212 3660 28218
rect 3608 28154 3660 28160
rect 3516 27396 3568 27402
rect 3516 27338 3568 27344
rect 3528 26042 3556 27338
rect 3620 27062 3648 28154
rect 3712 27946 3740 28358
rect 3988 28098 4016 28562
rect 4264 28558 4292 28630
rect 4724 28558 4752 29242
rect 4908 29170 4936 29260
rect 4804 29164 4856 29170
rect 4804 29106 4856 29112
rect 4896 29164 4948 29170
rect 4896 29106 4948 29112
rect 4816 28762 4844 29106
rect 4804 28756 4856 28762
rect 4804 28698 4856 28704
rect 4068 28552 4120 28558
rect 4068 28494 4120 28500
rect 4252 28552 4304 28558
rect 4252 28494 4304 28500
rect 4344 28552 4396 28558
rect 4344 28494 4396 28500
rect 4712 28552 4764 28558
rect 4712 28494 4764 28500
rect 4080 28218 4108 28494
rect 4068 28212 4120 28218
rect 4068 28154 4120 28160
rect 4264 28150 4292 28494
rect 3896 28082 4016 28098
rect 4252 28144 4304 28150
rect 4252 28086 4304 28092
rect 4356 28082 4384 28494
rect 4804 28416 4856 28422
rect 4804 28358 4856 28364
rect 3884 28076 4016 28082
rect 3936 28070 4016 28076
rect 3884 28018 3936 28024
rect 3792 28008 3844 28014
rect 3792 27950 3844 27956
rect 3700 27940 3752 27946
rect 3700 27882 3752 27888
rect 3608 27056 3660 27062
rect 3608 26998 3660 27004
rect 3712 26858 3740 27882
rect 3804 26994 3832 27950
rect 3988 27878 4016 28070
rect 4344 28076 4396 28082
rect 4344 28018 4396 28024
rect 4620 28008 4672 28014
rect 4620 27950 4672 27956
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3976 27872 4028 27878
rect 3976 27814 4028 27820
rect 3792 26988 3844 26994
rect 3792 26930 3844 26936
rect 3700 26852 3752 26858
rect 3700 26794 3752 26800
rect 3896 26790 3924 27814
rect 3988 27674 4016 27814
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 3976 27668 4028 27674
rect 3976 27610 4028 27616
rect 4068 27600 4120 27606
rect 4068 27542 4120 27548
rect 4080 27334 4108 27542
rect 4632 27470 4660 27950
rect 4712 27872 4764 27878
rect 4712 27814 4764 27820
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 27062 4108 27270
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4632 26994 4660 27406
rect 4620 26988 4672 26994
rect 4620 26930 4672 26936
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 3884 26784 3936 26790
rect 3884 26726 3936 26732
rect 4080 26466 4108 26862
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4080 26438 4200 26466
rect 3516 26036 3568 26042
rect 3516 25978 3568 25984
rect 4172 25786 4200 26438
rect 4632 26382 4660 26930
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 4724 26330 4752 27814
rect 4816 27334 4844 28358
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5276 28150 5304 32370
rect 5368 31890 5396 35430
rect 5736 35290 5764 35634
rect 5724 35284 5776 35290
rect 5724 35226 5776 35232
rect 5920 35222 5948 36110
rect 6000 35624 6052 35630
rect 6000 35566 6052 35572
rect 6012 35290 6040 35566
rect 6000 35284 6052 35290
rect 6000 35226 6052 35232
rect 5908 35216 5960 35222
rect 5908 35158 5960 35164
rect 6104 35086 6132 36722
rect 6932 36242 6960 37606
rect 7024 37262 7052 37878
rect 7576 37874 7604 38150
rect 7668 38010 7696 38150
rect 7656 38004 7708 38010
rect 7656 37946 7708 37952
rect 7654 37904 7710 37913
rect 7564 37868 7616 37874
rect 7760 37890 7788 38490
rect 8116 38344 8168 38350
rect 8116 38286 8168 38292
rect 7840 38208 7892 38214
rect 7840 38150 7892 38156
rect 7852 37942 7880 38150
rect 8128 38010 8156 38286
rect 8220 38282 8248 38898
rect 8300 38752 8352 38758
rect 8300 38694 8352 38700
rect 8208 38276 8260 38282
rect 8208 38218 8260 38224
rect 8116 38004 8168 38010
rect 8116 37946 8168 37952
rect 7710 37862 7788 37890
rect 7840 37936 7892 37942
rect 7840 37878 7892 37884
rect 7654 37839 7656 37848
rect 7564 37810 7616 37816
rect 7708 37839 7710 37848
rect 7656 37810 7708 37816
rect 7012 37256 7064 37262
rect 7012 37198 7064 37204
rect 7012 37120 7064 37126
rect 7012 37062 7064 37068
rect 7024 36378 7052 37062
rect 7288 36576 7340 36582
rect 7208 36524 7288 36530
rect 7208 36518 7340 36524
rect 7208 36502 7328 36518
rect 7012 36372 7064 36378
rect 7012 36314 7064 36320
rect 6920 36236 6972 36242
rect 6920 36178 6972 36184
rect 6736 35692 6788 35698
rect 6736 35634 6788 35640
rect 6092 35080 6144 35086
rect 6092 35022 6144 35028
rect 5540 35012 5592 35018
rect 5540 34954 5592 34960
rect 5448 33924 5500 33930
rect 5448 33866 5500 33872
rect 5460 32366 5488 33866
rect 5552 32910 5580 34954
rect 5908 34196 5960 34202
rect 5908 34138 5960 34144
rect 5920 33318 5948 34138
rect 6104 34066 6132 35022
rect 6748 35018 6776 35634
rect 6828 35216 6880 35222
rect 6828 35158 6880 35164
rect 6736 35012 6788 35018
rect 6736 34954 6788 34960
rect 6092 34060 6144 34066
rect 6092 34002 6144 34008
rect 6104 33590 6132 34002
rect 6092 33584 6144 33590
rect 6092 33526 6144 33532
rect 5908 33312 5960 33318
rect 5908 33254 5960 33260
rect 5540 32904 5592 32910
rect 5540 32846 5592 32852
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5448 31952 5500 31958
rect 5448 31894 5500 31900
rect 5356 31884 5408 31890
rect 5356 31826 5408 31832
rect 5356 31748 5408 31754
rect 5356 31690 5408 31696
rect 5368 30734 5396 31690
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 5356 30388 5408 30394
rect 5356 30330 5408 30336
rect 5368 29510 5396 30330
rect 5356 29504 5408 29510
rect 5356 29446 5408 29452
rect 5356 29164 5408 29170
rect 5356 29106 5408 29112
rect 5368 28694 5396 29106
rect 5460 29102 5488 31894
rect 5552 31754 5580 32846
rect 5816 32768 5868 32774
rect 5920 32722 5948 33254
rect 6104 32910 6132 33526
rect 6840 33522 6868 35158
rect 6932 33980 6960 36178
rect 7208 36174 7236 36502
rect 7196 36168 7248 36174
rect 7196 36110 7248 36116
rect 7104 36100 7156 36106
rect 7104 36042 7156 36048
rect 7012 33992 7064 33998
rect 6932 33952 7012 33980
rect 7012 33934 7064 33940
rect 6920 33856 6972 33862
rect 7116 33810 7144 36042
rect 7208 35698 7236 36110
rect 7472 36032 7524 36038
rect 7472 35974 7524 35980
rect 7484 35698 7512 35974
rect 7196 35692 7248 35698
rect 7196 35634 7248 35640
rect 7472 35692 7524 35698
rect 7472 35634 7524 35640
rect 7576 35086 7604 37810
rect 8220 36650 8248 38218
rect 8312 38214 8340 38694
rect 8680 38554 8708 39578
rect 10980 39438 11008 41200
rect 12912 39438 12940 41200
rect 10968 39432 11020 39438
rect 10968 39374 11020 39380
rect 12900 39432 12952 39438
rect 12900 39374 12952 39380
rect 10048 39296 10100 39302
rect 10048 39238 10100 39244
rect 10784 39296 10836 39302
rect 10784 39238 10836 39244
rect 11336 39296 11388 39302
rect 11336 39238 11388 39244
rect 12624 39296 12676 39302
rect 12624 39238 12676 39244
rect 10060 39098 10088 39238
rect 10048 39092 10100 39098
rect 10048 39034 10100 39040
rect 9772 38888 9824 38894
rect 9772 38830 9824 38836
rect 8668 38548 8720 38554
rect 8668 38490 8720 38496
rect 8484 38344 8536 38350
rect 8484 38286 8536 38292
rect 8300 38208 8352 38214
rect 8300 38150 8352 38156
rect 8312 37738 8340 38150
rect 8300 37732 8352 37738
rect 8300 37674 8352 37680
rect 7932 36644 7984 36650
rect 7932 36586 7984 36592
rect 8208 36644 8260 36650
rect 8208 36586 8260 36592
rect 7840 35556 7892 35562
rect 7840 35498 7892 35504
rect 7852 35086 7880 35498
rect 7564 35080 7616 35086
rect 7564 35022 7616 35028
rect 7840 35080 7892 35086
rect 7840 35022 7892 35028
rect 7472 34604 7524 34610
rect 7472 34546 7524 34552
rect 7288 34468 7340 34474
rect 7288 34410 7340 34416
rect 7196 34400 7248 34406
rect 7196 34342 7248 34348
rect 7208 33930 7236 34342
rect 7300 34202 7328 34410
rect 7288 34196 7340 34202
rect 7288 34138 7340 34144
rect 7380 34128 7432 34134
rect 7380 34070 7432 34076
rect 7392 33930 7420 34070
rect 7196 33924 7248 33930
rect 7196 33866 7248 33872
rect 7380 33924 7432 33930
rect 7380 33866 7432 33872
rect 6920 33798 6972 33804
rect 6828 33516 6880 33522
rect 6828 33458 6880 33464
rect 6840 33114 6868 33458
rect 6828 33108 6880 33114
rect 6828 33050 6880 33056
rect 6932 32910 6960 33798
rect 7024 33782 7144 33810
rect 6092 32904 6144 32910
rect 6092 32846 6144 32852
rect 6460 32904 6512 32910
rect 6460 32846 6512 32852
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 5868 32716 5948 32722
rect 5816 32710 5948 32716
rect 6276 32768 6328 32774
rect 6276 32710 6328 32716
rect 5828 32694 5948 32710
rect 5920 32434 5948 32694
rect 6288 32502 6316 32710
rect 6276 32496 6328 32502
rect 6276 32438 6328 32444
rect 5908 32428 5960 32434
rect 5908 32370 5960 32376
rect 5920 32026 5948 32370
rect 6000 32360 6052 32366
rect 6000 32302 6052 32308
rect 5908 32020 5960 32026
rect 5908 31962 5960 31968
rect 5920 31890 5948 31962
rect 5908 31884 5960 31890
rect 5908 31826 5960 31832
rect 6012 31822 6040 32302
rect 6184 31952 6236 31958
rect 6184 31894 6236 31900
rect 6000 31816 6052 31822
rect 6000 31758 6052 31764
rect 5552 31726 5672 31754
rect 5644 31278 5672 31726
rect 6196 31346 6224 31894
rect 6288 31822 6316 32438
rect 6276 31816 6328 31822
rect 6276 31758 6328 31764
rect 6184 31340 6236 31346
rect 6184 31282 6236 31288
rect 5632 31272 5684 31278
rect 5632 31214 5684 31220
rect 5540 31136 5592 31142
rect 5540 31078 5592 31084
rect 5552 30394 5580 31078
rect 5540 30388 5592 30394
rect 5540 30330 5592 30336
rect 5644 30122 5672 31214
rect 6288 30682 6316 31758
rect 6472 31346 6500 32846
rect 7024 32842 7052 33782
rect 7392 32910 7420 33866
rect 7484 33862 7512 34546
rect 7852 34202 7880 35022
rect 7840 34196 7892 34202
rect 7840 34138 7892 34144
rect 7852 33980 7880 34138
rect 7944 34134 7972 36586
rect 8208 36032 8260 36038
rect 8208 35974 8260 35980
rect 8024 35624 8076 35630
rect 8024 35566 8076 35572
rect 8036 35290 8064 35566
rect 8220 35494 8248 35974
rect 8116 35488 8168 35494
rect 8116 35430 8168 35436
rect 8208 35488 8260 35494
rect 8208 35430 8260 35436
rect 8024 35284 8076 35290
rect 8024 35226 8076 35232
rect 8128 35154 8156 35430
rect 8116 35148 8168 35154
rect 8116 35090 8168 35096
rect 7932 34128 7984 34134
rect 7932 34070 7984 34076
rect 8024 33992 8076 33998
rect 7852 33952 8024 33980
rect 8024 33934 8076 33940
rect 7472 33856 7524 33862
rect 7472 33798 7524 33804
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7484 32842 7512 33798
rect 7656 33380 7708 33386
rect 7656 33322 7708 33328
rect 7012 32836 7064 32842
rect 7012 32778 7064 32784
rect 7472 32836 7524 32842
rect 7472 32778 7524 32784
rect 7024 32026 7052 32778
rect 7668 32570 7696 33322
rect 8036 33114 8064 33934
rect 8128 33862 8156 35090
rect 8312 35018 8340 37674
rect 8392 35284 8444 35290
rect 8392 35226 8444 35232
rect 8300 35012 8352 35018
rect 8300 34954 8352 34960
rect 8404 34746 8432 35226
rect 8392 34740 8444 34746
rect 8392 34682 8444 34688
rect 8208 34604 8260 34610
rect 8208 34546 8260 34552
rect 8220 34202 8248 34546
rect 8208 34196 8260 34202
rect 8208 34138 8260 34144
rect 8116 33856 8168 33862
rect 8116 33798 8168 33804
rect 8496 33522 8524 38286
rect 8576 38208 8628 38214
rect 8576 38150 8628 38156
rect 8588 37806 8616 38150
rect 8576 37800 8628 37806
rect 8576 37742 8628 37748
rect 8680 37466 8708 38490
rect 9784 38350 9812 38830
rect 10796 38554 10824 39238
rect 11060 38752 11112 38758
rect 11060 38694 11112 38700
rect 10784 38548 10836 38554
rect 10784 38490 10836 38496
rect 11072 38350 11100 38694
rect 9772 38344 9824 38350
rect 9772 38286 9824 38292
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 11060 38344 11112 38350
rect 11060 38286 11112 38292
rect 10324 38208 10376 38214
rect 10324 38150 10376 38156
rect 10336 38010 10364 38150
rect 10612 38010 10640 38286
rect 8760 38004 8812 38010
rect 8760 37946 8812 37952
rect 9956 38004 10008 38010
rect 9956 37946 10008 37952
rect 10324 38004 10376 38010
rect 10324 37946 10376 37952
rect 10600 38004 10652 38010
rect 10600 37946 10652 37952
rect 8772 37913 8800 37946
rect 8758 37904 8814 37913
rect 8758 37839 8760 37848
rect 8812 37839 8814 37848
rect 8760 37810 8812 37816
rect 8668 37460 8720 37466
rect 8668 37402 8720 37408
rect 8576 36100 8628 36106
rect 8576 36042 8628 36048
rect 8588 35834 8616 36042
rect 8576 35828 8628 35834
rect 8576 35770 8628 35776
rect 8680 34474 8708 37402
rect 9968 37262 9996 37946
rect 11072 37874 11100 38286
rect 11060 37868 11112 37874
rect 11060 37810 11112 37816
rect 10876 37664 10928 37670
rect 10876 37606 10928 37612
rect 10888 37398 10916 37606
rect 10600 37392 10652 37398
rect 10600 37334 10652 37340
rect 10876 37392 10928 37398
rect 10876 37334 10928 37340
rect 9864 37256 9916 37262
rect 9864 37198 9916 37204
rect 9956 37256 10008 37262
rect 9956 37198 10008 37204
rect 9036 36848 9088 36854
rect 9036 36790 9088 36796
rect 9048 36038 9076 36790
rect 9876 36718 9904 37198
rect 9968 36922 9996 37198
rect 10048 37120 10100 37126
rect 10048 37062 10100 37068
rect 9956 36916 10008 36922
rect 9956 36858 10008 36864
rect 10060 36786 10088 37062
rect 10048 36780 10100 36786
rect 10048 36722 10100 36728
rect 10416 36780 10468 36786
rect 10416 36722 10468 36728
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 10060 36378 10088 36722
rect 10232 36712 10284 36718
rect 10232 36654 10284 36660
rect 10048 36372 10100 36378
rect 10048 36314 10100 36320
rect 9128 36168 9180 36174
rect 9128 36110 9180 36116
rect 9956 36168 10008 36174
rect 9956 36110 10008 36116
rect 9036 36032 9088 36038
rect 9036 35974 9088 35980
rect 8944 35624 8996 35630
rect 8944 35566 8996 35572
rect 8956 35290 8984 35566
rect 8944 35284 8996 35290
rect 8944 35226 8996 35232
rect 8668 34468 8720 34474
rect 8668 34410 8720 34416
rect 9048 34406 9076 35974
rect 9140 35834 9168 36110
rect 9968 35834 9996 36110
rect 10244 35834 10272 36654
rect 9128 35828 9180 35834
rect 9128 35770 9180 35776
rect 9956 35828 10008 35834
rect 9956 35770 10008 35776
rect 10232 35828 10284 35834
rect 10232 35770 10284 35776
rect 10324 35760 10376 35766
rect 10324 35702 10376 35708
rect 9496 35692 9548 35698
rect 9496 35634 9548 35640
rect 9956 35692 10008 35698
rect 9956 35634 10008 35640
rect 10232 35692 10284 35698
rect 10232 35634 10284 35640
rect 9312 35216 9364 35222
rect 9312 35158 9364 35164
rect 9220 34468 9272 34474
rect 9220 34410 9272 34416
rect 9036 34400 9088 34406
rect 9036 34342 9088 34348
rect 9048 33998 9076 34342
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 9232 33930 9260 34410
rect 9220 33924 9272 33930
rect 9220 33866 9272 33872
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 8484 33516 8536 33522
rect 8484 33458 8536 33464
rect 8668 33516 8720 33522
rect 8668 33458 8720 33464
rect 8024 33108 8076 33114
rect 8024 33050 8076 33056
rect 8312 33046 8340 33458
rect 8680 33114 8708 33458
rect 8760 33312 8812 33318
rect 8760 33254 8812 33260
rect 8668 33108 8720 33114
rect 8668 33050 8720 33056
rect 8300 33040 8352 33046
rect 8300 32982 8352 32988
rect 8772 32910 8800 33254
rect 8300 32904 8352 32910
rect 8760 32904 8812 32910
rect 8352 32852 8616 32858
rect 8300 32846 8616 32852
rect 8760 32846 8812 32852
rect 9036 32904 9088 32910
rect 9232 32858 9260 33866
rect 9324 33114 9352 35158
rect 9508 35086 9536 35634
rect 9680 35624 9732 35630
rect 9680 35566 9732 35572
rect 9772 35624 9824 35630
rect 9772 35566 9824 35572
rect 9692 35086 9720 35566
rect 9784 35290 9812 35566
rect 9864 35488 9916 35494
rect 9864 35430 9916 35436
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9876 35170 9904 35430
rect 9968 35290 9996 35634
rect 10244 35290 10272 35634
rect 9956 35284 10008 35290
rect 9956 35226 10008 35232
rect 10232 35284 10284 35290
rect 10232 35226 10284 35232
rect 9876 35154 9996 35170
rect 9876 35148 10008 35154
rect 9876 35142 9956 35148
rect 9496 35080 9548 35086
rect 9496 35022 9548 35028
rect 9680 35080 9732 35086
rect 9680 35022 9732 35028
rect 9508 33318 9536 35022
rect 9876 33998 9904 35142
rect 9956 35090 10008 35096
rect 10336 35018 10364 35702
rect 10428 35222 10456 36722
rect 10508 36576 10560 36582
rect 10508 36518 10560 36524
rect 10520 35698 10548 36518
rect 10612 36174 10640 37334
rect 10784 37256 10836 37262
rect 10888 37244 10916 37334
rect 11072 37262 11100 37810
rect 11244 37800 11296 37806
rect 11244 37742 11296 37748
rect 11152 37664 11204 37670
rect 11152 37606 11204 37612
rect 10836 37216 10916 37244
rect 10784 37198 10836 37204
rect 10784 36576 10836 36582
rect 10784 36518 10836 36524
rect 10796 36310 10824 36518
rect 10784 36304 10836 36310
rect 10784 36246 10836 36252
rect 10600 36168 10652 36174
rect 10598 36136 10600 36145
rect 10652 36136 10654 36145
rect 10598 36071 10654 36080
rect 10600 36032 10652 36038
rect 10600 35974 10652 35980
rect 10612 35698 10640 35974
rect 10508 35692 10560 35698
rect 10508 35634 10560 35640
rect 10600 35692 10652 35698
rect 10600 35634 10652 35640
rect 10796 35222 10824 36246
rect 10888 35562 10916 37216
rect 11060 37256 11112 37262
rect 11060 37198 11112 37204
rect 11164 36854 11192 37606
rect 11256 37262 11284 37742
rect 11244 37256 11296 37262
rect 11244 37198 11296 37204
rect 11256 37126 11284 37198
rect 11244 37120 11296 37126
rect 11244 37062 11296 37068
rect 11152 36848 11204 36854
rect 11152 36790 11204 36796
rect 11256 36786 11284 37062
rect 11244 36780 11296 36786
rect 11244 36722 11296 36728
rect 11348 36258 11376 39238
rect 12072 38752 12124 38758
rect 12072 38694 12124 38700
rect 11520 38344 11572 38350
rect 11520 38286 11572 38292
rect 11532 37466 11560 38286
rect 11888 38276 11940 38282
rect 11888 38218 11940 38224
rect 11704 37732 11756 37738
rect 11704 37674 11756 37680
rect 11716 37466 11744 37674
rect 11900 37670 11928 38218
rect 12084 37874 12112 38694
rect 12164 38548 12216 38554
rect 12216 38508 12296 38536
rect 12164 38490 12216 38496
rect 12164 38344 12216 38350
rect 12164 38286 12216 38292
rect 12072 37868 12124 37874
rect 12072 37810 12124 37816
rect 11888 37664 11940 37670
rect 11888 37606 11940 37612
rect 11520 37460 11572 37466
rect 11520 37402 11572 37408
rect 11704 37460 11756 37466
rect 11704 37402 11756 37408
rect 11716 37330 11744 37402
rect 11704 37324 11756 37330
rect 11704 37266 11756 37272
rect 11716 36718 11744 37266
rect 12084 37194 12112 37810
rect 12176 37738 12204 38286
rect 12268 38010 12296 38508
rect 12348 38208 12400 38214
rect 12348 38150 12400 38156
rect 12256 38004 12308 38010
rect 12256 37946 12308 37952
rect 12164 37732 12216 37738
rect 12164 37674 12216 37680
rect 12072 37188 12124 37194
rect 12072 37130 12124 37136
rect 11704 36712 11756 36718
rect 11704 36654 11756 36660
rect 12164 36644 12216 36650
rect 12164 36586 12216 36592
rect 12176 36378 12204 36586
rect 11428 36372 11480 36378
rect 11428 36314 11480 36320
rect 12164 36372 12216 36378
rect 12164 36314 12216 36320
rect 11256 36230 11376 36258
rect 11440 36242 11468 36314
rect 12072 36304 12124 36310
rect 12072 36246 12124 36252
rect 11428 36236 11480 36242
rect 11152 36168 11204 36174
rect 11150 36136 11152 36145
rect 11204 36136 11206 36145
rect 11150 36071 11206 36080
rect 11060 36032 11112 36038
rect 11060 35974 11112 35980
rect 11072 35766 11100 35974
rect 11060 35760 11112 35766
rect 11060 35702 11112 35708
rect 10968 35624 11020 35630
rect 11256 35612 11284 36230
rect 11428 36178 11480 36184
rect 11520 36168 11572 36174
rect 11520 36110 11572 36116
rect 11336 36100 11388 36106
rect 11336 36042 11388 36048
rect 11020 35584 11284 35612
rect 10968 35566 11020 35572
rect 10876 35556 10928 35562
rect 10876 35498 10928 35504
rect 10416 35216 10468 35222
rect 10416 35158 10468 35164
rect 10784 35216 10836 35222
rect 10784 35158 10836 35164
rect 10508 35080 10560 35086
rect 10888 35034 10916 35498
rect 10508 35022 10560 35028
rect 10232 35012 10284 35018
rect 10232 34954 10284 34960
rect 10324 35012 10376 35018
rect 10324 34954 10376 34960
rect 10416 35012 10468 35018
rect 10416 34954 10468 34960
rect 10048 34060 10100 34066
rect 10048 34002 10100 34008
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 9956 33992 10008 33998
rect 9956 33934 10008 33940
rect 9968 33658 9996 33934
rect 9956 33652 10008 33658
rect 9956 33594 10008 33600
rect 9956 33516 10008 33522
rect 9956 33458 10008 33464
rect 9496 33312 9548 33318
rect 9496 33254 9548 33260
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9864 33108 9916 33114
rect 9864 33050 9916 33056
rect 9404 33040 9456 33046
rect 9404 32982 9456 32988
rect 9088 32852 9260 32858
rect 9036 32846 9260 32852
rect 8312 32842 8616 32846
rect 8312 32836 8628 32842
rect 8312 32830 8576 32836
rect 9048 32830 9260 32846
rect 8576 32778 8628 32784
rect 9232 32774 9260 32830
rect 9128 32768 9180 32774
rect 9128 32710 9180 32716
rect 9220 32768 9272 32774
rect 9220 32710 9272 32716
rect 7656 32564 7708 32570
rect 7656 32506 7708 32512
rect 7012 32020 7064 32026
rect 7012 31962 7064 31968
rect 7012 31884 7064 31890
rect 7012 31826 7064 31832
rect 6920 31816 6972 31822
rect 6920 31758 6972 31764
rect 6828 31748 6880 31754
rect 6828 31690 6880 31696
rect 6552 31680 6604 31686
rect 6552 31622 6604 31628
rect 6368 31340 6420 31346
rect 6368 31282 6420 31288
rect 6460 31340 6512 31346
rect 6460 31282 6512 31288
rect 6196 30654 6316 30682
rect 5632 30116 5684 30122
rect 5632 30058 5684 30064
rect 5816 29708 5868 29714
rect 5816 29650 5868 29656
rect 5540 29504 5592 29510
rect 5540 29446 5592 29452
rect 5552 29238 5580 29446
rect 5540 29232 5592 29238
rect 5540 29174 5592 29180
rect 5448 29096 5500 29102
rect 5448 29038 5500 29044
rect 5828 28762 5856 29650
rect 6196 29646 6224 30654
rect 6380 30326 6408 31282
rect 6564 30802 6592 31622
rect 6840 31414 6868 31690
rect 6932 31414 6960 31758
rect 7024 31482 7052 31826
rect 8484 31816 8536 31822
rect 8484 31758 8536 31764
rect 7932 31680 7984 31686
rect 7932 31622 7984 31628
rect 8116 31680 8168 31686
rect 8116 31622 8168 31628
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 6828 31408 6880 31414
rect 6828 31350 6880 31356
rect 6920 31408 6972 31414
rect 6920 31350 6972 31356
rect 6736 31340 6788 31346
rect 6736 31282 6788 31288
rect 6748 30938 6776 31282
rect 6736 30932 6788 30938
rect 6736 30874 6788 30880
rect 6552 30796 6604 30802
rect 6552 30738 6604 30744
rect 6368 30320 6420 30326
rect 6368 30262 6420 30268
rect 6276 30116 6328 30122
rect 6276 30058 6328 30064
rect 6288 29646 6316 30058
rect 6380 29646 6408 30262
rect 6840 29646 6868 31350
rect 7944 30598 7972 31622
rect 8024 30728 8076 30734
rect 8128 30716 8156 31622
rect 8496 31482 8524 31758
rect 9140 31754 9168 32710
rect 9312 31816 9364 31822
rect 9312 31758 9364 31764
rect 9140 31726 9260 31754
rect 9128 31680 9180 31686
rect 9128 31622 9180 31628
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8220 30938 8248 31282
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 8076 30688 8156 30716
rect 8024 30670 8076 30676
rect 8392 30660 8444 30666
rect 8392 30602 8444 30608
rect 7012 30592 7064 30598
rect 7012 30534 7064 30540
rect 7932 30592 7984 30598
rect 7932 30534 7984 30540
rect 7024 29866 7052 30534
rect 8300 30252 8352 30258
rect 8300 30194 8352 30200
rect 6932 29838 7052 29866
rect 6184 29640 6236 29646
rect 6184 29582 6236 29588
rect 6276 29640 6328 29646
rect 6276 29582 6328 29588
rect 6368 29640 6420 29646
rect 6368 29582 6420 29588
rect 6828 29640 6880 29646
rect 6828 29582 6880 29588
rect 6380 29306 6408 29582
rect 6368 29300 6420 29306
rect 6368 29242 6420 29248
rect 6736 29028 6788 29034
rect 6736 28970 6788 28976
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5356 28688 5408 28694
rect 5356 28630 5408 28636
rect 6276 28416 6328 28422
rect 6276 28358 6328 28364
rect 6288 28150 6316 28358
rect 5264 28144 5316 28150
rect 6276 28144 6328 28150
rect 5316 28092 5580 28098
rect 5264 28086 5580 28092
rect 6276 28086 6328 28092
rect 5276 28070 5580 28086
rect 6748 28082 6776 28970
rect 6932 28626 6960 29838
rect 7012 29708 7064 29714
rect 7012 29650 7064 29656
rect 7024 28626 7052 29650
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7196 29164 7248 29170
rect 7196 29106 7248 29112
rect 7208 28762 7236 29106
rect 7196 28756 7248 28762
rect 7196 28698 7248 28704
rect 6920 28620 6972 28626
rect 6920 28562 6972 28568
rect 7012 28620 7064 28626
rect 7012 28562 7064 28568
rect 7392 28082 7420 29582
rect 8312 29170 8340 30194
rect 8300 29164 8352 29170
rect 8300 29106 8352 29112
rect 7748 29096 7800 29102
rect 7748 29038 7800 29044
rect 7760 28150 7788 29038
rect 7840 28688 7892 28694
rect 7840 28630 7892 28636
rect 7748 28144 7800 28150
rect 7748 28086 7800 28092
rect 4804 27328 4856 27334
rect 4804 27270 4856 27276
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 5552 27062 5580 28070
rect 6368 28076 6420 28082
rect 6368 28018 6420 28024
rect 6736 28076 6788 28082
rect 6736 28018 6788 28024
rect 7380 28076 7432 28082
rect 7380 28018 7432 28024
rect 5724 28008 5776 28014
rect 5724 27950 5776 27956
rect 5736 27674 5764 27950
rect 6276 27872 6328 27878
rect 6276 27814 6328 27820
rect 5724 27668 5776 27674
rect 5724 27610 5776 27616
rect 6288 27470 6316 27814
rect 6380 27538 6408 28018
rect 6920 27872 6972 27878
rect 6920 27814 6972 27820
rect 7564 27872 7616 27878
rect 7564 27814 7616 27820
rect 6368 27532 6420 27538
rect 6368 27474 6420 27480
rect 5816 27464 5868 27470
rect 5816 27406 5868 27412
rect 6276 27464 6328 27470
rect 6276 27406 6328 27412
rect 5540 27056 5592 27062
rect 5540 26998 5592 27004
rect 5828 26926 5856 27406
rect 5816 26920 5868 26926
rect 5816 26862 5868 26868
rect 5264 26512 5316 26518
rect 5264 26454 5316 26460
rect 4804 26376 4856 26382
rect 4724 26324 4804 26330
rect 4724 26318 4856 26324
rect 4724 26302 4844 26318
rect 4252 26240 4304 26246
rect 4252 26182 4304 26188
rect 4080 25758 4200 25786
rect 4080 25412 4108 25758
rect 4264 25702 4292 26182
rect 4724 26042 4752 26302
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4620 25832 4672 25838
rect 4620 25774 4672 25780
rect 4252 25696 4304 25702
rect 4252 25638 4304 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4080 25384 4200 25412
rect 4172 25226 4200 25384
rect 4160 25220 4212 25226
rect 4160 25162 4212 25168
rect 3792 25152 3844 25158
rect 3792 25094 3844 25100
rect 3804 24274 3832 25094
rect 4172 24954 4200 25162
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 3792 24268 3844 24274
rect 3792 24210 3844 24216
rect 4632 23866 4660 25774
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4620 23860 4672 23866
rect 4620 23802 4672 23808
rect 3056 23724 3108 23730
rect 3056 23666 3108 23672
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 3068 23186 3096 23666
rect 3160 23322 3188 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4724 23322 4752 25638
rect 5276 25362 5304 26454
rect 5828 26382 5856 26862
rect 6932 26382 6960 27814
rect 7472 27396 7524 27402
rect 7472 27338 7524 27344
rect 7484 27130 7512 27338
rect 7472 27124 7524 27130
rect 7472 27066 7524 27072
rect 7576 26994 7604 27814
rect 7852 27130 7880 28630
rect 8208 28552 8260 28558
rect 8208 28494 8260 28500
rect 7932 28484 7984 28490
rect 7932 28426 7984 28432
rect 7944 27878 7972 28426
rect 7932 27872 7984 27878
rect 7932 27814 7984 27820
rect 7944 27130 7972 27814
rect 8220 27334 8248 28494
rect 8404 28490 8432 30602
rect 8496 30394 8524 31418
rect 9140 31346 9168 31622
rect 9128 31340 9180 31346
rect 9128 31282 9180 31288
rect 8944 31204 8996 31210
rect 8944 31146 8996 31152
rect 8956 30870 8984 31146
rect 8944 30864 8996 30870
rect 8944 30806 8996 30812
rect 8484 30388 8536 30394
rect 8536 30348 8616 30376
rect 8484 30330 8536 30336
rect 8484 30048 8536 30054
rect 8484 29990 8536 29996
rect 8496 29850 8524 29990
rect 8484 29844 8536 29850
rect 8484 29786 8536 29792
rect 8588 29646 8616 30348
rect 9140 30258 9168 31282
rect 9128 30252 9180 30258
rect 9128 30194 9180 30200
rect 8760 30048 8812 30054
rect 8760 29990 8812 29996
rect 8772 29714 8800 29990
rect 8760 29708 8812 29714
rect 8760 29650 8812 29656
rect 8576 29640 8628 29646
rect 8576 29582 8628 29588
rect 8668 29572 8720 29578
rect 8668 29514 8720 29520
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 8496 28150 8524 29106
rect 8680 28218 8708 29514
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 8484 28144 8536 28150
rect 8484 28086 8536 28092
rect 8300 28076 8352 28082
rect 8300 28018 8352 28024
rect 8312 27606 8340 28018
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 8300 27600 8352 27606
rect 8300 27542 8352 27548
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7932 27124 7984 27130
rect 7932 27066 7984 27072
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 7852 26586 7880 27066
rect 8220 26926 8248 27270
rect 8404 27130 8432 27882
rect 8496 27674 8524 28086
rect 8484 27668 8536 27674
rect 8484 27610 8536 27616
rect 8496 27130 8524 27610
rect 8680 27538 8708 28154
rect 9128 27872 9180 27878
rect 9128 27814 9180 27820
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 8668 27532 8720 27538
rect 8668 27474 8720 27480
rect 8576 27396 8628 27402
rect 8576 27338 8628 27344
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8484 27124 8536 27130
rect 8484 27066 8536 27072
rect 8588 27010 8616 27338
rect 8496 26994 8616 27010
rect 8680 26994 8708 27474
rect 8956 26994 8984 27542
rect 9140 27470 9168 27814
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9036 27396 9088 27402
rect 9036 27338 9088 27344
rect 9048 27130 9076 27338
rect 9036 27124 9088 27130
rect 9036 27066 9088 27072
rect 9140 27010 9168 27406
rect 8484 26988 8616 26994
rect 8536 26982 8616 26988
rect 8668 26988 8720 26994
rect 8484 26930 8536 26936
rect 8668 26930 8720 26936
rect 8944 26988 8996 26994
rect 8944 26930 8996 26936
rect 9048 26982 9168 27010
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 7012 26580 7064 26586
rect 7012 26522 7064 26528
rect 7840 26580 7892 26586
rect 7840 26522 7892 26528
rect 5816 26376 5868 26382
rect 5816 26318 5868 26324
rect 6920 26376 6972 26382
rect 6920 26318 6972 26324
rect 5356 26308 5408 26314
rect 5356 26250 5408 26256
rect 5368 25702 5396 26250
rect 5632 25832 5684 25838
rect 5632 25774 5684 25780
rect 5356 25696 5408 25702
rect 5356 25638 5408 25644
rect 5264 25356 5316 25362
rect 5264 25298 5316 25304
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 5644 24954 5672 25774
rect 5828 25294 5856 26318
rect 6368 26308 6420 26314
rect 6368 26250 6420 26256
rect 6380 25770 6408 26250
rect 7024 25906 7052 26522
rect 8220 26450 8248 26862
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8208 26444 8260 26450
rect 8208 26386 8260 26392
rect 7932 26240 7984 26246
rect 7932 26182 7984 26188
rect 7944 25906 7972 26182
rect 8220 25974 8248 26386
rect 8208 25968 8260 25974
rect 8208 25910 8260 25916
rect 7012 25900 7064 25906
rect 7012 25842 7064 25848
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7932 25900 7984 25906
rect 7932 25842 7984 25848
rect 6368 25764 6420 25770
rect 6368 25706 6420 25712
rect 6000 25696 6052 25702
rect 6000 25638 6052 25644
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 7564 25696 7616 25702
rect 7564 25638 7616 25644
rect 6012 25294 6040 25638
rect 6920 25424 6972 25430
rect 6920 25366 6972 25372
rect 5816 25288 5868 25294
rect 5816 25230 5868 25236
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 6552 25288 6604 25294
rect 6604 25236 6684 25242
rect 6552 25230 6684 25236
rect 5632 24948 5684 24954
rect 5632 24890 5684 24896
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5460 24410 5488 24754
rect 5828 24682 5856 25230
rect 6564 25214 6684 25230
rect 6552 25152 6604 25158
rect 6552 25094 6604 25100
rect 5908 24744 5960 24750
rect 5908 24686 5960 24692
rect 6460 24744 6512 24750
rect 6460 24686 6512 24692
rect 5816 24676 5868 24682
rect 5816 24618 5868 24624
rect 5920 24426 5948 24686
rect 6368 24608 6420 24614
rect 6368 24550 6420 24556
rect 5448 24404 5500 24410
rect 5448 24346 5500 24352
rect 5828 24398 5948 24426
rect 5828 24274 5856 24398
rect 5908 24336 5960 24342
rect 6380 24290 6408 24550
rect 6472 24410 6500 24686
rect 6460 24404 6512 24410
rect 6460 24346 6512 24352
rect 5908 24278 5960 24284
rect 5816 24268 5868 24274
rect 5816 24210 5868 24216
rect 4804 24064 4856 24070
rect 4804 24006 4856 24012
rect 3148 23316 3200 23322
rect 3148 23258 3200 23264
rect 3332 23316 3384 23322
rect 3332 23258 3384 23264
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 3056 23180 3108 23186
rect 3056 23122 3108 23128
rect 2044 22976 2096 22982
rect 2044 22918 2096 22924
rect 846 22672 902 22681
rect 846 22607 848 22616
rect 900 22607 902 22616
rect 848 22578 900 22584
rect 1768 22500 1820 22506
rect 1768 22442 1820 22448
rect 848 22024 900 22030
rect 846 21992 848 22001
rect 900 21992 902 22001
rect 112 21956 164 21962
rect 846 21927 902 21936
rect 112 21898 164 21904
rect 1780 21554 1808 22442
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1306 21176 1362 21185
rect 1306 21111 1362 21120
rect 1320 20330 1348 21111
rect 1780 20874 1808 21490
rect 1492 20868 1544 20874
rect 1492 20810 1544 20816
rect 1768 20868 1820 20874
rect 1768 20810 1820 20816
rect 1504 20602 1532 20810
rect 1492 20596 1544 20602
rect 1492 20538 1544 20544
rect 1780 20534 1808 20810
rect 1872 20534 1900 21966
rect 2056 21554 2084 22918
rect 3068 22030 3096 23122
rect 3344 23118 3372 23258
rect 3332 23112 3384 23118
rect 3332 23054 3384 23060
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3240 23044 3292 23050
rect 3240 22986 3292 22992
rect 3252 22710 3280 22986
rect 3332 22976 3384 22982
rect 3332 22918 3384 22924
rect 3240 22704 3292 22710
rect 3240 22646 3292 22652
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 1952 21480 2004 21486
rect 1952 21422 2004 21428
rect 1768 20528 1820 20534
rect 1768 20470 1820 20476
rect 1860 20528 1912 20534
rect 1860 20470 1912 20476
rect 1964 20398 1992 21422
rect 1952 20392 2004 20398
rect 1952 20334 2004 20340
rect 1308 20324 1360 20330
rect 1308 20266 1360 20272
rect 846 19952 902 19961
rect 846 19887 902 19896
rect 860 19854 888 19887
rect 2056 19854 2084 21490
rect 2136 21344 2188 21350
rect 2136 21286 2188 21292
rect 2148 20466 2176 21286
rect 2332 20534 2360 21830
rect 2792 21672 2820 21966
rect 3068 21690 3096 21966
rect 2700 21644 2820 21672
rect 2872 21684 2924 21690
rect 2700 21146 2728 21644
rect 2872 21626 2924 21632
rect 3056 21684 3108 21690
rect 3056 21626 3108 21632
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2688 21140 2740 21146
rect 2688 21082 2740 21088
rect 2320 20528 2372 20534
rect 2320 20470 2372 20476
rect 2700 20466 2728 21082
rect 2792 20942 2820 21490
rect 2780 20936 2832 20942
rect 2780 20878 2832 20884
rect 2884 20534 2912 21626
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3068 21146 3096 21490
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 3148 21004 3200 21010
rect 3148 20946 3200 20952
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2872 20528 2924 20534
rect 2872 20470 2924 20476
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2976 20058 3004 20878
rect 3160 20602 3188 20946
rect 3344 20942 3372 22918
rect 3436 22642 3464 23054
rect 3700 23044 3752 23050
rect 3700 22986 3752 22992
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 3712 22506 3740 22986
rect 4620 22976 4672 22982
rect 4620 22918 4672 22924
rect 3884 22704 3936 22710
rect 3884 22646 3936 22652
rect 3896 22574 3924 22646
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 3700 22500 3752 22506
rect 3700 22442 3752 22448
rect 3792 21956 3844 21962
rect 3792 21898 3844 21904
rect 3700 21072 3752 21078
rect 3700 21014 3752 21020
rect 3332 20936 3384 20942
rect 3332 20878 3384 20884
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3620 20618 3648 20878
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 3252 20590 3648 20618
rect 3054 20496 3110 20505
rect 3054 20431 3056 20440
rect 3108 20431 3110 20440
rect 3056 20402 3108 20408
rect 3148 20392 3200 20398
rect 3148 20334 3200 20340
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2964 20052 3016 20058
rect 2964 19994 3016 20000
rect 848 19848 900 19854
rect 848 19790 900 19796
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 2320 19848 2372 19854
rect 2320 19790 2372 19796
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 17746 1440 19314
rect 2148 18970 2176 19654
rect 2332 18970 2360 19790
rect 2792 19258 2820 19994
rect 3160 19922 3188 20334
rect 3252 19990 3280 20590
rect 3516 20528 3568 20534
rect 3516 20470 3568 20476
rect 3332 20324 3384 20330
rect 3332 20266 3384 20272
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3148 19780 3200 19786
rect 3148 19722 3200 19728
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2884 19378 2912 19654
rect 3160 19514 3188 19722
rect 3252 19514 3280 19926
rect 3148 19508 3200 19514
rect 3148 19450 3200 19456
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 2872 19372 2924 19378
rect 3344 19334 3372 20266
rect 2872 19314 2924 19320
rect 2700 19230 2820 19258
rect 3252 19306 3372 19334
rect 3528 19310 3556 20470
rect 3620 20398 3648 20590
rect 3712 20466 3740 21014
rect 3804 20874 3832 21898
rect 3896 21554 3924 22510
rect 4632 22506 4660 22918
rect 4816 22642 4844 24006
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5264 22976 5316 22982
rect 5264 22918 5316 22924
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 5276 22710 5304 22918
rect 5264 22704 5316 22710
rect 5264 22646 5316 22652
rect 4804 22636 4856 22642
rect 4804 22578 4856 22584
rect 4620 22500 4672 22506
rect 4620 22442 4672 22448
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4632 21554 4660 22442
rect 4816 22438 4844 22578
rect 5816 22568 5868 22574
rect 5816 22510 5868 22516
rect 5920 22522 5948 24278
rect 6104 24262 6408 24290
rect 6000 24200 6052 24206
rect 6104 24188 6132 24262
rect 6380 24206 6408 24262
rect 6052 24160 6132 24188
rect 6000 24142 6052 24148
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 6012 22642 6040 22918
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 4804 22432 4856 22438
rect 4804 22374 4856 22380
rect 5632 22432 5684 22438
rect 5632 22374 5684 22380
rect 4712 22024 4764 22030
rect 4712 21966 4764 21972
rect 4724 21554 4752 21966
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5644 21622 5672 22374
rect 5828 21978 5856 22510
rect 5920 22494 6040 22522
rect 5908 22432 5960 22438
rect 5908 22374 5960 22380
rect 5736 21950 5856 21978
rect 5632 21616 5684 21622
rect 5632 21558 5684 21564
rect 5736 21554 5764 21950
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 3884 21548 3936 21554
rect 3884 21490 3936 21496
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 3896 21146 3924 21490
rect 3976 21344 4028 21350
rect 3976 21286 4028 21292
rect 4068 21344 4120 21350
rect 4068 21286 4120 21292
rect 3988 21146 4016 21286
rect 3884 21140 3936 21146
rect 3884 21082 3936 21088
rect 3976 21140 4028 21146
rect 3976 21082 4028 21088
rect 4080 21078 4108 21286
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4068 21072 4120 21078
rect 4068 21014 4120 21020
rect 4632 20942 4660 21490
rect 5736 21146 5764 21490
rect 5724 21140 5776 21146
rect 5724 21082 5776 21088
rect 5828 21010 5856 21830
rect 5816 21004 5868 21010
rect 5816 20946 5868 20952
rect 5920 20942 5948 22374
rect 4620 20936 4672 20942
rect 4620 20878 4672 20884
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 3792 20868 3844 20874
rect 3792 20810 3844 20816
rect 4712 20868 4764 20874
rect 4712 20810 4764 20816
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3792 20460 3844 20466
rect 3792 20402 3844 20408
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 3608 20256 3660 20262
rect 3608 20198 3660 20204
rect 3700 20256 3752 20262
rect 3700 20198 3752 20204
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2320 18964 2372 18970
rect 2320 18906 2372 18912
rect 2148 18358 2176 18906
rect 2136 18352 2188 18358
rect 2136 18294 2188 18300
rect 2700 18222 2728 19230
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2872 19168 2924 19174
rect 2872 19110 2924 19116
rect 2792 18766 2820 19110
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2228 18216 2280 18222
rect 2228 18158 2280 18164
rect 2688 18216 2740 18222
rect 2688 18158 2740 18164
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1400 17740 1452 17746
rect 1400 17682 1452 17688
rect 1688 17610 1716 18022
rect 2240 17762 2268 18158
rect 2792 18086 2820 18702
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2148 17734 2268 17762
rect 1676 17604 1728 17610
rect 1676 17546 1728 17552
rect 2148 17338 2176 17734
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2228 17604 2280 17610
rect 2228 17546 2280 17552
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2240 17202 2268 17546
rect 2792 17270 2820 17614
rect 2884 17542 2912 19110
rect 2964 18692 3016 18698
rect 2964 18634 3016 18640
rect 2976 18290 3004 18634
rect 3056 18420 3108 18426
rect 3056 18362 3108 18368
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2964 18148 3016 18154
rect 2964 18090 3016 18096
rect 2976 17882 3004 18090
rect 2964 17876 3016 17882
rect 2964 17818 3016 17824
rect 3068 17762 3096 18362
rect 3068 17746 3188 17762
rect 3056 17740 3188 17746
rect 3108 17734 3188 17740
rect 3056 17682 3108 17688
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 2872 17536 2924 17542
rect 2924 17496 3004 17524
rect 2872 17478 2924 17484
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2504 16448 2556 16454
rect 2504 16390 2556 16396
rect 2516 15502 2544 16390
rect 2504 15496 2556 15502
rect 2556 15456 2636 15484
rect 2504 15438 2556 15444
rect 2608 15366 2636 15456
rect 2688 15428 2740 15434
rect 2688 15370 2740 15376
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1872 14618 1900 14962
rect 1860 14612 1912 14618
rect 1860 14554 1912 14560
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 2056 13870 2084 14418
rect 2148 14414 2176 15302
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2608 14346 2636 15302
rect 2700 14482 2728 15370
rect 2792 15094 2820 17206
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16794 2912 17138
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 2884 16266 2912 16458
rect 2976 16454 3004 17496
rect 3068 16998 3096 17546
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 2964 16448 3016 16454
rect 2964 16390 3016 16396
rect 3068 16266 3096 16934
rect 3160 16726 3188 17734
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 2884 16238 3096 16266
rect 2884 15638 2912 16238
rect 2964 15700 3016 15706
rect 2964 15642 3016 15648
rect 2872 15632 2924 15638
rect 2872 15574 2924 15580
rect 2976 15502 3004 15642
rect 3160 15570 3188 16526
rect 3148 15564 3200 15570
rect 3148 15506 3200 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2976 15162 3004 15438
rect 3148 15428 3200 15434
rect 3148 15370 3200 15376
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2596 14340 2648 14346
rect 2596 14282 2648 14288
rect 2792 14006 2820 15030
rect 2976 14618 3004 15098
rect 3160 15026 3188 15370
rect 3148 15020 3200 15026
rect 3148 14962 3200 14968
rect 3160 14618 3188 14962
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3148 14612 3200 14618
rect 3148 14554 3200 14560
rect 2976 14414 3004 14554
rect 2964 14408 3016 14414
rect 2964 14350 3016 14356
rect 2872 14272 2924 14278
rect 2872 14214 2924 14220
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2596 13796 2648 13802
rect 2596 13738 2648 13744
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 2228 13728 2280 13734
rect 2228 13670 2280 13676
rect 1504 13258 1532 13670
rect 1492 13252 1544 13258
rect 1492 13194 1544 13200
rect 1306 13016 1362 13025
rect 1306 12951 1308 12960
rect 1360 12951 1362 12960
rect 1308 12922 1360 12928
rect 2240 12850 2268 13670
rect 2608 13530 2636 13738
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2332 12646 2360 13466
rect 2700 13462 2728 13874
rect 2688 13456 2740 13462
rect 2688 13398 2740 13404
rect 2700 12730 2728 13398
rect 2792 13326 2820 13942
rect 2884 13870 2912 14214
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2976 13938 3004 14010
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2792 12918 2820 13262
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2608 12702 2728 12730
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 1676 12232 1728 12238
rect 846 12200 902 12209
rect 1676 12174 1728 12180
rect 846 12135 902 12144
rect 860 12102 888 12135
rect 848 12096 900 12102
rect 848 12038 900 12044
rect 1122 11656 1178 11665
rect 1688 11626 1716 12174
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1122 11591 1178 11600
rect 1676 11620 1728 11626
rect 1136 11354 1164 11591
rect 1676 11562 1728 11568
rect 1124 11348 1176 11354
rect 1124 11290 1176 11296
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1306 10296 1362 10305
rect 1306 10231 1362 10240
rect 1030 9616 1086 9625
rect 1030 9551 1086 9560
rect 1044 9450 1072 9551
rect 1032 9444 1084 9450
rect 1032 9386 1084 9392
rect 1320 9382 1348 10231
rect 1780 10130 1808 11086
rect 1872 10985 1900 12038
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1858 10976 1914 10985
rect 1858 10911 1914 10920
rect 2056 10810 2084 11018
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2148 10674 2176 11494
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 2240 10674 2268 11018
rect 2320 11008 2372 11014
rect 2320 10950 2372 10956
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 1768 10124 1820 10130
rect 1768 10066 1820 10072
rect 1400 9988 1452 9994
rect 1400 9930 1452 9936
rect 1308 9376 1360 9382
rect 1308 9318 1360 9324
rect 848 9104 900 9110
rect 846 9072 848 9081
rect 900 9072 902 9081
rect 846 9007 902 9016
rect 1412 8566 1440 9930
rect 1676 9920 1728 9926
rect 1676 9862 1728 9868
rect 1688 9586 1716 9862
rect 1676 9580 1728 9586
rect 1676 9522 1728 9528
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1688 8974 1716 9318
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 1780 8430 1808 10066
rect 2332 8974 2360 10950
rect 2608 10826 2636 12702
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 11014 2728 12582
rect 2792 11762 2820 12854
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2884 11286 2912 11766
rect 2976 11694 3004 12174
rect 3056 12096 3108 12102
rect 3056 12038 3108 12044
rect 2964 11688 3016 11694
rect 2964 11630 3016 11636
rect 2976 11354 3004 11630
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2884 11150 2912 11222
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 3068 11082 3096 12038
rect 3252 11694 3280 19306
rect 3516 19304 3568 19310
rect 3516 19246 3568 19252
rect 3528 18698 3556 19246
rect 3516 18692 3568 18698
rect 3516 18634 3568 18640
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3344 17338 3372 17818
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3344 17066 3372 17274
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3344 15706 3372 17002
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 15008 3464 18090
rect 3528 17678 3556 18158
rect 3620 17882 3648 20198
rect 3712 19854 3740 20198
rect 3804 19922 3832 20402
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3700 19304 3752 19310
rect 3700 19246 3752 19252
rect 3712 18426 3740 19246
rect 3804 18834 3832 19858
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 3700 18420 3752 18426
rect 3700 18362 3752 18368
rect 3804 18290 3832 18770
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 3976 18284 4028 18290
rect 3976 18226 4028 18232
rect 3608 17876 3660 17882
rect 3608 17818 3660 17824
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3700 17332 3752 17338
rect 3700 17274 3752 17280
rect 3712 16998 3740 17274
rect 3804 17134 3832 18226
rect 3988 17882 4016 18226
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3700 16992 3752 16998
rect 3700 16934 3752 16940
rect 3804 16658 3832 17070
rect 3896 16794 3924 17206
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 3516 16652 3568 16658
rect 3516 16594 3568 16600
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3344 14980 3464 15008
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2424 10798 2728 10826
rect 2424 10674 2452 10798
rect 2596 10736 2648 10742
rect 2594 10704 2596 10713
rect 2648 10704 2650 10713
rect 2412 10668 2464 10674
rect 2594 10639 2650 10648
rect 2412 10610 2464 10616
rect 2412 10464 2464 10470
rect 2412 10406 2464 10412
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2424 9994 2452 10406
rect 2412 9988 2464 9994
rect 2412 9930 2464 9936
rect 2516 9874 2544 10406
rect 2424 9846 2544 9874
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2320 8968 2372 8974
rect 2320 8910 2372 8916
rect 2056 8634 2084 8910
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1768 8424 1820 8430
rect 1768 8366 1820 8372
rect 1780 8090 1808 8366
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7546 1716 7754
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1780 6866 1808 8026
rect 1952 7404 2004 7410
rect 1872 7364 1952 7392
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1768 5704 1820 5710
rect 1688 5652 1768 5658
rect 1688 5646 1820 5652
rect 1688 5630 1808 5646
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1492 5024 1544 5030
rect 1492 4966 1544 4972
rect 1504 4554 1532 4966
rect 1492 4548 1544 4554
rect 1492 4490 1544 4496
rect 1400 3936 1452 3942
rect 1400 3878 1452 3884
rect 20 1352 72 1358
rect 1412 1306 1440 3878
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1504 2378 1532 3334
rect 1492 2372 1544 2378
rect 1492 2314 1544 2320
rect 1596 1358 1624 5510
rect 1688 3126 1716 5630
rect 1872 5234 1900 7364
rect 1952 7346 2004 7352
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1964 5234 1992 5510
rect 1860 5228 1912 5234
rect 1860 5170 1912 5176
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1872 3534 1900 5170
rect 2056 5166 2084 6802
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2240 5710 2268 5782
rect 2332 5710 2360 8910
rect 2424 7313 2452 9846
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2516 8090 2544 9522
rect 2608 9042 2636 10639
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2596 8832 2648 8838
rect 2596 8774 2648 8780
rect 2608 8566 2636 8774
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2516 7478 2544 8026
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2596 7404 2648 7410
rect 2596 7346 2648 7352
rect 2410 7304 2466 7313
rect 2410 7239 2466 7248
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2320 5704 2372 5710
rect 2320 5646 2372 5652
rect 2136 5636 2188 5642
rect 2136 5578 2188 5584
rect 2044 5160 2096 5166
rect 2044 5102 2096 5108
rect 2056 4622 2084 5102
rect 2148 4826 2176 5578
rect 2332 5370 2360 5646
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1952 3528 2004 3534
rect 1952 3470 2004 3476
rect 1964 3194 1992 3470
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1676 3120 1728 3126
rect 1676 3062 1728 3068
rect 2056 3058 2084 4558
rect 2148 4146 2176 4762
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2148 2774 2176 3878
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2056 2746 2176 2774
rect 2056 1986 2084 2746
rect 2240 2446 2268 2994
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 1964 1958 2084 1986
rect 20 1294 72 1300
rect 32 800 60 1294
rect 664 1284 716 1290
rect 664 1226 716 1232
rect 1320 1278 1440 1306
rect 1584 1352 1636 1358
rect 1584 1294 1636 1300
rect 676 800 704 1226
rect 1320 800 1348 1278
rect 1964 800 1992 1958
rect 2332 1290 2360 3878
rect 2424 3602 2452 7239
rect 2608 5846 2636 7346
rect 2700 7206 2728 10798
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2792 10713 2820 10746
rect 2778 10704 2834 10713
rect 2777 10668 2778 10674
rect 3068 10674 3096 11018
rect 3344 10826 3372 14980
rect 3424 14884 3476 14890
rect 3424 14826 3476 14832
rect 3436 13870 3464 14826
rect 3528 14822 3556 16594
rect 3988 16182 4016 17614
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16516 4120 16522
rect 4068 16458 4120 16464
rect 4080 16250 4108 16458
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3988 15502 4016 16118
rect 4632 16046 4660 16934
rect 4724 16674 4752 20810
rect 5724 20800 5776 20806
rect 5724 20742 5776 20748
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5736 20534 5764 20742
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 5276 18426 5304 19110
rect 6012 18970 6040 22494
rect 6000 18964 6052 18970
rect 6000 18906 6052 18912
rect 5540 18692 5592 18698
rect 5540 18634 5592 18640
rect 5552 18426 5580 18634
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5540 18420 5592 18426
rect 5540 18362 5592 18368
rect 5276 17610 5304 18362
rect 6012 18358 6040 18906
rect 6000 18352 6052 18358
rect 6000 18294 6052 18300
rect 6104 18222 6132 24160
rect 6276 24200 6328 24206
rect 6276 24142 6328 24148
rect 6368 24200 6420 24206
rect 6368 24142 6420 24148
rect 6288 22778 6316 24142
rect 6564 24138 6592 25094
rect 6552 24132 6604 24138
rect 6552 24074 6604 24080
rect 6656 23594 6684 25214
rect 6828 24744 6880 24750
rect 6828 24686 6880 24692
rect 6840 24614 6868 24686
rect 6828 24608 6880 24614
rect 6828 24550 6880 24556
rect 6736 24336 6788 24342
rect 6932 24290 6960 25366
rect 7024 24410 7052 25638
rect 7576 25294 7604 25638
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7012 24404 7064 24410
rect 7012 24346 7064 24352
rect 6788 24284 6960 24290
rect 6736 24278 6960 24284
rect 6748 24262 6960 24278
rect 6644 23588 6696 23594
rect 6644 23530 6696 23536
rect 6656 23202 6684 23530
rect 6564 23174 6684 23202
rect 6276 22772 6328 22778
rect 6276 22714 6328 22720
rect 6564 22642 6592 23174
rect 6644 23112 6696 23118
rect 6644 23054 6696 23060
rect 6552 22636 6604 22642
rect 6552 22578 6604 22584
rect 6552 21888 6604 21894
rect 6552 21830 6604 21836
rect 6564 21350 6592 21830
rect 6656 21554 6684 23054
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6736 22568 6788 22574
rect 6736 22510 6788 22516
rect 6748 21894 6776 22510
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 21622 6776 21830
rect 6736 21616 6788 21622
rect 6736 21558 6788 21564
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6460 21344 6512 21350
rect 6460 21286 6512 21292
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6368 21072 6420 21078
rect 6472 21060 6500 21286
rect 6552 21072 6604 21078
rect 6472 21032 6552 21060
rect 6368 21014 6420 21020
rect 6840 21026 6868 22578
rect 7012 22500 7064 22506
rect 7012 22442 7064 22448
rect 7024 22030 7052 22442
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 7024 21690 7052 21966
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6932 21146 6960 21490
rect 6920 21140 6972 21146
rect 6920 21082 6972 21088
rect 6552 21014 6604 21020
rect 6184 20868 6236 20874
rect 6184 20810 6236 20816
rect 6196 20602 6224 20810
rect 6380 20602 6408 21014
rect 6748 20998 6868 21026
rect 6184 20596 6236 20602
rect 6184 20538 6236 20544
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6380 20058 6408 20402
rect 6368 20052 6420 20058
rect 6368 19994 6420 20000
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6656 19514 6684 19790
rect 6748 19718 6776 20998
rect 6828 20936 6880 20942
rect 6828 20878 6880 20884
rect 6840 20602 6868 20878
rect 6828 20596 6880 20602
rect 6828 20538 6880 20544
rect 6840 19854 6868 20538
rect 7012 20460 7064 20466
rect 7012 20402 7064 20408
rect 7024 19938 7052 20402
rect 7116 20058 7144 25230
rect 7472 25220 7524 25226
rect 7472 25162 7524 25168
rect 7484 24818 7512 25162
rect 7576 24886 7604 25230
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7564 24880 7616 24886
rect 7564 24822 7616 24828
rect 7668 24818 7696 25094
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7288 24744 7340 24750
rect 7564 24744 7616 24750
rect 7340 24692 7512 24698
rect 7288 24686 7512 24692
rect 7564 24686 7616 24692
rect 7748 24744 7800 24750
rect 7748 24686 7800 24692
rect 7300 24670 7512 24686
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7208 24138 7236 24550
rect 7392 24206 7420 24550
rect 7484 24410 7512 24670
rect 7576 24614 7604 24686
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7196 24132 7248 24138
rect 7196 24074 7248 24080
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7208 22030 7236 22374
rect 7300 22030 7328 22578
rect 7392 22098 7420 24142
rect 7760 24070 7788 24686
rect 7852 24410 7880 25842
rect 7944 25362 7972 25842
rect 8220 25770 8248 25910
rect 8404 25906 8432 26726
rect 8392 25900 8444 25906
rect 8392 25842 8444 25848
rect 8496 25838 8524 26930
rect 9048 25974 9076 26982
rect 9128 26852 9180 26858
rect 9128 26794 9180 26800
rect 9140 26382 9168 26794
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9036 25968 9088 25974
rect 9036 25910 9088 25916
rect 8484 25832 8536 25838
rect 8484 25774 8536 25780
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 7932 25356 7984 25362
rect 7932 25298 7984 25304
rect 8220 24614 8248 25706
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8208 24608 8260 24614
rect 8208 24550 8260 24556
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 8116 24404 8168 24410
rect 8116 24346 8168 24352
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7760 23866 7788 24006
rect 7748 23860 7800 23866
rect 7748 23802 7800 23808
rect 8128 23730 8156 24346
rect 8312 24274 8340 25230
rect 8392 25152 8444 25158
rect 8392 25094 8444 25100
rect 8300 24268 8352 24274
rect 8300 24210 8352 24216
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8220 23866 8248 24142
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8404 23730 8432 25094
rect 9140 24682 9168 26318
rect 9128 24676 9180 24682
rect 9128 24618 9180 24624
rect 8668 24064 8720 24070
rect 8668 24006 8720 24012
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8392 23724 8444 23730
rect 8392 23666 8444 23672
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7484 22642 7512 23462
rect 8484 23112 8536 23118
rect 8484 23054 8536 23060
rect 8496 22642 8524 23054
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 8484 22636 8536 22642
rect 8484 22578 8536 22584
rect 8392 22568 8444 22574
rect 8392 22510 8444 22516
rect 7472 22500 7524 22506
rect 7472 22442 7524 22448
rect 7380 22092 7432 22098
rect 7380 22034 7432 22040
rect 7196 22024 7248 22030
rect 7196 21966 7248 21972
rect 7288 22024 7340 22030
rect 7288 21966 7340 21972
rect 7300 21554 7328 21966
rect 7380 21956 7432 21962
rect 7380 21898 7432 21904
rect 7288 21548 7340 21554
rect 7288 21490 7340 21496
rect 7392 21434 7420 21898
rect 7484 21554 7512 22442
rect 7564 22432 7616 22438
rect 7564 22374 7616 22380
rect 7472 21548 7524 21554
rect 7472 21490 7524 21496
rect 7576 21486 7604 22374
rect 8404 22166 8432 22510
rect 8392 22160 8444 22166
rect 8392 22102 8444 22108
rect 7656 21956 7708 21962
rect 7656 21898 7708 21904
rect 7668 21690 7696 21898
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7300 21406 7420 21434
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7300 20942 7328 21406
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7288 20936 7340 20942
rect 7288 20878 7340 20884
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7024 19910 7144 19938
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 7012 19848 7064 19854
rect 7012 19790 7064 19796
rect 6736 19712 6788 19718
rect 6736 19654 6788 19660
rect 6644 19508 6696 19514
rect 6644 19450 6696 19456
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4724 16646 4844 16674
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3528 14414 3556 14758
rect 3516 14408 3568 14414
rect 3516 14350 3568 14356
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3424 13456 3476 13462
rect 3424 13398 3476 13404
rect 3436 12918 3464 13398
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 3620 12782 3648 14214
rect 3988 14074 4016 15438
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 4264 15026 4292 15302
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14340 4120 14346
rect 4068 14282 4120 14288
rect 4080 14074 4108 14282
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4068 14068 4120 14074
rect 4068 14010 4120 14016
rect 3792 14000 3844 14006
rect 3792 13942 3844 13948
rect 3804 13394 3832 13942
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3988 12986 4016 14010
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4252 13252 4304 13258
rect 4252 13194 4304 13200
rect 4264 12986 4292 13194
rect 3976 12980 4028 12986
rect 3976 12922 4028 12928
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4724 12866 4752 16050
rect 4632 12838 4752 12866
rect 3608 12776 3660 12782
rect 3608 12718 3660 12724
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 4080 12442 4108 12718
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12436 4120 12442
rect 3896 12406 4068 12434
rect 3896 12306 3924 12406
rect 4068 12378 4120 12384
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 4436 12232 4488 12238
rect 4436 12174 4488 12180
rect 3884 12164 3936 12170
rect 3884 12106 3936 12112
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11762 3648 12038
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3252 10798 3372 10826
rect 2829 10639 2834 10648
rect 3056 10668 3108 10674
rect 2777 10610 2829 10616
rect 3056 10610 3108 10616
rect 2964 10532 3016 10538
rect 2964 10474 3016 10480
rect 2976 10266 3004 10474
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 3068 9674 3096 10610
rect 3252 10470 3280 10798
rect 3436 10674 3464 11222
rect 3712 10674 3740 11290
rect 3804 11150 3832 11834
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 2792 9646 3096 9674
rect 2792 9110 2820 9646
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8265 2820 8774
rect 2976 8566 3004 8910
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 2964 8560 3016 8566
rect 2964 8502 3016 8508
rect 3056 8288 3108 8294
rect 2778 8256 2834 8265
rect 3056 8230 3108 8236
rect 2778 8191 2834 8200
rect 2964 7744 3016 7750
rect 2964 7686 3016 7692
rect 2976 7585 3004 7686
rect 2962 7576 3018 7585
rect 2962 7511 3018 7520
rect 2872 7472 2924 7478
rect 2872 7414 2924 7420
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2780 6996 2832 7002
rect 2780 6938 2832 6944
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 2700 6458 2728 6666
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2596 5840 2648 5846
rect 2596 5782 2648 5788
rect 2792 5658 2820 6938
rect 2884 6662 2912 7414
rect 2964 7404 3016 7410
rect 3068 7392 3096 8230
rect 3160 7886 3188 8570
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3016 7364 3096 7392
rect 2964 7346 3016 7352
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2872 6656 2924 6662
rect 2872 6598 2924 6604
rect 2884 5778 2912 6598
rect 2976 6322 3004 7142
rect 3068 7002 3096 7364
rect 3056 6996 3108 7002
rect 3056 6938 3108 6944
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3068 5846 3096 6258
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 2872 5772 2924 5778
rect 2872 5714 2924 5720
rect 2792 5630 2912 5658
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5302 2820 5510
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2884 4486 2912 5630
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4622 3004 4966
rect 2964 4616 3016 4622
rect 2964 4558 3016 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2884 4214 2912 4422
rect 2872 4208 2924 4214
rect 2872 4150 2924 4156
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2412 3596 2464 3602
rect 2412 3538 2464 3544
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2516 1714 2544 3334
rect 2608 3058 2636 3334
rect 2792 3194 2820 4082
rect 2976 3534 3004 4558
rect 3068 3670 3096 5782
rect 3240 5704 3292 5710
rect 3240 5646 3292 5652
rect 3252 5370 3280 5646
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3344 4162 3372 10610
rect 3424 10532 3476 10538
rect 3424 10474 3476 10480
rect 3436 7970 3464 10474
rect 3528 10062 3556 10610
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3528 9674 3556 9998
rect 3528 9646 3648 9674
rect 3516 9104 3568 9110
rect 3516 9046 3568 9052
rect 3528 8430 3556 9046
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3620 8022 3648 9646
rect 3712 8974 3740 10610
rect 3804 9654 3832 11086
rect 3896 10742 3924 12106
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11150 4016 11494
rect 4080 11354 4108 12038
rect 4356 11898 4384 12038
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4448 11540 4476 12174
rect 4632 11608 4660 12838
rect 4712 12776 4764 12782
rect 4712 12718 4764 12724
rect 4724 12238 4752 12718
rect 4816 12434 4844 16646
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5276 15722 5304 17546
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5368 16114 5396 16390
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5368 15910 5396 16050
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5276 15694 5396 15722
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 5276 12442 5304 13126
rect 5264 12436 5316 12442
rect 4816 12406 5212 12434
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11898 4752 12174
rect 5184 12152 5212 12406
rect 5368 12434 5396 15694
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5552 15366 5580 15574
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 15162 5580 15302
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5368 12406 5488 12434
rect 5264 12378 5316 12384
rect 5356 12368 5408 12374
rect 5356 12310 5408 12316
rect 5184 12124 5304 12152
rect 4804 12096 4856 12102
rect 4804 12038 4856 12044
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4632 11580 4752 11608
rect 4448 11512 4660 11540
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4632 11286 4660 11512
rect 4620 11280 4672 11286
rect 4620 11222 4672 11228
rect 3976 11144 4028 11150
rect 3976 11086 4028 11092
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 4172 10674 4200 10950
rect 4264 10742 4292 11018
rect 4724 11014 4752 11580
rect 4816 11218 4844 12038
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4896 11824 4948 11830
rect 4896 11766 4948 11772
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4908 11150 4936 11766
rect 5080 11756 5132 11762
rect 5080 11698 5132 11704
rect 5092 11354 5120 11698
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 4896 11144 4948 11150
rect 4896 11086 4948 11092
rect 4712 11008 4764 11014
rect 4712 10950 4764 10956
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4160 10668 4212 10674
rect 4080 10628 4160 10656
rect 4080 9722 4108 10628
rect 4160 10610 4212 10616
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 3792 9648 3844 9654
rect 3792 9590 3844 9596
rect 3804 9058 3832 9590
rect 4172 9518 4200 9930
rect 4632 9518 4660 10610
rect 4712 10464 4764 10470
rect 4712 10406 4764 10412
rect 4724 9518 4752 10406
rect 4896 10056 4948 10062
rect 4816 10004 4896 10010
rect 4816 9998 4948 10004
rect 4816 9982 4936 9998
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3804 9030 3924 9058
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3608 8016 3660 8022
rect 3436 7942 3556 7970
rect 3608 7958 3660 7964
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3436 4826 3464 7822
rect 3528 5794 3556 7942
rect 3712 7342 3740 8910
rect 3896 8498 3924 9030
rect 4080 8974 4108 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4436 9172 4488 9178
rect 4436 9114 4488 9120
rect 4344 9036 4396 9042
rect 4344 8978 4396 8984
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4356 8498 4384 8978
rect 4448 8498 4476 9114
rect 4632 9042 4660 9454
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3804 6798 3832 8366
rect 3896 8072 3924 8434
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 8090 4660 8366
rect 4620 8084 4672 8090
rect 3896 8044 4200 8072
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3792 6792 3844 6798
rect 3792 6734 3844 6740
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6390 3832 6598
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 3528 5766 3648 5794
rect 3516 5704 3568 5710
rect 3516 5646 3568 5652
rect 3528 5234 3556 5646
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3528 4185 3556 4558
rect 3514 4176 3570 4185
rect 3344 4134 3464 4162
rect 3148 4004 3200 4010
rect 3148 3946 3200 3952
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2792 2650 2820 3130
rect 3160 3058 3188 3946
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3252 2650 3280 3470
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3240 2644 3292 2650
rect 3240 2586 3292 2592
rect 3344 1986 3372 3946
rect 3436 3942 3464 4134
rect 3514 4111 3516 4120
rect 3568 4111 3570 4120
rect 3516 4082 3568 4088
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3620 3738 3648 5766
rect 3896 5710 3924 6054
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3896 5370 3924 5646
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3712 2854 3740 4082
rect 3896 3534 3924 5306
rect 3988 4826 4016 7822
rect 4172 7478 4200 8044
rect 4620 8026 4672 8032
rect 4528 7948 4580 7954
rect 4528 7890 4580 7896
rect 4252 7880 4304 7886
rect 4252 7822 4304 7828
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4264 7410 4292 7822
rect 4540 7478 4568 7890
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4632 7410 4660 7754
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4436 6792 4488 6798
rect 4436 6734 4488 6740
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 4172 6322 4200 6666
rect 4448 6390 4476 6734
rect 4540 6458 4568 6734
rect 4632 6662 4660 7142
rect 4724 6780 4752 8910
rect 4816 7546 4844 9982
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5092 8906 5120 9658
rect 5184 8945 5212 9658
rect 5170 8936 5226 8945
rect 5080 8900 5132 8906
rect 5170 8871 5226 8880
rect 5080 8842 5132 8848
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 7886 5304 12124
rect 5368 10452 5396 12310
rect 5460 10554 5488 12406
rect 5552 11830 5580 15098
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5736 12170 5764 13126
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5540 11824 5592 11830
rect 5592 11784 5672 11812
rect 5540 11766 5592 11772
rect 5540 11552 5592 11558
rect 5540 11494 5592 11500
rect 5552 10742 5580 11494
rect 5540 10736 5592 10742
rect 5540 10678 5592 10684
rect 5460 10526 5580 10554
rect 5448 10464 5500 10470
rect 5368 10424 5448 10452
rect 5368 9994 5396 10424
rect 5448 10406 5500 10412
rect 5552 10282 5580 10526
rect 5460 10254 5580 10282
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5368 9586 5396 9930
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5460 8974 5488 10254
rect 5644 9722 5672 11784
rect 5828 10810 5856 17070
rect 6104 15570 6132 18158
rect 6840 17746 6868 18226
rect 6184 17740 6236 17746
rect 6184 17682 6236 17688
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6196 17338 6224 17682
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6748 17338 6776 17478
rect 7024 17338 7052 19790
rect 7116 19334 7144 19910
rect 7208 19446 7236 20334
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7300 19334 7328 20878
rect 7392 19922 7420 21286
rect 7472 20936 7524 20942
rect 7472 20878 7524 20884
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7484 20602 7512 20878
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7380 19916 7432 19922
rect 7380 19858 7432 19864
rect 7484 19854 7512 20538
rect 7576 19854 7604 20878
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7760 20058 7788 20402
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7564 19848 7616 19854
rect 7564 19790 7616 19796
rect 7484 19334 7512 19790
rect 7116 19306 7328 19334
rect 7300 18358 7328 19306
rect 7392 19306 7512 19334
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7288 18352 7340 18358
rect 7288 18294 7340 18300
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7300 17202 7328 18294
rect 7392 18068 7420 19306
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7484 18426 7512 18770
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7472 18080 7524 18086
rect 7392 18040 7472 18068
rect 7472 18022 7524 18028
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7300 16726 7328 17138
rect 7484 16794 7512 18022
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 7288 16720 7340 16726
rect 7288 16662 7340 16668
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6472 15570 6500 16390
rect 7576 16250 7604 16458
rect 7564 16244 7616 16250
rect 7564 16186 7616 16192
rect 6920 16176 6972 16182
rect 6920 16118 6972 16124
rect 6644 16108 6696 16114
rect 6644 16050 6696 16056
rect 6656 15706 6684 16050
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6092 15564 6144 15570
rect 6092 15506 6144 15512
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 6828 15496 6880 15502
rect 6828 15438 6880 15444
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6656 14618 6684 14962
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6840 14550 6868 15438
rect 6932 15094 6960 16118
rect 7668 15570 7696 19314
rect 7852 19242 7880 20810
rect 8404 20262 8432 20810
rect 8576 20800 8628 20806
rect 8576 20742 8628 20748
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8588 20058 8616 20742
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8208 19440 8260 19446
rect 8208 19382 8260 19388
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 7840 19236 7892 19242
rect 7840 19178 7892 19184
rect 7852 17610 7880 19178
rect 8128 18970 8156 19314
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 8128 17678 8156 18022
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 7840 17604 7892 17610
rect 7840 17546 7892 17552
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 16046 7788 16390
rect 7852 16114 7880 17546
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8036 16250 8064 17138
rect 8116 16720 8168 16726
rect 8116 16662 8168 16668
rect 8024 16244 8076 16250
rect 8024 16186 8076 16192
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7748 16040 7800 16046
rect 7748 15982 7800 15988
rect 8128 15570 8156 16662
rect 8220 16182 8248 19382
rect 8576 18896 8628 18902
rect 8576 18838 8628 18844
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8312 17338 8340 17818
rect 8392 17536 8444 17542
rect 8392 17478 8444 17484
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8404 17202 8432 17478
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 8300 17060 8352 17066
rect 8300 17002 8352 17008
rect 8312 16726 8340 17002
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16794 8524 16934
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8300 16720 8352 16726
rect 8300 16662 8352 16668
rect 8496 16522 8524 16730
rect 8484 16516 8536 16522
rect 8484 16458 8536 16464
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8312 16182 8340 16390
rect 8208 16176 8260 16182
rect 8208 16118 8260 16124
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8220 16046 8248 16118
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8300 15904 8352 15910
rect 8300 15846 8352 15852
rect 8312 15706 8340 15846
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 7656 15564 7708 15570
rect 7656 15506 7708 15512
rect 8116 15564 8168 15570
rect 8116 15506 8168 15512
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6932 14414 6960 15030
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 6012 13870 6040 14282
rect 6932 14006 6960 14350
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5632 9716 5684 9722
rect 5632 9658 5684 9664
rect 5908 9172 5960 9178
rect 6012 9160 6040 13806
rect 6092 13184 6144 13190
rect 6092 13126 6144 13132
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6104 12986 6132 13126
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6196 12434 6224 13126
rect 5960 9132 6040 9160
rect 5908 9114 5960 9120
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 8072 5396 8842
rect 5368 8044 5488 8072
rect 5356 7948 5408 7954
rect 5356 7890 5408 7896
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 5368 7410 5396 7890
rect 5460 7426 5488 8044
rect 6012 7886 6040 9132
rect 6104 12406 6224 12434
rect 6104 8022 6132 12406
rect 6276 11076 6328 11082
rect 6276 11018 6328 11024
rect 6288 10810 6316 11018
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6380 9654 6408 13942
rect 6656 13326 6684 13942
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 6564 11286 6592 12378
rect 6656 12238 6684 13262
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 11762 6684 12174
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6656 11150 6684 11698
rect 7024 11354 7052 15302
rect 7392 14482 7420 15302
rect 7668 15162 7696 15506
rect 8128 15162 8156 15506
rect 7656 15156 7708 15162
rect 7656 15098 7708 15104
rect 8116 15156 8168 15162
rect 8116 15098 8168 15104
rect 7380 14476 7432 14482
rect 7380 14418 7432 14424
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7116 12850 7144 12922
rect 7104 12844 7156 12850
rect 7104 12786 7156 12792
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 7116 12442 7144 12786
rect 7208 12617 7236 12786
rect 7194 12608 7250 12617
rect 7194 12543 7250 12552
rect 7104 12436 7156 12442
rect 7392 12434 7420 12786
rect 7944 12646 7972 14350
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8128 12986 8156 14214
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8116 12776 8168 12782
rect 8116 12718 8168 12724
rect 7932 12640 7984 12646
rect 7932 12582 7984 12588
rect 7392 12406 7788 12434
rect 7104 12378 7156 12384
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11830 7420 12038
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7012 11348 7064 11354
rect 7012 11290 7064 11296
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10674 7328 10950
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6840 10266 6868 10542
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6196 8362 6224 8570
rect 6380 8566 6408 9590
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6920 9580 6972 9586
rect 7288 9580 7340 9586
rect 6972 9540 7052 9568
rect 6920 9522 6972 9528
rect 6460 8900 6512 8906
rect 6460 8842 6512 8848
rect 6368 8560 6420 8566
rect 6368 8502 6420 8508
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6092 8016 6144 8022
rect 6092 7958 6144 7964
rect 6000 7880 6052 7886
rect 5920 7840 6000 7868
rect 5356 7404 5408 7410
rect 5460 7398 5580 7426
rect 5356 7346 5408 7352
rect 5368 6882 5396 7346
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5276 6854 5396 6882
rect 5276 6798 5304 6854
rect 5460 6798 5488 7278
rect 4804 6792 4856 6798
rect 4724 6752 4804 6780
rect 4804 6734 4856 6740
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4436 6384 4488 6390
rect 4632 6338 4660 6394
rect 4488 6332 4660 6338
rect 4436 6326 4660 6332
rect 4160 6316 4212 6322
rect 4448 6310 4660 6326
rect 4724 6322 4752 6598
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 4712 6316 4764 6322
rect 4160 6258 4212 6264
rect 4712 6258 4764 6264
rect 4172 6202 4200 6258
rect 4080 6174 4200 6202
rect 4080 5234 4108 6174
rect 4804 6112 4856 6118
rect 4804 6054 4856 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 4080 4706 4108 5170
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3988 4678 4108 4706
rect 3988 4214 4016 4678
rect 4632 4622 4660 4966
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 3976 4208 4028 4214
rect 3976 4150 4028 4156
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3896 2938 3924 2994
rect 3988 2938 4016 4150
rect 4080 3058 4108 4558
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4632 4214 4660 4422
rect 4724 4282 4752 5170
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4620 4208 4672 4214
rect 4816 4162 4844 6054
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5172 5228 5224 5234
rect 5276 5216 5304 6394
rect 5368 5778 5396 6734
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5356 5772 5408 5778
rect 5356 5714 5408 5720
rect 5368 5234 5396 5714
rect 5224 5188 5304 5216
rect 5172 5170 5224 5176
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4620 4150 4672 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4250 3632 4306 3641
rect 4250 3567 4306 3576
rect 4264 3534 4292 3567
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4172 3194 4200 3334
rect 4160 3188 4212 3194
rect 4160 3130 4212 3136
rect 4540 3126 4568 3334
rect 4528 3120 4580 3126
rect 4528 3062 4580 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 3896 2922 4108 2938
rect 3896 2916 4120 2922
rect 3896 2910 4068 2916
rect 3700 2848 3752 2854
rect 3700 2790 3752 2796
rect 3712 2446 3740 2790
rect 3896 2774 3924 2910
rect 4068 2858 4120 2864
rect 3804 2746 3924 2774
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 3700 2440 3752 2446
rect 3700 2382 3752 2388
rect 3804 2378 3832 2746
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2446 4660 4150
rect 4724 4134 4844 4162
rect 4724 2446 4752 4134
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 4816 3194 4844 3470
rect 5000 3398 5028 3470
rect 5172 3460 5224 3466
rect 5276 3448 5304 5188
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5460 4978 5488 6326
rect 5552 5234 5580 7398
rect 5540 5228 5592 5234
rect 5816 5228 5868 5234
rect 5592 5188 5672 5216
rect 5540 5170 5592 5176
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5552 4978 5580 5034
rect 5460 4950 5580 4978
rect 5460 4570 5488 4950
rect 5540 4616 5592 4622
rect 5460 4564 5540 4570
rect 5460 4558 5592 4564
rect 5460 4542 5580 4558
rect 5460 3534 5488 4542
rect 5644 4486 5672 5188
rect 5816 5170 5868 5176
rect 5724 5024 5776 5030
rect 5724 4966 5776 4972
rect 5736 4554 5764 4966
rect 5724 4548 5776 4554
rect 5724 4490 5776 4496
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5448 3528 5500 3534
rect 5448 3470 5500 3476
rect 5224 3420 5304 3448
rect 5172 3402 5224 3408
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5460 2446 5488 3062
rect 5828 2990 5856 5170
rect 5920 5098 5948 7840
rect 6000 7822 6052 7828
rect 6196 7478 6224 8298
rect 6472 8090 6500 8842
rect 6656 8838 6684 9522
rect 6748 9450 6776 9522
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 6748 9178 6776 9386
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6932 8974 6960 9386
rect 6920 8968 6972 8974
rect 6920 8910 6972 8916
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6748 7886 6776 8502
rect 6932 8498 6960 8910
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 6736 7880 6788 7886
rect 6736 7822 6788 7828
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6552 6792 6604 6798
rect 6552 6734 6604 6740
rect 6000 6656 6052 6662
rect 6000 6598 6052 6604
rect 6012 6390 6040 6598
rect 6000 6384 6052 6390
rect 6000 6326 6052 6332
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 5920 4554 5948 5034
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5816 2576 5868 2582
rect 5816 2518 5868 2524
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 3792 2372 3844 2378
rect 3792 2314 3844 2320
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 4528 2304 4580 2310
rect 4528 2246 4580 2252
rect 5172 2304 5224 2310
rect 5224 2264 5304 2292
rect 5172 2246 5224 2252
rect 3252 1958 3372 1986
rect 2516 1686 2636 1714
rect 2320 1284 2372 1290
rect 2320 1226 2372 1232
rect 2608 800 2636 1686
rect 3252 800 3280 1958
rect 3896 800 3924 2246
rect 4540 800 4568 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1170 5304 2264
rect 5184 1142 5304 1170
rect 5184 800 5212 1142
rect 5828 800 5856 2518
rect 6012 2446 6040 6326
rect 6564 6322 6592 6734
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6564 4214 6592 6258
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6840 4554 6868 5238
rect 6932 5166 6960 6666
rect 7024 6458 7052 9540
rect 7288 9522 7340 9528
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7300 9110 7328 9522
rect 7484 9178 7512 9522
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8498 7512 8774
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 7886 7420 8366
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7196 7404 7248 7410
rect 7248 7364 7328 7392
rect 7196 7346 7248 7352
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 7024 5846 7052 6258
rect 7104 6248 7156 6254
rect 7104 6190 7156 6196
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7024 5234 7052 5646
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 7024 4826 7052 5170
rect 7012 4820 7064 4826
rect 7012 4762 7064 4768
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6552 4208 6604 4214
rect 6550 4176 6552 4185
rect 6604 4176 6606 4185
rect 6606 4134 6684 4162
rect 6550 4111 6606 4120
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6196 2446 6224 2790
rect 6564 2446 6592 2858
rect 6656 2446 6684 4134
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6840 3738 6868 4014
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6840 3126 6868 3674
rect 7024 3584 7052 4762
rect 7116 4264 7144 6190
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7208 4826 7236 5170
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7196 4276 7248 4282
rect 7116 4236 7196 4264
rect 7196 4218 7248 4224
rect 7208 4146 7236 4218
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 6932 3556 7052 3584
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6932 2650 6960 3556
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7024 3126 7052 3334
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 6644 2440 6696 2446
rect 7208 2428 7236 4082
rect 7300 4010 7328 7364
rect 7392 6798 7420 7822
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7576 5030 7604 5578
rect 7656 5568 7708 5574
rect 7656 5510 7708 5516
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7576 4214 7604 4966
rect 7668 4622 7696 5510
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7300 3641 7328 3674
rect 7286 3632 7342 3641
rect 7286 3567 7342 3576
rect 7300 3534 7328 3567
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7484 2650 7512 3470
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7576 2446 7604 4150
rect 7760 2774 7788 12406
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 10810 7880 12038
rect 7944 11218 7972 12582
rect 8128 12238 8156 12718
rect 8220 12322 8248 13262
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8312 12442 8340 12786
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8220 12306 8340 12322
rect 8208 12300 8340 12306
rect 8260 12294 8340 12300
rect 8208 12242 8260 12248
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8312 12102 8340 12294
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8404 11354 8432 13126
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8496 11234 8524 12378
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8404 11206 8524 11234
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8128 10062 8156 10610
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8312 9382 8340 10542
rect 8404 10062 8432 11206
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 7944 9042 7972 9318
rect 8312 9042 8340 9318
rect 7932 9036 7984 9042
rect 7932 8978 7984 8984
rect 8300 9036 8352 9042
rect 8300 8978 8352 8984
rect 8312 7818 8340 8978
rect 8404 8498 8432 9998
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8036 7546 8064 7754
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8392 7336 8444 7342
rect 8390 7304 8392 7313
rect 8444 7304 8446 7313
rect 8390 7239 8446 7248
rect 8404 6934 8432 7239
rect 8392 6928 8444 6934
rect 8392 6870 8444 6876
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7852 4758 7880 6734
rect 7944 6458 7972 6734
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 8036 5370 8064 6734
rect 8392 5772 8444 5778
rect 8392 5714 8444 5720
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 7840 4752 7892 4758
rect 7840 4694 7892 4700
rect 8036 4622 8064 5306
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7840 4208 7892 4214
rect 7838 4176 7840 4185
rect 7892 4176 7894 4185
rect 7838 4111 7894 4120
rect 8036 3534 8064 4558
rect 8220 3602 8248 4626
rect 8404 4554 8432 5714
rect 8392 4548 8444 4554
rect 8392 4490 8444 4496
rect 8404 4282 8432 4490
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 8116 3392 8168 3398
rect 8116 3334 8168 3340
rect 8128 3058 8156 3334
rect 8312 3194 8340 4014
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7760 2746 8064 2774
rect 8036 2582 8064 2746
rect 8024 2576 8076 2582
rect 8024 2518 8076 2524
rect 8312 2446 8340 3130
rect 7288 2440 7340 2446
rect 7208 2400 7288 2428
rect 6644 2382 6696 2388
rect 7288 2382 7340 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8404 2378 8432 4218
rect 8496 4010 8524 10610
rect 8588 9450 8616 18838
rect 8680 18834 8708 24006
rect 9232 23050 9260 31726
rect 9324 31482 9352 31758
rect 9416 31754 9444 32982
rect 9416 31726 9628 31754
rect 9404 31680 9456 31686
rect 9404 31622 9456 31628
rect 9496 31680 9548 31686
rect 9496 31622 9548 31628
rect 9312 31476 9364 31482
rect 9312 31418 9364 31424
rect 9324 30734 9352 31418
rect 9416 31278 9444 31622
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30938 9444 31214
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9312 30728 9364 30734
rect 9312 30670 9364 30676
rect 9508 30598 9536 31622
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 9496 30592 9548 30598
rect 9496 30534 9548 30540
rect 9324 30122 9352 30534
rect 9404 30252 9456 30258
rect 9404 30194 9456 30200
rect 9312 30116 9364 30122
rect 9312 30058 9364 30064
rect 9416 29782 9444 30194
rect 9600 30122 9628 31726
rect 9876 30258 9904 33050
rect 9968 32978 9996 33458
rect 9956 32972 10008 32978
rect 9956 32914 10008 32920
rect 9968 31346 9996 32914
rect 10060 32910 10088 34002
rect 10244 33980 10272 34954
rect 10428 34202 10456 34954
rect 10416 34196 10468 34202
rect 10416 34138 10468 34144
rect 10416 33992 10468 33998
rect 10244 33952 10416 33980
rect 10416 33934 10468 33940
rect 10140 33584 10192 33590
rect 10140 33526 10192 33532
rect 10152 32978 10180 33526
rect 10428 33386 10456 33934
rect 10416 33380 10468 33386
rect 10416 33322 10468 33328
rect 10520 33318 10548 35022
rect 10796 35006 10916 35034
rect 10692 34672 10744 34678
rect 10692 34614 10744 34620
rect 10508 33312 10560 33318
rect 10508 33254 10560 33260
rect 10600 33312 10652 33318
rect 10600 33254 10652 33260
rect 10140 32972 10192 32978
rect 10140 32914 10192 32920
rect 10048 32904 10100 32910
rect 10048 32846 10100 32852
rect 10060 32502 10088 32846
rect 10048 32496 10100 32502
rect 10048 32438 10100 32444
rect 10152 32434 10180 32914
rect 10612 32910 10640 33254
rect 10600 32904 10652 32910
rect 10600 32846 10652 32852
rect 10232 32836 10284 32842
rect 10232 32778 10284 32784
rect 10244 32434 10272 32778
rect 10704 32722 10732 34614
rect 10796 33658 10824 35006
rect 11164 34746 11192 35584
rect 11348 35562 11376 36042
rect 11532 35834 11560 36110
rect 11520 35828 11572 35834
rect 11520 35770 11572 35776
rect 11428 35760 11480 35766
rect 11428 35702 11480 35708
rect 11336 35556 11388 35562
rect 11336 35498 11388 35504
rect 11440 35442 11468 35702
rect 11348 35414 11468 35442
rect 11348 35086 11376 35414
rect 11532 35086 11560 35770
rect 12084 35698 12112 36246
rect 12176 35766 12204 36314
rect 12268 36038 12296 37946
rect 12360 37874 12388 38150
rect 12636 37942 12664 39238
rect 12716 38956 12768 38962
rect 12716 38898 12768 38904
rect 12728 38554 12756 38898
rect 13912 38888 13964 38894
rect 13912 38830 13964 38836
rect 12716 38548 12768 38554
rect 12716 38490 12768 38496
rect 13924 38418 13952 38830
rect 13912 38412 13964 38418
rect 13912 38354 13964 38360
rect 13084 38276 13136 38282
rect 13084 38218 13136 38224
rect 13096 38010 13124 38218
rect 13084 38004 13136 38010
rect 13084 37946 13136 37952
rect 12624 37936 12676 37942
rect 12624 37878 12676 37884
rect 12348 37868 12400 37874
rect 12348 37810 12400 37816
rect 12808 37868 12860 37874
rect 12808 37810 12860 37816
rect 13360 37868 13412 37874
rect 13360 37810 13412 37816
rect 12360 37330 12388 37810
rect 12624 37800 12676 37806
rect 12624 37742 12676 37748
rect 12348 37324 12400 37330
rect 12348 37266 12400 37272
rect 12636 37262 12664 37742
rect 12820 37466 12848 37810
rect 12808 37460 12860 37466
rect 12808 37402 12860 37408
rect 13372 37262 13400 37810
rect 12624 37256 12676 37262
rect 12624 37198 12676 37204
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 12992 37188 13044 37194
rect 12992 37130 13044 37136
rect 12808 36100 12860 36106
rect 12808 36042 12860 36048
rect 12256 36032 12308 36038
rect 12256 35974 12308 35980
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12164 35760 12216 35766
rect 12164 35702 12216 35708
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 11612 35080 11664 35086
rect 11612 35022 11664 35028
rect 11152 34740 11204 34746
rect 11152 34682 11204 34688
rect 11164 33998 11192 34682
rect 11348 34678 11376 35022
rect 11336 34672 11388 34678
rect 11336 34614 11388 34620
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 11244 33992 11296 33998
rect 11244 33934 11296 33940
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10796 33522 10824 33594
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10796 33318 10824 33458
rect 10784 33312 10836 33318
rect 10784 33254 10836 33260
rect 11164 33096 11192 33934
rect 11256 33454 11284 33934
rect 11624 33658 11652 35022
rect 12084 35018 12112 35634
rect 12268 35494 12296 35974
rect 12348 35760 12400 35766
rect 12452 35748 12480 35974
rect 12532 35760 12584 35766
rect 12452 35720 12532 35748
rect 12348 35702 12400 35708
rect 12532 35702 12584 35708
rect 12256 35488 12308 35494
rect 12256 35430 12308 35436
rect 12268 35154 12296 35430
rect 12360 35290 12388 35702
rect 12440 35624 12492 35630
rect 12440 35566 12492 35572
rect 12624 35624 12676 35630
rect 12624 35566 12676 35572
rect 12348 35284 12400 35290
rect 12348 35226 12400 35232
rect 12256 35148 12308 35154
rect 12256 35090 12308 35096
rect 12072 35012 12124 35018
rect 12072 34954 12124 34960
rect 12084 33862 12112 34954
rect 12452 34950 12480 35566
rect 12440 34944 12492 34950
rect 12440 34886 12492 34892
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12268 33998 12296 34546
rect 12452 34542 12480 34886
rect 12532 34604 12584 34610
rect 12532 34546 12584 34552
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12348 34400 12400 34406
rect 12348 34342 12400 34348
rect 12256 33992 12308 33998
rect 12256 33934 12308 33940
rect 12072 33856 12124 33862
rect 12072 33798 12124 33804
rect 11612 33652 11664 33658
rect 11612 33594 11664 33600
rect 11704 33652 11756 33658
rect 11704 33594 11756 33600
rect 11244 33448 11296 33454
rect 11244 33390 11296 33396
rect 11164 33068 11284 33096
rect 10876 32972 10928 32978
rect 10876 32914 10928 32920
rect 11152 32972 11204 32978
rect 11152 32914 11204 32920
rect 10520 32694 10732 32722
rect 10520 32570 10548 32694
rect 10508 32564 10560 32570
rect 10508 32506 10560 32512
rect 10140 32428 10192 32434
rect 10140 32370 10192 32376
rect 10232 32428 10284 32434
rect 10232 32370 10284 32376
rect 10244 31822 10272 32370
rect 10232 31816 10284 31822
rect 10232 31758 10284 31764
rect 9956 31340 10008 31346
rect 9956 31282 10008 31288
rect 10244 30818 10272 31758
rect 10244 30790 10364 30818
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 10232 30728 10284 30734
rect 10232 30670 10284 30676
rect 9968 30394 9996 30670
rect 9956 30388 10008 30394
rect 9956 30330 10008 30336
rect 9864 30252 9916 30258
rect 9864 30194 9916 30200
rect 9588 30116 9640 30122
rect 9588 30058 9640 30064
rect 9496 30048 9548 30054
rect 9496 29990 9548 29996
rect 9404 29776 9456 29782
rect 9404 29718 9456 29724
rect 9416 29306 9444 29718
rect 9508 29646 9536 29990
rect 9496 29640 9548 29646
rect 9496 29582 9548 29588
rect 10244 29578 10272 30670
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 9404 29300 9456 29306
rect 9404 29242 9456 29248
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 10244 28762 10272 29106
rect 10232 28756 10284 28762
rect 10232 28698 10284 28704
rect 10336 28150 10364 30790
rect 10416 29844 10468 29850
rect 10416 29786 10468 29792
rect 10428 29714 10456 29786
rect 10416 29708 10468 29714
rect 10416 29650 10468 29656
rect 10324 28144 10376 28150
rect 10324 28086 10376 28092
rect 10428 28082 10456 29650
rect 10520 28558 10548 32506
rect 10888 31414 10916 32914
rect 11164 32434 11192 32914
rect 11256 32434 11284 33068
rect 11716 32570 11744 33594
rect 11980 33516 12032 33522
rect 12084 33504 12112 33798
rect 12268 33522 12296 33934
rect 12360 33930 12388 34342
rect 12544 34202 12572 34546
rect 12532 34196 12584 34202
rect 12532 34138 12584 34144
rect 12438 34096 12494 34105
rect 12438 34031 12440 34040
rect 12492 34031 12494 34040
rect 12440 34002 12492 34008
rect 12348 33924 12400 33930
rect 12348 33866 12400 33872
rect 12636 33590 12664 35566
rect 12820 35494 12848 36042
rect 12808 35488 12860 35494
rect 12808 35430 12860 35436
rect 13004 35086 13032 37130
rect 13924 36242 13952 38354
rect 13912 36236 13964 36242
rect 13912 36178 13964 36184
rect 13084 36168 13136 36174
rect 13084 36110 13136 36116
rect 13096 35834 13124 36110
rect 13084 35828 13136 35834
rect 13084 35770 13136 35776
rect 12992 35080 13044 35086
rect 12992 35022 13044 35028
rect 12716 34944 12768 34950
rect 12716 34886 12768 34892
rect 12728 34610 12756 34886
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 12808 34604 12860 34610
rect 12808 34546 12860 34552
rect 12820 34474 12848 34546
rect 12900 34536 12952 34542
rect 12900 34478 12952 34484
rect 12808 34468 12860 34474
rect 12808 34410 12860 34416
rect 12716 34400 12768 34406
rect 12716 34342 12768 34348
rect 12728 34134 12756 34342
rect 12716 34128 12768 34134
rect 12716 34070 12768 34076
rect 12820 33998 12848 34410
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12624 33584 12676 33590
rect 12624 33526 12676 33532
rect 12032 33476 12112 33504
rect 12256 33516 12308 33522
rect 11980 33458 12032 33464
rect 12256 33458 12308 33464
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 12164 33448 12216 33454
rect 12164 33390 12216 33396
rect 12176 32978 12204 33390
rect 12716 33312 12768 33318
rect 12716 33254 12768 33260
rect 12164 32972 12216 32978
rect 12164 32914 12216 32920
rect 11704 32564 11756 32570
rect 11704 32506 11756 32512
rect 11152 32428 11204 32434
rect 11152 32370 11204 32376
rect 11244 32428 11296 32434
rect 11244 32370 11296 32376
rect 11428 32224 11480 32230
rect 11428 32166 11480 32172
rect 11440 31822 11468 32166
rect 11428 31816 11480 31822
rect 11428 31758 11480 31764
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11060 31680 11112 31686
rect 11060 31622 11112 31628
rect 10876 31408 10928 31414
rect 10876 31350 10928 31356
rect 10692 31136 10744 31142
rect 10692 31078 10744 31084
rect 10784 31136 10836 31142
rect 10784 31078 10836 31084
rect 10704 30734 10732 31078
rect 10796 30870 10824 31078
rect 11072 30938 11100 31622
rect 11532 31346 11560 31758
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 11060 30932 11112 30938
rect 11060 30874 11112 30880
rect 10784 30864 10836 30870
rect 10784 30806 10836 30812
rect 10692 30728 10744 30734
rect 10692 30670 10744 30676
rect 10968 30728 11020 30734
rect 11072 30716 11100 30874
rect 11716 30802 11744 32506
rect 11888 32496 11940 32502
rect 11888 32438 11940 32444
rect 11152 30796 11204 30802
rect 11152 30738 11204 30744
rect 11704 30796 11756 30802
rect 11704 30738 11756 30744
rect 11020 30688 11100 30716
rect 10968 30670 11020 30676
rect 10784 30592 10836 30598
rect 10784 30534 10836 30540
rect 10796 29646 10824 30534
rect 11060 30252 11112 30258
rect 11060 30194 11112 30200
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 10600 29504 10652 29510
rect 10600 29446 10652 29452
rect 10612 29306 10640 29446
rect 10704 29306 10732 29582
rect 10876 29572 10928 29578
rect 11072 29560 11100 30194
rect 11164 29866 11192 30738
rect 11336 30728 11388 30734
rect 11336 30670 11388 30676
rect 11244 30592 11296 30598
rect 11244 30534 11296 30540
rect 11256 30054 11284 30534
rect 11348 30258 11376 30670
rect 11336 30252 11388 30258
rect 11336 30194 11388 30200
rect 11244 30048 11296 30054
rect 11244 29990 11296 29996
rect 11428 30048 11480 30054
rect 11428 29990 11480 29996
rect 11164 29850 11284 29866
rect 11164 29844 11296 29850
rect 11164 29838 11244 29844
rect 11244 29786 11296 29792
rect 10928 29532 11100 29560
rect 10876 29514 10928 29520
rect 10600 29300 10652 29306
rect 10600 29242 10652 29248
rect 10692 29300 10744 29306
rect 10692 29242 10744 29248
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10612 28558 10640 29106
rect 11072 28762 11100 29532
rect 11440 29238 11468 29990
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11428 29232 11480 29238
rect 11428 29174 11480 29180
rect 11060 28756 11112 28762
rect 11060 28698 11112 28704
rect 10508 28552 10560 28558
rect 10508 28494 10560 28500
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 11520 28552 11572 28558
rect 11520 28494 11572 28500
rect 10520 28082 10548 28494
rect 10612 28218 10640 28494
rect 10692 28484 10744 28490
rect 10692 28426 10744 28432
rect 11428 28484 11480 28490
rect 11428 28426 11480 28432
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 10704 28082 10732 28426
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 10416 28076 10468 28082
rect 10416 28018 10468 28024
rect 10508 28076 10560 28082
rect 10508 28018 10560 28024
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 9508 27674 9812 27690
rect 9876 27674 9904 28018
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 9496 27668 9812 27674
rect 9548 27662 9812 27668
rect 9496 27610 9548 27616
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9312 27464 9364 27470
rect 9310 27432 9312 27441
rect 9364 27432 9366 27441
rect 9310 27367 9366 27376
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 9312 27328 9364 27334
rect 9312 27270 9364 27276
rect 9324 26586 9352 27270
rect 9600 26926 9628 27338
rect 9692 26994 9720 27542
rect 9784 27334 9812 27662
rect 9864 27668 9916 27674
rect 9864 27610 9916 27616
rect 10152 27538 10180 27950
rect 10428 27826 10456 28018
rect 10336 27798 10456 27826
rect 10140 27532 10192 27538
rect 10140 27474 10192 27480
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9784 26790 9812 27270
rect 10152 26994 10180 27474
rect 10232 27396 10284 27402
rect 10232 27338 10284 27344
rect 10244 27062 10272 27338
rect 10232 27056 10284 27062
rect 10232 26998 10284 27004
rect 10140 26988 10192 26994
rect 10140 26930 10192 26936
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9312 26580 9364 26586
rect 9312 26522 9364 26528
rect 9324 26042 9352 26522
rect 9312 26036 9364 26042
rect 9312 25978 9364 25984
rect 9324 25158 9352 25978
rect 10152 25922 10180 26930
rect 10060 25906 10180 25922
rect 10048 25900 10180 25906
rect 10100 25894 10180 25900
rect 10048 25842 10100 25848
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 9508 25226 9536 25638
rect 10060 25294 10088 25842
rect 10048 25288 10100 25294
rect 10048 25230 10100 25236
rect 9496 25220 9548 25226
rect 9496 25162 9548 25168
rect 9312 25152 9364 25158
rect 9312 25094 9364 25100
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9784 23730 9812 24006
rect 10060 23798 10088 25230
rect 10048 23792 10100 23798
rect 10048 23734 10100 23740
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 10060 23118 10088 23734
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 9220 23044 9272 23050
rect 9220 22986 9272 22992
rect 9864 22976 9916 22982
rect 9864 22918 9916 22924
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8772 20806 8800 22578
rect 9876 21962 9904 22918
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9692 21554 9720 21830
rect 9876 21554 9904 21898
rect 9968 21554 9996 22170
rect 10060 22098 10088 23054
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9864 21548 9916 21554
rect 9864 21490 9916 21496
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 8760 20800 8812 20806
rect 8760 20742 8812 20748
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8772 18068 8800 20742
rect 9692 20534 9720 21490
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9784 20874 9812 21422
rect 10244 21146 10272 26998
rect 10336 26450 10364 27798
rect 10600 27328 10652 27334
rect 10704 27282 10732 28018
rect 10784 27532 10836 27538
rect 10784 27474 10836 27480
rect 10652 27276 10732 27282
rect 10600 27270 10732 27276
rect 10612 27254 10732 27270
rect 10416 27124 10468 27130
rect 10416 27066 10468 27072
rect 10428 26450 10456 27066
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10416 26444 10468 26450
rect 10416 26386 10468 26392
rect 10612 25498 10640 27254
rect 10692 27056 10744 27062
rect 10692 26998 10744 27004
rect 10704 26382 10732 26998
rect 10796 26382 10824 27474
rect 11152 27464 11204 27470
rect 11152 27406 11204 27412
rect 11164 26382 11192 27406
rect 11440 27402 11468 28426
rect 11532 28218 11560 28494
rect 11520 28212 11572 28218
rect 11520 28154 11572 28160
rect 11428 27396 11480 27402
rect 11428 27338 11480 27344
rect 11624 27334 11652 29514
rect 11716 29238 11744 30738
rect 11796 30728 11848 30734
rect 11796 30670 11848 30676
rect 11808 30258 11836 30670
rect 11796 30252 11848 30258
rect 11796 30194 11848 30200
rect 11704 29232 11756 29238
rect 11704 29174 11756 29180
rect 11808 29170 11836 30194
rect 11796 29164 11848 29170
rect 11796 29106 11848 29112
rect 11900 28490 11928 32438
rect 12176 30802 12204 32914
rect 12440 31816 12492 31822
rect 12440 31758 12492 31764
rect 12624 31816 12676 31822
rect 12624 31758 12676 31764
rect 12452 30818 12480 31758
rect 12636 31210 12664 31758
rect 12624 31204 12676 31210
rect 12624 31146 12676 31152
rect 12164 30796 12216 30802
rect 12452 30790 12664 30818
rect 12164 30738 12216 30744
rect 12176 30258 12204 30738
rect 12440 30728 12492 30734
rect 12440 30670 12492 30676
rect 12452 30258 12480 30670
rect 12636 30326 12664 30790
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 12452 30122 12480 30194
rect 12440 30116 12492 30122
rect 12440 30058 12492 30064
rect 12636 30054 12664 30262
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12624 30048 12676 30054
rect 12624 29990 12676 29996
rect 12360 29646 12388 29990
rect 11980 29640 12032 29646
rect 11980 29582 12032 29588
rect 12348 29640 12400 29646
rect 12348 29582 12400 29588
rect 11992 29170 12020 29582
rect 12164 29572 12216 29578
rect 12164 29514 12216 29520
rect 12176 29170 12204 29514
rect 11980 29164 12032 29170
rect 11980 29106 12032 29112
rect 12164 29164 12216 29170
rect 12164 29106 12216 29112
rect 12072 29096 12124 29102
rect 12072 29038 12124 29044
rect 11888 28484 11940 28490
rect 11888 28426 11940 28432
rect 12084 28082 12112 29038
rect 12360 28642 12388 29582
rect 12728 29238 12756 33254
rect 12820 33114 12848 33458
rect 12808 33108 12860 33114
rect 12808 33050 12860 33056
rect 12912 32842 12940 34478
rect 13004 34406 13032 35022
rect 13096 34610 13124 35770
rect 13176 34672 13228 34678
rect 13176 34614 13228 34620
rect 13084 34604 13136 34610
rect 13084 34546 13136 34552
rect 12992 34400 13044 34406
rect 12992 34342 13044 34348
rect 13096 34202 13124 34546
rect 13084 34196 13136 34202
rect 13084 34138 13136 34144
rect 12992 34128 13044 34134
rect 13096 34105 13124 34138
rect 12992 34070 13044 34076
rect 13082 34096 13138 34105
rect 13004 33862 13032 34070
rect 13082 34031 13138 34040
rect 13188 33998 13216 34614
rect 13360 34604 13412 34610
rect 13360 34546 13412 34552
rect 13372 34134 13400 34546
rect 13728 34196 13780 34202
rect 13728 34138 13780 34144
rect 13360 34128 13412 34134
rect 13360 34070 13412 34076
rect 13176 33992 13228 33998
rect 13176 33934 13228 33940
rect 13372 33862 13400 34070
rect 13740 33930 13768 34138
rect 13924 34066 13952 36178
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 13728 33924 13780 33930
rect 13728 33866 13780 33872
rect 12992 33856 13044 33862
rect 12992 33798 13044 33804
rect 13084 33856 13136 33862
rect 13084 33798 13136 33804
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 13360 33856 13412 33862
rect 13360 33798 13412 33804
rect 13096 33114 13124 33798
rect 13084 33108 13136 33114
rect 13084 33050 13136 33056
rect 13188 32842 13216 33798
rect 13924 33522 13952 34002
rect 13912 33516 13964 33522
rect 13912 33458 13964 33464
rect 13924 32910 13952 33458
rect 13912 32904 13964 32910
rect 13912 32846 13964 32852
rect 12900 32836 12952 32842
rect 12900 32778 12952 32784
rect 13176 32836 13228 32842
rect 13176 32778 13228 32784
rect 13924 32502 13952 32846
rect 13912 32496 13964 32502
rect 13912 32438 13964 32444
rect 12900 31816 12952 31822
rect 12900 31758 12952 31764
rect 12992 31816 13044 31822
rect 12992 31758 13044 31764
rect 12808 31204 12860 31210
rect 12808 31146 12860 31152
rect 12820 30938 12848 31146
rect 12808 30932 12860 30938
rect 12808 30874 12860 30880
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12820 30394 12848 30670
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 12912 29782 12940 31758
rect 13004 31278 13032 31758
rect 13924 31754 13952 32438
rect 13924 31726 14136 31754
rect 13360 31680 13412 31686
rect 13360 31622 13412 31628
rect 13372 31414 13400 31622
rect 13176 31408 13228 31414
rect 13176 31350 13228 31356
rect 13360 31408 13412 31414
rect 13360 31350 13412 31356
rect 13544 31408 13596 31414
rect 13544 31350 13596 31356
rect 12992 31272 13044 31278
rect 12992 31214 13044 31220
rect 12992 31136 13044 31142
rect 12992 31078 13044 31084
rect 13004 30870 13032 31078
rect 12992 30864 13044 30870
rect 12992 30806 13044 30812
rect 12900 29776 12952 29782
rect 12900 29718 12952 29724
rect 12900 29504 12952 29510
rect 12900 29446 12952 29452
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12268 28614 12388 28642
rect 11704 28076 11756 28082
rect 11704 28018 11756 28024
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 11716 27470 11744 28018
rect 11704 27464 11756 27470
rect 11704 27406 11756 27412
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11624 27112 11652 27270
rect 11624 27084 11744 27112
rect 11612 26988 11664 26994
rect 11612 26930 11664 26936
rect 11624 26586 11652 26930
rect 11716 26858 11744 27084
rect 11704 26852 11756 26858
rect 11704 26794 11756 26800
rect 11716 26586 11744 26794
rect 11612 26580 11664 26586
rect 11612 26522 11664 26528
rect 11704 26580 11756 26586
rect 11704 26522 11756 26528
rect 11428 26512 11480 26518
rect 11428 26454 11480 26460
rect 10692 26376 10744 26382
rect 10692 26318 10744 26324
rect 10784 26376 10836 26382
rect 10784 26318 10836 26324
rect 11152 26376 11204 26382
rect 11152 26318 11204 26324
rect 10692 26240 10744 26246
rect 10692 26182 10744 26188
rect 10704 25974 10732 26182
rect 11164 26042 11192 26318
rect 11152 26036 11204 26042
rect 11152 25978 11204 25984
rect 10692 25968 10744 25974
rect 10692 25910 10744 25916
rect 10600 25492 10652 25498
rect 10600 25434 10652 25440
rect 11440 25294 11468 26454
rect 11808 26314 11836 27338
rect 12084 27334 12112 28018
rect 12268 27402 12296 28614
rect 12348 28484 12400 28490
rect 12348 28426 12400 28432
rect 12624 28484 12676 28490
rect 12624 28426 12676 28432
rect 12360 28014 12388 28426
rect 12348 28008 12400 28014
rect 12348 27950 12400 27956
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 12072 27328 12124 27334
rect 11992 27288 12072 27316
rect 11992 26314 12020 27288
rect 12072 27270 12124 27276
rect 12072 26988 12124 26994
rect 12072 26930 12124 26936
rect 12084 26586 12112 26930
rect 12164 26784 12216 26790
rect 12164 26726 12216 26732
rect 12072 26580 12124 26586
rect 12072 26522 12124 26528
rect 11796 26308 11848 26314
rect 11796 26250 11848 26256
rect 11980 26308 12032 26314
rect 11980 26250 12032 26256
rect 11992 26042 12020 26250
rect 11980 26036 12032 26042
rect 11980 25978 12032 25984
rect 11980 25900 12032 25906
rect 11980 25842 12032 25848
rect 11992 25498 12020 25842
rect 11980 25492 12032 25498
rect 11980 25434 12032 25440
rect 12176 25362 12204 26726
rect 12268 26586 12296 27338
rect 12256 26580 12308 26586
rect 12256 26522 12308 26528
rect 12360 25974 12388 27950
rect 12636 27130 12664 28426
rect 12624 27124 12676 27130
rect 12624 27066 12676 27072
rect 12728 27062 12756 29038
rect 12820 27441 12848 29106
rect 12912 29102 12940 29446
rect 13004 29306 13032 30806
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 12992 29300 13044 29306
rect 12992 29242 13044 29248
rect 13096 29170 13124 30534
rect 13188 30326 13216 31350
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 13280 30734 13308 30874
rect 13452 30864 13504 30870
rect 13452 30806 13504 30812
rect 13464 30734 13492 30806
rect 13268 30728 13320 30734
rect 13268 30670 13320 30676
rect 13452 30728 13504 30734
rect 13452 30670 13504 30676
rect 13176 30320 13228 30326
rect 13176 30262 13228 30268
rect 13188 30190 13216 30262
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13176 29776 13228 29782
rect 13176 29718 13228 29724
rect 13084 29164 13136 29170
rect 13084 29106 13136 29112
rect 12900 29096 12952 29102
rect 12900 29038 12952 29044
rect 13188 28558 13216 29718
rect 13280 29594 13308 30670
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 13372 30138 13400 30330
rect 13372 30110 13492 30138
rect 13464 29646 13492 30110
rect 13452 29640 13504 29646
rect 13280 29566 13400 29594
rect 13452 29582 13504 29588
rect 13372 28694 13400 29566
rect 13452 29096 13504 29102
rect 13452 29038 13504 29044
rect 13360 28688 13412 28694
rect 13360 28630 13412 28636
rect 13464 28626 13492 29038
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 13176 28552 13228 28558
rect 13176 28494 13228 28500
rect 13556 28490 13584 31350
rect 14108 31142 14136 31726
rect 14096 31136 14148 31142
rect 14096 31078 14148 31084
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14108 30802 14136 31078
rect 14004 30796 14056 30802
rect 14004 30738 14056 30744
rect 14096 30796 14148 30802
rect 14096 30738 14148 30744
rect 13728 30184 13780 30190
rect 13728 30126 13780 30132
rect 13636 30116 13688 30122
rect 13636 30058 13688 30064
rect 13648 29646 13676 30058
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 13740 28490 13768 30126
rect 14016 30122 14044 30738
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14108 30326 14136 30534
rect 14096 30320 14148 30326
rect 14096 30262 14148 30268
rect 14476 30258 14504 31078
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14004 30116 14056 30122
rect 14004 30058 14056 30064
rect 14832 29640 14884 29646
rect 14832 29582 14884 29588
rect 14844 29306 14872 29582
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 13820 28552 13872 28558
rect 13820 28494 13872 28500
rect 13544 28484 13596 28490
rect 13544 28426 13596 28432
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 12900 28416 12952 28422
rect 12900 28358 12952 28364
rect 12912 28150 12940 28358
rect 13740 28218 13768 28426
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 12900 28144 12952 28150
rect 12900 28086 12952 28092
rect 12806 27432 12862 27441
rect 12806 27367 12862 27376
rect 12440 27056 12492 27062
rect 12440 26998 12492 27004
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12452 26926 12480 26998
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12716 26920 12768 26926
rect 12820 26874 12848 27367
rect 13832 26994 13860 28494
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 12768 26868 12848 26874
rect 12716 26862 12848 26868
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 12348 25968 12400 25974
rect 12348 25910 12400 25916
rect 12452 25430 12480 26862
rect 12728 26846 12848 26862
rect 13096 26586 13124 26862
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 13924 26296 13952 26930
rect 13740 26268 13952 26296
rect 13740 25974 13768 26268
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 13728 25968 13780 25974
rect 13728 25910 13780 25916
rect 12440 25424 12492 25430
rect 12440 25366 12492 25372
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 11428 25288 11480 25294
rect 11428 25230 11480 25236
rect 10416 24200 10468 24206
rect 10416 24142 10468 24148
rect 11980 24200 12032 24206
rect 11980 24142 12032 24148
rect 12072 24200 12124 24206
rect 12256 24200 12308 24206
rect 12072 24142 12124 24148
rect 12176 24160 12256 24188
rect 10428 22778 10456 24142
rect 11612 24132 11664 24138
rect 11612 24074 11664 24080
rect 10784 24064 10836 24070
rect 10784 24006 10836 24012
rect 10796 23118 10824 24006
rect 10784 23112 10836 23118
rect 10784 23054 10836 23060
rect 10416 22772 10468 22778
rect 10416 22714 10468 22720
rect 11624 22642 11652 24074
rect 11888 23724 11940 23730
rect 11888 23666 11940 23672
rect 11900 23322 11928 23666
rect 11992 23322 12020 24142
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 11704 23044 11756 23050
rect 11704 22986 11756 22992
rect 11716 22778 11744 22986
rect 12084 22778 12112 24142
rect 12176 23526 12204 24160
rect 12256 24142 12308 24148
rect 13280 23730 13308 25910
rect 13176 23724 13228 23730
rect 13176 23666 13228 23672
rect 13268 23724 13320 23730
rect 13268 23666 13320 23672
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12176 23118 12204 23462
rect 13188 23322 13216 23666
rect 13176 23316 13228 23322
rect 13176 23258 13228 23264
rect 12164 23112 12216 23118
rect 12164 23054 12216 23060
rect 12808 23112 12860 23118
rect 12808 23054 12860 23060
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 12072 22772 12124 22778
rect 12072 22714 12124 22720
rect 11612 22636 11664 22642
rect 11612 22578 11664 22584
rect 12164 22636 12216 22642
rect 12164 22578 12216 22584
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 11624 22094 11652 22578
rect 11440 22066 11652 22094
rect 11336 22024 11388 22030
rect 11336 21966 11388 21972
rect 11348 21690 11376 21966
rect 11440 21894 11468 22066
rect 12176 21894 12204 22578
rect 12452 22166 12480 22578
rect 12820 22574 12848 23054
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 12808 22568 12860 22574
rect 12808 22510 12860 22516
rect 12440 22160 12492 22166
rect 12440 22102 12492 22108
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 11440 21690 11468 21830
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11152 21548 11204 21554
rect 11152 21490 11204 21496
rect 11164 21146 11192 21490
rect 11808 21486 11836 21830
rect 11796 21480 11848 21486
rect 11796 21422 11848 21428
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 11244 21412 11296 21418
rect 11244 21354 11296 21360
rect 10232 21140 10284 21146
rect 10232 21082 10284 21088
rect 11152 21140 11204 21146
rect 11152 21082 11204 21088
rect 9864 21072 9916 21078
rect 9864 21014 9916 21020
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9680 20528 9732 20534
rect 9680 20470 9732 20476
rect 9220 20392 9272 20398
rect 9220 20334 9272 20340
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8864 18766 8892 20198
rect 9232 19514 9260 20334
rect 9508 20058 9536 20334
rect 9496 20052 9548 20058
rect 9496 19994 9548 20000
rect 9220 19508 9272 19514
rect 9220 19450 9272 19456
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 9508 18698 9536 19994
rect 9588 19780 9640 19786
rect 9588 19722 9640 19728
rect 9600 19174 9628 19722
rect 9692 19378 9720 20470
rect 9784 20262 9812 20810
rect 9876 20602 9904 21014
rect 9864 20596 9916 20602
rect 9864 20538 9916 20544
rect 9772 20256 9824 20262
rect 9772 20198 9824 20204
rect 9784 19446 9812 20198
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 9876 19242 9904 19790
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9600 18834 9628 19110
rect 9588 18828 9640 18834
rect 9588 18770 9640 18776
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9600 18222 9628 18770
rect 9588 18216 9640 18222
rect 9588 18158 9640 18164
rect 9876 18086 9904 19178
rect 10140 18828 10192 18834
rect 10140 18770 10192 18776
rect 8680 18040 8800 18068
rect 9864 18080 9916 18086
rect 8680 16726 8708 18040
rect 9864 18022 9916 18028
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8956 17338 8984 17546
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8864 17202 8892 17274
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8668 16720 8720 16726
rect 8668 16662 8720 16668
rect 8680 14362 8708 16662
rect 8864 15434 8892 17138
rect 9128 17060 9180 17066
rect 9128 17002 9180 17008
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 16182 8984 16390
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 9048 15706 9076 16458
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 8852 15428 8904 15434
rect 8852 15370 8904 15376
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8772 14482 8800 15302
rect 8852 15088 8904 15094
rect 8852 15030 8904 15036
rect 8864 14618 8892 15030
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8680 14334 8800 14362
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8680 11898 8708 12718
rect 8772 12238 8800 14334
rect 8864 13394 8892 14554
rect 8956 14414 8984 14758
rect 9048 14618 9076 14962
rect 9036 14612 9088 14618
rect 9036 14554 9088 14560
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 8852 13388 8904 13394
rect 8852 13330 8904 13336
rect 8956 12306 8984 14350
rect 9140 14006 9168 17002
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 15706 9352 16390
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9128 14000 9180 14006
rect 9128 13942 9180 13948
rect 9140 13870 9168 13942
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9324 12986 9352 14214
rect 9508 13394 9536 15302
rect 9600 15094 9628 16594
rect 9784 16250 9812 17206
rect 9876 17134 9904 18022
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9876 16658 9904 17070
rect 9864 16652 9916 16658
rect 9864 16594 9916 16600
rect 9772 16244 9824 16250
rect 9772 16186 9824 16192
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9600 14482 9628 15030
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9600 13784 9628 14418
rect 9876 14414 9904 16594
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 16250 9996 16390
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 10152 15570 10180 18770
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10060 15162 10088 15438
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9680 13796 9732 13802
rect 9600 13756 9680 13784
rect 9680 13738 9732 13744
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9876 12986 9904 13194
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8680 11150 8708 11834
rect 8956 11694 8984 12038
rect 9048 11898 9076 12650
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9508 11898 9536 12106
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 8944 11688 8996 11694
rect 8944 11630 8996 11636
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 8668 11144 8720 11150
rect 8668 11086 8720 11092
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9508 10742 9536 11018
rect 9496 10736 9548 10742
rect 9496 10678 9548 10684
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 8944 10464 8996 10470
rect 8944 10406 8996 10412
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8588 9042 8616 9386
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8668 7812 8720 7818
rect 8668 7754 8720 7760
rect 8680 7342 8708 7754
rect 8668 7336 8720 7342
rect 8668 7278 8720 7284
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8588 5658 8616 7142
rect 8680 6866 8708 7278
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8680 5794 8708 6394
rect 8772 5914 8800 9998
rect 8956 9654 8984 10406
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9048 8498 9076 9114
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8864 7886 8892 8434
rect 9048 8090 9076 8434
rect 9036 8084 9088 8090
rect 9036 8026 9088 8032
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8864 6322 8892 7822
rect 9048 7546 9076 8026
rect 9036 7540 9088 7546
rect 9036 7482 9088 7488
rect 9048 7206 9076 7482
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8852 6316 8904 6322
rect 8852 6258 8904 6264
rect 8956 6186 8984 7142
rect 9048 6322 9076 7142
rect 9036 6316 9088 6322
rect 9036 6258 9088 6264
rect 8944 6180 8996 6186
rect 8944 6122 8996 6128
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8680 5766 8800 5794
rect 8772 5710 8800 5766
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5704 8812 5710
rect 8588 5642 8708 5658
rect 8760 5646 8812 5652
rect 8588 5636 8720 5642
rect 8588 5630 8668 5636
rect 8668 5578 8720 5584
rect 8772 4214 8800 5646
rect 8864 4486 8892 5714
rect 8956 5574 8984 6122
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 4758 8984 5170
rect 8944 4752 8996 4758
rect 8944 4694 8996 4700
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8576 3528 8628 3534
rect 8576 3470 8628 3476
rect 8588 2650 8616 3470
rect 9140 2854 9168 10542
rect 9416 10266 9444 10542
rect 9508 10266 9536 10678
rect 9600 10606 9628 11630
rect 9968 11354 9996 13874
rect 10152 12646 10180 15506
rect 10244 14074 10272 21082
rect 11256 20602 11284 21354
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11244 20596 11296 20602
rect 11244 20538 11296 20544
rect 11532 20466 11560 21082
rect 11520 20460 11572 20466
rect 11520 20402 11572 20408
rect 11624 20346 11652 21286
rect 11808 20942 11836 21422
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11532 20318 11652 20346
rect 11532 20262 11560 20318
rect 10784 20256 10836 20262
rect 10784 20198 10836 20204
rect 11520 20256 11572 20262
rect 11520 20198 11572 20204
rect 10796 19922 10824 20198
rect 10784 19916 10836 19922
rect 10784 19858 10836 19864
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11440 19514 11468 19790
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10796 18426 10824 18702
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 11440 16998 11468 19450
rect 11532 18834 11560 20198
rect 11808 19854 11836 20470
rect 11900 19854 11928 20538
rect 11992 20534 12020 21422
rect 12164 21412 12216 21418
rect 12164 21354 12216 21360
rect 12176 21078 12204 21354
rect 12268 21146 12296 21830
rect 12348 21548 12400 21554
rect 12348 21490 12400 21496
rect 12256 21140 12308 21146
rect 12256 21082 12308 21088
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12360 20890 12388 21490
rect 12452 21434 12480 22102
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12544 21690 12572 21966
rect 12624 21956 12676 21962
rect 12624 21898 12676 21904
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12636 21622 12664 21898
rect 12624 21616 12676 21622
rect 12624 21558 12676 21564
rect 12452 21418 12572 21434
rect 12452 21412 12584 21418
rect 12452 21406 12532 21412
rect 12532 21354 12584 21360
rect 12820 21078 12848 22510
rect 13004 22030 13032 22986
rect 12992 22024 13044 22030
rect 12992 21966 13044 21972
rect 13096 21622 13124 23054
rect 13832 22030 13860 23666
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 13820 22024 13872 22030
rect 13820 21966 13872 21972
rect 13360 21956 13412 21962
rect 13360 21898 13412 21904
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13084 21616 13136 21622
rect 13084 21558 13136 21564
rect 13280 21486 13308 21830
rect 13268 21480 13320 21486
rect 13268 21422 13320 21428
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12912 21146 12940 21354
rect 13372 21350 13400 21898
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13360 21344 13412 21350
rect 13360 21286 13412 21292
rect 13464 21146 13492 21490
rect 14188 21412 14240 21418
rect 14188 21354 14240 21360
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13452 21140 13504 21146
rect 13452 21082 13504 21088
rect 12808 21072 12860 21078
rect 12808 21014 12860 21020
rect 11980 20528 12032 20534
rect 11980 20470 12032 20476
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11624 17134 11652 19450
rect 11716 19378 11744 19654
rect 11992 19514 12020 20198
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11704 19372 11756 19378
rect 11704 19314 11756 19320
rect 11716 17202 11744 19314
rect 12084 19310 12112 19926
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 11888 18624 11940 18630
rect 11940 18584 12020 18612
rect 11888 18566 11940 18572
rect 11794 18456 11850 18465
rect 11794 18391 11850 18400
rect 11808 18358 11836 18391
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17610 11928 18022
rect 11888 17604 11940 17610
rect 11888 17546 11940 17552
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11612 17128 11664 17134
rect 11612 17070 11664 17076
rect 11428 16992 11480 16998
rect 11428 16934 11480 16940
rect 11624 16674 11652 17070
rect 11532 16646 11652 16674
rect 11532 16590 11560 16646
rect 11520 16584 11572 16590
rect 11520 16526 11572 16532
rect 11704 16584 11756 16590
rect 11704 16526 11756 16532
rect 11612 16448 11664 16454
rect 11612 16390 11664 16396
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10244 13326 10272 14010
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10060 11898 10088 12174
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 10060 11218 10088 11834
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10244 10606 10272 12786
rect 10336 12442 10364 15302
rect 11244 15020 11296 15026
rect 11244 14962 11296 14968
rect 11256 14414 11284 14962
rect 11624 14414 11652 16390
rect 11716 16114 11744 16526
rect 11808 16250 11836 17138
rect 11796 16244 11848 16250
rect 11796 16186 11848 16192
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11716 15434 11744 16050
rect 11704 15428 11756 15434
rect 11704 15370 11756 15376
rect 11900 15026 11928 17546
rect 11992 16590 12020 18584
rect 12084 18290 12112 18702
rect 12176 18698 12204 20878
rect 12360 20862 12480 20890
rect 12452 20806 12480 20862
rect 12256 20800 12308 20806
rect 12256 20742 12308 20748
rect 12440 20800 12492 20806
rect 12440 20742 12492 20748
rect 12268 20466 12296 20742
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12268 19378 12296 20402
rect 12256 19372 12308 19378
rect 12256 19314 12308 19320
rect 12268 18970 12296 19314
rect 12532 19304 12584 19310
rect 13096 19281 13124 21082
rect 13544 21072 13596 21078
rect 13544 21014 13596 21020
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13188 20262 13216 20334
rect 13464 20262 13492 20402
rect 13176 20256 13228 20262
rect 13176 20198 13228 20204
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 12532 19246 12584 19252
rect 13082 19272 13138 19281
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12268 18822 12480 18850
rect 12164 18692 12216 18698
rect 12164 18634 12216 18640
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12268 18222 12296 18822
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12360 18086 12388 18702
rect 12452 18630 12480 18822
rect 12544 18766 12572 19246
rect 12992 19236 13044 19242
rect 13082 19207 13138 19216
rect 12992 19178 13044 19184
rect 13004 18766 13032 19178
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12992 18760 13044 18766
rect 12992 18702 13044 18708
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12544 18290 12572 18702
rect 12900 18692 12952 18698
rect 12900 18634 12952 18640
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12348 18080 12400 18086
rect 12348 18022 12400 18028
rect 12164 17740 12216 17746
rect 12164 17682 12216 17688
rect 12176 17338 12204 17682
rect 12452 17542 12480 18226
rect 12544 17610 12572 18226
rect 12820 18086 12848 18226
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12532 17604 12584 17610
rect 12584 17564 12664 17592
rect 12532 17546 12584 17552
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12176 17202 12204 17274
rect 12348 17264 12400 17270
rect 12348 17206 12400 17212
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11888 14884 11940 14890
rect 11888 14826 11940 14832
rect 11900 14550 11928 14826
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11256 13938 11284 14350
rect 11900 14074 11928 14486
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11704 14000 11756 14006
rect 11704 13942 11756 13948
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 11256 13394 11284 13874
rect 11244 13388 11296 13394
rect 11244 13330 11296 13336
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11830 10456 12038
rect 10416 11824 10468 11830
rect 10416 11766 10468 11772
rect 10520 11218 10548 12582
rect 11348 11762 11376 12718
rect 11532 12170 11560 13262
rect 11612 12232 11664 12238
rect 11612 12174 11664 12180
rect 11520 12164 11572 12170
rect 11520 12106 11572 12112
rect 11624 11762 11652 12174
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11612 11756 11664 11762
rect 11716 11744 11744 13942
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13258 11836 13670
rect 11796 13252 11848 13258
rect 11796 13194 11848 13200
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11900 12986 11928 13126
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 12306 12020 16526
rect 12084 15910 12112 16730
rect 12176 16590 12204 16934
rect 12360 16794 12388 17206
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12544 16590 12572 17138
rect 12164 16584 12216 16590
rect 12532 16584 12584 16590
rect 12164 16526 12216 16532
rect 12452 16544 12532 16572
rect 12256 16244 12308 16250
rect 12256 16186 12308 16192
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12084 15706 12112 15846
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12268 15434 12296 16186
rect 12452 15978 12480 16544
rect 12532 16526 12584 16532
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12544 16250 12572 16390
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12440 15972 12492 15978
rect 12440 15914 12492 15920
rect 12438 15872 12494 15881
rect 12360 15830 12438 15858
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12162 13968 12218 13977
rect 12162 13903 12164 13912
rect 12216 13903 12218 13912
rect 12164 13874 12216 13880
rect 12268 13841 12296 14350
rect 12254 13832 12310 13841
rect 12254 13767 12310 13776
rect 12072 13388 12124 13394
rect 12072 13330 12124 13336
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 12084 12238 12112 13330
rect 12164 12844 12216 12850
rect 12164 12786 12216 12792
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11796 12096 11848 12102
rect 11796 12038 11848 12044
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11808 11898 11836 12038
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11900 11830 11928 12038
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11796 11756 11848 11762
rect 11716 11716 11796 11744
rect 11612 11698 11664 11704
rect 11796 11698 11848 11704
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 10508 11008 10560 11014
rect 10508 10950 10560 10956
rect 10520 10606 10548 10950
rect 9588 10600 9640 10606
rect 9588 10542 9640 10548
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9232 9586 9260 9930
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 9232 8498 9260 9522
rect 9600 9382 9628 10542
rect 10140 9988 10192 9994
rect 10140 9930 10192 9936
rect 10152 9722 10180 9930
rect 10140 9716 10192 9722
rect 10140 9658 10192 9664
rect 10244 9450 10272 10542
rect 10520 10266 10548 10542
rect 10600 10464 10652 10470
rect 10600 10406 10652 10412
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10612 9722 10640 10406
rect 11348 10266 11376 11086
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10704 9722 10732 9998
rect 10876 9920 10928 9926
rect 10876 9862 10928 9868
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10692 9716 10744 9722
rect 10692 9658 10744 9664
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9600 8566 9628 8978
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9324 7478 9352 7686
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9416 6322 9444 7482
rect 9508 7002 9536 7754
rect 9692 7750 9720 8842
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9784 7886 9812 8434
rect 9876 8362 9904 8774
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9876 7410 9904 8298
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 10152 7342 10180 7754
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9588 6384 9640 6390
rect 9588 6326 9640 6332
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9600 5710 9628 6326
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9876 5914 9904 6258
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9588 5704 9640 5710
rect 9588 5646 9640 5652
rect 9232 5234 9260 5646
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9600 5114 9628 5646
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9232 5086 9628 5114
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9232 4622 9260 5086
rect 9588 5024 9640 5030
rect 9508 4972 9588 4978
rect 9508 4966 9640 4972
rect 9508 4950 9628 4966
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9508 4486 9536 4950
rect 9692 4842 9720 5102
rect 9600 4814 9720 4842
rect 9600 4486 9628 4814
rect 9680 4548 9732 4554
rect 9680 4490 9732 4496
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9588 4480 9640 4486
rect 9588 4422 9640 4428
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8576 2644 8628 2650
rect 8576 2586 8628 2592
rect 9508 2514 9536 4422
rect 9600 4214 9628 4422
rect 9692 4282 9720 4490
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9600 3534 9628 4150
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9692 3534 9720 3946
rect 9784 3534 9812 4014
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9600 3058 9628 3334
rect 9876 3194 9904 3470
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9968 2446 9996 5578
rect 10060 4146 10088 6598
rect 10152 6118 10180 7278
rect 10520 7206 10548 8366
rect 10612 7274 10640 9454
rect 10888 9178 10916 9862
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11072 8974 11100 9114
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11428 8968 11480 8974
rect 11428 8910 11480 8916
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8498 11008 8842
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 10704 8090 10732 8434
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10704 7342 10732 8026
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7410 10916 7686
rect 10980 7410 11008 8434
rect 11336 7540 11388 7546
rect 11336 7482 11388 7488
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10600 7268 10652 7274
rect 10600 7210 10652 7216
rect 10508 7200 10560 7206
rect 10508 7142 10560 7148
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10152 5778 10180 6054
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10152 5302 10180 5714
rect 10244 5642 10272 6054
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10060 3738 10088 4082
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 3398 10088 3674
rect 10152 3534 10180 5238
rect 10428 5098 10456 5578
rect 10520 5574 10548 7142
rect 10888 6866 10916 7346
rect 10876 6860 10928 6866
rect 10876 6802 10928 6808
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10520 5216 10548 5510
rect 10600 5228 10652 5234
rect 10520 5188 10600 5216
rect 10600 5170 10652 5176
rect 10416 5092 10468 5098
rect 10416 5034 10468 5040
rect 10612 4146 10640 5170
rect 10980 5098 11008 7346
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 5710 11100 7142
rect 11152 6724 11204 6730
rect 11152 6666 11204 6672
rect 11164 6458 11192 6666
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11256 6322 11284 6598
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11244 5704 11296 5710
rect 11244 5646 11296 5652
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5234 11100 5510
rect 11256 5234 11284 5646
rect 11348 5370 11376 7482
rect 11440 6118 11468 8910
rect 11532 7970 11560 11222
rect 11624 10606 11652 11698
rect 11808 11354 11836 11698
rect 11992 11642 12020 12106
rect 12176 11762 12204 12786
rect 12360 12782 12388 15830
rect 12438 15807 12494 15816
rect 12636 15586 12664 17564
rect 12912 17338 12940 18634
rect 13004 18290 13032 18702
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 17882 13032 18226
rect 13096 18222 13124 19207
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 12900 17332 12952 17338
rect 12820 17292 12900 17320
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12544 15558 12664 15586
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12452 15094 12480 15302
rect 12544 15162 12572 15558
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12636 15026 12664 15438
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12728 14958 12756 16186
rect 12820 15026 12848 17292
rect 12900 17274 12952 17280
rect 13004 17202 13032 17614
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 13004 16590 13032 17138
rect 13096 16658 13124 18158
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13004 16182 13032 16526
rect 12992 16176 13044 16182
rect 12992 16118 13044 16124
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12532 14952 12584 14958
rect 12452 14912 12532 14940
rect 12452 14074 12480 14912
rect 12532 14894 12584 14900
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12820 14804 12848 14962
rect 12636 14776 12848 14804
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12544 14346 12572 14418
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12544 14074 12572 14282
rect 12636 14074 12664 14776
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 12532 14068 12584 14074
rect 12532 14010 12584 14016
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12440 13932 12492 13938
rect 12492 13892 12664 13920
rect 12440 13874 12492 13880
rect 12532 13796 12584 13802
rect 12532 13738 12584 13744
rect 12544 13326 12572 13738
rect 12636 13326 12664 13892
rect 12532 13320 12584 13326
rect 12532 13262 12584 13268
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 12850 12664 13262
rect 12728 13258 12756 14418
rect 12912 14414 12940 15982
rect 12992 15904 13044 15910
rect 12990 15872 12992 15881
rect 13044 15872 13046 15881
rect 12990 15807 13046 15816
rect 13188 15638 13216 20198
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13372 19514 13400 19722
rect 13464 19718 13492 19858
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13280 18902 13308 19314
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13372 18970 13400 19246
rect 13464 18970 13492 19654
rect 13556 19378 13584 21014
rect 14200 20942 14228 21354
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13648 19378 13676 20538
rect 13832 20466 13860 20742
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13740 19514 13768 20402
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13832 19922 13860 20198
rect 13912 19984 13964 19990
rect 13912 19926 13964 19932
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13728 19508 13780 19514
rect 13728 19450 13780 19456
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13268 18896 13320 18902
rect 13268 18838 13320 18844
rect 13280 17134 13308 18838
rect 13360 18760 13412 18766
rect 13360 18702 13412 18708
rect 13372 17338 13400 18702
rect 13556 18465 13584 19178
rect 13740 18630 13768 19178
rect 13728 18624 13780 18630
rect 13728 18566 13780 18572
rect 13542 18456 13598 18465
rect 13542 18391 13598 18400
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13268 16992 13320 16998
rect 13268 16934 13320 16940
rect 13280 16250 13308 16934
rect 13372 16590 13400 17274
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13268 16244 13320 16250
rect 13268 16186 13320 16192
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13176 15632 13228 15638
rect 13176 15574 13228 15580
rect 13188 15502 13216 15574
rect 13176 15496 13228 15502
rect 13176 15438 13228 15444
rect 13174 15192 13230 15201
rect 13084 15156 13136 15162
rect 13174 15127 13230 15136
rect 13084 15098 13136 15104
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 12900 14408 12952 14414
rect 12820 14368 12900 14396
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12348 12776 12400 12782
rect 12348 12718 12400 12724
rect 12820 12714 12848 14368
rect 12900 14350 12952 14356
rect 12898 13832 12954 13841
rect 12898 13767 12954 13776
rect 12912 13734 12940 13767
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12912 12850 12940 13398
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12808 12708 12860 12714
rect 12808 12650 12860 12656
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 11900 11614 12020 11642
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11808 11150 11836 11290
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11612 10600 11664 10606
rect 11612 10542 11664 10548
rect 11716 10062 11744 10950
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11704 8900 11756 8906
rect 11704 8842 11756 8848
rect 11716 8498 11744 8842
rect 11900 8566 11928 11614
rect 12440 11552 12492 11558
rect 11978 11520 12034 11529
rect 12440 11494 12492 11500
rect 11978 11455 12034 11464
rect 11992 11218 12020 11455
rect 11980 11212 12032 11218
rect 11980 11154 12032 11160
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12256 11144 12308 11150
rect 12452 11098 12480 11494
rect 12544 11150 12572 12242
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 12636 11150 12664 11834
rect 12308 11092 12480 11098
rect 12256 11086 12480 11092
rect 12532 11144 12584 11150
rect 12532 11086 12584 11092
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11992 10538 12020 11018
rect 12176 10810 12204 11086
rect 12268 11070 12480 11086
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12164 10804 12216 10810
rect 12164 10746 12216 10752
rect 12268 10674 12296 10950
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 11980 10532 12032 10538
rect 11980 10474 12032 10480
rect 12452 10470 12480 11070
rect 12728 11014 12756 11086
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12636 10606 12664 10950
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12624 10600 12676 10606
rect 12624 10542 12676 10548
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12728 9994 12756 10678
rect 12820 10674 12848 12650
rect 13004 12646 13032 14554
rect 13096 14482 13124 15098
rect 13188 15094 13216 15127
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13280 14890 13308 14962
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13372 14414 13400 15914
rect 13464 14414 13492 17070
rect 13556 16998 13584 18391
rect 13740 18290 13768 18566
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13832 18222 13860 19858
rect 13924 19242 13952 19926
rect 14292 19360 14320 22374
rect 16132 22234 16160 22578
rect 16394 22536 16450 22545
rect 16394 22471 16396 22480
rect 16448 22471 16450 22480
rect 16396 22442 16448 22448
rect 16120 22228 16172 22234
rect 16120 22170 16172 22176
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 16120 22024 16172 22030
rect 16120 21966 16172 21972
rect 14384 21554 14412 21966
rect 14372 21548 14424 21554
rect 14372 21490 14424 21496
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14660 21146 14688 21490
rect 15948 21486 15976 21966
rect 15936 21480 15988 21486
rect 15936 21422 15988 21428
rect 15844 21344 15896 21350
rect 15844 21286 15896 21292
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 14372 19372 14424 19378
rect 14200 19332 14372 19360
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 13912 19236 13964 19242
rect 13912 19178 13964 19184
rect 14004 19168 14056 19174
rect 14004 19110 14056 19116
rect 14016 18902 14044 19110
rect 14108 18970 14136 19246
rect 14096 18964 14148 18970
rect 14096 18906 14148 18912
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 14004 18284 14056 18290
rect 14004 18226 14056 18232
rect 13820 18216 13872 18222
rect 13820 18158 13872 18164
rect 14016 18154 14044 18226
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 14016 17542 14044 18090
rect 14200 18086 14228 19332
rect 14372 19314 14424 19320
rect 14278 19272 14334 19281
rect 14278 19207 14334 19216
rect 14292 19174 14320 19207
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 14476 18834 14504 20266
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14280 18216 14332 18222
rect 14280 18158 14332 18164
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17678 14228 18022
rect 14292 17678 14320 18158
rect 14476 17746 14504 18226
rect 14464 17740 14516 17746
rect 14464 17682 14516 17688
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13556 15586 13584 16730
rect 14016 16726 14044 17478
rect 14292 17320 14320 17614
rect 14292 17292 14412 17320
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13636 16448 13688 16454
rect 13636 16390 13688 16396
rect 13648 15910 13676 16390
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13556 15558 13676 15586
rect 13648 15502 13676 15558
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13556 15201 13584 15438
rect 13542 15192 13598 15201
rect 13542 15127 13598 15136
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13084 14340 13136 14346
rect 13084 14282 13136 14288
rect 13096 13326 13124 14282
rect 13176 14272 13228 14278
rect 13176 14214 13228 14220
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13188 14074 13216 14214
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13188 13530 13216 13874
rect 13280 13870 13308 14214
rect 13268 13864 13320 13870
rect 13268 13806 13320 13812
rect 13176 13524 13228 13530
rect 13176 13466 13228 13472
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13188 12850 13216 13194
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12238 13032 12582
rect 13188 12306 13216 12786
rect 13176 12300 13228 12306
rect 13176 12242 13228 12248
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11529 13032 12174
rect 13188 11694 13216 12242
rect 13176 11688 13228 11694
rect 13176 11630 13228 11636
rect 13176 11552 13228 11558
rect 12990 11520 13046 11529
rect 13176 11494 13228 11500
rect 12990 11455 13046 11464
rect 12900 11348 12952 11354
rect 12900 11290 12952 11296
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12912 11150 12940 11290
rect 13004 11150 13032 11290
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12912 10810 12940 11086
rect 13096 11082 13124 11222
rect 13188 11150 13216 11494
rect 13280 11218 13308 13398
rect 13372 11830 13400 14350
rect 13556 14278 13584 14826
rect 13544 14272 13596 14278
rect 13464 14232 13544 14260
rect 13464 13977 13492 14232
rect 13544 14214 13596 14220
rect 13648 14090 13676 15438
rect 13740 14618 13768 16458
rect 13832 16182 13860 16594
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 13820 16176 13872 16182
rect 13820 16118 13872 16124
rect 13820 15632 13872 15638
rect 13924 15586 13952 16458
rect 13872 15580 13952 15586
rect 13820 15574 13952 15580
rect 13832 15558 13952 15574
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13832 14226 13860 14418
rect 13556 14062 13676 14090
rect 13740 14198 13860 14226
rect 13450 13968 13506 13977
rect 13450 13903 13506 13912
rect 13464 13394 13492 13903
rect 13556 13734 13584 14062
rect 13636 14000 13688 14006
rect 13740 13954 13768 14198
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13688 13948 13768 13954
rect 13636 13942 13768 13948
rect 13648 13926 13768 13942
rect 13636 13864 13688 13870
rect 13832 13852 13860 14010
rect 13924 13938 13952 15558
rect 14016 15042 14044 16662
rect 14200 15502 14228 17206
rect 14384 17202 14412 17292
rect 14476 17270 14504 17682
rect 14464 17264 14516 17270
rect 14464 17206 14516 17212
rect 14568 17202 14596 19790
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14936 19514 14964 19722
rect 14924 19508 14976 19514
rect 14924 19450 14976 19456
rect 14740 19236 14792 19242
rect 14740 19178 14792 19184
rect 14648 18624 14700 18630
rect 14648 18566 14700 18572
rect 14660 18426 14688 18566
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14292 16114 14320 17138
rect 14384 16504 14412 17138
rect 14384 16476 14504 16504
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14476 15502 14504 16476
rect 14568 15570 14596 17138
rect 14752 16590 14780 19178
rect 15028 18426 15056 20742
rect 15396 20602 15424 20946
rect 15856 20942 15884 21286
rect 16132 21146 16160 21966
rect 16396 21888 16448 21894
rect 16394 21856 16396 21865
rect 16448 21856 16450 21865
rect 16394 21791 16450 21800
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15948 20398 15976 20878
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15292 20256 15344 20262
rect 15292 20198 15344 20204
rect 15304 19514 15332 20198
rect 15948 20058 15976 20334
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 15488 19310 15516 19654
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15396 18970 15424 19246
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 14832 17672 14884 17678
rect 14832 17614 14884 17620
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14108 15162 14136 15438
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14016 15026 14136 15042
rect 14016 15020 14148 15026
rect 14016 15014 14096 15020
rect 14096 14962 14148 14968
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13688 13824 13860 13852
rect 13636 13806 13688 13812
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13556 13530 13584 13670
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13452 13388 13504 13394
rect 13452 13330 13504 13336
rect 13832 12850 13860 13398
rect 13924 12918 13952 13874
rect 14016 13530 14044 13874
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14108 13410 14136 14962
rect 14200 14482 14228 15438
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14016 13382 14136 13410
rect 13912 12912 13964 12918
rect 13912 12854 13964 12860
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13740 12714 13768 12786
rect 13728 12708 13780 12714
rect 13728 12650 13780 12656
rect 13832 12434 13860 12786
rect 13924 12714 13952 12854
rect 13912 12708 13964 12714
rect 13912 12650 13964 12656
rect 13740 12406 13860 12434
rect 13360 11824 13412 11830
rect 13360 11766 13412 11772
rect 13268 11212 13320 11218
rect 13372 11200 13400 11766
rect 13544 11212 13596 11218
rect 13372 11172 13544 11200
rect 13268 11154 13320 11160
rect 13544 11154 13596 11160
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13084 11076 13136 11082
rect 13084 11018 13136 11024
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12808 10668 12860 10674
rect 12912 10656 12940 10746
rect 13280 10742 13308 11154
rect 13740 11150 13768 12406
rect 13820 12300 13872 12306
rect 13820 12242 13872 12248
rect 13832 11762 13860 12242
rect 14016 12238 14044 13382
rect 14200 13258 14228 14418
rect 14292 13938 14320 15302
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14292 13462 14320 13874
rect 14384 13870 14412 14894
rect 14476 14074 14504 15438
rect 14568 14482 14596 15506
rect 14752 15434 14780 16526
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14476 13394 14504 14010
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 14200 13138 14228 13194
rect 14108 13110 14228 13138
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13912 11620 13964 11626
rect 13912 11562 13964 11568
rect 13924 11354 13952 11562
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13648 11014 13676 11086
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 12992 10668 13044 10674
rect 12912 10628 12992 10656
rect 12808 10610 12860 10616
rect 12992 10610 13044 10616
rect 13544 10464 13596 10470
rect 13544 10406 13596 10412
rect 13556 10062 13584 10406
rect 13648 10198 13676 10950
rect 13740 10674 13768 11086
rect 13832 10826 13860 11290
rect 13832 10798 13952 10826
rect 14016 10810 14044 11698
rect 14108 11132 14136 13110
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14200 12442 14228 12786
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14292 11898 14320 13262
rect 14372 13252 14424 13258
rect 14372 13194 14424 13200
rect 14384 12918 14412 13194
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14476 12832 14504 13330
rect 14556 12844 14608 12850
rect 14476 12804 14556 12832
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14280 11892 14332 11898
rect 14280 11834 14332 11840
rect 14188 11144 14240 11150
rect 14108 11104 14188 11132
rect 14188 11086 14240 11092
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13636 10192 13688 10198
rect 13636 10134 13688 10140
rect 13832 10062 13860 10678
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 12716 9988 12768 9994
rect 12716 9930 12768 9936
rect 13924 9654 13952 10798
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 14384 10742 14412 12174
rect 14476 11150 14504 12804
rect 14556 12786 14608 12792
rect 14556 12708 14608 12714
rect 14556 12650 14608 12656
rect 14568 11558 14596 12650
rect 14660 11762 14688 14282
rect 14752 12850 14780 14418
rect 14844 14278 14872 17614
rect 15844 17536 15896 17542
rect 15844 17478 15896 17484
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15028 16794 15056 17138
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15016 16788 15068 16794
rect 15016 16730 15068 16736
rect 15396 16522 15424 16934
rect 15856 16590 15884 17478
rect 16408 17338 16436 17614
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 15948 16590 15976 17274
rect 16212 17196 16264 17202
rect 16212 17138 16264 17144
rect 16224 16794 16252 17138
rect 16394 17096 16450 17105
rect 16394 17031 16396 17040
rect 16448 17031 16450 17040
rect 16396 17002 16448 17008
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15384 16516 15436 16522
rect 15384 16458 15436 16464
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15660 15700 15712 15706
rect 15660 15642 15712 15648
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15120 15162 15148 15370
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15580 15094 15608 15302
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15672 14958 15700 15642
rect 15764 15502 15792 15846
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15856 15162 15884 15846
rect 16132 15706 16160 16050
rect 16394 15736 16450 15745
rect 16120 15700 16172 15706
rect 16394 15671 16396 15680
rect 16120 15642 16172 15648
rect 16448 15671 16450 15680
rect 16396 15642 16448 15648
rect 15844 15156 15896 15162
rect 15844 15098 15896 15104
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 16132 14618 16160 14962
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16120 14612 16172 14618
rect 16120 14554 16172 14560
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 15028 14074 15056 14282
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15016 13252 15068 13258
rect 15016 13194 15068 13200
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14752 12306 14780 12786
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14464 10600 14516 10606
rect 14568 10588 14596 11494
rect 14752 11218 14780 12242
rect 14740 11212 14792 11218
rect 14660 11172 14740 11200
rect 14660 10674 14688 11172
rect 14740 11154 14792 11160
rect 14648 10668 14700 10674
rect 14648 10610 14700 10616
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14516 10560 14596 10588
rect 14464 10542 14516 10548
rect 14660 10198 14688 10610
rect 14844 10266 14872 10610
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14648 10192 14700 10198
rect 14648 10134 14700 10140
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13912 9648 13964 9654
rect 13912 9590 13964 9596
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12820 8974 12848 9114
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12532 8968 12584 8974
rect 12808 8968 12860 8974
rect 12584 8928 12664 8956
rect 12532 8910 12584 8916
rect 12176 8838 12204 8910
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 11888 8560 11940 8566
rect 11888 8502 11940 8508
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11532 7942 11652 7970
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 11532 7546 11560 7754
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11060 5228 11112 5234
rect 11060 5170 11112 5176
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10232 3936 10284 3942
rect 10232 3878 10284 3884
rect 10244 3534 10272 3878
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10152 3126 10180 3470
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10980 2922 11008 3334
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 11072 2378 11100 5170
rect 11256 4146 11284 5170
rect 11624 4282 11652 7942
rect 11900 7886 11928 8366
rect 12176 7886 12204 8774
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12176 7410 12204 7822
rect 12268 7478 12296 8434
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 12164 7404 12216 7410
rect 12164 7346 12216 7352
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 11808 7206 11836 7346
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11808 6798 11836 7142
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11900 5234 11928 6394
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5302 12020 5646
rect 11980 5296 12032 5302
rect 11980 5238 12032 5244
rect 11888 5228 11940 5234
rect 11716 5188 11888 5216
rect 11612 4276 11664 4282
rect 11612 4218 11664 4224
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11256 3126 11284 4082
rect 11624 4078 11652 4218
rect 11716 4146 11744 5188
rect 11888 5170 11940 5176
rect 12072 5228 12124 5234
rect 12072 5170 12124 5176
rect 12084 5114 12112 5170
rect 11900 5098 12112 5114
rect 11888 5092 12112 5098
rect 11940 5086 12112 5092
rect 11888 5034 11940 5040
rect 11900 4146 11928 5034
rect 12176 4622 12204 7346
rect 12360 7274 12388 7346
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12360 5930 12388 6326
rect 12452 5930 12480 7754
rect 12636 7750 12664 8928
rect 12728 8928 12808 8956
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12636 7410 12664 7686
rect 12728 7478 12756 8928
rect 12808 8910 12860 8916
rect 13280 8906 13308 8978
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 13268 8900 13320 8906
rect 13268 8842 13320 8848
rect 13452 8900 13504 8906
rect 13452 8842 13504 8848
rect 12912 8242 12940 8842
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12912 8214 13032 8242
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7750 12848 7822
rect 12808 7744 12860 7750
rect 12808 7686 12860 7692
rect 12716 7472 12768 7478
rect 12716 7414 12768 7420
rect 12912 7410 12940 8026
rect 13004 7886 13032 8214
rect 13096 7954 13124 8774
rect 13280 8634 13308 8842
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13188 8090 13216 8434
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13360 7744 13412 7750
rect 13464 7732 13492 8842
rect 13412 7704 13492 7732
rect 13360 7686 13412 7692
rect 12624 7404 12676 7410
rect 12900 7404 12952 7410
rect 12624 7346 12676 7352
rect 12820 7364 12900 7392
rect 12360 5902 12480 5930
rect 12440 5568 12492 5574
rect 12440 5510 12492 5516
rect 12348 5364 12400 5370
rect 12348 5306 12400 5312
rect 12360 5098 12388 5306
rect 12452 5234 12480 5510
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12164 4616 12216 4622
rect 12164 4558 12216 4564
rect 11704 4140 11756 4146
rect 11888 4140 11940 4146
rect 11704 4082 11756 4088
rect 11808 4100 11888 4128
rect 11612 4072 11664 4078
rect 11518 4040 11574 4049
rect 11612 4014 11664 4020
rect 11518 3975 11520 3984
rect 11572 3975 11574 3984
rect 11520 3946 11572 3952
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11716 3058 11744 4082
rect 11808 3108 11836 4100
rect 11888 4082 11940 4088
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3466 11928 3878
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 11992 3398 12020 4082
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11888 3120 11940 3126
rect 11808 3080 11888 3108
rect 11888 3062 11940 3068
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11428 2984 11480 2990
rect 11428 2926 11480 2932
rect 11440 2446 11468 2926
rect 11992 2446 12020 3334
rect 12268 2514 12296 4014
rect 12532 4004 12584 4010
rect 12360 3964 12532 3992
rect 12360 3738 12388 3964
rect 12532 3946 12584 3952
rect 12348 3732 12400 3738
rect 12348 3674 12400 3680
rect 12440 3528 12492 3534
rect 12440 3470 12492 3476
rect 12452 2990 12480 3470
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12256 2508 12308 2514
rect 12256 2450 12308 2456
rect 12636 2446 12664 7346
rect 12820 6254 12848 7364
rect 12900 7346 12952 7352
rect 13096 7342 13124 7686
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12900 7200 12952 7206
rect 13096 7188 13124 7278
rect 13464 7206 13492 7704
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 12952 7160 13124 7188
rect 13452 7200 13504 7206
rect 12900 7142 12952 7148
rect 13452 7142 13504 7148
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12808 5296 12860 5302
rect 12912 5284 12940 7142
rect 13360 6928 13412 6934
rect 13360 6870 13412 6876
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13280 6254 13308 6598
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13084 5704 13136 5710
rect 13084 5646 13136 5652
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 13004 5370 13032 5578
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 13096 5302 13124 5646
rect 12860 5256 12940 5284
rect 13084 5296 13136 5302
rect 12808 5238 12860 5244
rect 13084 5238 13136 5244
rect 12820 4282 12848 5238
rect 13280 4690 13308 6190
rect 13268 4684 13320 4690
rect 13268 4626 13320 4632
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13096 3738 13124 4082
rect 13084 3732 13136 3738
rect 13004 3692 13084 3720
rect 13004 3194 13032 3692
rect 13084 3674 13136 3680
rect 13280 3602 13308 4626
rect 13372 3738 13400 6870
rect 13464 6730 13492 7142
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13464 5642 13492 6666
rect 13556 6390 13584 7346
rect 13544 6384 13596 6390
rect 13544 6326 13596 6332
rect 13910 6352 13966 6361
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13464 4214 13492 5578
rect 13556 4214 13584 6326
rect 13910 6287 13912 6296
rect 13964 6287 13966 6296
rect 13912 6258 13964 6264
rect 14016 6186 14044 9658
rect 14108 9586 14136 9862
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 14108 7886 14136 8502
rect 14292 8090 14320 8910
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14292 6798 14320 7346
rect 14384 7342 14412 8910
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14476 7274 14504 8910
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 7818 14780 8774
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14936 7410 14964 12786
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 14924 7404 14976 7410
rect 14924 7346 14976 7352
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14660 7002 14688 7346
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14936 6866 14964 7346
rect 14924 6860 14976 6866
rect 14924 6802 14976 6808
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 13820 6180 13872 6186
rect 13820 6122 13872 6128
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 13832 4604 13860 6122
rect 14292 5250 14320 6734
rect 14372 6724 14424 6730
rect 14372 6666 14424 6672
rect 14384 6390 14412 6666
rect 14476 6458 14504 6734
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14830 6352 14886 6361
rect 14464 6316 14516 6322
rect 14464 6258 14516 6264
rect 14648 6316 14700 6322
rect 14830 6287 14832 6296
rect 14648 6258 14700 6264
rect 14884 6287 14886 6296
rect 14832 6258 14884 6264
rect 14476 6186 14504 6258
rect 14464 6180 14516 6186
rect 14464 6122 14516 6128
rect 14660 6118 14688 6258
rect 14924 6180 14976 6186
rect 14924 6122 14976 6128
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14384 5370 14412 5578
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14188 5228 14240 5234
rect 14292 5222 14504 5250
rect 14188 5170 14240 5176
rect 14108 4826 14136 5170
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13912 4616 13964 4622
rect 13832 4576 13912 4604
rect 13912 4558 13964 4564
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13544 4208 13596 4214
rect 13544 4150 13596 4156
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13268 3596 13320 3602
rect 13268 3538 13320 3544
rect 13372 3534 13400 3674
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 12992 3188 13044 3194
rect 12992 3130 13044 3136
rect 13004 2446 13032 3130
rect 13096 3058 13124 3334
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13464 2774 13492 4150
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13832 3602 13860 4082
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 3194 13584 3470
rect 13544 3188 13596 3194
rect 13544 3130 13596 3136
rect 13924 3058 13952 4558
rect 14108 4282 14136 4626
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14108 3942 14136 4218
rect 14200 4146 14228 5170
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14292 4282 14320 4558
rect 14384 4282 14412 4558
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14372 4276 14424 4282
rect 14372 4218 14424 4224
rect 14476 4146 14504 5222
rect 14568 4622 14596 5510
rect 14660 5166 14688 6054
rect 14936 5234 14964 6122
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14648 5160 14700 5166
rect 15028 5114 15056 13194
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15844 13184 15896 13190
rect 15844 13126 15896 13132
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15212 12442 15240 12854
rect 15200 12436 15252 12442
rect 15200 12378 15252 12384
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11150 15148 11494
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15212 8634 15240 10610
rect 15396 10130 15424 13126
rect 15580 13025 15608 13126
rect 15566 13016 15622 13025
rect 15566 12951 15622 12960
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15580 12306 15608 12582
rect 15764 12306 15792 12922
rect 15568 12300 15620 12306
rect 15568 12242 15620 12248
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15856 12170 15884 13126
rect 15844 12164 15896 12170
rect 15844 12106 15896 12112
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15488 11898 15516 12038
rect 15948 11898 15976 13262
rect 16040 12714 16068 14350
rect 16132 13938 16160 14554
rect 16224 14414 16252 14758
rect 16212 14408 16264 14414
rect 16212 14350 16264 14356
rect 16394 14376 16450 14385
rect 16394 14311 16450 14320
rect 16408 14278 16436 14311
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16486 13696 16542 13705
rect 16486 13631 16542 13640
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16408 12986 16436 13262
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15580 11354 15608 11630
rect 16040 11354 16068 12174
rect 16132 11762 16160 12922
rect 16500 12850 16528 13631
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16396 12368 16448 12374
rect 16394 12336 16396 12345
rect 16448 12336 16450 12345
rect 16394 12271 16450 12280
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15936 10464 15988 10470
rect 15936 10406 15988 10412
rect 15488 10130 15516 10406
rect 15948 10130 15976 10406
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 15476 10124 15528 10130
rect 15476 10066 15528 10072
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 16224 9450 16252 11698
rect 16316 11354 16344 12174
rect 16394 11656 16450 11665
rect 16394 11591 16396 11600
rect 16448 11591 16450 11600
rect 16396 11562 16448 11568
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16408 10305 16436 10406
rect 16394 10296 16450 10305
rect 16394 10231 16450 10240
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 16500 9586 16528 10066
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15120 6798 15148 7822
rect 15396 7410 15424 8842
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 16224 7750 16252 8434
rect 16580 8356 16632 8362
rect 16580 8298 16632 8304
rect 16592 8265 16620 8298
rect 16578 8256 16634 8265
rect 16578 8191 16634 8200
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15108 6792 15160 6798
rect 15108 6734 15160 6740
rect 15120 6254 15148 6734
rect 15396 6390 15424 7210
rect 15844 6656 15896 6662
rect 15844 6598 15896 6604
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15856 6322 15884 6598
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 5302 15148 6190
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 14648 5102 14700 5108
rect 14936 5086 15056 5114
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 4146 14596 4422
rect 14188 4140 14240 4146
rect 14188 4082 14240 4088
rect 14280 4140 14332 4146
rect 14464 4140 14516 4146
rect 14280 4082 14332 4088
rect 14384 4100 14464 4128
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 3398 14228 3470
rect 14188 3392 14240 3398
rect 14188 3334 14240 3340
rect 14292 3058 14320 4082
rect 14384 3670 14412 4100
rect 14464 4082 14516 4088
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14476 3534 14504 3878
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14556 3528 14608 3534
rect 14556 3470 14608 3476
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13280 2746 13492 2774
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13280 2378 13308 2746
rect 13924 2446 13952 2858
rect 14384 2650 14412 3470
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14476 2514 14504 3130
rect 14568 2854 14596 3470
rect 14660 3126 14688 4626
rect 14752 4622 14780 4966
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14752 3534 14780 4558
rect 14936 4214 14964 5086
rect 15016 5024 15068 5030
rect 15016 4966 15068 4972
rect 15028 4758 15056 4966
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 15120 4690 15148 5238
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 15120 4078 15148 4490
rect 15108 4072 15160 4078
rect 15108 4014 15160 4020
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 3398 14780 3470
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 14648 3120 14700 3126
rect 14648 3062 14700 3068
rect 14660 2990 14688 3062
rect 14936 3058 14964 3334
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14556 2848 14608 2854
rect 14556 2790 14608 2796
rect 14660 2514 14688 2926
rect 15120 2650 15148 3334
rect 15212 3058 15240 5782
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15568 5228 15620 5234
rect 15568 5170 15620 5176
rect 15580 4486 15608 5170
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 14464 2508 14516 2514
rect 14464 2450 14516 2456
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 15396 2446 15424 3334
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 6460 2372 6512 2378
rect 6460 2314 6512 2320
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 6472 800 6500 2314
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7748 2304 7800 2310
rect 7748 2246 7800 2252
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 7024 1034 7052 2246
rect 7024 1006 7144 1034
rect 7116 800 7144 1006
rect 7760 800 7788 2246
rect 8312 1170 8340 2246
rect 8312 1142 8432 1170
rect 8404 800 8432 1142
rect 9048 800 9076 2246
rect 9692 800 9720 2246
rect 10336 800 10364 2246
rect 10980 800 11008 2246
rect 11624 800 11652 2246
rect 12268 800 12296 2246
rect 12912 800 12940 2246
rect 13556 800 13584 2246
rect 14188 1352 14240 1358
rect 14188 1294 14240 1300
rect 14200 800 14228 1294
rect 14832 1148 14884 1154
rect 14832 1090 14884 1096
rect 14844 800 14872 1090
rect 15488 800 15516 3606
rect 15580 2378 15608 4082
rect 15672 3534 15700 5238
rect 15856 4146 15884 6258
rect 16224 5710 16252 6394
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16580 5568 16632 5574
rect 16578 5536 16580 5545
rect 16632 5536 16634 5545
rect 16578 5471 16634 5480
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16500 4146 16528 4422
rect 15844 4140 15896 4146
rect 15844 4082 15896 4088
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 17408 4072 17460 4078
rect 17408 4014 17460 4020
rect 16764 4004 16816 4010
rect 16764 3946 16816 3952
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15568 2372 15620 2378
rect 15568 2314 15620 2320
rect 15856 1154 15884 3334
rect 16040 3194 16068 3470
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15844 1148 15896 1154
rect 15844 1090 15896 1096
rect 16132 800 16160 3878
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 16316 1358 16344 2790
rect 16304 1352 16356 1358
rect 16304 1294 16356 1300
rect 16776 800 16804 3946
rect 17420 800 17448 4014
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
<< via2 >>
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 110 39072 166 39128
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 846 26732 848 26752
rect 848 26732 900 26752
rect 900 26732 902 26752
rect 846 26696 902 26732
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 7654 37868 7710 37904
rect 7654 37848 7656 37868
rect 7656 37848 7708 37868
rect 7708 37848 7710 37868
rect 8758 37868 8814 37904
rect 8758 37848 8760 37868
rect 8760 37848 8812 37868
rect 8812 37848 8814 37868
rect 10598 36116 10600 36136
rect 10600 36116 10652 36136
rect 10652 36116 10654 36136
rect 10598 36080 10654 36116
rect 11150 36116 11152 36136
rect 11152 36116 11204 36136
rect 11204 36116 11206 36136
rect 11150 36080 11206 36116
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 846 22636 902 22672
rect 846 22616 848 22636
rect 848 22616 900 22636
rect 900 22616 902 22636
rect 846 21972 848 21992
rect 848 21972 900 21992
rect 900 21972 902 21992
rect 846 21936 902 21972
rect 1306 21120 1362 21176
rect 846 19896 902 19952
rect 3054 20460 3110 20496
rect 3054 20440 3056 20460
rect 3056 20440 3108 20460
rect 3108 20440 3110 20460
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 1306 12980 1362 13016
rect 1306 12960 1308 12980
rect 1308 12960 1360 12980
rect 1360 12960 1362 12980
rect 846 12144 902 12200
rect 1122 11600 1178 11656
rect 1306 10240 1362 10296
rect 1030 9560 1086 9616
rect 1858 10920 1914 10976
rect 846 9052 848 9072
rect 848 9052 900 9072
rect 900 9052 902 9072
rect 846 9016 902 9052
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 2594 10684 2596 10704
rect 2596 10684 2648 10704
rect 2648 10684 2650 10704
rect 2594 10648 2650 10684
rect 2410 7248 2466 7304
rect 2778 10668 2834 10704
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 2778 10648 2829 10668
rect 2829 10648 2834 10668
rect 2778 8200 2834 8256
rect 2962 7520 3018 7576
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 3514 4140 3570 4176
rect 3514 4120 3516 4140
rect 3516 4120 3568 4140
rect 3568 4120 3570 4140
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 5170 8880 5226 8936
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 7194 12552 7250 12608
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4250 3576 4306 3632
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 6550 4156 6552 4176
rect 6552 4156 6604 4176
rect 6604 4156 6606 4176
rect 6550 4120 6606 4156
rect 7286 3576 7342 3632
rect 8390 7284 8392 7304
rect 8392 7284 8444 7304
rect 8444 7284 8446 7304
rect 8390 7248 8446 7284
rect 7838 4156 7840 4176
rect 7840 4156 7892 4176
rect 7892 4156 7894 4176
rect 7838 4120 7894 4156
rect 12438 34060 12494 34096
rect 12438 34040 12440 34060
rect 12440 34040 12492 34060
rect 12492 34040 12494 34060
rect 9310 27412 9312 27432
rect 9312 27412 9364 27432
rect 9364 27412 9366 27432
rect 9310 27376 9366 27412
rect 13082 34040 13138 34096
rect 12806 27376 12862 27432
rect 11794 18400 11850 18456
rect 13082 19216 13138 19272
rect 12162 13932 12218 13968
rect 12162 13912 12164 13932
rect 12164 13912 12216 13932
rect 12216 13912 12218 13932
rect 12254 13776 12310 13832
rect 12438 15816 12494 15872
rect 12990 15852 12992 15872
rect 12992 15852 13044 15872
rect 13044 15852 13046 15872
rect 12990 15816 13046 15852
rect 13542 18400 13598 18456
rect 13174 15136 13230 15192
rect 12898 13776 12954 13832
rect 11978 11464 12034 11520
rect 16394 22500 16450 22536
rect 16394 22480 16396 22500
rect 16396 22480 16448 22500
rect 16448 22480 16450 22500
rect 14278 19216 14334 19272
rect 13542 15136 13598 15192
rect 12990 11464 13046 11520
rect 13450 13912 13506 13968
rect 16394 21836 16396 21856
rect 16396 21836 16448 21856
rect 16448 21836 16450 21856
rect 16394 21800 16450 21836
rect 16394 17060 16450 17096
rect 16394 17040 16396 17060
rect 16396 17040 16448 17060
rect 16448 17040 16450 17060
rect 16394 15700 16450 15736
rect 16394 15680 16396 15700
rect 16396 15680 16448 15700
rect 16448 15680 16450 15700
rect 11518 4004 11574 4040
rect 11518 3984 11520 4004
rect 11520 3984 11572 4004
rect 11572 3984 11574 4004
rect 13910 6316 13966 6352
rect 13910 6296 13912 6316
rect 13912 6296 13964 6316
rect 13964 6296 13966 6316
rect 14830 6316 14886 6352
rect 14830 6296 14832 6316
rect 14832 6296 14884 6316
rect 14884 6296 14886 6316
rect 15566 12960 15622 13016
rect 16394 14320 16450 14376
rect 16486 13640 16542 13696
rect 16394 12316 16396 12336
rect 16396 12316 16448 12336
rect 16448 12316 16450 12336
rect 16394 12280 16450 12316
rect 16394 11620 16450 11656
rect 16394 11600 16396 11620
rect 16396 11600 16448 11620
rect 16448 11600 16450 11620
rect 16394 10240 16450 10296
rect 16578 8200 16634 8256
rect 16578 5516 16580 5536
rect 16580 5516 16632 5536
rect 16632 5516 16634 5536
rect 16578 5480 16634 5516
<< metal3 >>
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 105 39130 171 39133
rect 105 39128 1042 39130
rect 105 39072 110 39128
rect 166 39072 1042 39128
rect 105 39070 1042 39072
rect 105 39067 171 39070
rect 0 38858 800 38888
rect 982 38858 1042 39070
rect 0 38798 1042 38858
rect 0 38768 800 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 7649 37906 7715 37909
rect 8753 37906 8819 37909
rect 7649 37904 8819 37906
rect 7649 37848 7654 37904
rect 7710 37848 8758 37904
rect 8814 37848 8819 37904
rect 7649 37846 8819 37848
rect 7649 37843 7715 37846
rect 8753 37843 8819 37846
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 10593 36138 10659 36141
rect 11145 36138 11211 36141
rect 10593 36136 11211 36138
rect 10593 36080 10598 36136
rect 10654 36080 11150 36136
rect 11206 36080 11211 36136
rect 10593 36078 11211 36080
rect 10593 36075 10659 36078
rect 11145 36075 11211 36078
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 12433 34098 12499 34101
rect 13077 34098 13143 34101
rect 12433 34096 13143 34098
rect 12433 34040 12438 34096
rect 12494 34040 13082 34096
rect 13138 34040 13143 34096
rect 12433 34038 13143 34040
rect 12433 34035 12499 34038
rect 13077 34035 13143 34038
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 9305 27434 9371 27437
rect 12801 27434 12867 27437
rect 9305 27432 12867 27434
rect 9305 27376 9310 27432
rect 9366 27376 12806 27432
rect 12862 27376 12867 27432
rect 9305 27374 12867 27376
rect 9305 27371 9371 27374
rect 12801 27371 12867 27374
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 841 26754 907 26757
rect 798 26752 907 26754
rect 798 26696 846 26752
rect 902 26696 907 26752
rect 798 26691 907 26696
rect 798 26648 858 26691
rect 0 26558 858 26648
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 0 26528 800 26558
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 841 22674 907 22677
rect 798 22672 907 22674
rect 798 22616 846 22672
rect 902 22616 907 22672
rect 798 22611 907 22616
rect 798 22568 858 22611
rect 0 22478 858 22568
rect 16389 22538 16455 22541
rect 17200 22538 18000 22568
rect 16389 22536 18000 22538
rect 16389 22480 16394 22536
rect 16450 22480 18000 22536
rect 16389 22478 18000 22480
rect 0 22448 800 22478
rect 16389 22475 16455 22478
rect 17200 22448 18000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 841 21994 907 21997
rect 798 21992 907 21994
rect 798 21936 846 21992
rect 902 21936 907 21992
rect 798 21931 907 21936
rect 798 21888 858 21931
rect 0 21798 858 21888
rect 16389 21858 16455 21861
rect 17200 21858 18000 21888
rect 16389 21856 18000 21858
rect 16389 21800 16394 21856
rect 16450 21800 18000 21856
rect 16389 21798 18000 21800
rect 0 21768 800 21798
rect 16389 21795 16455 21798
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 17200 21768 18000 21798
rect 4870 21727 5186 21728
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 1301 21178 1367 21181
rect 0 21176 1367 21178
rect 0 21120 1306 21176
rect 1362 21120 1367 21176
rect 0 21118 1367 21120
rect 0 21088 800 21118
rect 1301 21115 1367 21118
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 0 20498 800 20528
rect 3049 20498 3115 20501
rect 0 20496 3115 20498
rect 0 20440 3054 20496
rect 3110 20440 3115 20496
rect 0 20438 3115 20440
rect 0 20408 800 20438
rect 3049 20435 3115 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 841 19954 907 19957
rect 798 19952 907 19954
rect 798 19896 846 19952
rect 902 19896 907 19952
rect 798 19891 907 19896
rect 798 19848 858 19891
rect 0 19758 858 19848
rect 0 19728 800 19758
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 13077 19274 13143 19277
rect 14273 19274 14339 19277
rect 13077 19272 14339 19274
rect 13077 19216 13082 19272
rect 13138 19216 14278 19272
rect 14334 19216 14339 19272
rect 13077 19214 14339 19216
rect 13077 19211 13143 19214
rect 14273 19211 14339 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 11789 18458 11855 18461
rect 13537 18458 13603 18461
rect 11789 18456 13603 18458
rect 11789 18400 11794 18456
rect 11850 18400 13542 18456
rect 13598 18400 13603 18456
rect 11789 18398 13603 18400
rect 11789 18395 11855 18398
rect 13537 18395 13603 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 16389 17098 16455 17101
rect 17200 17098 18000 17128
rect 16389 17096 18000 17098
rect 16389 17040 16394 17096
rect 16450 17040 18000 17096
rect 16389 17038 18000 17040
rect 16389 17035 16455 17038
rect 17200 17008 18000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 12433 15874 12499 15877
rect 12985 15874 13051 15877
rect 12433 15872 13051 15874
rect 12433 15816 12438 15872
rect 12494 15816 12990 15872
rect 13046 15816 13051 15872
rect 12433 15814 13051 15816
rect 12433 15811 12499 15814
rect 12985 15811 13051 15814
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 16389 15738 16455 15741
rect 17200 15738 18000 15768
rect 16389 15736 18000 15738
rect 16389 15680 16394 15736
rect 16450 15680 18000 15736
rect 16389 15678 18000 15680
rect 16389 15675 16455 15678
rect 17200 15648 18000 15678
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 13169 15194 13235 15197
rect 13537 15194 13603 15197
rect 13169 15192 13603 15194
rect 13169 15136 13174 15192
rect 13230 15136 13542 15192
rect 13598 15136 13603 15192
rect 13169 15134 13603 15136
rect 13169 15131 13235 15134
rect 13537 15131 13603 15134
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 16389 14378 16455 14381
rect 17200 14378 18000 14408
rect 16389 14376 18000 14378
rect 16389 14320 16394 14376
rect 16450 14320 18000 14376
rect 16389 14318 18000 14320
rect 16389 14315 16455 14318
rect 17200 14288 18000 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 12157 13970 12223 13973
rect 13445 13970 13511 13973
rect 12157 13968 13511 13970
rect 12157 13912 12162 13968
rect 12218 13912 13450 13968
rect 13506 13912 13511 13968
rect 12157 13910 13511 13912
rect 12157 13907 12223 13910
rect 13445 13907 13511 13910
rect 12249 13834 12315 13837
rect 12893 13834 12959 13837
rect 12249 13832 12959 13834
rect 12249 13776 12254 13832
rect 12310 13776 12898 13832
rect 12954 13776 12959 13832
rect 12249 13774 12959 13776
rect 12249 13771 12315 13774
rect 12893 13771 12959 13774
rect 16481 13698 16547 13701
rect 17200 13698 18000 13728
rect 16481 13696 18000 13698
rect 16481 13640 16486 13696
rect 16542 13640 18000 13696
rect 16481 13638 18000 13640
rect 16481 13635 16547 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 17200 13608 18000 13638
rect 4210 13567 4526 13568
rect 4870 13088 5186 13089
rect 0 13018 800 13048
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 1301 13018 1367 13021
rect 0 13016 1367 13018
rect 0 12960 1306 13016
rect 1362 12960 1367 13016
rect 0 12958 1367 12960
rect 0 12928 800 12958
rect 1301 12955 1367 12958
rect 15561 13018 15627 13021
rect 17200 13018 18000 13048
rect 15561 13016 18000 13018
rect 15561 12960 15566 13016
rect 15622 12960 18000 13016
rect 15561 12958 18000 12960
rect 15561 12955 15627 12958
rect 17200 12928 18000 12958
rect 7189 12612 7255 12613
rect 7189 12608 7236 12612
rect 7300 12610 7306 12612
rect 7189 12552 7194 12608
rect 7189 12548 7236 12552
rect 7300 12550 7346 12610
rect 7300 12548 7306 12550
rect 7189 12547 7255 12548
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 0 12338 800 12368
rect 16389 12338 16455 12341
rect 17200 12338 18000 12368
rect 0 12248 858 12338
rect 16389 12336 18000 12338
rect 16389 12280 16394 12336
rect 16450 12280 18000 12336
rect 16389 12278 18000 12280
rect 16389 12275 16455 12278
rect 17200 12248 18000 12278
rect 798 12205 858 12248
rect 798 12200 907 12205
rect 798 12144 846 12200
rect 902 12144 907 12200
rect 798 12142 907 12144
rect 841 12139 907 12142
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 0 11658 800 11688
rect 1117 11658 1183 11661
rect 0 11656 1183 11658
rect 0 11600 1122 11656
rect 1178 11600 1183 11656
rect 0 11598 1183 11600
rect 0 11568 800 11598
rect 1117 11595 1183 11598
rect 16389 11658 16455 11661
rect 17200 11658 18000 11688
rect 16389 11656 18000 11658
rect 16389 11600 16394 11656
rect 16450 11600 18000 11656
rect 16389 11598 18000 11600
rect 16389 11595 16455 11598
rect 17200 11568 18000 11598
rect 11973 11522 12039 11525
rect 12985 11522 13051 11525
rect 11973 11520 13051 11522
rect 11973 11464 11978 11520
rect 12034 11464 12990 11520
rect 13046 11464 13051 11520
rect 11973 11462 13051 11464
rect 11973 11459 12039 11462
rect 12985 11459 13051 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 0 10978 800 11008
rect 1853 10978 1919 10981
rect 0 10976 1919 10978
rect 0 10920 1858 10976
rect 1914 10920 1919 10976
rect 0 10918 1919 10920
rect 0 10888 800 10918
rect 1853 10915 1919 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 2589 10706 2655 10709
rect 2773 10706 2839 10709
rect 2589 10704 2839 10706
rect 2589 10648 2594 10704
rect 2650 10648 2778 10704
rect 2834 10648 2839 10704
rect 2589 10646 2839 10648
rect 2589 10643 2655 10646
rect 2773 10643 2839 10646
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 1301 10298 1367 10301
rect 0 10296 1367 10298
rect 0 10240 1306 10296
rect 1362 10240 1367 10296
rect 0 10238 1367 10240
rect 0 10208 800 10238
rect 1301 10235 1367 10238
rect 16389 10298 16455 10301
rect 17200 10298 18000 10328
rect 16389 10296 18000 10298
rect 16389 10240 16394 10296
rect 16450 10240 18000 10296
rect 16389 10238 18000 10240
rect 16389 10235 16455 10238
rect 17200 10208 18000 10238
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 0 9618 800 9648
rect 1025 9618 1091 9621
rect 0 9616 1091 9618
rect 0 9560 1030 9616
rect 1086 9560 1091 9616
rect 0 9558 1091 9560
rect 0 9528 800 9558
rect 1025 9555 1091 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 841 9074 907 9077
rect 798 9072 907 9074
rect 798 9016 846 9072
rect 902 9016 907 9072
rect 798 9011 907 9016
rect 798 8968 858 9011
rect 0 8878 858 8968
rect 0 8848 800 8878
rect 4654 8876 4660 8940
rect 4724 8938 4730 8940
rect 5165 8938 5231 8941
rect 4724 8936 5231 8938
rect 4724 8880 5170 8936
rect 5226 8880 5231 8936
rect 4724 8878 5231 8880
rect 4724 8876 4730 8878
rect 5165 8875 5231 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 0 8258 800 8288
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8168 800 8198
rect 2773 8195 2839 8198
rect 16573 8258 16639 8261
rect 17200 8258 18000 8288
rect 16573 8256 18000 8258
rect 16573 8200 16578 8256
rect 16634 8200 18000 8256
rect 16573 8198 18000 8200
rect 16573 8195 16639 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 17200 8168 18000 8198
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 2957 7578 3023 7581
rect 0 7576 3023 7578
rect 0 7520 2962 7576
rect 3018 7520 3023 7576
rect 0 7518 3023 7520
rect 0 7488 800 7518
rect 2957 7515 3023 7518
rect 2405 7306 2471 7309
rect 8385 7306 8451 7309
rect 2405 7304 8451 7306
rect 2405 7248 2410 7304
rect 2466 7248 8390 7304
rect 8446 7248 8451 7304
rect 2405 7246 8451 7248
rect 2405 7243 2471 7246
rect 8385 7243 8451 7246
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 13905 6354 13971 6357
rect 14825 6354 14891 6357
rect 13905 6352 14891 6354
rect 13905 6296 13910 6352
rect 13966 6296 14830 6352
rect 14886 6296 14891 6352
rect 13905 6294 14891 6296
rect 13905 6291 13971 6294
rect 14825 6291 14891 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 16573 5538 16639 5541
rect 17200 5538 18000 5568
rect 16573 5536 18000 5538
rect 16573 5480 16578 5536
rect 16634 5480 18000 5536
rect 16573 5478 18000 5480
rect 16573 5475 16639 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 17200 5448 18000 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 3509 4178 3575 4181
rect 6545 4178 6611 4181
rect 7833 4178 7899 4181
rect 3509 4176 7899 4178
rect 3509 4120 3514 4176
rect 3570 4120 6550 4176
rect 6606 4120 7838 4176
rect 7894 4120 7899 4176
rect 3509 4118 7899 4120
rect 3509 4115 3575 4118
rect 6545 4115 6611 4118
rect 7833 4115 7899 4118
rect 7230 3980 7236 4044
rect 7300 4042 7306 4044
rect 11513 4042 11579 4045
rect 7300 4040 11579 4042
rect 7300 3984 11518 4040
rect 11574 3984 11579 4040
rect 7300 3982 11579 3984
rect 7300 3980 7306 3982
rect 11513 3979 11579 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 4245 3634 4311 3637
rect 4654 3634 4660 3636
rect 4245 3632 4660 3634
rect 4245 3576 4250 3632
rect 4306 3576 4660 3632
rect 4245 3574 4660 3576
rect 4245 3571 4311 3574
rect 4654 3572 4660 3574
rect 4724 3634 4730 3636
rect 7281 3634 7347 3637
rect 4724 3632 7347 3634
rect 4724 3576 7286 3632
rect 7342 3576 7347 3632
rect 4724 3574 7347 3576
rect 4724 3572 4730 3574
rect 7281 3571 7347 3574
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
<< via3 >>
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 7236 12608 7300 12612
rect 7236 12552 7250 12608
rect 7250 12552 7300 12608
rect 7236 12548 7300 12552
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4660 8876 4724 8940
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 7236 3980 7300 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4660 3572 4724 3636
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 39744 4528 39760
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4868 39200 5188 39760
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 35936 5188 36960
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 7235 12612 7301 12613
rect 7235 12548 7236 12612
rect 7300 12548 7301 12612
rect 7235 12547 7301 12548
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4659 8940 4725 8941
rect 4659 8876 4660 8940
rect 4724 8876 4725 8940
rect 4659 8875 4725 8876
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4662 3637 4722 8875
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4659 3636 4725 3637
rect 4659 3572 4660 3636
rect 4724 3572 4725 3636
rect 4659 3571 4725 3572
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 3296 5188 4320
rect 7238 4045 7298 12547
rect 7235 4044 7301 4045
rect 7235 3980 7236 4044
rect 7300 3980 7301 4044
rect 7235 3979 7301 3980
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__inv_2  _0527_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 8188 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0528_
timestamp 1730493024
transform -1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0529_
timestamp 1730493024
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0530_
timestamp 1730493024
transform -1 0 9752 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0531_
timestamp 1730493024
transform -1 0 12420 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0532_
timestamp 1730493024
transform 1 0 11684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0533_
timestamp 1730493024
transform -1 0 14812 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0534_
timestamp 1730493024
transform 1 0 9200 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0535_
timestamp 1730493024
transform 1 0 6256 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0536_
timestamp 1730493024
transform 1 0 14076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0537_
timestamp 1730493024
transform -1 0 12328 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0538_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 2760 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0539_
timestamp 1730493024
transform 1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0540_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3588 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0541_
timestamp 1730493024
transform -1 0 2576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0542_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 3128 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0543_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 3772 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0544_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 3680 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0545_
timestamp 1730493024
transform 1 0 2852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0546_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 3036 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0547_
timestamp 1730493024
transform 1 0 5520 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0548_
timestamp 1730493024
transform -1 0 7452 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0549_
timestamp 1730493024
transform 1 0 7636 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0550_
timestamp 1730493024
transform 1 0 7452 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _0551_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 6532 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0552_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 6348 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0553_
timestamp 1730493024
transform 1 0 6532 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0554_
timestamp 1704896540
transform 1 0 7912 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0555_
timestamp 1730493024
transform 1 0 9476 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0556_
timestamp 1730493024
transform 1 0 10948 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0557_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 6348 0 -1 33728
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _0558_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 11040 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0559_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 10212 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0560_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 10856 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0561_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 10212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0562_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 11500 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0563_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 10764 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0564_
timestamp 1730493024
transform 1 0 11500 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _0565_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 11500 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0566_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 10948 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_1  _0567_
timestamp 1730493024
transform -1 0 11316 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0568_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 10212 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0569_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 10856 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0570_
timestamp 1730493024
transform -1 0 9936 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0571_
timestamp 1730493024
transform -1 0 10120 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__and3b_1  _0572_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 12144 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0573_
timestamp 1730493024
transform 1 0 10580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__o311a_1  _0574_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 11040 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _0575_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 9936 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0576_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _0577_
timestamp 1730493024
transform 1 0 8924 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0578_
timestamp 1730493024
transform 1 0 8648 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0579_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _0580_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 10304 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0581_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 10764 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0582_
timestamp 1730493024
transform -1 0 10396 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a22oi_2  _0583_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9936 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0584_
timestamp 1730493024
transform 1 0 8924 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0585_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 2576 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0586_
timestamp 1730493024
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0587_
timestamp 1730493024
transform 1 0 3772 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0588_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 4048 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _0589_
timestamp 1730493024
transform 1 0 9476 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_2  _0590_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9568 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0591_
timestamp 1730493024
transform 1 0 12144 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0592_
timestamp 1730493024
transform 1 0 12880 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_2  _0593_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 14352 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0594_
timestamp 1730493024
transform -1 0 12420 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0595_
timestamp 1730493024
transform -1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _0596_
timestamp 1730493024
transform 1 0 11684 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0597_
timestamp 1730493024
transform 1 0 12696 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0598_
timestamp 1730493024
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0599_
timestamp 1730493024
transform 1 0 13524 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0600_
timestamp 1730493024
transform 1 0 13524 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0601_
timestamp 1730493024
transform 1 0 4232 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0602_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 5060 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0603_
timestamp 1730493024
transform 1 0 9660 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0604_
timestamp 1730493024
transform -1 0 12880 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _0605_
timestamp 1730493024
transform 1 0 13064 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0606_
timestamp 1730493024
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0607_
timestamp 1730493024
transform 1 0 12880 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0608_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 13892 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0609_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 13340 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0610_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 14076 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _0611_
timestamp 1730493024
transform 1 0 14076 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0612_
timestamp 1730493024
transform 1 0 13984 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0613_
timestamp 1730493024
transform 1 0 15088 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0614_
timestamp 1730493024
transform 1 0 8464 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0615_
timestamp 1730493024
transform -1 0 8832 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0616_
timestamp 1730493024
transform 1 0 7360 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0617_
timestamp 1730493024
transform 1 0 8280 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _0618_
timestamp 1730493024
transform -1 0 11592 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0619_
timestamp 1730493024
transform -1 0 10488 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0620_
timestamp 1730493024
transform 1 0 10488 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _0621_
timestamp 1730493024
transform 1 0 10396 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0622_
timestamp 1730493024
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0623_
timestamp 1730493024
transform 1 0 10120 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0624_
timestamp 1730493024
transform 1 0 10580 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0625_
timestamp 1730493024
transform -1 0 12052 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0626_
timestamp 1730493024
transform -1 0 12696 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0627_
timestamp 1730493024
transform -1 0 11316 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0628_
timestamp 1730493024
transform 1 0 10212 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0629_
timestamp 1730493024
transform -1 0 12144 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _0630_
timestamp 1730493024
transform -1 0 12696 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0631_
timestamp 1730493024
transform -1 0 11500 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0632_
timestamp 1730493024
transform 1 0 11500 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0633_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 10764 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0634_
timestamp 1730493024
transform 1 0 10672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0635_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 10488 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0636_
timestamp 1730493024
transform 1 0 9384 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0637_
timestamp 1730493024
transform -1 0 9660 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0638_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 8740 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _0639_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_1  _0640_
timestamp 1730493024
transform 1 0 9660 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0641_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 10764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2a_1  _0642_
timestamp 1730493024
transform 1 0 9292 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_1  _0643_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 13800 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _0644_
timestamp 1730493024
transform 1 0 11960 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0645_
timestamp 1704896540
transform 1 0 12604 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0646_
timestamp 1730493024
transform -1 0 13800 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0647_
timestamp 1730493024
transform -1 0 14168 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0648_
timestamp 1730493024
transform -1 0 13064 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0649_
timestamp 1704896540
transform 1 0 13064 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0650_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 12972 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0651_
timestamp 1730493024
transform 1 0 13432 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0652_
timestamp 1730493024
transform -1 0 13432 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0653_
timestamp 1704896540
transform 1 0 12696 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0654_
timestamp 1730493024
transform 1 0 12604 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0655_
timestamp 1704896540
transform 1 0 12420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0656_
timestamp 1730493024
transform -1 0 12052 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0657_
timestamp 1730493024
transform 1 0 12052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0658_
timestamp 1730493024
transform -1 0 12144 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0659_
timestamp 1704896540
transform 1 0 11500 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0660_
timestamp 1730493024
transform -1 0 11960 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0661_
timestamp 1730493024
transform -1 0 11408 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0662_
timestamp 1730493024
transform -1 0 11040 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0663_
timestamp 1704896540
transform 1 0 10028 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0664_
timestamp 1730493024
transform 1 0 8188 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0665_
timestamp 1704896540
transform 1 0 8832 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0666_
timestamp 1730493024
transform 1 0 8372 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0667_
timestamp 1730493024
transform 1 0 9660 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0668_
timestamp 1730493024
transform -1 0 9200 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0669_
timestamp 1704896540
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0670_
timestamp 1730493024
transform -1 0 8924 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0671_
timestamp 1730493024
transform -1 0 8372 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0672_
timestamp 1730493024
transform -1 0 7636 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _0673_
timestamp 1704896540
transform -1 0 8280 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1730493024
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0675_
timestamp 1730493024
transform 1 0 6440 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0676_
timestamp 1704896540
transform 1 0 6532 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0677_
timestamp 1730493024
transform -1 0 7176 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0678_
timestamp 1704896540
transform -1 0 7268 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _0679_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 8188 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _0680_
timestamp 1704896540
transform 1 0 7544 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _0681_
timestamp 1730493024
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0682_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 1472 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _0683_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 9936 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0684_
timestamp 1730493024
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0685_
timestamp 1730493024
transform 1 0 8372 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _0686_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 4600 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1730493024
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0688_
timestamp 1730493024
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _0689_
timestamp 1730493024
transform -1 0 4876 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0690_
timestamp 1730493024
transform 1 0 1656 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0691_
timestamp 1730493024
transform 1 0 1656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0692_
timestamp 1730493024
transform 1 0 4508 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0693_
timestamp 1730493024
transform -1 0 5060 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0694_
timestamp 1730493024
transform 1 0 3588 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0695_
timestamp 1730493024
transform -1 0 4784 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0696_
timestamp 1730493024
transform 1 0 1656 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0697_
timestamp 1730493024
transform -1 0 2668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0698_
timestamp 1730493024
transform 1 0 3772 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0699_
timestamp 1730493024
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0700_
timestamp 1730493024
transform 1 0 1380 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0701_
timestamp 1730493024
transform 1 0 2392 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0702_
timestamp 1730493024
transform 1 0 4784 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0703_
timestamp 1730493024
transform -1 0 4508 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0704_
timestamp 1730493024
transform 1 0 3312 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0705_
timestamp 1730493024
transform -1 0 4600 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0706_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9660 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0707_
timestamp 1730493024
transform 1 0 13248 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0708_
timestamp 1704896540
transform 1 0 12788 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0709_
timestamp 1730493024
transform 1 0 14536 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0710_
timestamp 1730493024
transform -1 0 15640 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0711_
timestamp 1730493024
transform 1 0 14076 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0712_
timestamp 1730493024
transform -1 0 14904 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0713_
timestamp 1730493024
transform -1 0 12328 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0714_
timestamp 1730493024
transform -1 0 13064 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0715_
timestamp 1730493024
transform 1 0 14168 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0716_
timestamp 1730493024
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0717_
timestamp 1730493024
transform -1 0 13340 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0718_
timestamp 1730493024
transform 1 0 12144 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0719_
timestamp 1730493024
transform 1 0 13524 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0720_
timestamp 1730493024
transform -1 0 15180 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0721_
timestamp 1730493024
transform -1 0 13524 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0722_
timestamp 1730493024
transform -1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0723_
timestamp 1730493024
transform 1 0 13248 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0724_
timestamp 1730493024
transform -1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _0725_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0726_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 12880 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0727_
timestamp 1704896540
transform 1 0 12880 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0728_
timestamp 1730493024
transform 1 0 13892 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0729_
timestamp 1730493024
transform 1 0 13064 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0730_
timestamp 1730493024
transform 1 0 7176 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0731_
timestamp 1730493024
transform 1 0 6992 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0732_
timestamp 1730493024
transform 1 0 7268 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0733_
timestamp 1730493024
transform 1 0 7176 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0734_
timestamp 1730493024
transform 1 0 13524 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0735_
timestamp 1730493024
transform -1 0 15180 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0736_
timestamp 1730493024
transform 1 0 8372 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0737_
timestamp 1730493024
transform 1 0 8096 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0738_
timestamp 1730493024
transform 1 0 13800 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0739_
timestamp 1730493024
transform -1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0740_
timestamp 1730493024
transform 1 0 8372 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0741_
timestamp 1730493024
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0742_
timestamp 1730493024
transform 1 0 6992 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0743_
timestamp 1730493024
transform 1 0 7452 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _0744_
timestamp 1704896540
transform -1 0 9384 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0745_
timestamp 1730493024
transform -1 0 5244 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0746_
timestamp 1704896540
transform -1 0 5612 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0747_
timestamp 1730493024
transform -1 0 3496 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0748_
timestamp 1730493024
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0749_
timestamp 1730493024
transform 1 0 3772 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0750_
timestamp 1730493024
transform -1 0 4600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0751_
timestamp 1730493024
transform 1 0 4140 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0752_
timestamp 1730493024
transform 1 0 4232 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0753_
timestamp 1730493024
transform -1 0 4140 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0754_
timestamp 1730493024
transform 1 0 2760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0755_
timestamp 1730493024
transform -1 0 6164 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0756_
timestamp 1730493024
transform -1 0 5336 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0757_
timestamp 1730493024
transform -1 0 4232 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0758_
timestamp 1730493024
transform 1 0 2668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0759_
timestamp 1730493024
transform 1 0 5796 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0760_
timestamp 1730493024
transform -1 0 5796 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0761_
timestamp 1730493024
transform 1 0 4140 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0762_
timestamp 1730493024
transform -1 0 5152 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _0763_
timestamp 1704896540
transform 1 0 8648 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _0764_
timestamp 1704896540
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0765_
timestamp 1704896540
transform -1 0 10948 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0766_
timestamp 1730493024
transform 1 0 1564 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0767_
timestamp 1730493024
transform 1 0 1472 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0768_
timestamp 1730493024
transform -1 0 11408 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0769_
timestamp 1730493024
transform 1 0 10212 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0770_
timestamp 1730493024
transform -1 0 11408 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0771_
timestamp 1730493024
transform 1 0 10212 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0772_
timestamp 1730493024
transform -1 0 2300 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0773_
timestamp 1730493024
transform 1 0 1472 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0774_
timestamp 1730493024
transform -1 0 11408 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0775_
timestamp 1730493024
transform 1 0 9384 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0776_
timestamp 1730493024
transform -1 0 2760 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0777_
timestamp 1730493024
transform 1 0 1564 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0778_
timestamp 1730493024
transform -1 0 10396 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0779_
timestamp 1730493024
transform -1 0 9936 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0780_
timestamp 1730493024
transform 1 0 12328 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0781_
timestamp 1730493024
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0782_
timestamp 1730493024
transform 1 0 2944 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0783_
timestamp 1730493024
transform -1 0 14444 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0784_
timestamp 1730493024
transform -1 0 3772 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0785_
timestamp 1730493024
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0786_
timestamp 1730493024
transform 1 0 6532 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0787_
timestamp 1730493024
transform -1 0 12144 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0788_
timestamp 1730493024
transform -1 0 7820 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0789_
timestamp 1730493024
transform -1 0 9568 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0790_
timestamp 1730493024
transform 1 0 6716 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0791_
timestamp 1730493024
transform -1 0 12328 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0792_
timestamp 1730493024
transform 1 0 6716 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0793_
timestamp 1730493024
transform 1 0 10120 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0794_
timestamp 1730493024
transform -1 0 15640 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0795_
timestamp 1730493024
transform 1 0 2852 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0796_
timestamp 1730493024
transform -1 0 4416 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0797_
timestamp 1730493024
transform 1 0 5704 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0798_
timestamp 1730493024
transform -1 0 12144 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0799_
timestamp 1730493024
transform 1 0 7636 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0800_
timestamp 1730493024
transform 1 0 7912 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0801_
timestamp 1730493024
transform 1 0 7360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0802_
timestamp 1730493024
transform 1 0 2760 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0803_
timestamp 1730493024
transform -1 0 14904 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0804_
timestamp 1730493024
transform -1 0 5428 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0805_
timestamp 1730493024
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0806_
timestamp 1730493024
transform -1 0 11500 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0807_
timestamp 1730493024
transform 1 0 8188 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0808_
timestamp 1730493024
transform 1 0 8188 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0809_
timestamp 1730493024
transform 1 0 8924 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0810_
timestamp 1730493024
transform 1 0 6348 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0811_
timestamp 1730493024
transform 1 0 12420 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0812_
timestamp 1730493024
transform 1 0 6440 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0813_
timestamp 1730493024
transform 1 0 7544 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0814_
timestamp 1730493024
transform 1 0 8004 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0815_
timestamp 1730493024
transform 1 0 9476 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1730493024
transform 1 0 6348 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0817_
timestamp 1730493024
transform 1 0 3036 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0818_
timestamp 1730493024
transform -1 0 4324 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _0819_
timestamp 1730493024
transform 1 0 3404 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0820_
timestamp 1730493024
transform -1 0 4140 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0821_
timestamp 1730493024
transform 1 0 6348 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1730493024
transform -1 0 9200 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0823_
timestamp 1730493024
transform -1 0 8004 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0824_
timestamp 1730493024
transform 1 0 10948 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0825_
timestamp 1730493024
transform 1 0 8188 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _0826_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 8004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0827_
timestamp 1730493024
transform -1 0 8464 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1730493024
transform -1 0 7912 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0829_
timestamp 1730493024
transform -1 0 5704 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0830_
timestamp 1730493024
transform 1 0 7176 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0831_
timestamp 1730493024
transform -1 0 9384 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0832_
timestamp 1730493024
transform 1 0 7176 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0833_
timestamp 1730493024
transform -1 0 8556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0834_
timestamp 1730493024
transform -1 0 8372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1730493024
transform -1 0 7176 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0836_
timestamp 1730493024
transform 1 0 7268 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0837_
timestamp 1730493024
transform -1 0 8924 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0838_
timestamp 1730493024
transform -1 0 9476 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _0839_
timestamp 1730493024
transform 1 0 7728 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _0840_
timestamp 1730493024
transform 1 0 7544 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1730493024
transform 1 0 6900 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0842_
timestamp 1730493024
transform 1 0 6992 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _0843_
timestamp 1730493024
transform 1 0 6440 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _0844_
timestamp 1730493024
transform -1 0 7912 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _0845_
timestamp 1730493024
transform 1 0 5428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0846_
timestamp 1730493024
transform -1 0 6716 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0847_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6716 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0848_
timestamp 1730493024
transform -1 0 6256 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0849_
timestamp 1730493024
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0850_
timestamp 1730493024
transform 1 0 8004 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0851_
timestamp 1730493024
transform 1 0 9016 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0852_
timestamp 1730493024
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0853_
timestamp 1730493024
transform 1 0 6900 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0854_
timestamp 1730493024
transform -1 0 6992 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0855_
timestamp 1730493024
transform -1 0 8648 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0856_
timestamp 1730493024
transform 1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0857_
timestamp 1730493024
transform 1 0 7728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0858_
timestamp 1730493024
transform 1 0 6900 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0859_
timestamp 1730493024
transform 1 0 9660 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0860_
timestamp 1730493024
transform 1 0 9568 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0861_
timestamp 1730493024
transform 1 0 9384 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0862_
timestamp 1730493024
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0863_
timestamp 1730493024
transform 1 0 6440 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0864_
timestamp 1730493024
transform 1 0 5428 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _0865_
timestamp 1730493024
transform 1 0 5796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0866_
timestamp 1730493024
transform 1 0 1932 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0867_
timestamp 1730493024
transform 1 0 5060 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0868_
timestamp 1730493024
transform -1 0 6072 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _0869_
timestamp 1730493024
transform 1 0 5244 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0870_
timestamp 1730493024
transform 1 0 5336 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0871_
timestamp 1730493024
transform 1 0 4968 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0872_
timestamp 1730493024
transform 1 0 4968 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0873_
timestamp 1730493024
transform 1 0 5796 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0874_
timestamp 1730493024
transform 1 0 4876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0875_
timestamp 1730493024
transform -1 0 5520 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0876_
timestamp 1730493024
transform 1 0 4508 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o41ai_1  _0877_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_1  _0878_
timestamp 1730493024
transform 1 0 3956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0879_
timestamp 1730493024
transform -1 0 4508 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0880_
timestamp 1730493024
transform 1 0 2576 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0881_
timestamp 1730493024
transform -1 0 3312 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0882_
timestamp 1730493024
transform -1 0 3220 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _0883_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 6440 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0884_
timestamp 1730493024
transform -1 0 4416 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0885_
timestamp 1730493024
transform -1 0 5152 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0886_
timestamp 1730493024
transform 1 0 4416 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0887_
timestamp 1730493024
transform 1 0 3772 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0888_
timestamp 1730493024
transform 1 0 4324 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0889_
timestamp 1730493024
transform 1 0 4416 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0890_
timestamp 1730493024
transform 1 0 4416 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0891_
timestamp 1730493024
transform -1 0 5336 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0892_
timestamp 1730493024
transform 1 0 3772 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0893_
timestamp 1730493024
transform -1 0 3588 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0894_
timestamp 1730493024
transform -1 0 4324 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0895_
timestamp 1730493024
transform 1 0 3220 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0896_
timestamp 1730493024
transform 1 0 3772 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0897_
timestamp 1730493024
transform -1 0 4048 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0898_
timestamp 1730493024
transform -1 0 3864 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0899_
timestamp 1730493024
transform 1 0 2944 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0900_
timestamp 1730493024
transform -1 0 3680 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0901_
timestamp 1730493024
transform 1 0 3772 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0902_
timestamp 1730493024
transform -1 0 3128 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0903_
timestamp 1730493024
transform -1 0 3496 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0904_
timestamp 1730493024
transform 1 0 3496 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _0905_
timestamp 1730493024
transform -1 0 3312 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1730493024
transform 1 0 4048 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0907_
timestamp 1730493024
transform 1 0 3588 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0908_
timestamp 1730493024
transform 1 0 4048 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _0909_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 5704 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0910_
timestamp 1730493024
transform -1 0 4048 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0911_
timestamp 1730493024
transform 1 0 5244 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0912_
timestamp 1730493024
transform 1 0 4784 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0913_
timestamp 1730493024
transform 1 0 3220 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0914_
timestamp 1730493024
transform 1 0 3128 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0915_
timestamp 1730493024
transform 1 0 7452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0916_
timestamp 1730493024
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _0917_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 1730493024
transform -1 0 6348 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0919_
timestamp 1730493024
transform -1 0 6440 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0920_
timestamp 1730493024
transform 1 0 5520 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0921_
timestamp 1730493024
transform -1 0 6900 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0922_
timestamp 1730493024
transform 1 0 6348 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1730493024
transform 1 0 7728 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0924_
timestamp 1730493024
transform 1 0 5612 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0925_
timestamp 1730493024
transform 1 0 6808 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _0926_
timestamp 1730493024
transform 1 0 11868 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0927_
timestamp 1730493024
transform -1 0 13340 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0928_
timestamp 1730493024
transform -1 0 13984 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0929_
timestamp 1730493024
transform 1 0 12880 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1730493024
transform -1 0 13064 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1730493024
transform -1 0 12880 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1730493024
transform 1 0 12512 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0933_
timestamp 1730493024
transform -1 0 13248 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0934_
timestamp 1730493024
transform -1 0 12420 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0935_
timestamp 1730493024
transform -1 0 12696 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1730493024
transform 1 0 12696 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0937_
timestamp 1730493024
transform 1 0 12144 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0938_
timestamp 1730493024
transform 1 0 12604 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0939_
timestamp 1730493024
transform 1 0 13156 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0940_
timestamp 1730493024
transform 1 0 12512 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0941_
timestamp 1730493024
transform -1 0 11960 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0942_
timestamp 1730493024
transform 1 0 12144 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0943_
timestamp 1730493024
transform -1 0 11868 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1730493024
transform 1 0 11868 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0945_
timestamp 1730493024
transform 1 0 11500 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0946_
timestamp 1730493024
transform -1 0 11316 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1730493024
transform -1 0 10856 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0948_
timestamp 1730493024
transform -1 0 10488 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0949_
timestamp 1730493024
transform -1 0 9016 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0950_
timestamp 1730493024
transform 1 0 8372 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0951_
timestamp 1730493024
transform -1 0 8096 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0952_
timestamp 1730493024
transform 1 0 8004 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1730493024
transform 1 0 8096 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0954_
timestamp 1730493024
transform 1 0 7176 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0955_
timestamp 1730493024
transform 1 0 7360 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0956_
timestamp 1730493024
transform 1 0 7084 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1730493024
transform -1 0 7176 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0958_
timestamp 1730493024
transform -1 0 7084 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0959_
timestamp 1730493024
transform 1 0 6440 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0960_
timestamp 1730493024
transform -1 0 7176 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0961_
timestamp 1730493024
transform -1 0 8280 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0962_
timestamp 1730493024
transform -1 0 7912 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0963_
timestamp 1730493024
transform 1 0 7360 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0964_
timestamp 1730493024
transform -1 0 7452 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0965_
timestamp 1730493024
transform -1 0 8832 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _0966_
timestamp 1730493024
transform 1 0 12972 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0967_
timestamp 1730493024
transform -1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0968_
timestamp 1730493024
transform 1 0 14168 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _0969_
timestamp 1730493024
transform 1 0 15180 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0970_
timestamp 1730493024
transform 1 0 2576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0971_
timestamp 1730493024
transform 1 0 1472 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0972_
timestamp 1704896540
transform -1 0 12328 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0973_
timestamp 1730493024
transform 1 0 12328 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0974_
timestamp 1730493024
transform 1 0 12236 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0975_
timestamp 1730493024
transform -1 0 12144 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0976_
timestamp 1730493024
transform 1 0 12420 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0977_
timestamp 1730493024
transform -1 0 13524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0978_
timestamp 1730493024
transform 1 0 12052 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0979_
timestamp 1730493024
transform 1 0 12144 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0980_
timestamp 1730493024
transform -1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _0981_
timestamp 1730493024
transform 1 0 11500 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0982_
timestamp 1730493024
transform -1 0 12328 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1730493024
transform -1 0 12788 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0984_
timestamp 1730493024
transform -1 0 12696 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0985_
timestamp 1730493024
transform -1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1730493024
transform -1 0 12144 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0987_
timestamp 1730493024
transform -1 0 12880 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0988_
timestamp 1730493024
transform -1 0 13432 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0989_
timestamp 1730493024
transform -1 0 12972 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0990_
timestamp 1730493024
transform 1 0 12052 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1730493024
transform -1 0 12420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 1730493024
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0993_
timestamp 1730493024
transform 1 0 12512 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0994_
timestamp 1730493024
transform -1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _0995_
timestamp 1730493024
transform -1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0996_
timestamp 1730493024
transform -1 0 12236 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0997_
timestamp 1730493024
transform -1 0 13892 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0998_
timestamp 1730493024
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _0999_
timestamp 1730493024
transform -1 0 14352 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1000_
timestamp 1730493024
transform 1 0 14076 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1730493024
transform 1 0 11776 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1002_
timestamp 1730493024
transform -1 0 14260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1730493024
transform 1 0 13708 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1004_
timestamp 1730493024
transform 1 0 14352 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1005_
timestamp 1730493024
transform 1 0 14812 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o221a_1  _1006_
timestamp 1730493024
transform 1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1007_
timestamp 1730493024
transform -1 0 14076 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1008_
timestamp 1730493024
transform 1 0 14076 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1009_
timestamp 1730493024
transform 1 0 15088 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1010_
timestamp 1730493024
transform 1 0 13340 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1730493024
transform -1 0 14536 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1012_
timestamp 1730493024
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1013_
timestamp 1730493024
transform 1 0 13156 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1014_
timestamp 1730493024
transform 1 0 14996 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _1015_
timestamp 1730493024
transform -1 0 13892 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1016_
timestamp 1730493024
transform -1 0 14444 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1017_
timestamp 1730493024
transform 1 0 14628 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1018_
timestamp 1730493024
transform 1 0 14260 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1019_
timestamp 1730493024
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1020_
timestamp 1730493024
transform 1 0 12696 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1021_
timestamp 1730493024
transform 1 0 13248 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1022_
timestamp 1730493024
transform -1 0 13432 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1023_
timestamp 1730493024
transform -1 0 13892 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1024_
timestamp 1730493024
transform 1 0 13248 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1025_
timestamp 1730493024
transform -1 0 15088 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1026_
timestamp 1730493024
transform 1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1027_
timestamp 1730493024
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1028_
timestamp 1730493024
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a32o_1  _1029_
timestamp 1730493024
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1030_
timestamp 1730493024
transform 1 0 11316 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1031_
timestamp 1730493024
transform 1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1032_
timestamp 1730493024
transform 1 0 3588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1033_
timestamp 1730493024
transform 1 0 2392 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1034_
timestamp 1730493024
transform -1 0 3312 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1035_
timestamp 1730493024
transform -1 0 2300 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1036_
timestamp 1730493024
transform -1 0 2208 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1037_
timestamp 1730493024
transform -1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1038_
timestamp 1730493024
transform 1 0 10580 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1730493024
transform 1 0 11684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1040_
timestamp 1730493024
transform -1 0 2300 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1041_
timestamp 1730493024
transform 1 0 1656 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1042_
timestamp 1730493024
transform 1 0 3036 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1043_
timestamp 1730493024
transform 1 0 4048 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and4b_1  _1044_
timestamp 1704896540
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1045_
timestamp 1730493024
transform -1 0 11408 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1730493024
transform 1 0 11592 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22ai_1  _1047_
timestamp 1730493024
transform 1 0 13156 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1048_
timestamp 1730493024
transform 1 0 3864 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1049_
timestamp 1730493024
transform 1 0 2300 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1050_
timestamp 1730493024
transform 1 0 2300 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1730493024
transform -1 0 11868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1052_
timestamp 1730493024
transform 1 0 12696 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1053_
timestamp 1730493024
transform 1 0 13156 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1054_
timestamp 1730493024
transform 1 0 12236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1055_
timestamp 1730493024
transform 1 0 14076 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1056_
timestamp 1730493024
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_2  _1057_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 3956 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1058_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 14720 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1059_
timestamp 1730493024
transform 1 0 12420 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1060_
timestamp 1730493024
transform 1 0 13064 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1061_
timestamp 1730493024
transform 1 0 14076 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1062_
timestamp 1730493024
transform 1 0 13432 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1063_
timestamp 1730493024
transform -1 0 14628 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1064_
timestamp 1730493024
transform 1 0 11684 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1065_
timestamp 1730493024
transform 1 0 9936 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1066_
timestamp 1730493024
transform 1 0 9200 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1067_
timestamp 1730493024
transform -1 0 10212 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1068_
timestamp 1730493024
transform 1 0 6808 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1069_
timestamp 1730493024
transform -1 0 7820 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1070_
timestamp 1730493024
transform 1 0 6440 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1071_
timestamp 1730493024
transform 1 0 7912 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1072_
timestamp 1730493024
transform 1 0 1380 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1073_
timestamp 1730493024
transform 1 0 8464 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1074_
timestamp 1730493024
transform 1 0 1748 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1075_
timestamp 1730493024
transform 1 0 4784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1076_
timestamp 1730493024
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1077_
timestamp 1730493024
transform 1 0 2116 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1078_
timestamp 1730493024
transform 1 0 3312 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1079_
timestamp 1730493024
transform 1 0 1840 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1080_
timestamp 1730493024
transform 1 0 4508 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1081_
timestamp 1730493024
transform 1 0 4600 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1082_
timestamp 1730493024
transform 1 0 15088 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1083_
timestamp 1730493024
transform 1 0 14628 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1084_
timestamp 1730493024
transform 1 0 12328 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1085_
timestamp 1730493024
transform 1 0 13524 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1086_
timestamp 1730493024
transform 1 0 11592 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1087_
timestamp 1730493024
transform 1 0 15088 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1088_
timestamp 1730493024
transform 1 0 13248 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1089_
timestamp 1730493024
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1090_
timestamp 1730493024
transform 1 0 12420 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1091_
timestamp 1730493024
transform -1 0 7912 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1092_
timestamp 1730493024
transform 1 0 6900 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1093_
timestamp 1730493024
transform 1 0 15088 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1094_
timestamp 1730493024
transform 1 0 8004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1095_
timestamp 1730493024
transform 1 0 14996 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1096_
timestamp 1730493024
transform 1 0 8648 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1097_
timestamp 1730493024
transform -1 0 7452 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1098_
timestamp 1730493024
transform 1 0 2300 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1099_
timestamp 1730493024
transform 1 0 4232 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1100_
timestamp 1730493024
transform 1 0 4048 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1101_
timestamp 1730493024
transform 1 0 2208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1102_
timestamp 1730493024
transform 1 0 5336 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1103_
timestamp 1730493024
transform 1 0 2024 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1104_
timestamp 1730493024
transform 1 0 5520 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1105_
timestamp 1730493024
transform 1 0 4600 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1106_
timestamp 1730493024
transform 1 0 1380 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1107_
timestamp 1730493024
transform 1 0 10120 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1108_
timestamp 1730493024
transform 1 0 10396 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1109_
timestamp 1730493024
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1110_
timestamp 1730493024
transform 1 0 9476 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1111_
timestamp 1730493024
transform 1 0 1380 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1112_
timestamp 1730493024
transform 1 0 9936 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1113_
timestamp 1730493024
transform 1 0 10856 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1114_
timestamp 1730493024
transform 1 0 9476 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1115_
timestamp 1730493024
transform 1 0 4784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1116_
timestamp 1730493024
transform 1 0 8924 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1117_
timestamp 1730493024
transform 1 0 9108 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1118_
timestamp 1730493024
transform 1 0 5336 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1119_
timestamp 1730493024
transform 1 0 6900 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1120_
timestamp 1730493024
transform 1 0 5428 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1121_
timestamp 1730493024
transform 1 0 8648 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1122_
timestamp 1730493024
transform 1 0 7176 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1123_
timestamp 1730493024
transform 1 0 7360 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1124_
timestamp 1730493024
transform 1 0 9200 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1125_
timestamp 1730493024
transform 1 0 6072 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1126_
timestamp 1730493024
transform 1 0 3772 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1127_
timestamp 1730493024
transform 1 0 4232 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1128_
timestamp 1730493024
transform 1 0 6072 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1129_
timestamp 1730493024
transform 1 0 8004 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1130_
timestamp 1730493024
transform -1 0 5612 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1131_
timestamp 1730493024
transform 1 0 6716 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1132_
timestamp 1730493024
transform 1 0 5704 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1133_
timestamp 1730493024
transform 1 0 7820 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1134_
timestamp 1730493024
transform -1 0 9384 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1135_
timestamp 1730493024
transform 1 0 6348 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1136_
timestamp 1730493024
transform 1 0 6532 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1137_
timestamp 1730493024
transform 1 0 6348 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1138_
timestamp 1730493024
transform 1 0 8096 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1139_
timestamp 1730493024
transform 1 0 8464 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1140_
timestamp 1730493024
transform 1 0 5244 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1141_
timestamp 1730493024
transform -1 0 3680 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1142_
timestamp 1730493024
transform -1 0 3680 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1143_
timestamp 1730493024
transform 1 0 3956 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1144_
timestamp 1730493024
transform 1 0 4416 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1145_
timestamp 1730493024
transform 1 0 4600 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1146_
timestamp 1730493024
transform 1 0 2852 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1147_
timestamp 1730493024
transform -1 0 4784 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1148_
timestamp 1730493024
transform 1 0 3864 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1149_
timestamp 1730493024
transform 1 0 2208 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1150_
timestamp 1730493024
transform 1 0 2208 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1151_
timestamp 1730493024
transform 1 0 4508 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1152_
timestamp 1730493024
transform -1 0 5704 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1153_
timestamp 1730493024
transform -1 0 3128 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1154_
timestamp 1730493024
transform -1 0 5244 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1155_
timestamp 1730493024
transform 1 0 3772 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1156_
timestamp 1730493024
transform 1 0 3036 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1157_
timestamp 1730493024
transform 1 0 7360 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1158_
timestamp 1730493024
transform 1 0 7176 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1159_
timestamp 1730493024
transform 1 0 4784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1160_
timestamp 1730493024
transform 1 0 4692 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1161_
timestamp 1730493024
transform 1 0 5336 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1162_
timestamp 1730493024
transform 1 0 2760 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1163_
timestamp 1730493024
transform 1 0 3772 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1164_
timestamp 1730493024
transform 1 0 12604 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1165_
timestamp 1730493024
transform 1 0 14076 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1166_
timestamp 1730493024
transform -1 0 14076 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1167_
timestamp 1730493024
transform -1 0 13984 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1168_
timestamp 1730493024
transform -1 0 13984 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1169_
timestamp 1730493024
transform -1 0 13432 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1170_
timestamp 1730493024
transform 1 0 9844 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1171_
timestamp 1730493024
transform 1 0 8924 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1172_
timestamp 1730493024
transform 1 0 7636 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1173_
timestamp 1730493024
transform 1 0 6072 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1174_
timestamp 1730493024
transform 1 0 6348 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1175_
timestamp 1730493024
transform 1 0 6624 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1176_
timestamp 1730493024
transform 1 0 8372 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1177_
timestamp 1730493024
transform 1 0 14812 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1178_
timestamp 1730493024
transform 1 0 1380 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1179_
timestamp 1730493024
transform -1 0 10948 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1180_
timestamp 1730493024
transform -1 0 11408 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1181_
timestamp 1730493024
transform -1 0 11408 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1182_
timestamp 1730493024
transform -1 0 11316 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1183_
timestamp 1730493024
transform -1 0 13524 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1184_
timestamp 1730493024
transform -1 0 12052 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1185_
timestamp 1730493024
transform -1 0 11316 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1186_
timestamp 1730493024
transform 1 0 14352 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1187_
timestamp 1730493024
transform 1 0 14720 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1188_
timestamp 1730493024
transform 1 0 14720 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1189_
timestamp 1730493024
transform 1 0 14536 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1190_
timestamp 1730493024
transform 1 0 8924 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1191_
timestamp 1730493024
transform 1 0 14536 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1192_
timestamp 1730493024
transform 1 0 9936 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1193_
timestamp 1730493024
transform 1 0 9844 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1194_
timestamp 1730493024
transform 1 0 9844 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1195_
timestamp 1730493024
transform 1 0 1380 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1196_
timestamp 1730493024
transform 1 0 2300 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1197_
timestamp 1730493024
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1198_
timestamp 1730493024
transform -1 0 10580 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1199_
timestamp 1730493024
transform 1 0 10488 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1200_
timestamp 1730493024
transform 1 0 1380 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1201_
timestamp 1730493024
transform 1 0 4140 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1202_
timestamp 1730493024
transform 1 0 10120 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1203_
timestamp 1730493024
transform -1 0 13892 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1204_
timestamp 1730493024
transform 1 0 3680 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1205_
timestamp 1730493024
transform 1 0 1932 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1206_
timestamp 1730493024
transform -1 0 13340 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1207_
timestamp 1730493024
transform 1 0 14812 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _1208_ ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 16192 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1730493024
transform -1 0 15824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1210_
timestamp 1730493024
transform -1 0 16192 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1730493024
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1212_
timestamp 1730493024
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1730493024
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1214_
timestamp 1730493024
transform -1 0 16192 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1215_
timestamp 1730493024
transform -1 0 16192 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 8924 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_clk ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 4784 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_clk
timestamp 1730493024
transform 1 0 6348 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_clk
timestamp 1730493024
transform 1 0 4140 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_clk
timestamp 1730493024
transform 1 0 6532 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_clk
timestamp 1730493024
transform -1 0 10764 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_clk
timestamp 1730493024
transform 1 0 12236 0 -1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_clk
timestamp 1730493024
transform 1 0 10580 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_clk
timestamp 1730493024
transform 1 0 12420 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_clk
timestamp 1730493024
transform 1 0 4692 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_clk
timestamp 1730493024
transform 1 0 6532 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_clk
timestamp 1730493024
transform -1 0 5336 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_clk
timestamp 1730493024
transform -1 0 6992 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_clk
timestamp 1730493024
transform -1 0 11040 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_clk
timestamp 1730493024
transform 1 0 11868 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_clk
timestamp 1730493024
transform 1 0 10028 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_clk
timestamp 1730493024
transform 1 0 12144 0 -1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkload0
timestamp 1730493024
transform 1 0 3772 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_4  clkload1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 6256 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  clkload2 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 6532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkinvlp_4  clkload3 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 9752 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  clkload4
timestamp 1730493024
transform -1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_4  clkload5
timestamp 1730493024
transform 1 0 11500 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__bufinv_16  clkload6 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12420 0 -1 11968
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinvlp_4  clkload7
timestamp 1730493024
transform 1 0 4692 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_4  clkload8
timestamp 1730493024
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  clkload9 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 4324 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload10 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 5980 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload11
timestamp 1730493024
transform 1 0 10028 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_6  clkload12
timestamp 1730493024
transform -1 0 11868 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_8  clkload13
timestamp 1730493024
transform 1 0 10028 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  clkload14
timestamp 1730493024
transform 1 0 12144 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  fanout58 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 3864 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 1730493024
transform -1 0 8740 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout60
timestamp 1730493024
transform -1 0 9660 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 1730493024
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout63
timestamp 1730493024
transform -1 0 8188 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout64 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 8832 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout65 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout66
timestamp 1730493024
transform 1 0 8924 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout69
timestamp 1730493024
transform 1 0 11408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout70
timestamp 1730493024
transform -1 0 9292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  fanout71
timestamp 1730493024
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  fanout72
timestamp 1730493024
transform 1 0 8096 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout73
timestamp 1730493024
transform 1 0 9660 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout74
timestamp 1730493024
transform -1 0 8188 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout75
timestamp 1730493024
transform 1 0 3404 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout76
timestamp 1730493024
transform -1 0 2760 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout77
timestamp 1730493024
transform -1 0 10396 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout78 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 15456 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout79 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 11500 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout80
timestamp 1730493024
transform -1 0 3312 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  fanout81
timestamp 1730493024
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout82
timestamp 1730493024
transform -1 0 10856 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout83
timestamp 1730493024
transform -1 0 11408 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout84
timestamp 1730493024
transform 1 0 11500 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1730493024
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1730493024
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 4324 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1730493024
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1730493024
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_91 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_98
timestamp 1730493024
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_105
timestamp 1730493024
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1730493024
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp 1730493024
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_126
timestamp 1730493024
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_133
timestamp 1730493024
transform 1 0 13340 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_151
timestamp 1730493024
transform 1 0 14996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1730493024
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_10
timestamp 1730493024
transform 1 0 2024 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1730493024
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1730493024
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_74
timestamp 1730493024
transform 1 0 7912 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_120
timestamp 1730493024
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_144
timestamp 1730493024
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1730493024
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1730493024
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_12
timestamp 1730493024
transform 1 0 2208 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1730493024
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1730493024
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62
timestamp 1730493024
transform 1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_72 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 7728 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1730493024
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_89
timestamp 1730493024
transform 1 0 9292 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1730493024
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1730493024
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1730493024
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_7
timestamp 1730493024
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1730493024
transform 1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_31
timestamp 1730493024
transform 1 0 3956 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_38 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 4600 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_50 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 5704 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_57
timestamp 1730493024
transform 1 0 6348 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_68
timestamp 1730493024
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_78
timestamp 1730493024
transform 1 0 8280 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_90 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 9384 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_98
timestamp 1730493024
transform 1 0 10120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_133
timestamp 1730493024
transform 1 0 13340 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_137
timestamp 1730493024
transform 1 0 13708 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_153
timestamp 1730493024
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1730493024
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1730493024
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1730493024
transform 1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_74
timestamp 1730493024
transform 1 0 7912 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_78
timestamp 1730493024
transform 1 0 8280 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_93
timestamp 1730493024
transform 1 0 9660 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_101
timestamp 1730493024
transform 1 0 10396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_113
timestamp 1730493024
transform 1 0 11500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_125
timestamp 1730493024
transform 1 0 12604 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1730493024
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_149
timestamp 1730493024
transform 1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1730493024
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 1730493024
transform 1 0 4140 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_42
timestamp 1730493024
transform 1 0 4968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1730493024
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_5_79
timestamp 1730493024
transform 1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_98
timestamp 1730493024
transform 1 0 10120 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1730493024
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_130
timestamp 1730493024
transform 1 0 13064 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_134
timestamp 1730493024
transform 1 0 13432 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_158
timestamp 1730493024
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1730493024
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1730493024
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1730493024
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_17
timestamp 1730493024
transform 1 0 2668 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1730493024
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1730493024
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1730493024
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1730493024
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1730493024
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_72
timestamp 1730493024
transform 1 0 7728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_76
timestamp 1730493024
transform 1 0 8096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1730493024
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1730493024
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1730493024
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_147
timestamp 1730493024
transform 1 0 14628 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_159
timestamp 1730493024
transform 1 0 15732 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_163
timestamp 1730493024
transform 1 0 16100 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1730493024
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_15
timestamp 1730493024
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_29
timestamp 1730493024
transform 1 0 3772 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1730493024
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1730493024
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1730493024
transform 1 0 8556 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_93
timestamp 1730493024
transform 1 0 9660 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_113
timestamp 1730493024
transform 1 0 11500 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1730493024
transform 1 0 12236 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_133
timestamp 1730493024
transform 1 0 13340 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_137
timestamp 1730493024
transform 1 0 13708 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1730493024
transform 1 0 14904 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_8_3
timestamp 1730493024
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1730493024
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1730493024
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_34
timestamp 1730493024
transform 1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_49
timestamp 1730493024
transform 1 0 5612 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1730493024
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1730493024
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1730493024
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_112
timestamp 1730493024
transform 1 0 11408 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_124
timestamp 1730493024
transform 1 0 12512 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_132
timestamp 1730493024
transform 1 0 13248 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1730493024
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_167
timestamp 1730493024
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1730493024
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_25
timestamp 1730493024
transform 1 0 3404 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1730493024
transform 1 0 4140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_37
timestamp 1730493024
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_45
timestamp 1730493024
transform 1 0 5244 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1730493024
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_57
timestamp 1730493024
transform 1 0 6348 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_68
timestamp 1730493024
transform 1 0 7360 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_74
timestamp 1730493024
transform 1 0 7912 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_90
timestamp 1730493024
transform 1 0 9384 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1730493024
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1730493024
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_137
timestamp 1730493024
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_156
timestamp 1730493024
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1730493024
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1730493024
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_44
timestamp 1730493024
transform 1 0 5152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_56
timestamp 1730493024
transform 1 0 6256 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1730493024
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1730493024
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_122
timestamp 1730493024
transform 1 0 12328 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1730493024
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_157
timestamp 1730493024
transform 1 0 15548 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_165
timestamp 1730493024
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_3
timestamp 1730493024
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_90
timestamp 1730493024
transform 1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_100
timestamp 1730493024
transform 1 0 10304 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1730493024
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1730493024
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1730493024
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_148
timestamp 1730493024
transform 1 0 14720 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1730493024
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 1730493024
transform 1 0 1748 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_21
timestamp 1730493024
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1730493024
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 1730493024
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1730493024
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1730493024
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_103
timestamp 1730493024
transform 1 0 10580 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1730493024
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1730493024
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_149
timestamp 1730493024
transform 1 0 14812 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_161
timestamp 1730493024
transform 1 0 15916 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1730493024
transform 1 0 16468 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_11
timestamp 1730493024
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_23
timestamp 1730493024
transform 1 0 3220 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_45
timestamp 1730493024
transform 1 0 5244 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_57
timestamp 1730493024
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_65
timestamp 1730493024
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1730493024
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1730493024
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1730493024
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1730493024
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1730493024
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_144
timestamp 1730493024
transform 1 0 14352 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_156
timestamp 1730493024
transform 1 0 15456 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_164
timestamp 1730493024
transform 1 0 16192 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1730493024
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_47
timestamp 1730493024
transform 1 0 5428 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_59
timestamp 1730493024
transform 1 0 6532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_71
timestamp 1730493024
transform 1 0 7636 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1730493024
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1730493024
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_149
timestamp 1730493024
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_167
timestamp 1730493024
transform 1 0 16468 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1730493024
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1730493024
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_81
timestamp 1730493024
transform 1 0 8556 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_102
timestamp 1730493024
transform 1 0 10488 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1730493024
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_129
timestamp 1730493024
transform 1 0 12972 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_145
timestamp 1730493024
transform 1 0 14444 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1730493024
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1730493024
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1730493024
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_34
timestamp 1730493024
transform 1 0 4232 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_43
timestamp 1730493024
transform 1 0 5060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1730493024
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1730493024
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_85
timestamp 1730493024
transform 1 0 8924 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_102
timestamp 1730493024
transform 1 0 10488 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_148
timestamp 1730493024
transform 1 0 14720 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 1730493024
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_11
timestamp 1730493024
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1730493024
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_79
timestamp 1730493024
transform 1 0 8372 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_92
timestamp 1730493024
transform 1 0 9568 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1730493024
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_11
timestamp 1730493024
transform 1 0 2116 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_18
timestamp 1730493024
transform 1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1730493024
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_42
timestamp 1730493024
transform 1 0 4968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_62
timestamp 1730493024
transform 1 0 6808 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_77
timestamp 1730493024
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1730493024
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp 1730493024
transform 1 0 13432 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1730493024
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_162
timestamp 1730493024
transform 1 0 16008 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1730493024
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_35
timestamp 1730493024
transform 1 0 4324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_47
timestamp 1730493024
transform 1 0 5428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1730493024
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1730493024
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_73
timestamp 1730493024
transform 1 0 7820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_84
timestamp 1730493024
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1730493024
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_122
timestamp 1730493024
transform 1 0 12328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_128
timestamp 1730493024
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_20
timestamp 1730493024
transform 1 0 2944 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_46
timestamp 1730493024
transform 1 0 5336 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_93
timestamp 1730493024
transform 1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1730493024
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1730493024
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1730493024
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_150
timestamp 1730493024
transform 1 0 14904 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1730493024
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_22
timestamp 1730493024
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1730493024
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 1730493024
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_70
timestamp 1730493024
transform 1 0 7544 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 1730493024
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1730493024
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_146
timestamp 1730493024
transform 1 0 14536 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_150
timestamp 1730493024
transform 1 0 14904 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1730493024
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_12
timestamp 1730493024
transform 1 0 2208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_20
timestamp 1730493024
transform 1 0 2944 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_29
timestamp 1730493024
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1730493024
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_51
timestamp 1730493024
transform 1 0 5796 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1730493024
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_94
timestamp 1730493024
transform 1 0 9752 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_134
timestamp 1730493024
transform 1 0 13432 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1730493024
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1730493024
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 1730493024
transform 1 0 14628 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1730493024
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1730493024
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_32
timestamp 1730493024
transform 1 0 4048 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_50
timestamp 1730493024
transform 1 0 5704 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_73
timestamp 1730493024
transform 1 0 7820 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_90
timestamp 1730493024
transform 1 0 9384 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1730493024
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_141
timestamp 1730493024
transform 1 0 14076 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_149
timestamp 1730493024
transform 1 0 14812 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1730493024
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_3
timestamp 1730493024
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_7
timestamp 1730493024
transform 1 0 1748 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1730493024
transform 1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_29
timestamp 1730493024
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1730493024
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_53
timestamp 1730493024
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1730493024
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_99
timestamp 1730493024
transform 1 0 10212 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_124
timestamp 1730493024
transform 1 0 12512 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_130
timestamp 1730493024
transform 1 0 13064 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1730493024
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1730493024
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_27
timestamp 1730493024
transform 1 0 3588 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_31
timestamp 1730493024
transform 1 0 3956 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_41
timestamp 1730493024
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1730493024
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_79
timestamp 1730493024
transform 1 0 8372 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_104
timestamp 1730493024
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_113
timestamp 1730493024
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_128
timestamp 1730493024
transform 1 0 12880 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_139
timestamp 1730493024
transform 1 0 13892 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_151
timestamp 1730493024
transform 1 0 14996 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_3
timestamp 1730493024
transform 1 0 1380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_11
timestamp 1730493024
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_24
timestamp 1730493024
transform 1 0 3312 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1730493024
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_48
timestamp 1730493024
transform 1 0 5520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1730493024
transform 1 0 6256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_73
timestamp 1730493024
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_81
timestamp 1730493024
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_94
timestamp 1730493024
transform 1 0 9752 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_126
timestamp 1730493024
transform 1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1730493024
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_150
timestamp 1730493024
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_164
timestamp 1730493024
transform 1 0 16192 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1730493024
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_7
timestamp 1730493024
transform 1 0 1748 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_34
timestamp 1730493024
transform 1 0 4232 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_66
timestamp 1730493024
transform 1 0 7176 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_91
timestamp 1730493024
transform 1 0 9476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1730493024
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_121
timestamp 1730493024
transform 1 0 12236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_133
timestamp 1730493024
transform 1 0 13340 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1730493024
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_147
timestamp 1730493024
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_20
timestamp 1730493024
transform 1 0 2944 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1730493024
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_29
timestamp 1730493024
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_39
timestamp 1730493024
transform 1 0 4692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1730493024
transform 1 0 5796 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1730493024
transform 1 0 7268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_71
timestamp 1730493024
transform 1 0 7636 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1730493024
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1730493024
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1730493024
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_109
timestamp 1730493024
transform 1 0 11132 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_122
timestamp 1730493024
transform 1 0 12328 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1730493024
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1730493024
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_149
timestamp 1730493024
transform 1 0 14812 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_157
timestamp 1730493024
transform 1 0 15548 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1730493024
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1730493024
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_22
timestamp 1730493024
transform 1 0 3128 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_45
timestamp 1730493024
transform 1 0 5244 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1730493024
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_72
timestamp 1730493024
transform 1 0 7728 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_84
timestamp 1730493024
transform 1 0 8832 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_90
timestamp 1730493024
transform 1 0 9384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1730493024
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1730493024
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_120
timestamp 1730493024
transform 1 0 12144 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_128
timestamp 1730493024
transform 1 0 12880 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1730493024
transform 1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_151
timestamp 1730493024
transform 1 0 14996 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_163
timestamp 1730493024
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1730493024
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1730493024
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_23
timestamp 1730493024
transform 1 0 3220 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1730493024
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1730493024
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_41
timestamp 1730493024
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_69
timestamp 1730493024
transform 1 0 7452 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_94
timestamp 1730493024
transform 1 0 9752 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_102
timestamp 1730493024
transform 1 0 10488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_113
timestamp 1730493024
transform 1 0 11500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_125
timestamp 1730493024
transform 1 0 12604 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_131
timestamp 1730493024
transform 1 0 13156 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1730493024
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1730493024
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_152
timestamp 1730493024
transform 1 0 15088 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_164
timestamp 1730493024
transform 1 0 16192 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_30
timestamp 1730493024
transform 1 0 3864 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_42
timestamp 1730493024
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1730493024
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_57
timestamp 1730493024
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_63
timestamp 1730493024
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_122
timestamp 1730493024
transform 1 0 12328 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_126
timestamp 1730493024
transform 1 0 12696 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_149
timestamp 1730493024
transform 1 0 14812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_159
timestamp 1730493024
transform 1 0 15732 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1730493024
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1730493024
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_20
timestamp 1730493024
transform 1 0 2944 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_45
timestamp 1730493024
transform 1 0 5244 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_53
timestamp 1730493024
transform 1 0 5980 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_57
timestamp 1730493024
transform 1 0 6348 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_73
timestamp 1730493024
transform 1 0 7820 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_85
timestamp 1730493024
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_119
timestamp 1730493024
transform 1 0 12052 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp 1730493024
transform 1 0 12788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1730493024
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_141
timestamp 1730493024
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_145
timestamp 1730493024
transform 1 0 14444 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_162
timestamp 1730493024
transform 1 0 16008 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1730493024
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_16
timestamp 1730493024
transform 1 0 2576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_24
timestamp 1730493024
transform 1 0 3312 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_29
timestamp 1730493024
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1730493024
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_92
timestamp 1730493024
transform 1 0 9568 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1730493024
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_117
timestamp 1730493024
transform 1 0 11868 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_129
timestamp 1730493024
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_147
timestamp 1730493024
transform 1 0 14628 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_155
timestamp 1730493024
transform 1 0 15364 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1730493024
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1730493024
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_43
timestamp 1730493024
transform 1 0 5060 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_47
timestamp 1730493024
transform 1 0 5428 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_71
timestamp 1730493024
transform 1 0 7636 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_105
timestamp 1730493024
transform 1 0 10764 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_113
timestamp 1730493024
transform 1 0 11500 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_118
timestamp 1730493024
transform 1 0 11960 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1730493024
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_146
timestamp 1730493024
transform 1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_158
timestamp 1730493024
transform 1 0 15640 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_164
timestamp 1730493024
transform 1 0 16192 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_3
timestamp 1730493024
transform 1 0 1380 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_37
timestamp 1730493024
transform 1 0 4508 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1730493024
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_62
timestamp 1730493024
transform 1 0 6808 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_75
timestamp 1730493024
transform 1 0 8004 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_87
timestamp 1730493024
transform 1 0 9108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_91
timestamp 1730493024
transform 1 0 9476 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_101
timestamp 1730493024
transform 1 0 10396 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_105
timestamp 1730493024
transform 1 0 10764 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_121
timestamp 1730493024
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_136
timestamp 1730493024
transform 1 0 13616 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_21
timestamp 1730493024
transform 1 0 3036 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1730493024
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1730493024
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1730493024
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_45
timestamp 1730493024
transform 1 0 5244 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_85
timestamp 1730493024
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_36_117
timestamp 1730493024
transform 1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1730493024
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1730493024
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_153
timestamp 1730493024
transform 1 0 15180 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_7
timestamp 1730493024
transform 1 0 1748 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_19
timestamp 1730493024
transform 1 0 2852 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_43
timestamp 1730493024
transform 1 0 5060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_57
timestamp 1730493024
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_96
timestamp 1730493024
transform 1 0 9936 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1730493024
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_113
timestamp 1730493024
transform 1 0 11500 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_37_117
timestamp 1730493024
transform 1 0 11868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1730493024
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_127
timestamp 1730493024
transform 1 0 12788 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_134
timestamp 1730493024
transform 1 0 13432 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_146
timestamp 1730493024
transform 1 0 14536 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_158
timestamp 1730493024
transform 1 0 15640 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_38_3
timestamp 1730493024
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_38_53
timestamp 1730493024
transform 1 0 5980 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_62
timestamp 1730493024
transform 1 0 6808 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_74
timestamp 1730493024
transform 1 0 7912 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1730493024
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_101
timestamp 1730493024
transform 1 0 10396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1730493024
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1730493024
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1730493024
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1730493024
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_165
timestamp 1730493024
transform 1 0 16284 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1730493024
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_15
timestamp 1730493024
transform 1 0 2484 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_37
timestamp 1730493024
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1730493024
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1730493024
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1730493024
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_80
timestamp 1730493024
transform 1 0 8464 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_88
timestamp 1730493024
transform 1 0 9200 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1730493024
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_113
timestamp 1730493024
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_133
timestamp 1730493024
transform 1 0 13340 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_145
timestamp 1730493024
transform 1 0 14444 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_157
timestamp 1730493024
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1730493024
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1730493024
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1730493024
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1730493024
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_29
timestamp 1730493024
transform 1 0 3772 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_40
timestamp 1730493024
transform 1 0 4784 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_46
timestamp 1730493024
transform 1 0 5336 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1730493024
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_91
timestamp 1730493024
transform 1 0 9476 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_103
timestamp 1730493024
transform 1 0 10580 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_123
timestamp 1730493024
transform 1 0 12420 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_135
timestamp 1730493024
transform 1 0 13524 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1730493024
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1730493024
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1730493024
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_165
timestamp 1730493024
transform 1 0 16284 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1730493024
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1730493024
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_27
timestamp 1730493024
transform 1 0 3588 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1730493024
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_91
timestamp 1730493024
transform 1 0 9476 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_103
timestamp 1730493024
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1730493024
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1730493024
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1730493024
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1730493024
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1730493024
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1730493024
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1730493024
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1730493024
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1730493024
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1730493024
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_82
timestamp 1730493024
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_104
timestamp 1730493024
transform 1 0 10672 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_112
timestamp 1730493024
transform 1 0 11408 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1730493024
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1730493024
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1730493024
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1730493024
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1730493024
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_165
timestamp 1730493024
transform 1 0 16284 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1730493024
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1730493024
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_27
timestamp 1730493024
transform 1 0 3588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_43_37
timestamp 1730493024
transform 1 0 4508 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_46
timestamp 1730493024
transform 1 0 5336 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_61
timestamp 1730493024
transform 1 0 6716 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_75
timestamp 1730493024
transform 1 0 8004 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_92
timestamp 1730493024
transform 1 0 9568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_113
timestamp 1730493024
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_131
timestamp 1730493024
transform 1 0 13156 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_143
timestamp 1730493024
transform 1 0 14260 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_155
timestamp 1730493024
transform 1 0 15364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1730493024
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1730493024
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1730493024
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1730493024
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_29
timestamp 1730493024
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_37
timestamp 1730493024
transform 1 0 4508 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_49
timestamp 1730493024
transform 1 0 5612 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_53
timestamp 1730493024
transform 1 0 5980 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_70
timestamp 1730493024
transform 1 0 7544 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_82
timestamp 1730493024
transform 1 0 8648 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_89
timestamp 1730493024
transform 1 0 9292 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_108
timestamp 1730493024
transform 1 0 11040 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_112
timestamp 1730493024
transform 1 0 11408 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_123
timestamp 1730493024
transform 1 0 12420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_132
timestamp 1730493024
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1730493024
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1730493024
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_165
timestamp 1730493024
transform 1 0 16284 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_7
timestamp 1730493024
transform 1 0 1748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_15
timestamp 1730493024
transform 1 0 2484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_24
timestamp 1730493024
transform 1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_45_53
timestamp 1730493024
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1730493024
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_88
timestamp 1730493024
transform 1 0 9200 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_96
timestamp 1730493024
transform 1 0 9936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_104
timestamp 1730493024
transform 1 0 10672 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1730493024
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_45_120
timestamp 1730493024
transform 1 0 12144 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_147
timestamp 1730493024
transform 1 0 14628 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_159
timestamp 1730493024
transform 1 0 15732 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1730493024
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_3
timestamp 1730493024
transform 1 0 1380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_11
timestamp 1730493024
transform 1 0 2116 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_29
timestamp 1730493024
transform 1 0 3772 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_58
timestamp 1730493024
transform 1 0 6440 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_78
timestamp 1730493024
transform 1 0 8280 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_108
timestamp 1730493024
transform 1 0 11040 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_118
timestamp 1730493024
transform 1 0 11960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_130
timestamp 1730493024
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1730493024
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1730493024
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1730493024
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_165
timestamp 1730493024
transform 1 0 16284 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1730493024
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_15
timestamp 1730493024
transform 1 0 2484 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_66
timestamp 1730493024
transform 1 0 7176 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_71
timestamp 1730493024
transform 1 0 7636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_75
timestamp 1730493024
transform 1 0 8004 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_99
timestamp 1730493024
transform 1 0 10212 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1730493024
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_119
timestamp 1730493024
transform 1 0 12052 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_139
timestamp 1730493024
transform 1 0 13892 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_151
timestamp 1730493024
transform 1 0 14996 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_163
timestamp 1730493024
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1730493024
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1730493024
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1730493024
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1730493024
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_48_29
timestamp 1730493024
transform 1 0 3772 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_35
timestamp 1730493024
transform 1 0 4324 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_67
timestamp 1730493024
transform 1 0 7268 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_79
timestamp 1730493024
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1730493024
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1730493024
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_97
timestamp 1730493024
transform 1 0 10028 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_138
timestamp 1730493024
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_144
timestamp 1730493024
transform 1 0 14352 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_156
timestamp 1730493024
transform 1 0 15456 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1730493024
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_22
timestamp 1730493024
transform 1 0 3128 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_28
timestamp 1730493024
transform 1 0 3680 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1730493024
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1730493024
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_73
timestamp 1730493024
transform 1 0 7820 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_77
timestamp 1730493024
transform 1 0 8188 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_84
timestamp 1730493024
transform 1 0 8832 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_96
timestamp 1730493024
transform 1 0 9936 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_150
timestamp 1730493024
transform 1 0 14904 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_162
timestamp 1730493024
transform 1 0 16008 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1730493024
transform 1 0 1380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_11
timestamp 1730493024
transform 1 0 2116 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_35
timestamp 1730493024
transform 1 0 4324 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_50_49
timestamp 1730493024
transform 1 0 5612 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_50_57
timestamp 1730493024
transform 1 0 6348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_65
timestamp 1730493024
transform 1 0 7084 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_75
timestamp 1730493024
transform 1 0 8004 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_113
timestamp 1730493024
transform 1 0 11500 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_125
timestamp 1730493024
transform 1 0 12604 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_50_137
timestamp 1730493024
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1730493024
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1730493024
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_165
timestamp 1730493024
transform 1 0 16284 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1730493024
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_15
timestamp 1730493024
transform 1 0 2484 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_19
timestamp 1730493024
transform 1 0 2852 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_46
timestamp 1730493024
transform 1 0 5336 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1730493024
transform 1 0 6072 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1730493024
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_69
timestamp 1730493024
transform 1 0 7452 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_77
timestamp 1730493024
transform 1 0 8188 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_96
timestamp 1730493024
transform 1 0 9936 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_104
timestamp 1730493024
transform 1 0 10672 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1730493024
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_113
timestamp 1730493024
transform 1 0 11500 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_120
timestamp 1730493024
transform 1 0 12144 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_129
timestamp 1730493024
transform 1 0 12972 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_142
timestamp 1730493024
transform 1 0 14168 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_154
timestamp 1730493024
transform 1 0 15272 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1730493024
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1730493024
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1730493024
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1730493024
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_32
timestamp 1730493024
transform 1 0 4048 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_40
timestamp 1730493024
transform 1 0 4784 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_48
timestamp 1730493024
transform 1 0 5520 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_56
timestamp 1730493024
transform 1 0 6256 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_52_67
timestamp 1730493024
transform 1 0 7268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_78
timestamp 1730493024
transform 1 0 8280 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1730493024
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_126
timestamp 1730493024
transform 1 0 12696 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1730493024
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_157
timestamp 1730493024
transform 1 0 15548 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_165
timestamp 1730493024
transform 1 0 16284 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1730493024
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_15
timestamp 1730493024
transform 1 0 2484 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_23
timestamp 1730493024
transform 1 0 3220 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_40
timestamp 1730493024
transform 1 0 4784 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_48
timestamp 1730493024
transform 1 0 5520 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_52
timestamp 1730493024
transform 1 0 5888 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_57
timestamp 1730493024
transform 1 0 6348 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_90
timestamp 1730493024
transform 1 0 9384 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_99
timestamp 1730493024
transform 1 0 10212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1730493024
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1730493024
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_125
timestamp 1730493024
transform 1 0 12604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_129
timestamp 1730493024
transform 1 0 12972 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_146
timestamp 1730493024
transform 1 0 14536 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_158
timestamp 1730493024
transform 1 0 15640 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_166
timestamp 1730493024
transform 1 0 16376 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1730493024
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1730493024
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1730493024
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_41
timestamp 1730493024
transform 1 0 4876 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_57
timestamp 1730493024
transform 1 0 6348 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_66
timestamp 1730493024
transform 1 0 7176 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_72
timestamp 1730493024
transform 1 0 7728 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_85
timestamp 1730493024
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_97
timestamp 1730493024
transform 1 0 10028 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_114
timestamp 1730493024
transform 1 0 11592 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1730493024
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1730493024
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1730493024
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1730493024
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_165
timestamp 1730493024
transform 1 0 16284 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1730493024
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_15
timestamp 1730493024
transform 1 0 2484 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1730493024
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1730493024
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1730493024
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1730493024
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_93
timestamp 1730493024
transform 1 0 9660 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_106
timestamp 1730493024
transform 1 0 10856 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_119
timestamp 1730493024
transform 1 0 12052 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_131
timestamp 1730493024
transform 1 0 13156 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_143
timestamp 1730493024
transform 1 0 14260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_155
timestamp 1730493024
transform 1 0 15364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1730493024
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1730493024
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_15
timestamp 1730493024
transform 1 0 2484 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_19
timestamp 1730493024
transform 1 0 2852 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1730493024
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_44
timestamp 1730493024
transform 1 0 5152 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_115
timestamp 1730493024
transform 1 0 11684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_119
timestamp 1730493024
transform 1 0 12052 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_132
timestamp 1730493024
transform 1 0 13248 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1730493024
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1730493024
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_165
timestamp 1730493024
transform 1 0 16284 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1730493024
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_15
timestamp 1730493024
transform 1 0 2484 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_54
timestamp 1730493024
transform 1 0 6072 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_100
timestamp 1730493024
transform 1 0 10304 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_106
timestamp 1730493024
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_121
timestamp 1730493024
transform 1 0 12236 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_141
timestamp 1730493024
transform 1 0 14076 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_153
timestamp 1730493024
transform 1 0 15180 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1730493024
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1730493024
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1730493024
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1730493024
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_29
timestamp 1730493024
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_35
timestamp 1730493024
transform 1 0 4324 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_46
timestamp 1730493024
transform 1 0 5336 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_52
timestamp 1730493024
transform 1 0 5888 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_78
timestamp 1730493024
transform 1 0 8280 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_93
timestamp 1730493024
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_111
timestamp 1730493024
transform 1 0 11316 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_115
timestamp 1730493024
transform 1 0 11684 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_157
timestamp 1730493024
transform 1 0 15548 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_165
timestamp 1730493024
transform 1 0 16284 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1730493024
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_15
timestamp 1730493024
transform 1 0 2484 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_22
timestamp 1730493024
transform 1 0 3128 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_34
timestamp 1730493024
transform 1 0 4232 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_46
timestamp 1730493024
transform 1 0 5336 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_54
timestamp 1730493024
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_57
timestamp 1730493024
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_65
timestamp 1730493024
transform 1 0 7084 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_71
timestamp 1730493024
transform 1 0 7636 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_83
timestamp 1730493024
transform 1 0 8740 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_95
timestamp 1730493024
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1730493024
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1730493024
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_113
timestamp 1730493024
transform 1 0 11500 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_59_122
timestamp 1730493024
transform 1 0 12328 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_133
timestamp 1730493024
transform 1 0 13340 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_145
timestamp 1730493024
transform 1 0 14444 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_157
timestamp 1730493024
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_165
timestamp 1730493024
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_3
timestamp 1730493024
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_11
timestamp 1730493024
transform 1 0 2116 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_52
timestamp 1730493024
transform 1 0 5888 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_59
timestamp 1730493024
transform 1 0 6532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_76
timestamp 1730493024
transform 1 0 8096 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1730493024
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_92
timestamp 1730493024
transform 1 0 9568 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_105
timestamp 1730493024
transform 1 0 10764 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_115
timestamp 1730493024
transform 1 0 11684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_129
timestamp 1730493024
transform 1 0 12972 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_137
timestamp 1730493024
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1730493024
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1730493024
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_165
timestamp 1730493024
transform 1 0 16284 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1730493024
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_15
timestamp 1730493024
transform 1 0 2484 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_24
timestamp 1730493024
transform 1 0 3312 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_36
timestamp 1730493024
transform 1 0 4416 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_44
timestamp 1730493024
transform 1 0 5152 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_52
timestamp 1730493024
transform 1 0 5888 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1730493024
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_104
timestamp 1730493024
transform 1 0 10672 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_141
timestamp 1730493024
transform 1 0 14076 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_153
timestamp 1730493024
transform 1 0 15180 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_165
timestamp 1730493024
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_3
timestamp 1730493024
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_62_29
timestamp 1730493024
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_65
timestamp 1730493024
transform 1 0 7084 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1730493024
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1730493024
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_91
timestamp 1730493024
transform 1 0 9476 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_99
timestamp 1730493024
transform 1 0 10212 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_116
timestamp 1730493024
transform 1 0 11776 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1730493024
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1730493024
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_165
timestamp 1730493024
transform 1 0 16284 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1730493024
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_15
timestamp 1730493024
transform 1 0 2484 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_23
timestamp 1730493024
transform 1 0 3220 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_47
timestamp 1730493024
transform 1 0 5428 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1730493024
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_73
timestamp 1730493024
transform 1 0 7820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_85
timestamp 1730493024
transform 1 0 8924 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_93
timestamp 1730493024
transform 1 0 9660 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_98
timestamp 1730493024
transform 1 0 10120 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_102
timestamp 1730493024
transform 1 0 10488 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_107
timestamp 1730493024
transform 1 0 10948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1730493024
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1730493024
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1730493024
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1730493024
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1730493024
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1730493024
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1730493024
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1730493024
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1730493024
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1730493024
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1730493024
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1730493024
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_53
timestamp 1730493024
transform 1 0 5980 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_66
timestamp 1730493024
transform 1 0 7176 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_78
timestamp 1730493024
transform 1 0 8280 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_64_85
timestamp 1730493024
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_93
timestamp 1730493024
transform 1 0 9660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_112
timestamp 1730493024
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_118
timestamp 1730493024
transform 1 0 11960 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_124
timestamp 1730493024
transform 1 0 12512 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_128
timestamp 1730493024
transform 1 0 12880 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1730493024
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1730493024
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1730493024
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1730493024
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1730493024
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1730493024
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1730493024
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1730493024
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1730493024
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_57
timestamp 1730493024
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_65_86
timestamp 1730493024
transform 1 0 9016 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_98
timestamp 1730493024
transform 1 0 10120 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_136
timestamp 1730493024
transform 1 0 13616 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_148
timestamp 1730493024
transform 1 0 14720 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_160
timestamp 1730493024
transform 1 0 15824 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1730493024
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1730493024
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1730493024
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1730493024
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1730493024
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_53
timestamp 1730493024
transform 1 0 5980 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_70
timestamp 1730493024
transform 1 0 7544 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_101
timestamp 1730493024
transform 1 0 10396 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_106
timestamp 1730493024
transform 1 0 10856 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_111
timestamp 1730493024
transform 1 0 11316 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_122
timestamp 1730493024
transform 1 0 12328 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1730493024
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1730493024
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_165
timestamp 1730493024
transform 1 0 16284 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_67_3
timestamp 1730493024
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_15
timestamp 1730493024
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_27
timestamp 1730493024
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_39
timestamp 1730493024
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_51
timestamp 1730493024
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1730493024
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_57
timestamp 1730493024
transform 1 0 6348 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_67_87
timestamp 1730493024
transform 1 0 9108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1730493024
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_113
timestamp 1730493024
transform 1 0 11500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_117
timestamp 1730493024
transform 1 0 11868 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_134
timestamp 1730493024
transform 1 0 13432 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_146
timestamp 1730493024
transform 1 0 14536 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_158
timestamp 1730493024
transform 1 0 15640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1730493024
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1730493024
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1730493024
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1730493024
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1730493024
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1730493024
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_53
timestamp 1730493024
transform 1 0 5980 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_57
timestamp 1730493024
transform 1 0 6348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_69
timestamp 1730493024
transform 1 0 7452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_81
timestamp 1730493024
transform 1 0 8556 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1730493024
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_102
timestamp 1730493024
transform 1 0 10488 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_111
timestamp 1730493024
transform 1 0 11316 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_113
timestamp 1730493024
transform 1 0 11500 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_125
timestamp 1730493024
transform 1 0 12604 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_132
timestamp 1730493024
transform 1 0 13248 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1730493024
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1730493024
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_165
timestamp 1730493024
transform 1 0 16284 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform -1 0 10580 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1730493024
transform 1 0 4600 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1730493024
transform 1 0 11316 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1730493024
transform -1 0 3036 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1730493024
transform -1 0 7912 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1730493024
transform -1 0 8832 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1730493024
transform -1 0 11316 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1730493024
transform -1 0 16560 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1730493024
transform -1 0 16560 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1730493024
transform 1 0 14444 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1730493024
transform 1 0 6532 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1730493024
transform -1 0 16560 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1730493024
transform -1 0 16560 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1730493024
transform -1 0 3220 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1730493024
transform 1 0 2208 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1730493024
transform -1 0 16560 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1730493024
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1730493024
transform -1 0 16376 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1730493024
transform 1 0 11592 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1730493024
transform -1 0 16468 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1730493024
transform -1 0 7176 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1730493024
transform -1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1730493024
transform -1 0 9568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1730493024
transform -1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1730493024
transform -1 0 6808 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1730493024
transform -1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1730493024
transform -1 0 7176 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1730493024
transform -1 0 4784 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1730493024
transform 1 0 10120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1730493024
transform -1 0 9660 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1730493024
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1730493024
transform -1 0 11132 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1730493024
transform 1 0 10764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1730493024
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1730493024
transform -1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1730493024
transform -1 0 7728 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1730493024
transform 1 0 6532 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1730493024
transform 1 0 6716 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1730493024
transform 1 0 5060 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1730493024
transform -1 0 6440 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1730493024
transform -1 0 13156 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1730493024
transform -1 0 9660 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1730493024
transform -1 0 12696 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1730493024
transform -1 0 11684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1730493024
transform -1 0 8096 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1730493024
transform 1 0 4048 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1730493024
transform -1 0 4784 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1730493024
transform -1 0 7452 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1730493024
transform -1 0 5980 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1730493024
transform 1 0 2024 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1730493024
transform -1 0 8648 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1730493024
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1730493024
transform 1 0 11316 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1730493024
transform -1 0 7176 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1730493024
transform -1 0 14812 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1730493024
transform -1 0 8464 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1730493024
transform -1 0 11040 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1730493024
transform -1 0 11316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1730493024
transform 1 0 12972 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1730493024
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1730493024
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1730493024
transform 1 0 1380 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1730493024
transform 1 0 3036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1730493024
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap67
timestamp 1730493024
transform 1 0 11040 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  max_cap68
timestamp 1730493024
transform 1 0 10212 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1730493024
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1730493024
transform 1 0 16192 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1730493024
transform 1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1730493024
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1730493024
transform 1 0 16192 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1730493024
transform -1 0 15824 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1730493024
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1730493024
transform 1 0 16192 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1730493024
transform -1 0 2576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1730493024
transform -1 0 2760 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1730493024
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1730493024
transform -1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1730493024
transform -1 0 2392 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1730493024
transform -1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1730493024
transform -1 0 2116 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1730493024
transform -1 0 9476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1730493024
transform -1 0 12696 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1730493024
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1730493024
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1730493024
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1730493024
transform -1 0 2760 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1730493024
transform -1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output30
timestamp 1730493024
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1730493024
transform -1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1730493024
transform -1 0 4784 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1730493024
transform -1 0 13984 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1730493024
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1730493024
transform -1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output36
timestamp 1730493024
transform -1 0 16560 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output37
timestamp 1730493024
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1730493024
transform 1 0 15824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1730493024
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1730493024
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1730493024
transform 1 0 15456 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1730493024
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1730493024
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output44
timestamp 1730493024
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output45
timestamp 1730493024
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1730493024
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1730493024
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1730493024
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1730493024
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1730493024
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1730493024
transform -1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1730493024
transform -1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1730493024
transform -1 0 1748 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1730493024
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1730493024
transform -1 0 2116 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1730493024
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1730493024
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_69
timestamp 1730493024
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1730493024
transform -1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_70
timestamp 1730493024
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1730493024
transform -1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_71
timestamp 1730493024
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1730493024
transform -1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_72
timestamp 1730493024
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1730493024
transform -1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_73
timestamp 1730493024
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1730493024
transform -1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_74
timestamp 1730493024
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1730493024
transform -1 0 16836 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_75
timestamp 1730493024
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1730493024
transform -1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_76
timestamp 1730493024
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1730493024
transform -1 0 16836 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_77
timestamp 1730493024
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1730493024
transform -1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_78
timestamp 1730493024
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1730493024
transform -1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_79
timestamp 1730493024
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1730493024
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_80
timestamp 1730493024
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1730493024
transform -1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_81
timestamp 1730493024
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1730493024
transform -1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_82
timestamp 1730493024
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1730493024
transform -1 0 16836 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_83
timestamp 1730493024
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1730493024
transform -1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_84
timestamp 1730493024
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1730493024
transform -1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_85
timestamp 1730493024
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1730493024
transform -1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_86
timestamp 1730493024
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1730493024
transform -1 0 16836 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_87
timestamp 1730493024
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1730493024
transform -1 0 16836 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_88
timestamp 1730493024
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1730493024
transform -1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_89
timestamp 1730493024
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1730493024
transform -1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_90
timestamp 1730493024
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1730493024
transform -1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_91
timestamp 1730493024
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1730493024
transform -1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_92
timestamp 1730493024
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1730493024
transform -1 0 16836 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_93
timestamp 1730493024
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1730493024
transform -1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_94
timestamp 1730493024
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1730493024
transform -1 0 16836 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_95
timestamp 1730493024
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1730493024
transform -1 0 16836 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_96
timestamp 1730493024
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1730493024
transform -1 0 16836 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_97
timestamp 1730493024
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1730493024
transform -1 0 16836 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_98
timestamp 1730493024
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1730493024
transform -1 0 16836 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_99
timestamp 1730493024
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1730493024
transform -1 0 16836 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_100
timestamp 1730493024
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 1730493024
transform -1 0 16836 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Left_101
timestamp 1730493024
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_32_Right_32
timestamp 1730493024
transform -1 0 16836 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Left_102
timestamp 1730493024
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_33_Right_33
timestamp 1730493024
transform -1 0 16836 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Left_103
timestamp 1730493024
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_34_Right_34
timestamp 1730493024
transform -1 0 16836 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Left_104
timestamp 1730493024
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_35_Right_35
timestamp 1730493024
transform -1 0 16836 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Left_105
timestamp 1730493024
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_36_Right_36
timestamp 1730493024
transform -1 0 16836 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Left_106
timestamp 1730493024
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_37_Right_37
timestamp 1730493024
transform -1 0 16836 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Left_107
timestamp 1730493024
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_38_Right_38
timestamp 1730493024
transform -1 0 16836 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Left_108
timestamp 1730493024
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_39_Right_39
timestamp 1730493024
transform -1 0 16836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Left_109
timestamp 1730493024
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_40_Right_40
timestamp 1730493024
transform -1 0 16836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Left_110
timestamp 1730493024
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_41_Right_41
timestamp 1730493024
transform -1 0 16836 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Left_111
timestamp 1730493024
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_42_Right_42
timestamp 1730493024
transform -1 0 16836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Left_112
timestamp 1730493024
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_43_Right_43
timestamp 1730493024
transform -1 0 16836 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Left_113
timestamp 1730493024
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_44_Right_44
timestamp 1730493024
transform -1 0 16836 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Left_114
timestamp 1730493024
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_45_Right_45
timestamp 1730493024
transform -1 0 16836 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Left_115
timestamp 1730493024
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_46_Right_46
timestamp 1730493024
transform -1 0 16836 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Left_116
timestamp 1730493024
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_47_Right_47
timestamp 1730493024
transform -1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Left_117
timestamp 1730493024
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_48_Right_48
timestamp 1730493024
transform -1 0 16836 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Left_118
timestamp 1730493024
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_49_Right_49
timestamp 1730493024
transform -1 0 16836 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Left_119
timestamp 1730493024
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_50_Right_50
timestamp 1730493024
transform -1 0 16836 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Left_120
timestamp 1730493024
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_51_Right_51
timestamp 1730493024
transform -1 0 16836 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Left_121
timestamp 1730493024
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_52_Right_52
timestamp 1730493024
transform -1 0 16836 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Left_122
timestamp 1730493024
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_53_Right_53
timestamp 1730493024
transform -1 0 16836 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Left_123
timestamp 1730493024
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_54_Right_54
timestamp 1730493024
transform -1 0 16836 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Left_124
timestamp 1730493024
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_55_Right_55
timestamp 1730493024
transform -1 0 16836 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Left_125
timestamp 1730493024
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_56_Right_56
timestamp 1730493024
transform -1 0 16836 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Left_126
timestamp 1730493024
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_57_Right_57
timestamp 1730493024
transform -1 0 16836 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Left_127
timestamp 1730493024
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_58_Right_58
timestamp 1730493024
transform -1 0 16836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Left_128
timestamp 1730493024
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_59_Right_59
timestamp 1730493024
transform -1 0 16836 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Left_129
timestamp 1730493024
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_60_Right_60
timestamp 1730493024
transform -1 0 16836 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Left_130
timestamp 1730493024
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_61_Right_61
timestamp 1730493024
transform -1 0 16836 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Left_131
timestamp 1730493024
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_62_Right_62
timestamp 1730493024
transform -1 0 16836 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Left_132
timestamp 1730493024
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_63_Right_63
timestamp 1730493024
transform -1 0 16836 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Left_133
timestamp 1730493024
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_64_Right_64
timestamp 1730493024
transform -1 0 16836 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Left_134
timestamp 1730493024
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_65_Right_65
timestamp 1730493024
transform -1 0 16836 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Left_135
timestamp 1730493024
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_66_Right_66
timestamp 1730493024
transform -1 0 16836 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Left_136
timestamp 1730493024
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_67_Right_67
timestamp 1730493024
transform -1 0 16836 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Left_137
timestamp 1730493024
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_68_Right_68
timestamp 1730493024
transform -1 0 16836 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_138 ~/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730493024
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_139
timestamp 1730493024
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_140
timestamp 1730493024
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_141
timestamp 1730493024
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_142
timestamp 1730493024
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_143
timestamp 1730493024
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_144
timestamp 1730493024
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_145
timestamp 1730493024
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_146
timestamp 1730493024
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_147
timestamp 1730493024
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_148
timestamp 1730493024
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_149
timestamp 1730493024
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_150
timestamp 1730493024
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_151
timestamp 1730493024
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_152
timestamp 1730493024
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_153
timestamp 1730493024
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_154
timestamp 1730493024
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_155
timestamp 1730493024
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_156
timestamp 1730493024
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_157
timestamp 1730493024
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_158
timestamp 1730493024
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_159
timestamp 1730493024
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_160
timestamp 1730493024
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_161
timestamp 1730493024
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_162
timestamp 1730493024
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_163
timestamp 1730493024
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_164
timestamp 1730493024
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_165
timestamp 1730493024
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_166
timestamp 1730493024
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_167
timestamp 1730493024
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_168
timestamp 1730493024
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_169
timestamp 1730493024
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_170
timestamp 1730493024
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_171
timestamp 1730493024
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_172
timestamp 1730493024
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_173
timestamp 1730493024
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_174
timestamp 1730493024
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_175
timestamp 1730493024
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_176
timestamp 1730493024
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_177
timestamp 1730493024
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_178
timestamp 1730493024
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_179
timestamp 1730493024
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_180
timestamp 1730493024
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_181
timestamp 1730493024
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_182
timestamp 1730493024
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_183
timestamp 1730493024
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_184
timestamp 1730493024
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_185
timestamp 1730493024
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_186
timestamp 1730493024
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_187
timestamp 1730493024
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 1730493024
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 1730493024
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_190
timestamp 1730493024
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_191
timestamp 1730493024
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_192
timestamp 1730493024
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_193
timestamp 1730493024
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_194
timestamp 1730493024
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_195
timestamp 1730493024
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_196
timestamp 1730493024
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_197
timestamp 1730493024
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_198
timestamp 1730493024
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_199
timestamp 1730493024
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_200
timestamp 1730493024
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_201
timestamp 1730493024
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_202
timestamp 1730493024
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_203
timestamp 1730493024
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_204
timestamp 1730493024
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_205
timestamp 1730493024
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_206
timestamp 1730493024
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_207
timestamp 1730493024
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_208
timestamp 1730493024
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_209
timestamp 1730493024
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_210
timestamp 1730493024
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_211
timestamp 1730493024
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_212
timestamp 1730493024
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_213
timestamp 1730493024
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_214
timestamp 1730493024
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_215
timestamp 1730493024
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_216
timestamp 1730493024
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_217
timestamp 1730493024
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_218
timestamp 1730493024
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_219
timestamp 1730493024
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_220
timestamp 1730493024
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_221
timestamp 1730493024
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_32_222
timestamp 1730493024
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_223
timestamp 1730493024
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_33_224
timestamp 1730493024
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_225
timestamp 1730493024
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_226
timestamp 1730493024
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_34_227
timestamp 1730493024
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_228
timestamp 1730493024
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_35_229
timestamp 1730493024
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_230
timestamp 1730493024
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_231
timestamp 1730493024
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_36_232
timestamp 1730493024
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_233
timestamp 1730493024
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_37_234
timestamp 1730493024
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_235
timestamp 1730493024
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_236
timestamp 1730493024
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_38_237
timestamp 1730493024
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_238
timestamp 1730493024
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_39_239
timestamp 1730493024
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_240
timestamp 1730493024
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_241
timestamp 1730493024
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_40_242
timestamp 1730493024
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_243
timestamp 1730493024
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_41_244
timestamp 1730493024
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_245
timestamp 1730493024
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_246
timestamp 1730493024
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_42_247
timestamp 1730493024
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_248
timestamp 1730493024
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_43_249
timestamp 1730493024
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_250
timestamp 1730493024
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_251
timestamp 1730493024
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_44_252
timestamp 1730493024
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_253
timestamp 1730493024
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_45_254
timestamp 1730493024
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_255
timestamp 1730493024
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_256
timestamp 1730493024
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_46_257
timestamp 1730493024
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_258
timestamp 1730493024
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_47_259
timestamp 1730493024
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_260
timestamp 1730493024
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_261
timestamp 1730493024
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_48_262
timestamp 1730493024
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_263
timestamp 1730493024
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_49_264
timestamp 1730493024
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_265
timestamp 1730493024
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_266
timestamp 1730493024
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_50_267
timestamp 1730493024
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_268
timestamp 1730493024
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_51_269
timestamp 1730493024
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_270
timestamp 1730493024
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_271
timestamp 1730493024
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_52_272
timestamp 1730493024
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_273
timestamp 1730493024
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_53_274
timestamp 1730493024
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_275
timestamp 1730493024
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_276
timestamp 1730493024
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_54_277
timestamp 1730493024
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_278
timestamp 1730493024
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_55_279
timestamp 1730493024
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_280
timestamp 1730493024
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_281
timestamp 1730493024
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_56_282
timestamp 1730493024
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_283
timestamp 1730493024
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_57_284
timestamp 1730493024
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_285
timestamp 1730493024
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_286
timestamp 1730493024
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_58_287
timestamp 1730493024
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_288
timestamp 1730493024
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_59_289
timestamp 1730493024
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_290
timestamp 1730493024
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_291
timestamp 1730493024
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_60_292
timestamp 1730493024
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_293
timestamp 1730493024
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_61_294
timestamp 1730493024
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_295
timestamp 1730493024
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_296
timestamp 1730493024
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_62_297
timestamp 1730493024
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_298
timestamp 1730493024
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_63_299
timestamp 1730493024
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_300
timestamp 1730493024
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_301
timestamp 1730493024
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_64_302
timestamp 1730493024
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_303
timestamp 1730493024
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_65_304
timestamp 1730493024
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_305
timestamp 1730493024
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_306
timestamp 1730493024
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_66_307
timestamp 1730493024
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_308
timestamp 1730493024
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_67_309
timestamp 1730493024
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_310
timestamp 1730493024
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_311
timestamp 1730493024
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_312
timestamp 1730493024
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_313
timestamp 1730493024
transform 1 0 11408 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_68_314
timestamp 1730493024
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire62
timestamp 1730493024
transform 1 0 6900 0 -1 28288
box -38 -48 314 592
<< labels >>
flabel metal4 s 4868 2128 5188 39760 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 39760 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 10966 41200 11022 42000 0 FreeSans 224 90 0 0 b0
port 2 nsew signal input
flabel metal2 s 12898 41200 12954 42000 0 FreeSans 224 90 0 0 b1
port 3 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 clk
port 4 nsew signal input
flabel metal3 s 17200 13608 18000 13728 0 FreeSans 480 0 0 0 compr
port 5 nsew signal input
flabel metal3 s 17200 22448 18000 22568 0 FreeSans 480 0 0 0 dac[0]
port 6 nsew signal output
flabel metal3 s 17200 15648 18000 15768 0 FreeSans 480 0 0 0 dac[1]
port 7 nsew signal output
flabel metal3 s 17200 14288 18000 14408 0 FreeSans 480 0 0 0 dac[2]
port 8 nsew signal output
flabel metal3 s 17200 11568 18000 11688 0 FreeSans 480 0 0 0 dac[3]
port 9 nsew signal output
flabel metal3 s 17200 12248 18000 12368 0 FreeSans 480 0 0 0 dac[4]
port 10 nsew signal output
flabel metal3 s 17200 12928 18000 13048 0 FreeSans 480 0 0 0 dac[5]
port 11 nsew signal output
flabel metal3 s 17200 17008 18000 17128 0 FreeSans 480 0 0 0 dac[6]
port 12 nsew signal output
flabel metal3 s 17200 21768 18000 21888 0 FreeSans 480 0 0 0 dac[7]
port 13 nsew signal output
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 dac_coupl
port 14 nsew signal output
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 m0
port 15 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 m1
port 16 nsew signal input
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 reg0[0]
port 17 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 reg0[1]
port 18 nsew signal output
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 reg0[2]
port 19 nsew signal output
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 reg0[3]
port 20 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 reg0[4]
port 21 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 reg0[5]
port 22 nsew signal output
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 reg0[6]
port 23 nsew signal output
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 reg0[7]
port 24 nsew signal output
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 reg1[0]
port 25 nsew signal output
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 reg1[1]
port 26 nsew signal output
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 reg1[2]
port 27 nsew signal output
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 reg1[3]
port 28 nsew signal output
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 reg1[4]
port 29 nsew signal output
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 reg1[5]
port 30 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 reg1[6]
port 31 nsew signal output
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 reg1[7]
port 32 nsew signal output
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 reg2[0]
port 33 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 reg2[1]
port 34 nsew signal output
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 reg2[2]
port 35 nsew signal output
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 reg2[3]
port 36 nsew signal output
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 reg2[4]
port 37 nsew signal output
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 reg2[5]
port 38 nsew signal output
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 reg2[6]
port 39 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 reg2[7]
port 40 nsew signal output
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 reg3[0]
port 41 nsew signal output
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 reg3[1]
port 42 nsew signal output
flabel metal2 s 14186 0 14242 800 0 FreeSans 224 90 0 0 reg3[2]
port 43 nsew signal output
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 reg3[3]
port 44 nsew signal output
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 reg3[4]
port 45 nsew signal output
flabel metal3 s 17200 5448 18000 5568 0 FreeSans 480 0 0 0 reg3[5]
port 46 nsew signal output
flabel metal3 s 17200 10208 18000 10328 0 FreeSans 480 0 0 0 reg3[6]
port 47 nsew signal output
flabel metal3 s 17200 8168 18000 8288 0 FreeSans 480 0 0 0 reg3[7]
port 48 nsew signal output
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 reg4[0]
port 49 nsew signal output
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 reg4[1]
port 50 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 reg4[2]
port 51 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 reg4[3]
port 52 nsew signal output
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 reg4[4]
port 53 nsew signal output
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 reg4[5]
port 54 nsew signal output
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 reg4[6]
port 55 nsew signal output
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 reg4[7]
port 56 nsew signal output
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 rst
port 57 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 rx
port 58 nsew signal input
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 tx
port 59 nsew signal output
rlabel metal1 8970 39168 8970 39168 0 VGND
rlabel metal1 8970 39712 8970 39712 0 VPWR
rlabel metal2 4094 16354 4094 16354 0 _0000_
rlabel metal1 15088 16762 15088 16762 0 _0001_
rlabel metal1 12829 28118 12829 28118 0 _0002_
rlabel metal1 13340 31654 13340 31654 0 _0003_
rlabel metal1 14060 30634 14060 30634 0 _0004_
rlabel metal1 13554 29206 13554 29206 0 _0005_
rlabel metal1 13712 27030 13712 27030 0 _0006_
rlabel metal1 12098 25466 12098 25466 0 _0007_
rlabel metal1 10483 25942 10483 25942 0 _0008_
rlabel via1 9517 25194 9517 25194 0 _0009_
rlabel metal1 9614 27608 9614 27608 0 _0010_
rlabel metal1 7544 27098 7544 27098 0 _0011_
rlabel metal2 7222 28934 7222 28934 0 _0012_
rlabel metal1 6670 30906 6670 30906 0 _0013_
rlabel metal2 8234 31110 8234 31110 0 _0014_
rlabel metal2 1518 20706 1518 20706 0 _0015_
rlabel metal1 7038 17068 7038 17068 0 _0016_
rlabel metal1 1886 10778 1886 10778 0 _0017_
rlabel metal1 5060 11322 5060 11322 0 _0018_
rlabel metal1 5004 8466 5004 8466 0 _0019_
rlabel metal1 2525 8534 2525 8534 0 _0020_
rlabel via1 3629 11730 3629 11730 0 _0021_
rlabel metal1 2295 9962 2295 9962 0 _0022_
rlabel metal1 4630 10710 4630 10710 0 _0023_
rlabel metal1 4722 8874 4722 8874 0 _0024_
rlabel via1 15405 2414 15405 2414 0 _0025_
rlabel via1 14945 3026 14945 3026 0 _0026_
rlabel metal2 13018 5474 13018 5474 0 _0027_
rlabel metal2 14122 4998 14122 4998 0 _0028_
rlabel via1 11909 3434 11909 3434 0 _0029_
rlabel via1 15405 6358 15405 6358 0 _0030_
rlabel metal2 13202 8262 13202 8262 0 _0031_
rlabel metal1 14577 7786 14577 7786 0 _0032_
rlabel metal1 12921 3026 12921 3026 0 _0033_
rlabel metal1 7318 3094 7318 3094 0 _0034_
rlabel metal2 7222 4998 7222 4998 0 _0035_
rlabel metal2 15134 4284 15134 4284 0 _0036_
rlabel metal1 8224 3026 8224 3026 0 _0037_
rlabel metal1 15118 6698 15118 6698 0 _0038_
rlabel metal2 8970 4964 8970 4964 0 _0039_
rlabel metal1 7329 6698 7329 6698 0 _0040_
rlabel via1 2617 3026 2617 3026 0 _0041_
rlabel via1 4549 3094 4549 3094 0 _0042_
rlabel metal1 4503 4590 4503 4590 0 _0043_
rlabel metal2 2806 5406 2806 5406 0 _0044_
rlabel metal1 5458 3434 5458 3434 0 _0045_
rlabel metal2 2714 6562 2714 6562 0 _0046_
rlabel viali 5837 4590 5837 4590 0 _0047_
rlabel metal1 4820 6290 4820 6290 0 _0048_
rlabel metal1 1594 2346 1594 2346 0 _0049_
rlabel metal1 10340 3502 10340 3502 0 _0050_
rlabel metal1 10350 5066 10350 5066 0 _0051_
rlabel metal1 1594 4522 1594 4522 0 _0052_
rlabel metal1 9696 3026 9696 3026 0 _0053_
rlabel metal1 1656 7514 1656 7514 0 _0054_
rlabel metal2 9890 6086 9890 6086 0 _0055_
rlabel metal2 11546 7650 11546 7650 0 _0056_
rlabel metal1 5745 17238 5745 17238 0 _0057_
rlabel metal2 9522 12002 9522 12002 0 _0058_
rlabel metal2 10166 9826 10166 9826 0 _0059_
rlabel metal1 5699 12138 5699 12138 0 _0060_
rlabel metal1 7309 11798 7309 11798 0 _0061_
rlabel metal1 6348 10778 6348 10778 0 _0062_
rlabel via1 8965 9622 8965 9622 0 _0063_
rlabel metal1 7544 9146 7544 9146 0 _0064_
rlabel metal2 8050 7650 8050 7650 0 _0065_
rlabel metal2 9522 7378 9522 7378 0 _0066_
rlabel metal1 6440 8058 6440 8058 0 _0067_
rlabel metal2 4278 13090 4278 13090 0 _0068_
rlabel metal2 4094 14178 4094 14178 0 _0069_
rlabel metal2 6394 26010 6394 26010 0 _0070_
rlabel metal1 8132 24786 8132 24786 0 _0071_
rlabel metal2 5474 24582 5474 24582 0 _0072_
rlabel metal2 6486 24548 6486 24548 0 _0073_
rlabel metal2 5658 25364 5658 25364 0 _0074_
rlabel metal1 8096 18938 8096 18938 0 _0075_
rlabel metal1 9016 14586 9016 14586 0 _0076_
rlabel metal1 6808 15674 6808 15674 0 _0077_
rlabel metal1 7447 13226 7447 13226 0 _0078_
rlabel metal1 6808 14586 6808 14586 0 _0079_
rlabel metal1 9011 13906 9011 13906 0 _0080_
rlabel metal1 8873 16150 8873 16150 0 _0081_
rlabel metal1 5520 18394 5520 18394 0 _0082_
rlabel metal2 3082 34850 3082 34850 0 _0083_
rlabel metal1 3086 36142 3086 36142 0 _0084_
rlabel metal1 4048 36346 4048 36346 0 _0085_
rlabel metal1 4538 34986 4538 34986 0 _0086_
rlabel via1 4917 33490 4917 33490 0 _0087_
rlabel metal2 2990 33286 2990 33286 0 _0088_
rlabel metal2 4370 31518 4370 31518 0 _0089_
rlabel metal1 4084 30226 4084 30226 0 _0090_
rlabel metal2 2530 29410 2530 29410 0 _0091_
rlabel metal2 2714 27234 2714 27234 0 _0092_
rlabel metal1 4630 27030 4630 27030 0 _0093_
rlabel metal2 6302 27642 6302 27642 0 _0094_
rlabel metal2 3266 22848 3266 22848 0 _0095_
rlabel metal1 5024 25262 5024 25262 0 _0096_
rlabel metal1 3496 22474 3496 22474 0 _0097_
rlabel metal2 3174 23494 3174 23494 0 _0098_
rlabel metal2 7682 21794 7682 21794 0 _0099_
rlabel metal2 7774 20230 7774 20230 0 _0100_
rlabel metal1 5515 20434 5515 20434 0 _0101_
rlabel metal1 5331 21590 5331 21590 0 _0102_
rlabel metal1 6251 21930 6251 21930 0 _0103_
rlabel metal1 12726 35734 12726 35734 0 _0104_
rlabel metal1 13928 33966 13928 33966 0 _0105_
rlabel metal2 12834 33286 12834 33286 0 _0106_
rlabel metal1 12696 35462 12696 35462 0 _0107_
rlabel metal2 13110 38114 13110 38114 0 _0108_
rlabel metal2 12742 38726 12742 38726 0 _0109_
rlabel viali 10161 38998 10161 38998 0 _0110_
rlabel metal1 9000 38250 9000 38250 0 _0111_
rlabel metal1 7758 38998 7758 38998 0 _0112_
rlabel metal2 6670 38114 6670 38114 0 _0113_
rlabel metal1 6711 36822 6711 36822 0 _0114_
rlabel via1 6941 32878 6941 32878 0 _0115_
rlabel metal1 8740 33082 8740 33082 0 _0116_
rlabel metal1 15175 12886 15175 12886 0 _0117_
rlabel metal1 1594 13226 1594 13226 0 _0118_
rlabel metal1 11101 18326 11101 18326 0 _0119_
rlabel metal1 11331 15062 11331 15062 0 _0120_
rlabel metal1 11331 11798 11331 11798 0 _0121_
rlabel metal1 11561 14314 11561 14314 0 _0122_
rlabel metal1 12976 9962 12976 9962 0 _0123_
rlabel via1 11734 10030 11734 10030 0 _0124_
rlabel metal1 11285 12886 11285 12886 0 _0125_
rlabel metal1 14766 21114 14766 21114 0 _0126_
rlabel metal2 15134 15266 15134 15266 0 _0127_
rlabel metal2 15042 14178 15042 14178 0 _0128_
rlabel metal1 14904 10234 14904 10234 0 _0129_
rlabel metal2 14950 19618 14950 19618 0 _0130_
rlabel metal1 10897 19414 10897 19414 0 _0131_
rlabel metal1 10851 17170 10851 17170 0 _0132_
rlabel metal1 10529 16558 10529 16558 0 _0133_
rlabel metal1 2709 19414 2709 19414 0 _0134_
rlabel metal2 2898 16966 2898 16966 0 _0135_
rlabel metal1 1840 14586 1840 14586 0 _0136_
rlabel metal1 10457 19754 10457 19754 0 _0137_
rlabel metal1 11684 24242 11684 24242 0 _0138_
rlabel via1 1697 17578 1697 17578 0 _0139_
rlabel metal1 4360 14994 4360 14994 0 _0140_
rlabel metal1 11081 21930 11081 21930 0 _0141_
rlabel metal2 13386 21624 13386 21624 0 _0142_
rlabel metal1 3956 17850 3956 17850 0 _0143_
rlabel via1 2249 12818 2249 12818 0 _0144_
rlabel metal1 13248 23290 13248 23290 0 _0145_
rlabel via1 15129 11118 15129 11118 0 _0146_
rlabel metal2 7774 24276 7774 24276 0 _0147_
rlabel metal1 12098 12818 12098 12818 0 _0148_
rlabel metal2 4646 7582 4646 7582 0 _0149_
rlabel metal1 9384 7514 9384 7514 0 _0150_
rlabel metal1 12374 21114 12374 21114 0 _0151_
rlabel metal1 12926 20944 12926 20944 0 _0152_
rlabel metal1 13984 14994 13984 14994 0 _0153_
rlabel metal1 8556 35054 8556 35054 0 _0154_
rlabel metal1 5290 28050 5290 28050 0 _0155_
rlabel metal1 14076 9622 14076 9622 0 _0156_
rlabel metal2 12834 34272 12834 34272 0 _0157_
rlabel via1 3174 20366 3174 20366 0 _0158_
rlabel metal1 2208 18938 2208 18938 0 _0159_
rlabel metal2 2622 14824 2622 14824 0 _0160_
rlabel metal1 2622 15504 2622 15504 0 _0161_
rlabel metal1 3588 17850 3588 17850 0 _0162_
rlabel metal1 3312 20570 3312 20570 0 _0163_
rlabel metal1 4094 21522 4094 21522 0 _0164_
rlabel metal1 6486 32810 6486 32810 0 _0165_
rlabel metal1 7878 35734 7878 35734 0 _0166_
rlabel metal2 8050 35428 8050 35428 0 _0167_
rlabel metal1 8050 35666 8050 35666 0 _0168_
rlabel metal1 5474 35632 5474 35632 0 _0169_
rlabel metal1 6716 29750 6716 29750 0 _0170_
rlabel metal1 7728 35802 7728 35802 0 _0171_
rlabel metal1 8970 36074 8970 36074 0 _0172_
rlabel metal1 10120 33490 10120 33490 0 _0173_
rlabel metal1 11546 32538 11546 32538 0 _0174_
rlabel metal2 7682 32946 7682 32946 0 _0175_
rlabel metal1 11914 32946 11914 32946 0 _0176_
rlabel metal1 10350 36244 10350 36244 0 _0177_
rlabel metal1 10534 37162 10534 37162 0 _0178_
rlabel metal1 10580 36142 10580 36142 0 _0179_
rlabel metal1 10718 35734 10718 35734 0 _0180_
rlabel metal1 11454 35802 11454 35802 0 _0181_
rlabel viali 10810 36143 10810 36143 0 _0182_
rlabel metal1 11592 33626 11592 33626 0 _0183_
rlabel metal1 10580 35258 10580 35258 0 _0184_
rlabel metal1 10764 33898 10764 33898 0 _0185_
rlabel metal1 10810 34000 10810 34000 0 _0186_
rlabel metal2 10442 34578 10442 34578 0 _0187_
rlabel metal1 10166 35632 10166 35632 0 _0188_
rlabel metal2 10534 36108 10534 36108 0 _0189_
rlabel metal1 11454 35530 11454 35530 0 _0190_
rlabel metal1 10718 36278 10718 36278 0 _0191_
rlabel metal2 10626 35836 10626 35836 0 _0192_
rlabel metal2 9982 35972 9982 35972 0 _0193_
rlabel metal1 8924 35054 8924 35054 0 _0194_
rlabel metal2 8970 35428 8970 35428 0 _0195_
rlabel metal1 9062 35802 9062 35802 0 _0196_
rlabel metal1 13064 33898 13064 33898 0 _0197_
rlabel metal1 10304 33286 10304 33286 0 _0198_
rlabel metal1 10434 34918 10434 34918 0 _0199_
rlabel metal2 9982 35462 9982 35462 0 _0200_
rlabel metal2 9890 34714 9890 34714 0 _0201_
rlabel metal2 2254 17374 2254 17374 0 _0202_
rlabel metal1 3726 16762 3726 16762 0 _0203_
rlabel metal2 4646 16490 4646 16490 0 _0204_
rlabel metal2 12466 20825 12466 20825 0 _0205_
rlabel metal1 13938 20502 13938 20502 0 _0206_
rlabel metal1 12190 22746 12190 22746 0 _0207_
rlabel metal2 14352 19346 14352 19346 0 _0208_
rlabel metal1 14352 19210 14352 19210 0 _0209_
rlabel metal1 13110 17204 13110 17204 0 _0210_
rlabel metal2 12558 16320 12558 16320 0 _0211_
rlabel metal2 12926 15198 12926 15198 0 _0212_
rlabel metal1 13432 14586 13432 14586 0 _0213_
rlabel metal1 13340 17306 13340 17306 0 _0214_
rlabel metal1 14076 12410 14076 12410 0 _0215_
rlabel metal1 14214 16626 14214 16626 0 _0216_
rlabel metal1 8602 21080 8602 21080 0 _0217_
rlabel metal1 2277 21386 2277 21386 0 _0218_
rlabel metal1 14582 20366 14582 20366 0 _0219_
rlabel metal1 12742 20808 12742 20808 0 _0220_
rlabel metal1 13662 12852 13662 12852 0 _0221_
rlabel metal2 13662 16150 13662 16150 0 _0222_
rlabel metal1 13708 21046 13708 21046 0 _0223_
rlabel metal2 11822 18377 11822 18377 0 _0224_
rlabel metal2 13478 21318 13478 21318 0 _0225_
rlabel metal1 15272 16626 15272 16626 0 _0226_
rlabel metal2 14490 17986 14490 17986 0 _0227_
rlabel metal1 15502 16490 15502 16490 0 _0228_
rlabel metal2 8510 29920 8510 29920 0 _0229_
rlabel metal1 8510 29716 8510 29716 0 _0230_
rlabel metal1 8326 29512 8326 29512 0 _0231_
rlabel metal1 10534 29580 10534 29580 0 _0232_
rlabel metal1 10718 31824 10718 31824 0 _0233_
rlabel viali 10544 31790 10544 31790 0 _0234_
rlabel metal2 11040 30702 11040 30702 0 _0235_
rlabel metal2 10626 28356 10626 28356 0 _0236_
rlabel metal2 11546 28356 11546 28356 0 _0237_
rlabel metal1 10396 28730 10396 28730 0 _0238_
rlabel metal2 10994 29546 10994 29546 0 _0239_
rlabel metal1 11224 30702 11224 30702 0 _0240_
rlabel metal1 11362 30770 11362 30770 0 _0241_
rlabel metal1 10442 30362 10442 30362 0 _0242_
rlabel metal2 10626 29376 10626 29376 0 _0243_
rlabel metal1 11178 29172 11178 29172 0 _0244_
rlabel metal2 12006 29376 12006 29376 0 _0245_
rlabel metal1 11316 29818 11316 29818 0 _0246_
rlabel metal1 11454 29138 11454 29138 0 _0247_
rlabel metal2 10810 30090 10810 30090 0 _0248_
rlabel metal2 10718 29444 10718 29444 0 _0249_
rlabel metal1 10258 29614 10258 29614 0 _0250_
rlabel metal2 9522 29818 9522 29818 0 _0251_
rlabel metal1 9200 31654 9200 31654 0 _0252_
rlabel metal1 9292 29682 9292 29682 0 _0253_
rlabel metal2 13202 29138 13202 29138 0 _0254_
rlabel metal2 10718 30906 10718 30906 0 _0255_
rlabel metal1 9982 30838 9982 30838 0 _0256_
rlabel metal1 13340 28458 13340 28458 0 _0257_
rlabel metal1 12846 31858 12846 31858 0 _0258_
rlabel metal1 13110 30362 13110 30362 0 _0259_
rlabel metal1 14076 30090 14076 30090 0 _0260_
rlabel metal1 13260 30634 13260 30634 0 _0261_
rlabel metal1 12581 26418 12581 26418 0 _0262_
rlabel metal1 13386 29648 13386 29648 0 _0263_
rlabel metal1 13076 29070 13076 29070 0 _0264_
rlabel metal1 13156 26554 13156 26554 0 _0265_
rlabel metal2 11638 26758 11638 26758 0 _0266_
rlabel metal2 12098 26758 12098 26758 0 _0267_
rlabel metal1 12110 25330 12110 25330 0 _0268_
rlabel metal1 10120 27438 10120 27438 0 _0269_
rlabel metal1 10994 26316 10994 26316 0 _0270_
rlabel metal1 10730 26282 10730 26282 0 _0271_
rlabel metal1 8786 25840 8786 25840 0 _0272_
rlabel metal1 8556 27574 8556 27574 0 _0273_
rlabel metal1 9430 26962 9430 26962 0 _0274_
rlabel metal2 9062 27234 9062 27234 0 _0275_
rlabel metal1 7728 31790 7728 31790 0 _0276_
rlabel metal1 7590 28016 7590 28016 0 _0277_
rlabel metal1 7669 26962 7669 26962 0 _0278_
rlabel metal1 6624 31450 6624 31450 0 _0279_
rlabel via1 7050 28594 7050 28594 0 _0280_
rlabel metal2 6578 31212 6578 31212 0 _0281_
rlabel via1 8062 30702 8062 30702 0 _0282_
rlabel metal2 2162 20876 2162 20876 0 _0283_
rlabel metal1 9614 12682 9614 12682 0 _0284_
rlabel metal1 8648 20026 8648 20026 0 _0285_
rlabel metal2 4784 16660 4784 16660 0 _0286_
rlabel metal1 12972 7378 12972 7378 0 _0287_
rlabel metal1 1702 11832 1702 11832 0 _0288_
rlabel metal1 2254 8976 2254 8976 0 _0289_
rlabel metal2 2162 11084 2162 11084 0 _0290_
rlabel metal1 4554 11152 4554 11152 0 _0291_
rlabel metal1 4278 8500 4278 8500 0 _0292_
rlabel metal2 2070 8772 2070 8772 0 _0293_
rlabel metal1 4140 11322 4140 11322 0 _0294_
rlabel metal1 2392 10234 2392 10234 0 _0295_
rlabel metal1 4968 9486 4968 9486 0 _0296_
rlabel metal2 4094 9146 4094 9146 0 _0297_
rlabel metal1 10626 8942 10626 8942 0 _0298_
rlabel metal1 14352 2346 14352 2346 0 _0299_
rlabel via1 14491 3502 14491 3502 0 _0300_
rlabel metal1 15042 2618 15042 2618 0 _0301_
rlabel metal1 14444 2618 14444 2618 0 _0302_
rlabel metal2 12466 5372 12466 5372 0 _0303_
rlabel metal2 14582 5066 14582 5066 0 _0304_
rlabel metal1 12650 4080 12650 4080 0 _0305_
rlabel metal1 14306 6970 14306 6970 0 _0306_
rlabel metal1 12742 7888 12742 7888 0 _0307_
rlabel metal1 13984 8058 13984 8058 0 _0308_
rlabel metal2 11178 6562 11178 6562 0 _0309_
rlabel metal1 7820 2346 7820 2346 0 _0310_
rlabel metal1 9338 4624 9338 4624 0 _0311_
rlabel metal1 13938 3162 13938 3162 0 _0312_
rlabel metal1 7544 2618 7544 2618 0 _0313_
rlabel metal2 7682 5066 7682 5066 0 _0314_
rlabel metal1 14628 4114 14628 4114 0 _0315_
rlabel metal1 8694 2618 8694 2618 0 _0316_
rlabel metal1 14352 6426 14352 6426 0 _0317_
rlabel metal1 9430 4556 9430 4556 0 _0318_
rlabel metal1 7682 6426 7682 6426 0 _0319_
rlabel metal1 8418 5576 8418 5576 0 _0320_
rlabel metal1 3634 2346 3634 2346 0 _0321_
rlabel metal1 4738 6800 4738 6800 0 _0322_
rlabel metal1 3174 2618 3174 2618 0 _0323_
rlabel metal2 4186 3264 4186 3264 0 _0324_
rlabel metal1 4646 4250 4646 4250 0 _0325_
rlabel metal1 3496 5338 3496 5338 0 _0326_
rlabel metal1 5290 3162 5290 3162 0 _0327_
rlabel metal1 3174 6324 3174 6324 0 _0328_
rlabel metal1 5290 5236 5290 5236 0 _0329_
rlabel metal2 4554 6596 4554 6596 0 _0330_
rlabel metal1 9476 8534 9476 8534 0 _0331_
rlabel metal1 2024 5678 2024 5678 0 _0332_
rlabel metal2 1886 4352 1886 4352 0 _0333_
rlabel metal2 1978 3332 1978 3332 0 _0334_
rlabel metal1 10718 4080 10718 4080 0 _0335_
rlabel metal1 10718 5236 10718 5236 0 _0336_
rlabel metal2 1978 5372 1978 5372 0 _0337_
rlabel metal1 10442 3162 10442 3162 0 _0338_
rlabel metal1 2070 7412 2070 7412 0 _0339_
rlabel metal1 9430 5712 9430 5712 0 _0340_
rlabel metal1 12006 7344 12006 7344 0 _0341_
rlabel metal1 3496 3910 3496 3910 0 _0342_
rlabel metal1 13202 3978 13202 3978 0 _0343_
rlabel metal1 6348 17102 6348 17102 0 _0344_
rlabel metal1 7590 2550 7590 2550 0 _0345_
rlabel via3 7245 12580 7245 12580 0 _0346_
rlabel metal1 8418 12682 8418 12682 0 _0347_
rlabel metal2 7314 5678 7314 5678 0 _0348_
rlabel metal1 11546 5338 11546 5338 0 _0349_
rlabel metal1 8694 7242 8694 7242 0 _0350_
rlabel metal2 15042 4862 15042 4862 0 _0351_
rlabel metal2 3450 6324 3450 6324 0 _0352_
rlabel metal2 6210 12789 6210 12789 0 _0353_
rlabel metal1 10350 2822 10350 2822 0 _0354_
rlabel metal1 8372 3978 8372 3978 0 _0355_
rlabel metal1 7912 10778 7912 10778 0 _0356_
rlabel metal1 4094 7514 4094 7514 0 _0357_
rlabel metal1 14168 6154 14168 6154 0 _0358_
rlabel metal1 6118 10234 6118 10234 0 _0359_
rlabel metal2 10902 9520 10902 9520 0 _0360_
rlabel metal2 8786 7956 8786 7956 0 _0361_
rlabel metal1 8832 10234 8832 10234 0 _0362_
rlabel metal1 6992 6426 6992 6426 0 _0363_
rlabel metal2 7314 9316 7314 9316 0 _0364_
rlabel metal1 8004 9010 8004 9010 0 _0365_
rlabel metal2 3634 13498 3634 13498 0 _0366_
rlabel metal2 3450 14348 3450 14348 0 _0367_
rlabel metal2 7682 24956 7682 24956 0 _0368_
rlabel metal2 7590 25466 7590 25466 0 _0369_
rlabel metal1 9660 23834 9660 23834 0 _0370_
rlabel metal1 8648 24038 8648 24038 0 _0371_
rlabel metal1 7130 19788 7130 19788 0 _0372_
rlabel metal2 7498 23052 7498 23052 0 _0373_
rlabel metal1 6762 25194 6762 25194 0 _0374_
rlabel metal2 7590 20366 7590 20366 0 _0375_
rlabel metal1 8648 15674 8648 15674 0 _0376_
rlabel metal1 7958 16014 7958 16014 0 _0377_
rlabel metal2 8326 16286 8326 16286 0 _0378_
rlabel metal1 7958 16218 7958 16218 0 _0379_
rlabel metal1 6946 20570 6946 20570 0 _0380_
rlabel metal1 8188 17646 8188 17646 0 _0381_
rlabel metal2 8326 17578 8326 17578 0 _0382_
rlabel metal2 8970 17442 8970 17442 0 _0383_
rlabel metal1 8326 17170 8326 17170 0 _0384_
rlabel metal1 7314 17306 7314 17306 0 _0385_
rlabel via1 7406 21318 7406 21318 0 _0386_
rlabel metal1 6854 19482 6854 19482 0 _0387_
rlabel metal1 6808 20026 6808 20026 0 _0388_
rlabel metal1 6118 24208 6118 24208 0 _0389_
rlabel metal1 5842 20910 5842 20910 0 _0390_
rlabel metal1 8694 18666 8694 18666 0 _0391_
rlabel metal1 9200 12954 9200 12954 0 _0392_
rlabel metal1 6808 15334 6808 15334 0 _0393_
rlabel metal1 8510 11322 8510 11322 0 _0394_
rlabel metal1 7544 14246 7544 14246 0 _0395_
rlabel metal1 9844 11322 9844 11322 0 _0396_
rlabel metal1 9384 15674 9384 15674 0 _0397_
rlabel metal1 6164 18394 6164 18394 0 _0398_
rlabel metal1 5566 31824 5566 31824 0 _0399_
rlabel metal2 2070 36516 2070 36516 0 _0400_
rlabel metal1 4738 36074 4738 36074 0 _0401_
rlabel metal2 5658 35904 5658 35904 0 _0402_
rlabel metal2 5382 33660 5382 33660 0 _0403_
rlabel metal2 5014 31994 5014 31994 0 _0404_
rlabel metal1 4922 31450 4922 31450 0 _0405_
rlabel metal1 5612 31926 5612 31926 0 _0406_
rlabel metal1 6026 28730 6026 28730 0 _0407_
rlabel metal1 5106 29172 5106 29172 0 _0408_
rlabel metal1 4968 29138 4968 29138 0 _0409_
rlabel metal1 4692 28730 4692 28730 0 _0410_
rlabel metal1 6946 28050 6946 28050 0 _0411_
rlabel metal1 4416 26010 4416 26010 0 _0412_
rlabel metal1 3588 32742 3588 32742 0 _0413_
rlabel metal1 2944 35802 2944 35802 0 _0414_
rlabel metal1 4224 36074 4224 36074 0 _0415_
rlabel metal1 3956 35190 3956 35190 0 _0416_
rlabel metal1 4416 35258 4416 35258 0 _0417_
rlabel metal2 4554 33898 4554 33898 0 _0418_
rlabel metal1 4784 31994 4784 31994 0 _0419_
rlabel metal1 3818 33014 3818 33014 0 _0420_
rlabel metal1 3496 33082 3496 33082 0 _0421_
rlabel metal1 3772 31926 3772 31926 0 _0422_
rlabel metal1 3910 31994 3910 31994 0 _0423_
rlabel metal2 3174 30294 3174 30294 0 _0424_
rlabel metal1 3328 30294 3328 30294 0 _0425_
rlabel metal1 3174 29002 3174 29002 0 _0426_
rlabel metal1 3358 28968 3358 28968 0 _0427_
rlabel metal1 3588 28186 3588 28186 0 _0428_
rlabel metal1 3404 26758 3404 26758 0 _0429_
rlabel metal1 4278 26792 4278 26792 0 _0430_
rlabel metal1 4148 27098 4148 27098 0 _0431_
rlabel metal1 4830 22542 4830 22542 0 _0432_
rlabel metal1 7636 21454 7636 21454 0 _0433_
rlabel metal2 6394 20230 6394 20230 0 _0434_
rlabel metal1 5796 21114 5796 21114 0 _0435_
rlabel metal1 6670 20468 6670 20468 0 _0436_
rlabel metal1 7774 21454 7774 21454 0 _0437_
rlabel metal2 7038 21828 7038 21828 0 _0438_
rlabel metal1 13018 34612 13018 34612 0 _0439_
rlabel metal1 13432 33898 13432 33898 0 _0440_
rlabel metal2 12742 34748 12742 34748 0 _0441_
rlabel metal1 12512 34170 12512 34170 0 _0442_
rlabel metal1 12956 32810 12956 32810 0 _0443_
rlabel metal1 12972 35054 12972 35054 0 _0444_
rlabel metal1 12742 35088 12742 35088 0 _0445_
rlabel metal1 12834 35190 12834 35190 0 _0446_
rlabel metal1 12788 37434 12788 37434 0 _0447_
rlabel metal1 13248 37910 13248 37910 0 _0448_
rlabel metal1 11592 38318 11592 38318 0 _0449_
rlabel metal2 12190 38012 12190 38012 0 _0450_
rlabel metal1 11922 38182 11922 38182 0 _0451_
rlabel metal2 10626 38148 10626 38148 0 _0452_
rlabel metal1 10810 38352 10810 38352 0 _0453_
rlabel metal2 10810 38896 10810 38896 0 _0454_
rlabel metal1 8510 37774 8510 37774 0 _0455_
rlabel metal2 7682 38080 7682 38080 0 _0456_
rlabel via1 8145 37978 8145 37978 0 _0457_
rlabel metal1 7774 38454 7774 38454 0 _0458_
rlabel metal1 7452 37638 7452 37638 0 _0459_
rlabel metal2 7222 38454 7222 38454 0 _0460_
rlabel metal1 6984 37978 6984 37978 0 _0461_
rlabel metal2 7038 36720 7038 36720 0 _0462_
rlabel metal1 7912 34578 7912 34578 0 _0463_
rlabel metal2 7498 33320 7498 33320 0 _0464_
rlabel via1 7214 33898 7214 33898 0 _0465_
rlabel metal1 13432 12818 13432 12818 0 _0466_
rlabel metal1 14950 12954 14950 12954 0 _0467_
rlabel metal1 15180 12614 15180 12614 0 _0468_
rlabel metal1 1978 14416 1978 14416 0 _0469_
rlabel metal1 13386 21386 13386 21386 0 _0470_
rlabel metal1 14076 19346 14076 19346 0 _0471_
rlabel metal1 12098 18326 12098 18326 0 _0472_
rlabel metal2 12926 17986 12926 17986 0 _0473_
rlabel metal1 13340 15062 13340 15062 0 _0474_
rlabel metal1 12926 15334 12926 15334 0 _0475_
rlabel metal1 12006 14960 12006 14960 0 _0476_
rlabel metal1 12650 14450 12650 14450 0 _0477_
rlabel metal1 11960 16558 11960 16558 0 _0478_
rlabel metal1 13386 13328 13386 13328 0 _0479_
rlabel metal2 12558 14246 12558 14246 0 _0480_
rlabel metal2 11914 11934 11914 11934 0 _0481_
rlabel metal2 13386 15164 13386 15164 0 _0482_
rlabel metal1 12920 13940 12920 13940 0 _0483_
rlabel metal1 11960 14382 11960 14382 0 _0484_
rlabel metal1 13202 10438 13202 10438 0 _0485_
rlabel metal1 13524 11118 13524 11118 0 _0486_
rlabel metal2 12650 10778 12650 10778 0 _0487_
rlabel metal1 12144 10506 12144 10506 0 _0488_
rlabel metal3 12742 15844 12742 15844 0 _0489_
rlabel metal1 13846 19482 13846 19482 0 _0490_
rlabel metal2 13846 20604 13846 20604 0 _0491_
rlabel metal1 11822 19346 11822 19346 0 _0492_
rlabel metal1 14812 20570 14812 20570 0 _0493_
rlabel metal1 14260 18258 14260 18258 0 _0494_
rlabel metal1 14996 18394 14996 18394 0 _0495_
rlabel metal2 15686 15300 15686 15300 0 _0496_
rlabel metal1 14076 15130 14076 15130 0 _0497_
rlabel metal2 15594 15198 15594 15198 0 _0498_
rlabel metal1 13892 13498 13892 13498 0 _0499_
rlabel metal1 15594 13804 15594 13804 0 _0500_
rlabel metal2 13202 13702 13202 13702 0 _0501_
rlabel metal1 13754 14008 13754 14008 0 _0502_
rlabel metal1 13892 10642 13892 10642 0 _0503_
rlabel metal2 15502 10268 15502 10268 0 _0504_
rlabel metal1 14536 11866 14536 11866 0 _0505_
rlabel metal1 15134 13158 15134 13158 0 _0506_
rlabel metal1 13156 18734 13156 18734 0 _0507_
rlabel metal1 13432 19890 13432 19890 0 _0508_
rlabel metal1 13202 19788 13202 19788 0 _0509_
rlabel metal2 15502 19482 15502 19482 0 _0510_
rlabel metal1 14168 18394 14168 18394 0 _0511_
rlabel metal1 15226 18938 15226 18938 0 _0512_
rlabel metal2 12006 19856 12006 19856 0 _0513_
rlabel metal2 2346 19380 2346 19380 0 _0514_
rlabel metal1 3082 16592 3082 16592 0 _0515_
rlabel metal2 2162 14858 2162 14858 0 _0516_
rlabel metal1 12190 19890 12190 19890 0 _0517_
rlabel metal1 2024 17306 2024 17306 0 _0518_
rlabel metal1 4646 15572 4646 15572 0 _0519_
rlabel metal2 12650 21760 12650 21760 0 _0520_
rlabel metal2 11362 21828 11362 21828 0 _0521_
rlabel metal2 2898 14042 2898 14042 0 _0522_
rlabel metal2 11730 22882 11730 22882 0 _0523_
rlabel metal2 13938 11458 13938 11458 0 _0524_
rlabel metal1 13202 11220 13202 11220 0 _0525_
rlabel metal1 15134 11322 15134 11322 0 _0526_
rlabel metal1 11040 39406 11040 39406 0 b0
rlabel metal1 13064 39406 13064 39406 0 b1
rlabel metal1 1288 21930 1288 21930 0 clk
rlabel metal1 10442 13294 10442 13294 0 clknet_0_clk
rlabel metal1 1840 2414 1840 2414 0 clknet_4_0_0_clk
rlabel metal1 4600 32334 4600 32334 0 clknet_4_10_0_clk
rlabel metal1 6900 38862 6900 38862 0 clknet_4_11_0_clk
rlabel metal1 10120 22066 10120 22066 0 clknet_4_12_0_clk
rlabel metal1 14122 21998 14122 21998 0 clknet_4_13_0_clk
rlabel metal2 12650 34578 12650 34578 0 clknet_4_14_0_clk
rlabel metal2 13938 38624 13938 38624 0 clknet_4_15_0_clk
rlabel via1 5566 4573 5566 4573 0 clknet_4_1_0_clk
rlabel metal1 1610 15028 1610 15028 0 clknet_4_2_0_clk
rlabel metal1 7866 19380 7866 19380 0 clknet_4_3_0_clk
rlabel metal1 7958 3026 7958 3026 0 clknet_4_4_0_clk
rlabel metal2 14674 2720 14674 2720 0 clknet_4_5_0_clk
rlabel metal1 9338 14858 9338 14858 0 clknet_4_6_0_clk
rlabel metal1 14674 17170 14674 17170 0 clknet_4_7_0_clk
rlabel metal2 2254 28560 2254 28560 0 clknet_4_8_0_clk
rlabel metal1 7084 24174 7084 24174 0 clknet_4_9_0_clk
rlabel metal2 16514 13243 16514 13243 0 compr
rlabel metal2 9890 21726 9890 21726 0 control.baud_clk
rlabel metal2 13110 35360 13110 35360 0 control.baud_rate_gen.count\[0\]
rlabel metal2 7222 35904 7222 35904 0 control.baud_rate_gen.count\[10\]
rlabel metal2 7866 35292 7866 35292 0 control.baud_rate_gen.count\[11\]
rlabel metal1 9292 33286 9292 33286 0 control.baud_rate_gen.count\[12\]
rlabel metal1 13938 33864 13938 33864 0 control.baud_rate_gen.count\[1\]
rlabel metal1 12535 33354 12535 33354 0 control.baud_rate_gen.count\[2\]
rlabel metal2 12098 35972 12098 35972 0 control.baud_rate_gen.count\[3\]
rlabel metal1 13110 37230 13110 37230 0 control.baud_rate_gen.count\[4\]
rlabel metal2 11270 36992 11270 36992 0 control.baud_rate_gen.count\[5\]
rlabel metal2 11086 38522 11086 38522 0 control.baud_rate_gen.count\[6\]
rlabel metal2 10350 38080 10350 38080 0 control.baud_rate_gen.count\[7\]
rlabel metal2 6762 35326 6762 35326 0 control.baud_rate_gen.count\[8\]
rlabel metal2 7590 36448 7590 36448 0 control.baud_rate_gen.count\[9\]
rlabel metal2 9154 32241 9154 32241 0 control.baud_rate_gen.n805_o
rlabel metal1 12834 20876 12834 20876 0 control.n576_q\[0\]
rlabel metal1 13018 21420 13018 21420 0 control.n576_q\[1\]
rlabel metal1 11224 21454 11224 21454 0 control.n576_q\[2\]
rlabel metal2 11914 23494 11914 23494 0 control.n579_q
rlabel metal1 12466 16490 12466 16490 0 control.n588_o
rlabel metal1 15778 21420 15778 21420 0 control.n598_o
rlabel metal1 16008 16082 16008 16082 0 control.n600_o
rlabel metal2 16146 14790 16146 14790 0 control.n602_o
rlabel metal1 16146 10098 16146 10098 0 control.n604_o
rlabel metal1 16146 11322 16146 11322 0 control.n606_o
rlabel metal1 16330 12954 16330 12954 0 control.n608_o
rlabel metal1 16284 17306 16284 17306 0 control.n610_o
rlabel metal1 16100 20366 16100 20366 0 control.n612_o
rlabel metal1 10166 18394 10166 18394 0 control.n633_o
rlabel metal1 10626 15470 10626 15470 0 control.n635_o
rlabel metal1 10028 11866 10028 11866 0 control.n637_o
rlabel metal1 10626 14586 10626 14586 0 control.n639_o
rlabel metal1 14766 10166 14766 10166 0 control.n641_o
rlabel metal1 10350 10166 10350 10166 0 control.n643_o
rlabel metal2 9890 13090 9890 13090 0 control.n645_o
rlabel metal1 9338 20026 9338 20026 0 control.n647_o
rlabel metal2 13018 17408 13018 17408 0 control.n651_o
rlabel metal1 12098 17680 12098 17680 0 control.n653_o
rlabel via2 16422 22491 16422 22491 0 dac[0]
rlabel via2 16422 15691 16422 15691 0 dac[1]
rlabel metal2 16422 14297 16422 14297 0 dac[2]
rlabel via2 16422 11611 16422 11611 0 dac[3]
rlabel via2 16422 12325 16422 12325 0 dac[4]
rlabel metal2 15594 13073 15594 13073 0 dac[5]
rlabel via2 16422 17051 16422 17051 0 dac[6]
rlabel via2 16422 21845 16422 21845 0 dac[7]
rlabel metal1 1840 20298 1840 20298 0 dac_coupl
rlabel metal3 751 22508 751 22508 0 m0
rlabel metal3 751 21828 751 21828 0 m1
rlabel metal2 9062 8806 9062 8806 0 n119_q\[0\]
rlabel metal1 10764 7718 10764 7718 0 n119_q\[1\]
rlabel metal1 7084 8806 7084 8806 0 n119_q\[2\]
rlabel metal1 10948 23698 10948 23698 0 n120_q
rlabel metal1 6762 17714 6762 17714 0 n126_q\[0\]
rlabel metal1 10074 15334 10074 15334 0 n126_q\[1\]
rlabel metal2 10534 10608 10534 10608 0 n126_q\[2\]
rlabel metal2 7130 12886 7130 12886 0 n126_q\[3\]
rlabel metal1 8510 11866 8510 11866 0 n126_q\[4\]
rlabel metal1 7084 10982 7084 10982 0 n126_q\[5\]
rlabel metal1 9844 12818 9844 12818 0 n126_q\[6\]
rlabel metal1 8970 18870 8970 18870 0 n126_q\[7\]
rlabel metal1 10166 22746 10166 22746 0 n127_q
rlabel metal1 10902 35666 10902 35666 0 net1
rlabel metal2 16238 14586 16238 14586 0 net10
rlabel metal1 15548 20910 15548 20910 0 net100
rlabel metal1 12098 11798 12098 11798 0 net101
rlabel metal2 15318 19856 15318 19856 0 net102
rlabel metal2 11914 13056 11914 13056 0 net103
rlabel metal1 15548 9894 15548 9894 0 net104
rlabel metal2 6486 15980 6486 15980 0 net105
rlabel metal1 9568 10642 9568 10642 0 net106
rlabel metal1 8694 18734 8694 18734 0 net107
rlabel metal2 9982 16320 9982 16320 0 net108
rlabel metal2 6026 22780 6026 22780 0 net109
rlabel metal1 16284 9418 16284 9418 0 net11
rlabel metal1 9798 11798 9798 11798 0 net110
rlabel metal1 6302 12954 6302 12954 0 net111
rlabel metal1 3496 19822 3496 19822 0 net112
rlabel metal1 10948 19890 10948 19890 0 net113
rlabel metal1 8740 13158 8740 13158 0 net114
rlabel metal1 9108 14450 9108 14450 0 net115
rlabel metal1 10258 13906 10258 13906 0 net116
rlabel metal2 12098 18496 12098 18496 0 net117
rlabel metal2 12190 10948 12190 10948 0 net118
rlabel metal2 7406 14892 7406 14892 0 net119
rlabel metal2 16330 11764 16330 11764 0 net12
rlabel metal1 6808 24378 6808 24378 0 net120
rlabel metal1 7125 24106 7125 24106 0 net121
rlabel metal1 7314 22406 7314 22406 0 net122
rlabel metal1 6026 28526 6026 28526 0 net123
rlabel metal1 5581 27370 5581 27370 0 net124
rlabel metal1 12512 21658 12512 21658 0 net125
rlabel metal1 8464 8874 8464 8874 0 net126
rlabel metal2 12006 23732 12006 23732 0 net127
rlabel via1 10805 23086 10805 23086 0 net128
rlabel metal2 6762 8194 6762 8194 0 net129
rlabel metal1 15870 13294 15870 13294 0 net13
rlabel metal2 4830 23324 4830 23324 0 net130
rlabel metal1 3818 22610 3818 22610 0 net131
rlabel metal1 5980 18326 5980 18326 0 net132
rlabel metal1 4646 22678 4646 22678 0 net133
rlabel metal2 2898 21080 2898 21080 0 net134
rlabel metal1 6762 24786 6762 24786 0 net135
rlabel via1 6021 25262 6021 25262 0 net136
rlabel metal2 12650 15232 12650 15232 0 net137
rlabel metal1 6440 20570 6440 20570 0 net138
rlabel metal2 14122 9724 14122 9724 0 net139
rlabel metal1 16192 16762 16192 16762 0 net14
rlabel metal1 7452 21522 7452 21522 0 net140
rlabel metal1 10120 6698 10120 6698 0 net141
rlabel metal2 16146 21556 16146 21556 0 net15
rlabel metal2 2714 20774 2714 20774 0 net16
rlabel metal1 2070 3128 2070 3128 0 net17
rlabel metal1 11776 3366 11776 3366 0 net18
rlabel metal1 10580 2346 10580 2346 0 net19
rlabel metal2 12650 38590 12650 38590 0 net2
rlabel metal1 2254 4114 2254 4114 0 net20
rlabel metal1 11408 2414 11408 2414 0 net21
rlabel metal2 2530 8806 2530 8806 0 net22
rlabel metal1 9706 2414 9706 2414 0 net23
rlabel metal1 12604 7378 12604 7378 0 net24
rlabel metal1 3496 2414 3496 2414 0 net25
rlabel metal1 1702 4046 1702 4046 0 net26
rlabel metal1 4462 2414 4462 2414 0 net27
rlabel metal1 3082 4590 3082 4590 0 net28
rlabel metal1 6808 3706 6808 3706 0 net29
rlabel metal1 14812 14382 14812 14382 0 net3
rlabel metal1 1702 5712 1702 5712 0 net30
rlabel metal1 5106 2516 5106 2516 0 net31
rlabel metal1 4462 6290 4462 6290 0 net32
rlabel metal1 14214 3026 14214 3026 0 net33
rlabel metal1 6210 2448 6210 2448 0 net34
rlabel metal1 7774 2414 7774 2414 0 net35
rlabel metal2 15594 4828 15594 4828 0 net36
rlabel metal1 8188 2414 8188 2414 0 net37
rlabel metal1 16146 6630 16146 6630 0 net38
rlabel metal1 9982 2482 9982 2482 0 net39
rlabel metal1 1748 21522 1748 21522 0 net4
rlabel metal1 5934 2414 5934 2414 0 net40
rlabel metal1 15640 2346 15640 2346 0 net41
rlabel metal1 14306 2448 14306 2448 0 net42
rlabel metal1 14490 5814 14490 5814 0 net43
rlabel metal1 15502 5270 15502 5270 0 net44
rlabel metal1 13064 3706 13064 3706 0 net45
rlabel metal1 14490 6358 14490 6358 0 net46
rlabel metal1 14950 8602 14950 8602 0 net47
rlabel metal1 13248 7854 13248 7854 0 net48
rlabel metal1 1978 11084 1978 11084 0 net49
rlabel metal1 1794 21998 1794 21998 0 net5
rlabel metal2 4738 12478 4738 12478 0 net50
rlabel metal2 6210 7888 6210 7888 0 net51
rlabel metal1 2346 8568 2346 8568 0 net52
rlabel metal2 1702 11900 1702 11900 0 net53
rlabel metal1 1610 9928 1610 9928 0 net54
rlabel metal1 2070 12274 2070 12274 0 net55
rlabel metal2 1702 9146 1702 9146 0 net56
rlabel metal1 2231 26962 2231 26962 0 net57
rlabel metal1 3450 31790 3450 31790 0 net58
rlabel metal1 13064 29138 13064 29138 0 net59
rlabel metal2 3266 15491 3266 15491 0 net6
rlabel metal1 13064 33082 13064 33082 0 net60
rlabel metal1 8326 38250 8326 38250 0 net61
rlabel metal1 5842 26282 5842 26282 0 net62
rlabel metal2 13478 30770 13478 30770 0 net63
rlabel metal1 6440 13362 6440 13362 0 net64
rlabel metal1 13570 19856 13570 19856 0 net65
rlabel metal1 6210 15538 6210 15538 0 net66
rlabel metal2 14674 6188 14674 6188 0 net67
rlabel metal2 11868 4114 11868 4114 0 net68
rlabel metal2 12558 19006 12558 19006 0 net69
rlabel metal2 2714 18717 2714 18717 0 net7
rlabel metal2 12742 28050 12742 28050 0 net70
rlabel metal1 13892 28662 13892 28662 0 net71
rlabel metal1 7958 12818 7958 12818 0 net72
rlabel viali 10914 31790 10914 31790 0 net73
rlabel metal1 9246 35632 9246 35632 0 net74
rlabel metal1 2530 5203 2530 5203 0 net75
rlabel metal1 1978 9010 1978 9010 0 net76
rlabel metal2 14766 4794 14766 4794 0 net77
rlabel metal1 14490 7412 14490 7412 0 net78
rlabel metal1 14122 8908 14122 8908 0 net79
rlabel metal2 16146 22406 16146 22406 0 net8
rlabel metal1 3772 10642 3772 10642 0 net80
rlabel metal1 14306 14246 14306 14246 0 net81
rlabel metal1 6026 32470 6026 32470 0 net82
rlabel metal1 12650 29206 12650 29206 0 net83
rlabel metal2 5566 33932 5566 33932 0 net84
rlabel via1 9793 23698 9793 23698 0 net85
rlabel metal1 5014 25670 5014 25670 0 net86
rlabel metal1 12374 14416 12374 14416 0 net87
rlabel metal1 2185 20502 2185 20502 0 net88
rlabel metal1 6992 10642 6992 10642 0 net89
rlabel metal1 16008 15470 16008 15470 0 net9
rlabel metal1 7958 12206 7958 12206 0 net90
rlabel metal1 10580 9690 10580 9690 0 net91
rlabel metal1 15640 13906 15640 13906 0 net92
rlabel metal1 15686 16558 15686 16558 0 net93
rlabel metal2 15502 11968 15502 11968 0 net94
rlabel metal2 6762 17408 6762 17408 0 net95
rlabel metal1 15686 15130 15686 15130 0 net96
rlabel metal1 15732 12138 15732 12138 0 net97
rlabel metal1 2484 18802 2484 18802 0 net98
rlabel metal1 3266 19346 3266 19346 0 net99
rlabel metal2 690 1010 690 1010 0 reg0[0]
rlabel metal2 11638 1520 11638 1520 0 reg0[1]
rlabel metal2 9706 1520 9706 1520 0 reg0[2]
rlabel metal2 1978 1367 1978 1367 0 reg0[3]
rlabel metal2 10994 1520 10994 1520 0 reg0[4]
rlabel metal3 866 9588 866 9588 0 reg0[5]
rlabel metal2 9062 1520 9062 1520 0 reg0[6]
rlabel metal2 12282 1520 12282 1520 0 reg0[7]
rlabel metal2 3266 1367 3266 1367 0 reg1[0]
rlabel metal2 1334 1027 1334 1027 0 reg1[1]
rlabel metal2 3910 1520 3910 1520 0 reg1[2]
rlabel metal2 2622 1231 2622 1231 0 reg1[3]
rlabel metal2 5842 1656 5842 1656 0 reg1[4]
rlabel metal2 46 1044 46 1044 0 reg1[5]
rlabel metal2 5198 959 5198 959 0 reg1[6]
rlabel metal2 4554 1520 4554 1520 0 reg1[7]
rlabel metal2 13570 1520 13570 1520 0 reg2[0]
rlabel metal2 7130 891 7130 891 0 reg2[1]
rlabel metal2 7774 1520 7774 1520 0 reg2[2]
rlabel metal1 16238 3910 16238 3910 0 reg2[3]
rlabel metal2 8418 959 8418 959 0 reg2[4]
rlabel metal1 16422 3978 16422 3978 0 reg2[5]
rlabel metal2 10350 1520 10350 1520 0 reg2[6]
rlabel metal2 6486 1554 6486 1554 0 reg2[7]
rlabel metal1 16560 4046 16560 4046 0 reg3[0]
rlabel metal1 15870 3638 15870 3638 0 reg3[1]
rlabel metal2 14214 1044 14214 1044 0 reg3[2]
rlabel metal2 14858 942 14858 942 0 reg3[3]
rlabel metal2 12926 1520 12926 1520 0 reg3[4]
rlabel metal1 16514 5542 16514 5542 0 reg3[5]
rlabel metal2 16422 10353 16422 10353 0 reg3[6]
rlabel metal1 16514 8330 16514 8330 0 reg3[7]
rlabel metal1 1334 11322 1334 11322 0 reg4[0]
rlabel metal1 1426 12954 1426 12954 0 reg4[1]
rlabel metal2 2806 8517 2806 8517 0 reg4[2]
rlabel metal2 2990 7633 2990 7633 0 reg4[3]
rlabel metal3 751 12308 751 12308 0 reg4[4]
rlabel metal1 1426 9350 1426 9350 0 reg4[5]
rlabel metal3 1280 10948 1280 10948 0 reg4[6]
rlabel metal3 751 8908 751 8908 0 reg4[7]
rlabel via2 3082 20451 3082 20451 0 rst
rlabel metal3 751 19788 751 19788 0 rx
rlabel metal3 751 26588 751 26588 0 tx
rlabel metal1 3956 24242 3956 24242 0 uart_receive.baud_clk
rlabel metal1 4554 21522 4554 21522 0 uart_receive.baud_clk2
rlabel metal1 2024 19822 2024 19822 0 uart_receive.baud_clk3
rlabel metal1 2208 35258 2208 35258 0 uart_receive.baud_rate_gen.count\[0\]
rlabel metal1 4140 26962 4140 26962 0 uart_receive.baud_rate_gen.count\[10\]
rlabel metal1 4876 28390 4876 28390 0 uart_receive.baud_rate_gen.count\[11\]
rlabel metal1 1978 36108 1978 36108 0 uart_receive.baud_rate_gen.count\[1\]
rlabel metal1 5336 36142 5336 36142 0 uart_receive.baud_rate_gen.count\[2\]
rlabel metal2 5750 35462 5750 35462 0 uart_receive.baud_rate_gen.count\[3\]
rlabel metal1 5888 32402 5888 32402 0 uart_receive.baud_rate_gen.count\[4\]
rlabel metal1 5566 32368 5566 32368 0 uart_receive.baud_rate_gen.count\[5\]
rlabel metal1 4554 32266 4554 32266 0 uart_receive.baud_rate_gen.count\[6\]
rlabel metal1 5428 30362 5428 30362 0 uart_receive.baud_rate_gen.count\[7\]
rlabel metal1 4002 29580 4002 29580 0 uart_receive.baud_rate_gen.count\[8\]
rlabel metal1 5014 28560 5014 28560 0 uart_receive.baud_rate_gen.count\[9\]
rlabel metal2 3082 21318 3082 21318 0 uart_receive.n328_o\[0\]
rlabel metal1 3848 19754 3848 19754 0 uart_receive.n328_o\[1\]
rlabel metal2 4646 24820 4646 24820 0 uart_receive.n345_q
rlabel metal1 2162 18700 2162 18700 0 uart_receive.n346_q\[0\]
rlabel metal1 2162 19890 2162 19890 0 uart_receive.n346_q\[1\]
rlabel metal1 2254 15606 2254 15606 0 uart_receive.n352_o
rlabel metal1 2346 15538 2346 15538 0 uart_receive.n354_o
rlabel metal1 2944 18734 2944 18734 0 uart_receive.n360_o
rlabel metal1 2162 18156 2162 18156 0 uart_receive.n370_o
rlabel metal1 14398 15504 14398 15504 0 uart_receive.n372_o
rlabel metal1 12742 5134 12742 5134 0 uart_receive.n374_o
rlabel metal1 1886 13838 1886 13838 0 uart_receive.n376_o
rlabel metal1 13754 11050 13754 11050 0 uart_receive.n378_o
rlabel metal1 14490 12784 14490 12784 0 uart_receive.n380_o
rlabel metal2 14306 16626 14306 16626 0 uart_receive.n382_o
rlabel metal1 14582 18836 14582 18836 0 uart_receive.n384_o
rlabel metal2 7958 25602 7958 25602 0 uart_transmit.baud_clk
rlabel metal1 12558 30328 12558 30328 0 uart_transmit.baud_rate_gen.count\[0\]
rlabel metal1 7406 31926 7406 31926 0 uart_transmit.baud_rate_gen.count\[10\]
rlabel metal1 8188 31450 8188 31450 0 uart_transmit.baud_rate_gen.count\[11\]
rlabel metal1 9062 31790 9062 31790 0 uart_transmit.baud_rate_gen.count\[12\]
rlabel metal2 12650 30549 12650 30549 0 uart_transmit.baud_rate_gen.count\[1\]
rlabel metal2 14122 30430 14122 30430 0 uart_transmit.baud_rate_gen.count\[2\]
rlabel metal1 14260 29614 14260 29614 0 uart_transmit.baud_rate_gen.count\[3\]
rlabel metal1 12834 26316 12834 26316 0 uart_transmit.baud_rate_gen.count\[4\]
rlabel metal1 12650 29104 12650 29104 0 uart_transmit.baud_rate_gen.count\[5\]
rlabel metal2 11178 26180 11178 26180 0 uart_transmit.baud_rate_gen.count\[6\]
rlabel metal1 10258 27302 10258 27302 0 uart_transmit.baud_rate_gen.count\[7\]
rlabel metal1 8878 29614 8878 29614 0 uart_transmit.baud_rate_gen.count\[8\]
rlabel metal1 8142 28084 8142 28084 0 uart_transmit.baud_rate_gen.count\[9\]
rlabel metal1 7314 18836 7314 18836 0 uart_transmit.n167_o
rlabel metal2 13846 27744 13846 27744 0 uart_transmit.n224_q
rlabel metal1 8004 24378 8004 24378 0 uart_transmit.n226_q\[0\]
rlabel metal1 6854 25126 6854 25126 0 uart_transmit.n226_q\[1\]
rlabel metal1 7590 17170 7590 17170 0 uart_transmit.n227_q\[0\]
rlabel metal1 8786 16490 8786 16490 0 uart_transmit.n227_q\[1\]
rlabel metal1 7820 17578 7820 17578 0 uart_transmit.n227_q\[2\]
rlabel metal1 6624 21522 6624 21522 0 uart_transmit.n227_q\[3\]
rlabel metal1 6670 21862 6670 21862 0 uart_transmit.n227_q\[4\]
rlabel metal2 9246 19924 9246 19924 0 uart_transmit.n231_o
rlabel metal2 8142 16116 8142 16116 0 uart_transmit.n232_o
rlabel metal1 7360 16490 7360 16490 0 uart_transmit.n233_o
rlabel metal2 9522 14348 9522 14348 0 uart_transmit.n234_o
rlabel metal1 7820 15538 7820 15538 0 uart_transmit.n235_o
rlabel metal1 9522 13804 9522 13804 0 uart_transmit.n236_o
rlabel metal1 9844 16218 9844 16218 0 uart_transmit.n237_o
<< properties >>
string FIXED_BBOX 0 0 18000 42000
<< end >>
