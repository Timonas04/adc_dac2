VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.000000 ;
    ANTENNADIFFAREA 17.400000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 74.440 122.650 87.610 130.490 ;
      LAYER pwell ;
        RECT 74.450 118.150 87.620 121.940 ;
        RECT 74.450 110.660 88.300 117.880 ;
      LAYER nwell ;
        RECT 123.065 110.755 129.915 116.750 ;
      LAYER pwell ;
        RECT 74.450 104.670 85.340 110.660 ;
      LAYER nwell ;
        RECT 121.045 104.565 129.915 110.755 ;
        RECT 123.065 104.560 129.915 104.565 ;
      LAYER pwell ;
        RECT 121.040 104.260 123.150 104.265 ;
        RECT 121.040 101.165 129.915 104.260 ;
        RECT 123.065 97.160 129.915 101.165 ;
        RECT 149.600 94.520 159.010 100.510 ;
        RECT 125.920 88.000 159.010 94.520 ;
        RECT 75.535 64.505 79.635 86.665 ;
      LAYER nwell ;
        RECT 80.015 83.205 89.975 87.325 ;
        RECT 80.015 75.895 90.205 83.205 ;
        RECT 80.010 75.815 90.205 75.895 ;
        RECT 80.010 67.480 88.510 75.815 ;
        RECT 80.010 64.590 86.200 67.480 ;
        RECT 80.010 64.505 86.215 64.590 ;
      LAYER pwell ;
        RECT 75.535 64.415 79.640 64.505 ;
        RECT 76.540 62.480 79.640 64.415 ;
      LAYER nwell ;
        RECT 80.025 62.565 86.215 64.505 ;
      LAYER pwell ;
        RECT 92.535 64.505 96.635 86.665 ;
      LAYER nwell ;
        RECT 97.015 83.205 106.975 87.325 ;
        RECT 97.015 75.895 107.205 83.205 ;
        RECT 97.010 75.815 107.205 75.895 ;
        RECT 97.010 67.480 105.510 75.815 ;
        RECT 97.010 64.590 103.200 67.480 ;
        RECT 97.010 64.505 103.215 64.590 ;
      LAYER pwell ;
        RECT 92.535 64.415 96.640 64.505 ;
      LAYER nwell ;
        RECT 80.025 62.480 90.220 62.565 ;
      LAYER pwell ;
        RECT 93.540 62.480 96.640 64.415 ;
      LAYER nwell ;
        RECT 97.025 62.565 103.215 64.505 ;
      LAYER pwell ;
        RECT 109.535 64.505 113.635 86.665 ;
      LAYER nwell ;
        RECT 114.015 83.205 123.975 87.325 ;
        RECT 114.015 75.895 124.205 83.205 ;
        RECT 114.010 75.815 124.205 75.895 ;
        RECT 114.010 67.480 122.510 75.815 ;
        RECT 114.010 64.590 120.200 67.480 ;
        RECT 114.010 64.505 120.215 64.590 ;
      LAYER pwell ;
        RECT 109.535 64.415 113.640 64.505 ;
      LAYER nwell ;
        RECT 97.025 62.480 107.220 62.565 ;
      LAYER pwell ;
        RECT 110.540 62.480 113.640 64.415 ;
      LAYER nwell ;
        RECT 114.025 62.565 120.215 64.505 ;
      LAYER pwell ;
        RECT 126.535 64.505 130.635 86.665 ;
      LAYER nwell ;
        RECT 131.015 83.205 140.975 87.325 ;
        RECT 131.015 75.895 141.205 83.205 ;
        RECT 131.010 75.815 141.205 75.895 ;
        RECT 131.010 67.480 139.510 75.815 ;
        RECT 131.010 64.590 137.200 67.480 ;
        RECT 131.010 64.505 137.215 64.590 ;
      LAYER pwell ;
        RECT 126.535 64.415 130.640 64.505 ;
      LAYER nwell ;
        RECT 114.025 62.480 124.220 62.565 ;
      LAYER pwell ;
        RECT 127.540 62.480 130.640 64.415 ;
      LAYER nwell ;
        RECT 131.025 62.565 137.215 64.505 ;
      LAYER pwell ;
        RECT 143.535 64.505 147.635 86.665 ;
      LAYER nwell ;
        RECT 148.015 83.205 157.975 87.325 ;
        RECT 148.015 75.895 158.205 83.205 ;
        RECT 148.010 75.815 158.205 75.895 ;
        RECT 148.010 67.480 156.510 75.815 ;
        RECT 148.010 64.590 154.200 67.480 ;
        RECT 148.010 64.505 154.215 64.590 ;
      LAYER pwell ;
        RECT 143.535 64.415 147.640 64.505 ;
      LAYER nwell ;
        RECT 131.025 62.480 141.220 62.565 ;
      LAYER pwell ;
        RECT 144.540 62.480 147.640 64.415 ;
      LAYER nwell ;
        RECT 148.025 62.565 154.215 64.505 ;
        RECT 148.025 62.480 158.220 62.565 ;
      LAYER pwell ;
        RECT 75.545 60.370 79.645 62.480 ;
      LAYER nwell ;
        RECT 80.030 60.455 90.220 62.480 ;
      LAYER pwell ;
        RECT 92.545 60.370 96.645 62.480 ;
      LAYER nwell ;
        RECT 97.030 60.455 107.220 62.480 ;
      LAYER pwell ;
        RECT 109.545 60.370 113.645 62.480 ;
      LAYER nwell ;
        RECT 114.030 60.455 124.220 62.480 ;
      LAYER pwell ;
        RECT 126.545 60.370 130.645 62.480 ;
      LAYER nwell ;
        RECT 131.030 60.455 141.220 62.480 ;
      LAYER pwell ;
        RECT 143.545 60.370 147.645 62.480 ;
      LAYER nwell ;
        RECT 148.030 60.455 158.220 62.480 ;
        RECT 22.330 57.825 58.590 59.430 ;
      LAYER pwell ;
        RECT 22.525 56.625 23.895 57.435 ;
        RECT 23.905 56.625 29.415 57.435 ;
        RECT 30.830 57.305 32.175 57.535 ;
        RECT 30.345 56.625 32.175 57.305 ;
        RECT 32.315 56.625 35.315 57.535 ;
        RECT 35.415 56.710 35.845 57.495 ;
        RECT 39.440 57.305 40.360 57.535 ;
        RECT 36.895 56.625 40.360 57.305 ;
        RECT 41.385 57.305 42.730 57.535 ;
        RECT 45.880 57.305 46.800 57.535 ;
        RECT 41.385 56.625 43.215 57.305 ;
        RECT 43.335 56.625 46.800 57.305 ;
        RECT 46.905 56.625 48.275 57.405 ;
        RECT 48.295 56.710 48.725 57.495 ;
        RECT 49.665 57.305 51.010 57.535 ;
        RECT 49.665 56.625 51.495 57.305 ;
        RECT 51.505 56.625 52.875 57.435 ;
        RECT 52.885 56.625 54.255 57.405 ;
        RECT 54.265 56.625 55.635 57.405 ;
        RECT 55.645 56.625 57.015 57.405 ;
        RECT 57.025 56.625 58.395 57.435 ;
        RECT 22.665 56.415 22.835 56.625 ;
        RECT 24.045 56.415 24.215 56.625 ;
        RECT 27.720 56.465 27.840 56.575 ;
        RECT 29.575 56.470 29.735 56.580 ;
        RECT 30.485 56.435 30.655 56.625 ;
        RECT 35.085 56.415 35.255 56.625 ;
        RECT 35.545 56.415 35.715 56.605 ;
        RECT 36.015 56.470 36.175 56.580 ;
        RECT 36.925 56.435 37.095 56.625 ;
        RECT 40.615 56.470 40.775 56.580 ;
        RECT 42.905 56.435 43.075 56.625 ;
        RECT 43.365 56.435 43.535 56.625 ;
        RECT 47.055 56.605 47.225 56.625 ;
        RECT 44.745 56.435 44.915 56.605 ;
        RECT 44.745 56.415 44.910 56.435 ;
        RECT 45.205 56.415 45.375 56.605 ;
        RECT 47.045 56.435 47.225 56.605 ;
        RECT 47.045 56.415 47.215 56.435 ;
        RECT 48.885 56.415 49.055 56.605 ;
        RECT 51.185 56.435 51.355 56.625 ;
        RECT 51.645 56.435 51.815 56.625 ;
        RECT 52.105 56.415 52.275 56.605 ;
        RECT 53.945 56.435 54.115 56.625 ;
        RECT 55.325 56.435 55.495 56.625 ;
        RECT 56.695 56.415 56.865 56.625 ;
        RECT 58.085 56.415 58.255 56.625 ;
        RECT 22.525 55.605 23.895 56.415 ;
        RECT 23.905 55.605 27.575 56.415 ;
        RECT 28.085 55.735 35.395 56.415 ;
        RECT 35.405 55.735 42.715 56.415 ;
        RECT 28.085 55.505 29.435 55.735 ;
        RECT 30.970 55.515 31.880 55.735 ;
        RECT 38.920 55.515 39.830 55.735 ;
        RECT 41.365 55.505 42.715 55.735 ;
        RECT 43.075 55.735 44.910 56.415 ;
        RECT 45.065 55.735 46.895 56.415 ;
        RECT 43.075 55.505 44.005 55.735 ;
        RECT 45.550 55.505 46.895 55.735 ;
        RECT 46.915 55.505 48.265 56.415 ;
        RECT 48.295 55.545 48.725 56.330 ;
        RECT 48.825 55.505 51.825 56.415 ;
        RECT 52.075 55.735 55.540 56.415 ;
        RECT 54.620 55.505 55.540 55.735 ;
        RECT 55.645 55.635 57.015 56.415 ;
        RECT 57.025 55.605 58.395 56.415 ;
      LAYER nwell ;
        RECT 22.330 52.385 58.590 55.215 ;
      LAYER pwell ;
        RECT 22.525 51.185 23.895 51.995 ;
        RECT 27.420 51.865 28.330 52.085 ;
        RECT 29.865 51.865 31.215 52.095 ;
        RECT 23.905 51.185 31.215 51.865 ;
        RECT 31.360 51.865 32.280 52.095 ;
        RECT 31.360 51.185 34.825 51.865 ;
        RECT 35.415 51.270 35.845 52.055 ;
        RECT 35.865 51.865 36.795 52.095 ;
        RECT 41.515 51.865 42.445 52.095 ;
        RECT 35.865 51.185 39.765 51.865 ;
        RECT 40.610 51.185 42.445 51.865 ;
        RECT 42.775 51.185 44.125 52.095 ;
        RECT 47.660 51.865 48.570 52.085 ;
        RECT 50.105 51.865 51.455 52.095 ;
        RECT 53.015 51.865 53.945 52.095 ;
        RECT 44.145 51.185 51.455 51.865 ;
        RECT 52.110 51.185 53.945 51.865 ;
        RECT 54.265 51.185 55.635 51.965 ;
        RECT 55.645 51.185 57.015 51.965 ;
        RECT 57.025 51.185 58.395 51.995 ;
        RECT 22.665 50.975 22.835 51.185 ;
        RECT 24.045 50.995 24.215 51.185 ;
        RECT 25.425 50.975 25.595 51.165 ;
        RECT 26.160 50.975 26.330 51.165 ;
        RECT 30.025 50.975 30.195 51.165 ;
        RECT 34.625 50.995 34.795 51.185 ;
        RECT 35.080 51.025 35.200 51.135 ;
        RECT 36.280 50.995 36.450 51.185 ;
        RECT 40.610 51.165 40.775 51.185 ;
        RECT 40.145 51.135 40.315 51.165 ;
        RECT 40.140 51.025 40.315 51.135 ;
        RECT 40.145 50.975 40.315 51.025 ;
        RECT 40.605 50.995 40.775 51.165 ;
        RECT 43.825 50.975 43.995 51.185 ;
        RECT 44.285 50.975 44.455 51.185 ;
        RECT 52.110 51.165 52.275 51.185 ;
        RECT 22.525 50.165 23.895 50.975 ;
        RECT 23.905 50.295 25.735 50.975 ;
        RECT 25.745 50.295 29.645 50.975 ;
        RECT 23.905 50.065 25.250 50.295 ;
        RECT 25.745 50.065 26.675 50.295 ;
        RECT 29.885 50.165 31.255 50.975 ;
        RECT 31.350 50.295 40.455 50.975 ;
        RECT 40.560 50.295 44.025 50.975 ;
        RECT 40.560 50.065 41.480 50.295 ;
        RECT 44.145 50.165 45.515 50.975 ;
        RECT 45.670 50.945 45.840 51.165 ;
        RECT 48.885 50.975 49.055 51.165 ;
        RECT 51.640 51.025 51.760 51.135 ;
        RECT 52.105 50.995 52.275 51.165 ;
        RECT 52.565 50.975 52.735 51.165 ;
        RECT 54.405 50.995 54.575 51.185 ;
        RECT 56.255 51.020 56.415 51.130 ;
        RECT 56.695 50.995 56.865 51.185 ;
        RECT 58.085 50.975 58.255 51.185 ;
        RECT 47.330 50.945 48.275 50.975 ;
        RECT 45.525 50.265 48.275 50.945 ;
        RECT 47.330 50.065 48.275 50.265 ;
        RECT 48.295 50.105 48.725 50.890 ;
        RECT 48.825 50.065 52.275 50.975 ;
        RECT 52.505 50.065 55.955 50.975 ;
        RECT 57.025 50.165 58.395 50.975 ;
      LAYER nwell ;
        RECT 22.330 46.945 58.590 49.775 ;
      LAYER pwell ;
        RECT 22.525 45.745 23.895 46.555 ;
        RECT 23.905 46.425 24.835 46.655 ;
        RECT 31.560 46.425 32.470 46.645 ;
        RECT 34.005 46.425 35.355 46.655 ;
        RECT 23.905 45.745 27.805 46.425 ;
        RECT 28.045 45.745 35.355 46.425 ;
        RECT 35.415 45.830 35.845 46.615 ;
        RECT 39.380 46.425 40.290 46.645 ;
        RECT 41.825 46.425 43.175 46.655 ;
        RECT 35.865 45.745 43.175 46.425 ;
        RECT 43.685 46.425 45.050 46.655 ;
        RECT 43.685 45.745 46.895 46.425 ;
        RECT 47.905 45.745 50.905 46.655 ;
        RECT 51.045 45.745 52.395 46.655 ;
        RECT 52.965 45.745 56.415 46.655 ;
        RECT 57.025 45.745 58.395 46.555 ;
        RECT 22.665 45.535 22.835 45.745 ;
        RECT 24.320 45.555 24.490 45.745 ;
        RECT 28.185 45.555 28.355 45.745 ;
        RECT 30.945 45.535 31.115 45.725 ;
        RECT 31.405 45.535 31.575 45.725 ;
        RECT 34.160 45.585 34.280 45.695 ;
        RECT 34.625 45.535 34.795 45.725 ;
        RECT 36.005 45.555 36.175 45.745 ;
        RECT 43.360 45.585 43.480 45.695 ;
        RECT 46.580 45.555 46.750 45.745 ;
        RECT 47.045 45.535 47.215 45.725 ;
        RECT 47.515 45.580 47.675 45.690 ;
        RECT 47.965 45.555 48.135 45.745 ;
        RECT 51.190 45.725 51.360 45.745 ;
        RECT 22.525 44.725 23.895 45.535 ;
        RECT 23.945 44.855 31.255 45.535 ;
        RECT 23.945 44.625 25.295 44.855 ;
        RECT 26.830 44.635 27.740 44.855 ;
        RECT 31.265 44.725 34.015 45.535 ;
        RECT 34.485 44.855 43.590 45.535 ;
        RECT 43.780 44.855 47.245 45.535 ;
        RECT 48.880 45.505 49.050 45.725 ;
        RECT 51.185 45.555 51.360 45.725 ;
        RECT 52.560 45.585 52.680 45.695 ;
        RECT 53.025 45.555 53.195 45.745 ;
        RECT 53.940 45.585 54.060 45.695 ;
        RECT 51.185 45.535 51.355 45.555 ;
        RECT 55.320 45.535 55.490 45.725 ;
        RECT 56.705 45.695 56.875 45.725 ;
        RECT 56.700 45.585 56.875 45.695 ;
        RECT 56.705 45.535 56.875 45.585 ;
        RECT 58.085 45.535 58.255 45.745 ;
        RECT 50.080 45.505 51.035 45.535 ;
        RECT 43.780 44.625 44.700 44.855 ;
        RECT 48.295 44.665 48.725 45.450 ;
        RECT 48.755 44.825 51.035 45.505 ;
        RECT 50.080 44.625 51.035 44.825 ;
        RECT 51.045 44.725 53.795 45.535 ;
        RECT 54.285 44.625 55.635 45.535 ;
        RECT 55.645 44.755 57.015 45.535 ;
        RECT 57.025 44.725 58.395 45.535 ;
      LAYER nwell ;
        RECT 22.330 41.505 58.590 44.335 ;
      LAYER pwell ;
        RECT 22.525 40.305 23.895 41.115 ;
        RECT 23.905 40.305 25.275 41.115 ;
        RECT 27.940 40.985 28.860 41.215 ;
        RECT 25.395 40.305 28.860 40.985 ;
        RECT 29.060 40.985 29.980 41.215 ;
        RECT 29.060 40.305 32.525 40.985 ;
        RECT 32.645 40.305 35.395 41.115 ;
        RECT 35.415 40.390 35.845 41.175 ;
        RECT 35.885 40.305 37.235 41.215 ;
        RECT 37.315 40.305 41.375 41.215 ;
        RECT 41.480 40.985 42.400 41.215 ;
        RECT 41.480 40.305 44.945 40.985 ;
        RECT 45.065 40.305 46.435 41.115 ;
        RECT 46.445 41.015 47.395 41.215 ;
        RECT 46.445 40.335 50.115 41.015 ;
        RECT 46.445 40.305 47.395 40.335 ;
        RECT 22.665 40.095 22.835 40.305 ;
        RECT 24.045 40.115 24.215 40.305 ;
        RECT 25.425 40.095 25.595 40.305 ;
        RECT 25.880 40.145 26.000 40.255 ;
        RECT 26.620 40.095 26.790 40.285 ;
        RECT 30.485 40.095 30.655 40.285 ;
        RECT 32.325 40.115 32.495 40.305 ;
        RECT 32.785 40.115 32.955 40.305 ;
        RECT 36.920 40.115 37.090 40.305 ;
        RECT 38.120 40.095 38.290 40.285 ;
        RECT 41.065 40.115 41.235 40.305 ;
        RECT 44.745 40.115 44.915 40.305 ;
        RECT 45.205 40.095 45.375 40.305 ;
        RECT 45.665 40.095 45.835 40.285 ;
        RECT 49.800 40.115 49.970 40.335 ;
        RECT 50.125 40.305 51.475 41.215 ;
        RECT 51.505 40.305 52.875 41.085 ;
        RECT 53.025 40.305 56.475 41.215 ;
        RECT 57.025 40.305 58.395 41.115 ;
        RECT 50.270 40.115 50.440 40.305 ;
        RECT 51.655 40.285 51.825 40.305 ;
        RECT 51.640 40.115 51.825 40.285 ;
        RECT 52.115 40.140 52.275 40.250 ;
        RECT 51.640 40.095 51.810 40.115 ;
        RECT 56.245 40.095 56.415 40.305 ;
        RECT 56.700 40.145 56.820 40.255 ;
        RECT 58.085 40.095 58.255 40.305 ;
        RECT 22.525 39.285 23.895 40.095 ;
        RECT 23.905 39.415 25.735 40.095 ;
        RECT 26.205 39.415 30.105 40.095 ;
        RECT 30.345 39.415 37.655 40.095 ;
        RECT 23.905 39.185 25.250 39.415 ;
        RECT 26.205 39.185 27.135 39.415 ;
        RECT 33.860 39.195 34.770 39.415 ;
        RECT 36.305 39.185 37.655 39.415 ;
        RECT 37.705 39.415 41.605 40.095 ;
        RECT 41.940 39.415 45.405 40.095 ;
        RECT 37.705 39.185 38.635 39.415 ;
        RECT 41.940 39.185 42.860 39.415 ;
        RECT 45.525 39.285 48.275 40.095 ;
        RECT 48.295 39.225 48.725 40.010 ;
        RECT 49.035 39.185 51.955 40.095 ;
        RECT 53.025 39.185 56.475 40.095 ;
        RECT 57.025 39.285 58.395 40.095 ;
      LAYER nwell ;
        RECT 22.330 36.065 58.590 38.895 ;
      LAYER pwell ;
        RECT 22.525 34.865 23.895 35.675 ;
        RECT 27.420 35.545 28.330 35.765 ;
        RECT 29.865 35.545 31.215 35.775 ;
        RECT 23.905 34.865 31.215 35.545 ;
        RECT 31.265 34.865 34.935 35.675 ;
        RECT 35.415 34.950 35.845 35.735 ;
        RECT 39.380 35.545 40.290 35.765 ;
        RECT 41.825 35.545 43.175 35.775 ;
        RECT 45.070 35.545 46.435 35.775 ;
        RECT 35.865 34.865 43.175 35.545 ;
        RECT 43.225 34.865 46.435 35.545 ;
        RECT 46.445 34.865 49.195 35.675 ;
        RECT 52.320 35.545 53.240 35.775 ;
        RECT 49.775 34.865 53.240 35.545 ;
        RECT 53.425 34.865 56.425 35.775 ;
        RECT 57.025 34.865 58.395 35.675 ;
        RECT 75.535 35.505 79.635 57.665 ;
      LAYER nwell ;
        RECT 80.015 54.205 89.975 58.325 ;
        RECT 80.015 46.895 90.205 54.205 ;
        RECT 80.010 46.815 90.205 46.895 ;
        RECT 80.010 38.480 88.510 46.815 ;
        RECT 80.010 35.590 86.200 38.480 ;
        RECT 80.010 35.505 86.215 35.590 ;
      LAYER pwell ;
        RECT 75.535 35.415 79.640 35.505 ;
        RECT 22.665 34.655 22.835 34.865 ;
        RECT 24.045 34.675 24.215 34.865 ;
        RECT 25.425 34.655 25.595 34.845 ;
        RECT 25.895 34.700 26.055 34.810 ;
        RECT 26.805 34.655 26.975 34.845 ;
        RECT 30.495 34.700 30.655 34.810 ;
        RECT 31.405 34.655 31.575 34.865 ;
        RECT 35.080 34.705 35.200 34.815 ;
        RECT 36.005 34.675 36.175 34.865 ;
        RECT 38.490 34.655 38.660 34.845 ;
        RECT 39.225 34.655 39.395 34.845 ;
        RECT 41.065 34.655 41.235 34.845 ;
        RECT 43.370 34.675 43.540 34.865 ;
        RECT 46.585 34.675 46.755 34.865 ;
        RECT 49.160 34.655 49.330 34.845 ;
        RECT 49.340 34.705 49.460 34.815 ;
        RECT 49.805 34.675 49.975 34.865 ;
        RECT 53.025 34.655 53.195 34.845 ;
        RECT 53.485 34.675 53.655 34.865 ;
        RECT 22.525 33.845 23.895 34.655 ;
        RECT 23.905 33.975 25.735 34.655 ;
        RECT 26.775 33.975 30.240 34.655 ;
        RECT 31.375 33.975 34.840 34.655 ;
        RECT 35.175 33.975 39.075 34.655 ;
        RECT 23.905 33.745 25.250 33.975 ;
        RECT 29.320 33.745 30.240 33.975 ;
        RECT 33.920 33.745 34.840 33.975 ;
        RECT 38.145 33.745 39.075 33.975 ;
        RECT 39.085 33.845 40.915 34.655 ;
        RECT 40.925 33.975 48.235 34.655 ;
        RECT 44.440 33.755 45.350 33.975 ;
        RECT 46.885 33.745 48.235 33.975 ;
        RECT 48.295 33.785 48.725 34.570 ;
        RECT 48.745 33.975 52.645 34.655 ;
        RECT 48.745 33.745 49.675 33.975 ;
        RECT 52.885 33.875 54.255 34.655 ;
        RECT 54.265 34.625 55.210 34.655 ;
        RECT 56.700 34.625 56.870 34.845 ;
        RECT 58.085 34.655 58.255 34.865 ;
        RECT 54.265 33.945 57.015 34.625 ;
        RECT 54.265 33.745 55.210 33.945 ;
        RECT 57.025 33.845 58.395 34.655 ;
        RECT 76.540 33.480 79.640 35.415 ;
      LAYER nwell ;
        RECT 80.025 33.565 86.215 35.505 ;
      LAYER pwell ;
        RECT 92.535 35.505 96.635 57.665 ;
      LAYER nwell ;
        RECT 97.015 54.205 106.975 58.325 ;
        RECT 97.015 46.895 107.205 54.205 ;
        RECT 97.010 46.815 107.205 46.895 ;
        RECT 97.010 38.480 105.510 46.815 ;
        RECT 97.010 35.590 103.200 38.480 ;
        RECT 97.010 35.505 103.215 35.590 ;
      LAYER pwell ;
        RECT 92.535 35.415 96.640 35.505 ;
      LAYER nwell ;
        RECT 80.025 33.480 90.220 33.565 ;
      LAYER pwell ;
        RECT 93.540 33.480 96.640 35.415 ;
      LAYER nwell ;
        RECT 97.025 33.565 103.215 35.505 ;
      LAYER pwell ;
        RECT 109.535 35.505 113.635 57.665 ;
      LAYER nwell ;
        RECT 114.015 54.205 123.975 58.325 ;
        RECT 114.015 46.895 124.205 54.205 ;
        RECT 114.010 46.815 124.205 46.895 ;
        RECT 114.010 38.480 122.510 46.815 ;
        RECT 114.010 35.590 120.200 38.480 ;
        RECT 114.010 35.505 120.215 35.590 ;
      LAYER pwell ;
        RECT 109.535 35.415 113.640 35.505 ;
      LAYER nwell ;
        RECT 97.025 33.480 107.220 33.565 ;
      LAYER pwell ;
        RECT 110.540 33.480 113.640 35.415 ;
      LAYER nwell ;
        RECT 114.025 33.565 120.215 35.505 ;
      LAYER pwell ;
        RECT 126.535 35.505 130.635 57.665 ;
      LAYER nwell ;
        RECT 131.015 54.205 140.975 58.325 ;
        RECT 131.015 46.895 141.205 54.205 ;
        RECT 131.010 46.815 141.205 46.895 ;
        RECT 131.010 38.480 139.510 46.815 ;
        RECT 131.010 35.590 137.200 38.480 ;
        RECT 131.010 35.505 137.215 35.590 ;
      LAYER pwell ;
        RECT 126.535 35.415 130.640 35.505 ;
      LAYER nwell ;
        RECT 114.025 33.480 124.220 33.565 ;
      LAYER pwell ;
        RECT 127.540 33.480 130.640 35.415 ;
      LAYER nwell ;
        RECT 131.025 33.565 137.215 35.505 ;
      LAYER pwell ;
        RECT 143.535 35.505 147.635 57.665 ;
      LAYER nwell ;
        RECT 148.015 54.205 157.975 58.325 ;
        RECT 148.015 46.895 158.205 54.205 ;
        RECT 148.010 46.815 158.205 46.895 ;
        RECT 148.010 38.480 156.510 46.815 ;
        RECT 148.010 35.590 154.200 38.480 ;
        RECT 148.010 35.505 154.215 35.590 ;
      LAYER pwell ;
        RECT 143.535 35.415 147.640 35.505 ;
      LAYER nwell ;
        RECT 131.025 33.480 141.220 33.565 ;
      LAYER pwell ;
        RECT 144.540 33.480 147.640 35.415 ;
      LAYER nwell ;
        RECT 148.025 33.565 154.215 35.505 ;
        RECT 148.025 33.480 158.220 33.565 ;
        RECT 22.330 30.625 58.590 33.455 ;
      LAYER pwell ;
        RECT 75.545 31.370 79.645 33.480 ;
      LAYER nwell ;
        RECT 80.030 31.455 90.220 33.480 ;
      LAYER pwell ;
        RECT 92.545 31.370 96.645 33.480 ;
      LAYER nwell ;
        RECT 97.030 31.455 107.220 33.480 ;
      LAYER pwell ;
        RECT 109.545 31.370 113.645 33.480 ;
      LAYER nwell ;
        RECT 114.030 31.455 124.220 33.480 ;
      LAYER pwell ;
        RECT 126.545 31.370 130.645 33.480 ;
      LAYER nwell ;
        RECT 131.030 31.455 141.220 33.480 ;
      LAYER pwell ;
        RECT 143.545 31.370 147.645 33.480 ;
      LAYER nwell ;
        RECT 148.030 31.455 158.220 33.480 ;
      LAYER pwell ;
        RECT 22.525 29.425 23.895 30.235 ;
        RECT 23.945 30.105 25.295 30.335 ;
        RECT 26.830 30.105 27.740 30.325 ;
        RECT 23.945 29.425 31.255 30.105 ;
        RECT 31.265 29.425 34.935 30.235 ;
        RECT 35.415 29.510 35.845 30.295 ;
        RECT 35.865 29.425 44.970 30.105 ;
        RECT 45.065 29.425 46.435 30.235 ;
        RECT 46.445 29.425 47.815 30.205 ;
        RECT 47.825 29.425 49.195 30.205 ;
        RECT 49.205 29.425 50.575 30.205 ;
        RECT 50.585 29.425 51.955 30.205 ;
        RECT 51.985 29.425 53.335 30.335 ;
        RECT 53.425 29.425 56.875 30.335 ;
        RECT 57.025 29.425 58.395 30.235 ;
        RECT 22.665 29.215 22.835 29.425 ;
        RECT 25.425 29.215 25.595 29.405 ;
        RECT 25.895 29.260 26.055 29.370 ;
        RECT 27.080 29.215 27.250 29.405 ;
        RECT 30.945 29.215 31.115 29.425 ;
        RECT 31.405 29.235 31.575 29.425 ;
        RECT 34.625 29.215 34.795 29.405 ;
        RECT 35.080 29.265 35.200 29.375 ;
        RECT 36.005 29.235 36.175 29.425 ;
        RECT 42.905 29.215 43.075 29.405 ;
        RECT 43.640 29.215 43.810 29.405 ;
        RECT 45.205 29.235 45.375 29.425 ;
        RECT 46.585 29.235 46.755 29.425 ;
        RECT 47.515 29.260 47.675 29.370 ;
        RECT 47.965 29.235 48.135 29.425 ;
        RECT 49.345 29.235 49.515 29.425 ;
        RECT 50.725 29.235 50.895 29.425 ;
        RECT 52.105 29.215 52.275 29.405 ;
        RECT 52.575 29.260 52.735 29.370 ;
        RECT 53.020 29.235 53.190 29.425 ;
        RECT 53.485 29.235 53.655 29.425 ;
        RECT 55.785 29.215 55.955 29.405 ;
        RECT 56.255 29.260 56.415 29.370 ;
        RECT 58.085 29.215 58.255 29.425 ;
        RECT 22.525 28.405 23.895 29.215 ;
        RECT 23.905 28.535 25.735 29.215 ;
        RECT 26.665 28.535 30.565 29.215 ;
        RECT 23.905 28.305 25.250 28.535 ;
        RECT 26.665 28.305 27.595 28.535 ;
        RECT 30.805 28.405 34.475 29.215 ;
        RECT 34.485 28.405 35.855 29.215 ;
        RECT 35.905 28.535 43.215 29.215 ;
        RECT 43.225 28.535 47.125 29.215 ;
        RECT 35.905 28.305 37.255 28.535 ;
        RECT 38.790 28.315 39.700 28.535 ;
        RECT 43.225 28.305 44.155 28.535 ;
        RECT 48.295 28.345 48.725 29.130 ;
        RECT 48.840 28.535 52.305 29.215 ;
        RECT 48.840 28.305 49.760 28.535 ;
        RECT 53.345 28.305 56.095 29.215 ;
        RECT 57.025 28.405 58.395 29.215 ;
      LAYER nwell ;
        RECT 22.330 25.185 58.590 28.015 ;
      LAYER pwell ;
        RECT 22.525 23.985 23.895 24.795 ;
        RECT 23.905 23.985 29.415 24.795 ;
        RECT 29.425 23.985 33.095 24.795 ;
        RECT 34.050 24.665 35.395 24.895 ;
        RECT 33.565 23.985 35.395 24.665 ;
        RECT 35.415 24.070 35.845 24.855 ;
        RECT 36.325 24.665 37.670 24.895 ;
        RECT 41.680 24.665 42.590 24.885 ;
        RECT 44.125 24.665 45.475 24.895 ;
        RECT 36.325 23.985 38.155 24.665 ;
        RECT 38.165 23.985 45.475 24.665 ;
        RECT 45.525 24.665 46.870 24.895 ;
        RECT 45.525 23.985 47.355 24.665 ;
        RECT 48.295 24.070 48.725 24.855 ;
        RECT 50.150 24.665 51.495 24.895 ;
        RECT 49.665 23.985 51.495 24.665 ;
        RECT 51.505 23.985 52.875 24.765 ;
        RECT 55.625 24.665 56.555 24.895 ;
        RECT 53.805 23.985 56.555 24.665 ;
        RECT 57.025 23.985 58.395 24.795 ;
        RECT 22.665 23.795 22.835 23.985 ;
        RECT 24.045 23.795 24.215 23.985 ;
        RECT 29.565 23.795 29.735 23.985 ;
        RECT 33.240 23.825 33.360 23.935 ;
        RECT 33.705 23.795 33.875 23.985 ;
        RECT 36.000 23.825 36.120 23.935 ;
        RECT 37.845 23.795 38.015 23.985 ;
        RECT 38.305 23.795 38.475 23.985 ;
        RECT 47.045 23.795 47.215 23.985 ;
        RECT 47.515 23.830 47.675 23.940 ;
        RECT 48.895 23.830 49.055 23.940 ;
        RECT 49.805 23.795 49.975 23.985 ;
        RECT 52.555 23.795 52.725 23.985 ;
        RECT 53.035 23.830 53.195 23.940 ;
        RECT 53.945 23.795 54.115 23.985 ;
        RECT 56.700 23.825 56.820 23.935 ;
        RECT 58.085 23.795 58.255 23.985 ;
        RECT 75.535 6.505 79.635 28.665 ;
      LAYER nwell ;
        RECT 80.015 25.205 89.975 29.325 ;
        RECT 80.015 17.895 90.205 25.205 ;
        RECT 80.010 17.815 90.205 17.895 ;
        RECT 80.010 9.480 88.510 17.815 ;
        RECT 80.010 6.590 86.200 9.480 ;
        RECT 80.010 6.505 86.215 6.590 ;
      LAYER pwell ;
        RECT 75.535 6.415 79.640 6.505 ;
        RECT 76.540 4.480 79.640 6.415 ;
      LAYER nwell ;
        RECT 80.025 4.565 86.215 6.505 ;
      LAYER pwell ;
        RECT 92.535 6.505 96.635 28.665 ;
      LAYER nwell ;
        RECT 97.015 25.205 106.975 29.325 ;
        RECT 97.015 17.895 107.205 25.205 ;
        RECT 97.010 17.815 107.205 17.895 ;
        RECT 97.010 9.480 105.510 17.815 ;
        RECT 97.010 6.590 103.200 9.480 ;
        RECT 97.010 6.505 103.215 6.590 ;
      LAYER pwell ;
        RECT 92.535 6.415 96.640 6.505 ;
      LAYER nwell ;
        RECT 80.025 4.480 90.220 4.565 ;
      LAYER pwell ;
        RECT 93.540 4.480 96.640 6.415 ;
      LAYER nwell ;
        RECT 97.025 4.565 103.215 6.505 ;
      LAYER pwell ;
        RECT 109.535 6.505 113.635 28.665 ;
      LAYER nwell ;
        RECT 114.015 25.205 123.975 29.325 ;
        RECT 114.015 17.895 124.205 25.205 ;
        RECT 114.010 17.815 124.205 17.895 ;
        RECT 114.010 9.480 122.510 17.815 ;
        RECT 114.010 6.590 120.200 9.480 ;
        RECT 114.010 6.505 120.215 6.590 ;
      LAYER pwell ;
        RECT 109.535 6.415 113.640 6.505 ;
      LAYER nwell ;
        RECT 97.025 4.480 107.220 4.565 ;
      LAYER pwell ;
        RECT 110.540 4.480 113.640 6.415 ;
      LAYER nwell ;
        RECT 114.025 4.565 120.215 6.505 ;
      LAYER pwell ;
        RECT 126.535 6.505 130.635 28.665 ;
      LAYER nwell ;
        RECT 131.015 25.205 140.975 29.325 ;
        RECT 131.015 17.895 141.205 25.205 ;
        RECT 131.010 17.815 141.205 17.895 ;
        RECT 131.010 9.480 139.510 17.815 ;
        RECT 131.010 6.590 137.200 9.480 ;
        RECT 131.010 6.505 137.215 6.590 ;
      LAYER pwell ;
        RECT 126.535 6.415 130.640 6.505 ;
      LAYER nwell ;
        RECT 114.025 4.480 124.220 4.565 ;
      LAYER pwell ;
        RECT 127.540 4.480 130.640 6.415 ;
      LAYER nwell ;
        RECT 131.025 4.565 137.215 6.505 ;
      LAYER pwell ;
        RECT 143.535 6.505 147.635 28.665 ;
      LAYER nwell ;
        RECT 148.015 25.205 157.975 29.325 ;
        RECT 148.015 17.895 158.205 25.205 ;
        RECT 148.010 17.815 158.205 17.895 ;
        RECT 148.010 9.480 156.510 17.815 ;
        RECT 148.010 6.590 154.200 9.480 ;
        RECT 148.010 6.505 154.215 6.590 ;
      LAYER pwell ;
        RECT 143.535 6.415 147.640 6.505 ;
      LAYER nwell ;
        RECT 131.025 4.480 141.220 4.565 ;
      LAYER pwell ;
        RECT 144.540 4.480 147.640 6.415 ;
      LAYER nwell ;
        RECT 148.025 4.565 154.215 6.505 ;
        RECT 148.025 4.480 158.220 4.565 ;
      LAYER pwell ;
        RECT 75.545 2.370 79.645 4.480 ;
      LAYER nwell ;
        RECT 80.030 2.455 90.220 4.480 ;
      LAYER pwell ;
        RECT 92.545 2.370 96.645 4.480 ;
      LAYER nwell ;
        RECT 97.030 2.455 107.220 4.480 ;
      LAYER pwell ;
        RECT 109.545 2.370 113.645 4.480 ;
      LAYER nwell ;
        RECT 114.030 2.455 124.220 4.480 ;
      LAYER pwell ;
        RECT 126.545 2.370 130.645 4.480 ;
      LAYER nwell ;
        RECT 131.030 2.455 141.220 4.480 ;
      LAYER pwell ;
        RECT 143.545 2.370 147.645 4.480 ;
      LAYER nwell ;
        RECT 148.030 2.455 158.220 4.480 ;
      LAYER li1 ;
        RECT 74.670 130.310 87.380 130.920 ;
        RECT 74.620 130.110 87.430 130.310 ;
        RECT 74.620 123.000 74.790 130.110 ;
        RECT 75.190 123.730 75.360 129.770 ;
        RECT 75.630 123.730 75.800 129.770 ;
        RECT 75.330 123.345 75.660 123.515 ;
        RECT 76.200 123.000 76.370 130.110 ;
        RECT 76.770 123.730 76.940 129.770 ;
        RECT 77.210 123.730 77.380 129.770 ;
        RECT 76.910 123.345 77.240 123.515 ;
        RECT 77.780 123.000 77.950 130.110 ;
        RECT 78.350 123.730 78.520 129.770 ;
        RECT 78.790 123.730 78.960 129.770 ;
        RECT 78.490 123.345 78.820 123.515 ;
        RECT 79.360 123.000 79.530 130.110 ;
        RECT 79.930 123.730 80.100 129.770 ;
        RECT 80.370 123.730 80.540 129.770 ;
        RECT 80.070 123.345 80.400 123.515 ;
        RECT 80.940 123.000 81.110 130.110 ;
        RECT 81.510 123.730 81.680 129.770 ;
        RECT 81.950 123.730 82.120 129.770 ;
        RECT 81.650 123.345 81.980 123.515 ;
        RECT 82.520 123.000 82.690 130.110 ;
        RECT 83.090 123.730 83.260 129.770 ;
        RECT 83.530 123.730 83.700 129.770 ;
        RECT 83.230 123.345 83.560 123.515 ;
        RECT 84.100 123.000 84.270 130.110 ;
        RECT 84.670 123.730 84.840 129.770 ;
        RECT 85.110 123.730 85.280 129.770 ;
        RECT 84.810 123.345 85.140 123.515 ;
        RECT 85.680 123.000 85.850 130.110 ;
        RECT 86.250 123.730 86.420 129.770 ;
        RECT 86.690 123.730 86.860 129.770 ;
        RECT 86.390 123.345 86.720 123.515 ;
        RECT 87.260 123.000 87.430 130.110 ;
        RECT 74.620 122.830 87.430 123.000 ;
        RECT 74.630 121.590 87.440 121.760 ;
        RECT 74.630 118.520 74.800 121.590 ;
        RECT 75.340 121.080 75.670 121.250 ;
        RECT 75.200 118.870 75.370 120.910 ;
        RECT 75.640 118.870 75.810 120.910 ;
        RECT 76.210 118.520 76.380 121.590 ;
        RECT 76.920 121.080 77.250 121.250 ;
        RECT 76.780 118.870 76.950 120.910 ;
        RECT 77.220 118.870 77.390 120.910 ;
        RECT 77.790 118.520 77.960 121.590 ;
        RECT 78.500 121.080 78.830 121.250 ;
        RECT 78.360 118.870 78.530 120.910 ;
        RECT 78.800 118.870 78.970 120.910 ;
        RECT 79.370 118.520 79.540 121.590 ;
        RECT 80.080 121.080 80.410 121.250 ;
        RECT 79.940 118.870 80.110 120.910 ;
        RECT 80.380 118.870 80.550 120.910 ;
        RECT 80.950 118.520 81.120 121.590 ;
        RECT 81.660 121.080 81.990 121.250 ;
        RECT 81.520 118.870 81.690 120.910 ;
        RECT 81.960 118.870 82.130 120.910 ;
        RECT 82.530 118.520 82.700 121.590 ;
        RECT 83.240 121.080 83.570 121.250 ;
        RECT 83.100 118.870 83.270 120.910 ;
        RECT 83.540 118.870 83.710 120.910 ;
        RECT 84.110 118.520 84.280 121.590 ;
        RECT 84.820 121.080 85.150 121.250 ;
        RECT 84.680 118.870 84.850 120.910 ;
        RECT 85.120 118.870 85.290 120.910 ;
        RECT 85.690 118.520 85.860 121.590 ;
        RECT 86.400 121.080 86.730 121.250 ;
        RECT 86.260 118.870 86.430 120.910 ;
        RECT 86.700 118.870 86.870 120.910 ;
        RECT 87.270 118.520 87.440 121.590 ;
        RECT 74.630 118.330 87.440 118.520 ;
        RECT 74.710 117.700 87.400 118.330 ;
        RECT 74.630 117.530 88.120 117.700 ;
        RECT 74.630 111.010 74.800 117.530 ;
        RECT 75.280 114.890 75.630 117.050 ;
        RECT 75.280 111.490 75.630 113.650 ;
        RECT 76.110 111.010 76.280 117.530 ;
        RECT 76.760 114.890 77.110 117.050 ;
        RECT 76.760 111.490 77.110 113.650 ;
        RECT 77.590 111.010 77.760 117.530 ;
        RECT 78.240 114.890 78.590 117.050 ;
        RECT 78.240 111.490 78.590 113.650 ;
        RECT 79.070 111.010 79.240 117.530 ;
        RECT 79.720 114.890 80.070 117.050 ;
        RECT 79.720 111.490 80.070 113.650 ;
        RECT 80.550 111.010 80.720 117.530 ;
        RECT 81.200 114.890 81.550 117.050 ;
        RECT 81.200 111.490 81.550 113.650 ;
        RECT 82.030 111.010 82.200 117.530 ;
        RECT 82.680 114.890 83.030 117.050 ;
        RECT 82.680 111.490 83.030 113.650 ;
        RECT 83.510 111.010 83.680 117.530 ;
        RECT 84.160 114.890 84.510 117.050 ;
        RECT 84.160 111.490 84.510 113.650 ;
        RECT 84.990 111.010 85.160 117.530 ;
        RECT 85.640 114.890 85.990 117.050 ;
        RECT 85.640 111.490 85.990 113.650 ;
        RECT 86.470 111.010 86.640 117.530 ;
        RECT 87.120 114.890 87.470 117.050 ;
        RECT 87.120 111.490 87.470 113.650 ;
        RECT 87.950 111.010 88.120 117.530 ;
        RECT 121.335 116.975 123.280 117.010 ;
        RECT 121.210 116.435 129.735 116.975 ;
        RECT 74.630 110.840 88.120 111.010 ;
        RECT 121.215 116.400 129.735 116.435 ;
        RECT 74.630 105.020 74.800 110.840 ;
        RECT 75.280 108.200 75.630 110.360 ;
        RECT 75.280 105.500 75.630 107.660 ;
        RECT 76.110 105.020 76.280 110.840 ;
        RECT 76.760 108.200 77.110 110.360 ;
        RECT 76.760 105.500 77.110 107.660 ;
        RECT 77.590 105.020 77.760 110.840 ;
        RECT 78.240 108.200 78.590 110.360 ;
        RECT 78.240 105.500 78.590 107.660 ;
        RECT 79.070 105.020 79.240 110.840 ;
        RECT 79.720 108.200 80.070 110.360 ;
        RECT 79.720 105.500 80.070 107.660 ;
        RECT 80.550 105.020 80.720 110.840 ;
        RECT 81.200 108.200 81.550 110.360 ;
        RECT 81.200 105.500 81.550 107.660 ;
        RECT 82.030 105.020 82.200 110.840 ;
        RECT 82.680 108.200 83.030 110.360 ;
        RECT 82.680 105.500 83.030 107.660 ;
        RECT 83.510 105.020 83.680 110.840 ;
        RECT 84.160 108.200 84.510 110.360 ;
        RECT 84.160 105.500 84.510 107.660 ;
        RECT 84.990 105.020 85.160 110.840 ;
        RECT 121.215 110.435 123.415 116.400 ;
        RECT 123.955 115.890 124.285 116.060 ;
        RECT 74.630 104.850 85.160 105.020 ;
        RECT 121.225 110.405 122.975 110.435 ;
        RECT 121.225 104.915 121.395 110.405 ;
        RECT 121.935 109.895 122.265 110.065 ;
        RECT 121.795 105.640 121.965 109.680 ;
        RECT 122.235 105.640 122.405 109.680 ;
        RECT 121.935 105.255 122.265 105.425 ;
        RECT 122.805 104.915 122.975 110.405 ;
        RECT 121.225 104.745 122.975 104.915 ;
        RECT 123.245 104.910 123.415 110.435 ;
        RECT 123.815 105.635 123.985 115.675 ;
        RECT 124.255 105.635 124.425 115.675 ;
        RECT 123.955 105.250 124.285 105.420 ;
        RECT 124.825 104.910 124.995 116.400 ;
        RECT 125.535 115.890 125.865 116.060 ;
        RECT 125.395 105.635 125.565 115.675 ;
        RECT 125.835 105.635 126.005 115.675 ;
        RECT 125.535 105.250 125.865 105.420 ;
        RECT 126.405 104.910 126.575 116.400 ;
        RECT 127.115 115.890 127.445 116.060 ;
        RECT 126.975 105.635 127.145 115.675 ;
        RECT 127.415 105.635 127.585 115.675 ;
        RECT 127.115 105.250 127.445 105.420 ;
        RECT 127.985 104.910 128.155 116.400 ;
        RECT 128.695 115.890 129.025 116.060 ;
        RECT 128.555 105.635 128.725 115.675 ;
        RECT 128.995 105.635 129.165 115.675 ;
        RECT 128.695 105.250 129.025 105.420 ;
        RECT 129.565 104.910 129.735 116.400 ;
        RECT 123.245 104.740 129.735 104.910 ;
        RECT 122.030 104.305 124.595 104.490 ;
        RECT 121.220 103.915 122.970 104.085 ;
        RECT 121.220 101.515 121.390 103.915 ;
        RECT 121.930 103.405 122.260 103.575 ;
        RECT 121.790 102.195 121.960 103.235 ;
        RECT 122.230 102.195 122.400 103.235 ;
        RECT 121.930 101.855 122.260 102.025 ;
        RECT 122.800 101.515 122.970 103.915 ;
        RECT 121.220 101.485 122.970 101.515 ;
        RECT 123.245 103.910 129.735 104.080 ;
        RECT 123.245 101.485 123.415 103.910 ;
        RECT 123.955 103.400 124.285 103.570 ;
        RECT 121.220 97.510 123.415 101.485 ;
        RECT 123.815 98.190 123.985 103.230 ;
        RECT 124.255 98.190 124.425 103.230 ;
        RECT 123.955 97.850 124.285 98.020 ;
        RECT 124.825 97.510 124.995 103.910 ;
        RECT 125.535 103.400 125.865 103.570 ;
        RECT 125.395 98.190 125.565 103.230 ;
        RECT 125.835 98.190 126.005 103.230 ;
        RECT 125.535 97.850 125.865 98.020 ;
        RECT 126.405 97.510 126.575 103.910 ;
        RECT 127.115 103.400 127.445 103.570 ;
        RECT 126.975 98.190 127.145 103.230 ;
        RECT 127.415 98.190 127.585 103.230 ;
        RECT 127.115 97.850 127.445 98.020 ;
        RECT 127.985 97.510 128.155 103.910 ;
        RECT 128.695 103.400 129.025 103.570 ;
        RECT 128.555 98.190 128.725 103.230 ;
        RECT 128.995 98.190 129.165 103.230 ;
        RECT 128.695 97.850 129.025 98.020 ;
        RECT 129.565 97.510 129.735 103.910 ;
        RECT 121.220 97.455 129.735 97.510 ;
        RECT 149.780 100.160 158.830 100.330 ;
        RECT 121.220 97.335 129.750 97.455 ;
        RECT 121.230 97.000 129.750 97.335 ;
        RECT 149.780 94.340 149.950 100.160 ;
        RECT 150.430 97.520 150.780 99.680 ;
        RECT 150.430 94.820 150.780 96.980 ;
        RECT 151.260 94.340 151.430 100.160 ;
        RECT 151.910 97.520 152.260 99.680 ;
        RECT 151.910 94.820 152.260 96.980 ;
        RECT 152.740 94.340 152.910 100.160 ;
        RECT 153.390 97.520 153.740 99.680 ;
        RECT 153.390 94.820 153.740 96.980 ;
        RECT 154.220 94.340 154.390 100.160 ;
        RECT 154.870 97.520 155.220 99.680 ;
        RECT 154.870 94.820 155.220 96.980 ;
        RECT 155.700 94.340 155.870 100.160 ;
        RECT 156.350 97.520 156.700 99.680 ;
        RECT 156.350 94.820 156.700 96.980 ;
        RECT 157.180 94.340 157.350 100.160 ;
        RECT 157.830 97.520 158.180 99.680 ;
        RECT 157.830 94.820 158.180 96.980 ;
        RECT 158.660 94.340 158.830 100.160 ;
        RECT 126.100 94.170 158.830 94.340 ;
        RECT 126.100 88.350 126.270 94.170 ;
        RECT 126.750 91.530 127.100 93.690 ;
        RECT 126.750 88.830 127.100 90.990 ;
        RECT 127.580 88.350 127.750 94.170 ;
        RECT 128.230 91.530 128.580 93.690 ;
        RECT 128.230 88.830 128.580 90.990 ;
        RECT 129.060 88.350 129.230 94.170 ;
        RECT 129.710 91.530 130.060 93.690 ;
        RECT 129.710 88.830 130.060 90.990 ;
        RECT 130.540 88.350 130.710 94.170 ;
        RECT 131.190 91.530 131.540 93.690 ;
        RECT 131.190 88.830 131.540 90.990 ;
        RECT 132.020 88.350 132.190 94.170 ;
        RECT 132.670 91.530 133.020 93.690 ;
        RECT 132.670 88.830 133.020 90.990 ;
        RECT 133.500 88.350 133.670 94.170 ;
        RECT 134.150 91.530 134.500 93.690 ;
        RECT 134.150 88.830 134.500 90.990 ;
        RECT 134.980 88.350 135.150 94.170 ;
        RECT 135.630 91.530 135.980 93.690 ;
        RECT 135.630 88.830 135.980 90.990 ;
        RECT 136.460 88.350 136.630 94.170 ;
        RECT 137.110 91.530 137.460 93.690 ;
        RECT 137.110 88.830 137.460 90.990 ;
        RECT 137.940 88.350 138.110 94.170 ;
        RECT 138.590 91.530 138.940 93.690 ;
        RECT 138.590 88.830 138.940 90.990 ;
        RECT 139.420 88.350 139.590 94.170 ;
        RECT 140.070 91.530 140.420 93.690 ;
        RECT 140.070 88.830 140.420 90.990 ;
        RECT 140.900 88.350 141.070 94.170 ;
        RECT 141.550 91.530 141.900 93.690 ;
        RECT 141.550 88.830 141.900 90.990 ;
        RECT 142.380 88.350 142.550 94.170 ;
        RECT 143.030 91.530 143.380 93.690 ;
        RECT 143.030 88.830 143.380 90.990 ;
        RECT 143.860 88.350 144.030 94.170 ;
        RECT 144.510 91.530 144.860 93.690 ;
        RECT 144.510 88.830 144.860 90.990 ;
        RECT 145.340 88.350 145.510 94.170 ;
        RECT 145.990 91.530 146.340 93.690 ;
        RECT 145.990 88.830 146.340 90.990 ;
        RECT 146.820 88.350 146.990 94.170 ;
        RECT 147.470 91.530 147.820 93.690 ;
        RECT 147.470 88.830 147.820 90.990 ;
        RECT 148.300 88.350 148.470 94.170 ;
        RECT 148.950 91.530 149.300 93.690 ;
        RECT 148.950 88.830 149.300 90.990 ;
        RECT 149.780 88.350 149.950 94.170 ;
        RECT 150.430 91.530 150.780 93.690 ;
        RECT 150.430 88.830 150.780 90.990 ;
        RECT 151.260 88.350 151.430 94.170 ;
        RECT 151.910 91.530 152.260 93.690 ;
        RECT 151.910 88.830 152.260 90.990 ;
        RECT 152.740 88.350 152.910 94.170 ;
        RECT 153.390 91.530 153.740 93.690 ;
        RECT 153.390 88.830 153.740 90.990 ;
        RECT 154.220 88.350 154.390 94.170 ;
        RECT 154.870 91.530 155.220 93.690 ;
        RECT 154.870 88.830 155.220 90.990 ;
        RECT 155.700 88.350 155.870 94.170 ;
        RECT 156.350 91.530 156.700 93.690 ;
        RECT 156.350 88.830 156.700 90.990 ;
        RECT 157.180 88.350 157.350 94.170 ;
        RECT 157.830 91.530 158.180 93.690 ;
        RECT 157.830 88.830 158.180 90.990 ;
        RECT 158.660 88.350 158.830 94.170 ;
        RECT 126.100 88.260 158.830 88.350 ;
        RECT 126.050 88.180 158.830 88.260 ;
        RECT 89.625 87.165 90.100 87.180 ;
        RECT 106.625 87.165 107.100 87.180 ;
        RECT 123.625 87.165 124.100 87.180 ;
        RECT 89.625 87.145 90.580 87.165 ;
        RECT 106.625 87.145 107.580 87.165 ;
        RECT 123.625 87.145 124.580 87.165 ;
        RECT 75.000 86.485 75.865 87.140 ;
        RECT 80.195 86.975 90.580 87.145 ;
        RECT 75.000 86.315 79.455 86.485 ;
        RECT 75.000 81.055 75.885 86.315 ;
        RECT 76.565 85.745 78.605 85.915 ;
        RECT 76.225 81.685 76.395 85.685 ;
        RECT 78.775 81.685 78.945 85.685 ;
        RECT 76.565 81.455 78.605 81.625 ;
        RECT 79.285 81.055 79.455 86.315 ;
        RECT 80.195 83.485 80.365 86.975 ;
        RECT 80.995 86.465 88.995 86.635 ;
        RECT 80.765 84.210 80.935 86.250 ;
        RECT 89.055 84.210 89.225 86.250 ;
        RECT 80.995 83.825 88.995 83.995 ;
        RECT 89.625 83.485 90.580 86.975 ;
        RECT 80.195 83.315 90.580 83.485 ;
        RECT 89.625 83.025 90.580 83.315 ;
        RECT 75.000 80.885 79.455 81.055 ;
        RECT 75.000 75.625 75.885 80.885 ;
        RECT 76.565 80.315 78.605 80.485 ;
        RECT 76.225 76.255 76.395 80.255 ;
        RECT 78.775 76.255 78.945 80.255 ;
        RECT 76.565 76.025 78.605 76.195 ;
        RECT 79.285 75.625 79.455 80.885 ;
        RECT 80.195 82.855 90.580 83.025 ;
        RECT 80.195 79.595 80.365 82.855 ;
        RECT 81.090 82.285 89.130 82.455 ;
        RECT 80.705 80.225 80.875 82.225 ;
        RECT 89.345 80.225 89.515 82.225 ;
        RECT 81.090 79.995 89.130 80.165 ;
        RECT 89.855 79.595 90.580 82.855 ;
        RECT 80.195 79.425 90.580 79.595 ;
        RECT 80.195 76.165 80.365 79.425 ;
        RECT 81.090 78.855 89.130 79.025 ;
        RECT 80.705 76.795 80.875 78.795 ;
        RECT 89.345 76.795 89.515 78.795 ;
        RECT 81.090 76.565 89.130 76.735 ;
        RECT 89.855 76.165 90.580 79.425 ;
        RECT 80.195 75.995 90.580 76.165 ;
        RECT 85.905 75.715 90.580 75.995 ;
        RECT 75.000 75.455 79.455 75.625 ;
        RECT 75.000 70.195 75.885 75.455 ;
        RECT 76.565 74.885 78.605 75.055 ;
        RECT 76.225 70.825 76.395 74.825 ;
        RECT 78.775 70.825 78.945 74.825 ;
        RECT 76.565 70.595 78.605 70.765 ;
        RECT 79.285 70.195 79.455 75.455 ;
        RECT 75.000 70.025 79.455 70.195 ;
        RECT 75.000 64.765 75.885 70.025 ;
        RECT 76.565 69.455 78.605 69.625 ;
        RECT 76.225 65.395 76.395 69.395 ;
        RECT 78.775 65.395 78.945 69.395 ;
        RECT 76.565 65.165 78.605 65.335 ;
        RECT 79.285 64.765 79.455 70.025 ;
        RECT 75.000 64.595 79.455 64.765 ;
        RECT 80.190 75.545 90.580 75.715 ;
        RECT 80.190 70.285 80.360 75.545 ;
        RECT 81.085 74.975 85.125 75.145 ;
        RECT 80.700 70.915 80.870 74.915 ;
        RECT 85.340 70.915 85.510 74.915 ;
        RECT 85.850 74.435 90.580 75.545 ;
        RECT 81.085 70.685 85.125 70.855 ;
        RECT 85.850 70.285 86.020 74.435 ;
        RECT 80.190 70.115 86.020 70.285 ;
        RECT 80.190 64.855 80.360 70.115 ;
        RECT 81.085 69.545 85.125 69.715 ;
        RECT 80.700 65.485 80.870 69.485 ;
        RECT 85.340 65.485 85.510 69.485 ;
        RECT 81.085 65.255 85.125 65.425 ;
        RECT 85.850 64.855 86.020 70.115 ;
        RECT 86.535 74.360 88.285 74.435 ;
        RECT 86.535 67.870 86.705 74.360 ;
        RECT 87.245 73.850 87.575 74.020 ;
        RECT 87.105 68.595 87.275 73.635 ;
        RECT 87.545 68.595 87.715 73.635 ;
        RECT 87.245 68.210 87.575 68.380 ;
        RECT 88.115 67.870 88.285 74.360 ;
        RECT 86.535 67.700 88.285 67.870 ;
        RECT 80.190 64.685 86.020 64.855 ;
        RECT 75.000 64.325 76.860 64.595 ;
        RECT 75.000 64.155 79.460 64.325 ;
        RECT 75.000 62.745 76.890 64.155 ;
        RECT 77.230 63.285 77.400 63.615 ;
        RECT 77.570 63.585 78.610 63.755 ;
        RECT 77.570 63.145 78.610 63.315 ;
        RECT 78.780 63.285 78.950 63.615 ;
        RECT 79.290 62.745 79.460 64.155 ;
        RECT 75.000 62.575 79.460 62.745 ;
        RECT 80.205 64.240 86.035 64.410 ;
        RECT 80.205 62.830 80.375 64.240 ;
        RECT 80.715 63.370 80.885 63.700 ;
        RECT 81.100 63.670 85.140 63.840 ;
        RECT 81.100 63.230 85.140 63.400 ;
        RECT 85.355 63.370 85.525 63.700 ;
        RECT 85.865 62.830 86.035 64.240 ;
        RECT 80.205 62.660 86.035 62.830 ;
        RECT 75.000 62.300 76.860 62.575 ;
        RECT 89.880 62.385 90.580 74.435 ;
        RECT 75.000 62.130 79.465 62.300 ;
        RECT 75.000 60.720 75.895 62.130 ;
        RECT 76.235 61.260 76.405 61.590 ;
        RECT 76.575 61.560 78.615 61.730 ;
        RECT 76.575 61.120 78.615 61.290 ;
        RECT 78.785 61.260 78.955 61.590 ;
        RECT 79.295 60.720 79.465 62.130 ;
        RECT 75.000 60.560 79.465 60.720 ;
        RECT 80.210 62.215 90.580 62.385 ;
        RECT 80.210 60.805 80.380 62.215 ;
        RECT 80.720 61.345 80.890 61.675 ;
        RECT 81.105 61.645 89.145 61.815 ;
        RECT 81.105 61.205 89.145 61.375 ;
        RECT 89.360 61.345 89.530 61.675 ;
        RECT 89.870 60.805 90.580 62.215 ;
        RECT 80.210 60.690 90.580 60.805 ;
        RECT 92.000 86.485 92.865 87.140 ;
        RECT 97.195 86.975 107.580 87.145 ;
        RECT 92.000 86.315 96.455 86.485 ;
        RECT 92.000 81.055 92.885 86.315 ;
        RECT 93.565 85.745 95.605 85.915 ;
        RECT 93.225 81.685 93.395 85.685 ;
        RECT 95.775 81.685 95.945 85.685 ;
        RECT 93.565 81.455 95.605 81.625 ;
        RECT 96.285 81.055 96.455 86.315 ;
        RECT 97.195 83.485 97.365 86.975 ;
        RECT 97.995 86.465 105.995 86.635 ;
        RECT 97.765 84.210 97.935 86.250 ;
        RECT 106.055 84.210 106.225 86.250 ;
        RECT 97.995 83.825 105.995 83.995 ;
        RECT 106.625 83.485 107.580 86.975 ;
        RECT 97.195 83.315 107.580 83.485 ;
        RECT 106.625 83.025 107.580 83.315 ;
        RECT 92.000 80.885 96.455 81.055 ;
        RECT 92.000 75.625 92.885 80.885 ;
        RECT 93.565 80.315 95.605 80.485 ;
        RECT 93.225 76.255 93.395 80.255 ;
        RECT 95.775 76.255 95.945 80.255 ;
        RECT 93.565 76.025 95.605 76.195 ;
        RECT 96.285 75.625 96.455 80.885 ;
        RECT 97.195 82.855 107.580 83.025 ;
        RECT 97.195 79.595 97.365 82.855 ;
        RECT 98.090 82.285 106.130 82.455 ;
        RECT 97.705 80.225 97.875 82.225 ;
        RECT 106.345 80.225 106.515 82.225 ;
        RECT 98.090 79.995 106.130 80.165 ;
        RECT 106.855 79.595 107.580 82.855 ;
        RECT 97.195 79.425 107.580 79.595 ;
        RECT 97.195 76.165 97.365 79.425 ;
        RECT 98.090 78.855 106.130 79.025 ;
        RECT 97.705 76.795 97.875 78.795 ;
        RECT 106.345 76.795 106.515 78.795 ;
        RECT 98.090 76.565 106.130 76.735 ;
        RECT 106.855 76.165 107.580 79.425 ;
        RECT 97.195 75.995 107.580 76.165 ;
        RECT 102.905 75.715 107.580 75.995 ;
        RECT 92.000 75.455 96.455 75.625 ;
        RECT 92.000 70.195 92.885 75.455 ;
        RECT 93.565 74.885 95.605 75.055 ;
        RECT 93.225 70.825 93.395 74.825 ;
        RECT 95.775 70.825 95.945 74.825 ;
        RECT 93.565 70.595 95.605 70.765 ;
        RECT 96.285 70.195 96.455 75.455 ;
        RECT 92.000 70.025 96.455 70.195 ;
        RECT 92.000 64.765 92.885 70.025 ;
        RECT 93.565 69.455 95.605 69.625 ;
        RECT 93.225 65.395 93.395 69.395 ;
        RECT 95.775 65.395 95.945 69.395 ;
        RECT 93.565 65.165 95.605 65.335 ;
        RECT 96.285 64.765 96.455 70.025 ;
        RECT 92.000 64.595 96.455 64.765 ;
        RECT 97.190 75.545 107.580 75.715 ;
        RECT 97.190 70.285 97.360 75.545 ;
        RECT 98.085 74.975 102.125 75.145 ;
        RECT 97.700 70.915 97.870 74.915 ;
        RECT 102.340 70.915 102.510 74.915 ;
        RECT 102.850 74.435 107.580 75.545 ;
        RECT 98.085 70.685 102.125 70.855 ;
        RECT 102.850 70.285 103.020 74.435 ;
        RECT 97.190 70.115 103.020 70.285 ;
        RECT 97.190 64.855 97.360 70.115 ;
        RECT 98.085 69.545 102.125 69.715 ;
        RECT 97.700 65.485 97.870 69.485 ;
        RECT 102.340 65.485 102.510 69.485 ;
        RECT 98.085 65.255 102.125 65.425 ;
        RECT 102.850 64.855 103.020 70.115 ;
        RECT 103.535 74.360 105.285 74.435 ;
        RECT 103.535 67.870 103.705 74.360 ;
        RECT 104.245 73.850 104.575 74.020 ;
        RECT 104.105 68.595 104.275 73.635 ;
        RECT 104.545 68.595 104.715 73.635 ;
        RECT 104.245 68.210 104.575 68.380 ;
        RECT 105.115 67.870 105.285 74.360 ;
        RECT 103.535 67.700 105.285 67.870 ;
        RECT 97.190 64.685 103.020 64.855 ;
        RECT 92.000 64.325 93.860 64.595 ;
        RECT 92.000 64.155 96.460 64.325 ;
        RECT 92.000 62.745 93.890 64.155 ;
        RECT 94.230 63.285 94.400 63.615 ;
        RECT 94.570 63.585 95.610 63.755 ;
        RECT 94.570 63.145 95.610 63.315 ;
        RECT 95.780 63.285 95.950 63.615 ;
        RECT 96.290 62.745 96.460 64.155 ;
        RECT 92.000 62.575 96.460 62.745 ;
        RECT 97.205 64.240 103.035 64.410 ;
        RECT 97.205 62.830 97.375 64.240 ;
        RECT 97.715 63.370 97.885 63.700 ;
        RECT 98.100 63.670 102.140 63.840 ;
        RECT 98.100 63.230 102.140 63.400 ;
        RECT 102.355 63.370 102.525 63.700 ;
        RECT 102.865 62.830 103.035 64.240 ;
        RECT 97.205 62.660 103.035 62.830 ;
        RECT 92.000 62.300 93.860 62.575 ;
        RECT 106.880 62.385 107.580 74.435 ;
        RECT 92.000 62.130 96.465 62.300 ;
        RECT 92.000 60.720 92.895 62.130 ;
        RECT 93.235 61.260 93.405 61.590 ;
        RECT 93.575 61.560 95.615 61.730 ;
        RECT 93.575 61.120 95.615 61.290 ;
        RECT 95.785 61.260 95.955 61.590 ;
        RECT 96.295 60.720 96.465 62.130 ;
        RECT 80.210 60.635 90.040 60.690 ;
        RECT 92.000 60.560 96.465 60.720 ;
        RECT 97.210 62.215 107.580 62.385 ;
        RECT 97.210 60.805 97.380 62.215 ;
        RECT 97.720 61.345 97.890 61.675 ;
        RECT 98.105 61.645 106.145 61.815 ;
        RECT 98.105 61.205 106.145 61.375 ;
        RECT 106.360 61.345 106.530 61.675 ;
        RECT 106.870 60.805 107.580 62.215 ;
        RECT 97.210 60.690 107.580 60.805 ;
        RECT 109.000 86.485 109.865 87.140 ;
        RECT 114.195 86.975 124.580 87.145 ;
        RECT 126.050 87.140 126.945 88.180 ;
        RECT 140.625 87.165 141.100 87.180 ;
        RECT 157.625 87.165 158.100 87.180 ;
        RECT 140.625 87.145 141.580 87.165 ;
        RECT 157.625 87.145 158.580 87.165 ;
        RECT 109.000 86.315 113.455 86.485 ;
        RECT 109.000 81.055 109.885 86.315 ;
        RECT 110.565 85.745 112.605 85.915 ;
        RECT 110.225 81.685 110.395 85.685 ;
        RECT 112.775 81.685 112.945 85.685 ;
        RECT 110.565 81.455 112.605 81.625 ;
        RECT 113.285 81.055 113.455 86.315 ;
        RECT 114.195 83.485 114.365 86.975 ;
        RECT 114.995 86.465 122.995 86.635 ;
        RECT 114.765 84.210 114.935 86.250 ;
        RECT 123.055 84.210 123.225 86.250 ;
        RECT 114.995 83.825 122.995 83.995 ;
        RECT 123.625 83.485 124.580 86.975 ;
        RECT 114.195 83.315 124.580 83.485 ;
        RECT 123.625 83.025 124.580 83.315 ;
        RECT 109.000 80.885 113.455 81.055 ;
        RECT 109.000 75.625 109.885 80.885 ;
        RECT 110.565 80.315 112.605 80.485 ;
        RECT 110.225 76.255 110.395 80.255 ;
        RECT 112.775 76.255 112.945 80.255 ;
        RECT 110.565 76.025 112.605 76.195 ;
        RECT 113.285 75.625 113.455 80.885 ;
        RECT 114.195 82.855 124.580 83.025 ;
        RECT 114.195 79.595 114.365 82.855 ;
        RECT 115.090 82.285 123.130 82.455 ;
        RECT 114.705 80.225 114.875 82.225 ;
        RECT 123.345 80.225 123.515 82.225 ;
        RECT 115.090 79.995 123.130 80.165 ;
        RECT 123.855 79.595 124.580 82.855 ;
        RECT 114.195 79.425 124.580 79.595 ;
        RECT 114.195 76.165 114.365 79.425 ;
        RECT 115.090 78.855 123.130 79.025 ;
        RECT 114.705 76.795 114.875 78.795 ;
        RECT 123.345 76.795 123.515 78.795 ;
        RECT 115.090 76.565 123.130 76.735 ;
        RECT 123.855 76.165 124.580 79.425 ;
        RECT 114.195 75.995 124.580 76.165 ;
        RECT 119.905 75.715 124.580 75.995 ;
        RECT 109.000 75.455 113.455 75.625 ;
        RECT 109.000 70.195 109.885 75.455 ;
        RECT 110.565 74.885 112.605 75.055 ;
        RECT 110.225 70.825 110.395 74.825 ;
        RECT 112.775 70.825 112.945 74.825 ;
        RECT 110.565 70.595 112.605 70.765 ;
        RECT 113.285 70.195 113.455 75.455 ;
        RECT 109.000 70.025 113.455 70.195 ;
        RECT 109.000 64.765 109.885 70.025 ;
        RECT 110.565 69.455 112.605 69.625 ;
        RECT 110.225 65.395 110.395 69.395 ;
        RECT 112.775 65.395 112.945 69.395 ;
        RECT 110.565 65.165 112.605 65.335 ;
        RECT 113.285 64.765 113.455 70.025 ;
        RECT 109.000 64.595 113.455 64.765 ;
        RECT 114.190 75.545 124.580 75.715 ;
        RECT 114.190 70.285 114.360 75.545 ;
        RECT 115.085 74.975 119.125 75.145 ;
        RECT 114.700 70.915 114.870 74.915 ;
        RECT 119.340 70.915 119.510 74.915 ;
        RECT 119.850 74.435 124.580 75.545 ;
        RECT 115.085 70.685 119.125 70.855 ;
        RECT 119.850 70.285 120.020 74.435 ;
        RECT 114.190 70.115 120.020 70.285 ;
        RECT 114.190 64.855 114.360 70.115 ;
        RECT 115.085 69.545 119.125 69.715 ;
        RECT 114.700 65.485 114.870 69.485 ;
        RECT 119.340 65.485 119.510 69.485 ;
        RECT 115.085 65.255 119.125 65.425 ;
        RECT 119.850 64.855 120.020 70.115 ;
        RECT 120.535 74.360 122.285 74.435 ;
        RECT 120.535 67.870 120.705 74.360 ;
        RECT 121.245 73.850 121.575 74.020 ;
        RECT 121.105 68.595 121.275 73.635 ;
        RECT 121.545 68.595 121.715 73.635 ;
        RECT 121.245 68.210 121.575 68.380 ;
        RECT 122.115 67.870 122.285 74.360 ;
        RECT 120.535 67.700 122.285 67.870 ;
        RECT 114.190 64.685 120.020 64.855 ;
        RECT 109.000 64.325 110.860 64.595 ;
        RECT 109.000 64.155 113.460 64.325 ;
        RECT 109.000 62.745 110.890 64.155 ;
        RECT 111.230 63.285 111.400 63.615 ;
        RECT 111.570 63.585 112.610 63.755 ;
        RECT 111.570 63.145 112.610 63.315 ;
        RECT 112.780 63.285 112.950 63.615 ;
        RECT 113.290 62.745 113.460 64.155 ;
        RECT 109.000 62.575 113.460 62.745 ;
        RECT 114.205 64.240 120.035 64.410 ;
        RECT 114.205 62.830 114.375 64.240 ;
        RECT 114.715 63.370 114.885 63.700 ;
        RECT 115.100 63.670 119.140 63.840 ;
        RECT 115.100 63.230 119.140 63.400 ;
        RECT 119.355 63.370 119.525 63.700 ;
        RECT 119.865 62.830 120.035 64.240 ;
        RECT 114.205 62.660 120.035 62.830 ;
        RECT 109.000 62.300 110.860 62.575 ;
        RECT 123.880 62.385 124.580 74.435 ;
        RECT 109.000 62.130 113.465 62.300 ;
        RECT 109.000 60.720 109.895 62.130 ;
        RECT 110.235 61.260 110.405 61.590 ;
        RECT 110.575 61.560 112.615 61.730 ;
        RECT 110.575 61.120 112.615 61.290 ;
        RECT 112.785 61.260 112.955 61.590 ;
        RECT 113.295 60.720 113.465 62.130 ;
        RECT 97.210 60.635 107.040 60.690 ;
        RECT 109.000 60.560 113.465 60.720 ;
        RECT 114.210 62.215 124.580 62.385 ;
        RECT 114.210 60.805 114.380 62.215 ;
        RECT 114.720 61.345 114.890 61.675 ;
        RECT 115.105 61.645 123.145 61.815 ;
        RECT 115.105 61.205 123.145 61.375 ;
        RECT 123.360 61.345 123.530 61.675 ;
        RECT 123.870 60.805 124.580 62.215 ;
        RECT 114.210 60.690 124.580 60.805 ;
        RECT 126.000 86.485 126.945 87.140 ;
        RECT 131.195 86.975 141.580 87.145 ;
        RECT 126.000 86.315 130.455 86.485 ;
        RECT 126.000 81.055 126.885 86.315 ;
        RECT 127.565 85.745 129.605 85.915 ;
        RECT 127.225 81.685 127.395 85.685 ;
        RECT 129.775 81.685 129.945 85.685 ;
        RECT 127.565 81.455 129.605 81.625 ;
        RECT 130.285 81.055 130.455 86.315 ;
        RECT 131.195 83.485 131.365 86.975 ;
        RECT 131.995 86.465 139.995 86.635 ;
        RECT 131.765 84.210 131.935 86.250 ;
        RECT 140.055 84.210 140.225 86.250 ;
        RECT 131.995 83.825 139.995 83.995 ;
        RECT 140.625 83.485 141.580 86.975 ;
        RECT 131.195 83.315 141.580 83.485 ;
        RECT 140.625 83.025 141.580 83.315 ;
        RECT 126.000 80.885 130.455 81.055 ;
        RECT 126.000 75.625 126.885 80.885 ;
        RECT 127.565 80.315 129.605 80.485 ;
        RECT 127.225 76.255 127.395 80.255 ;
        RECT 129.775 76.255 129.945 80.255 ;
        RECT 127.565 76.025 129.605 76.195 ;
        RECT 130.285 75.625 130.455 80.885 ;
        RECT 131.195 82.855 141.580 83.025 ;
        RECT 131.195 79.595 131.365 82.855 ;
        RECT 132.090 82.285 140.130 82.455 ;
        RECT 131.705 80.225 131.875 82.225 ;
        RECT 140.345 80.225 140.515 82.225 ;
        RECT 132.090 79.995 140.130 80.165 ;
        RECT 140.855 79.595 141.580 82.855 ;
        RECT 131.195 79.425 141.580 79.595 ;
        RECT 131.195 76.165 131.365 79.425 ;
        RECT 132.090 78.855 140.130 79.025 ;
        RECT 131.705 76.795 131.875 78.795 ;
        RECT 140.345 76.795 140.515 78.795 ;
        RECT 132.090 76.565 140.130 76.735 ;
        RECT 140.855 76.165 141.580 79.425 ;
        RECT 131.195 75.995 141.580 76.165 ;
        RECT 136.905 75.715 141.580 75.995 ;
        RECT 126.000 75.455 130.455 75.625 ;
        RECT 126.000 70.195 126.885 75.455 ;
        RECT 127.565 74.885 129.605 75.055 ;
        RECT 127.225 70.825 127.395 74.825 ;
        RECT 129.775 70.825 129.945 74.825 ;
        RECT 127.565 70.595 129.605 70.765 ;
        RECT 130.285 70.195 130.455 75.455 ;
        RECT 126.000 70.025 130.455 70.195 ;
        RECT 126.000 64.765 126.885 70.025 ;
        RECT 127.565 69.455 129.605 69.625 ;
        RECT 127.225 65.395 127.395 69.395 ;
        RECT 129.775 65.395 129.945 69.395 ;
        RECT 127.565 65.165 129.605 65.335 ;
        RECT 130.285 64.765 130.455 70.025 ;
        RECT 126.000 64.595 130.455 64.765 ;
        RECT 131.190 75.545 141.580 75.715 ;
        RECT 131.190 70.285 131.360 75.545 ;
        RECT 132.085 74.975 136.125 75.145 ;
        RECT 131.700 70.915 131.870 74.915 ;
        RECT 136.340 70.915 136.510 74.915 ;
        RECT 136.850 74.435 141.580 75.545 ;
        RECT 132.085 70.685 136.125 70.855 ;
        RECT 136.850 70.285 137.020 74.435 ;
        RECT 131.190 70.115 137.020 70.285 ;
        RECT 131.190 64.855 131.360 70.115 ;
        RECT 132.085 69.545 136.125 69.715 ;
        RECT 131.700 65.485 131.870 69.485 ;
        RECT 136.340 65.485 136.510 69.485 ;
        RECT 132.085 65.255 136.125 65.425 ;
        RECT 136.850 64.855 137.020 70.115 ;
        RECT 137.535 74.360 139.285 74.435 ;
        RECT 137.535 67.870 137.705 74.360 ;
        RECT 138.245 73.850 138.575 74.020 ;
        RECT 138.105 68.595 138.275 73.635 ;
        RECT 138.545 68.595 138.715 73.635 ;
        RECT 138.245 68.210 138.575 68.380 ;
        RECT 139.115 67.870 139.285 74.360 ;
        RECT 137.535 67.700 139.285 67.870 ;
        RECT 131.190 64.685 137.020 64.855 ;
        RECT 126.000 64.325 127.860 64.595 ;
        RECT 126.000 64.155 130.460 64.325 ;
        RECT 126.000 62.745 127.890 64.155 ;
        RECT 128.230 63.285 128.400 63.615 ;
        RECT 128.570 63.585 129.610 63.755 ;
        RECT 128.570 63.145 129.610 63.315 ;
        RECT 129.780 63.285 129.950 63.615 ;
        RECT 130.290 62.745 130.460 64.155 ;
        RECT 126.000 62.575 130.460 62.745 ;
        RECT 131.205 64.240 137.035 64.410 ;
        RECT 131.205 62.830 131.375 64.240 ;
        RECT 131.715 63.370 131.885 63.700 ;
        RECT 132.100 63.670 136.140 63.840 ;
        RECT 132.100 63.230 136.140 63.400 ;
        RECT 136.355 63.370 136.525 63.700 ;
        RECT 136.865 62.830 137.035 64.240 ;
        RECT 131.205 62.660 137.035 62.830 ;
        RECT 126.000 62.300 127.860 62.575 ;
        RECT 140.880 62.385 141.580 74.435 ;
        RECT 126.000 62.130 130.465 62.300 ;
        RECT 126.000 60.720 126.895 62.130 ;
        RECT 127.235 61.260 127.405 61.590 ;
        RECT 127.575 61.560 129.615 61.730 ;
        RECT 127.575 61.120 129.615 61.290 ;
        RECT 129.785 61.260 129.955 61.590 ;
        RECT 130.295 60.720 130.465 62.130 ;
        RECT 114.210 60.635 124.040 60.690 ;
        RECT 126.000 60.560 130.465 60.720 ;
        RECT 131.210 62.215 141.580 62.385 ;
        RECT 131.210 60.805 131.380 62.215 ;
        RECT 131.720 61.345 131.890 61.675 ;
        RECT 132.105 61.645 140.145 61.815 ;
        RECT 132.105 61.205 140.145 61.375 ;
        RECT 140.360 61.345 140.530 61.675 ;
        RECT 140.870 60.805 141.580 62.215 ;
        RECT 131.210 60.690 141.580 60.805 ;
        RECT 143.000 86.485 143.865 87.140 ;
        RECT 148.195 86.975 158.580 87.145 ;
        RECT 143.000 86.315 147.455 86.485 ;
        RECT 143.000 81.055 143.885 86.315 ;
        RECT 144.565 85.745 146.605 85.915 ;
        RECT 144.225 81.685 144.395 85.685 ;
        RECT 146.775 81.685 146.945 85.685 ;
        RECT 144.565 81.455 146.605 81.625 ;
        RECT 147.285 81.055 147.455 86.315 ;
        RECT 148.195 83.485 148.365 86.975 ;
        RECT 148.995 86.465 156.995 86.635 ;
        RECT 148.765 84.210 148.935 86.250 ;
        RECT 157.055 84.210 157.225 86.250 ;
        RECT 148.995 83.825 156.995 83.995 ;
        RECT 157.625 83.485 158.580 86.975 ;
        RECT 148.195 83.315 158.580 83.485 ;
        RECT 157.625 83.025 158.580 83.315 ;
        RECT 143.000 80.885 147.455 81.055 ;
        RECT 143.000 75.625 143.885 80.885 ;
        RECT 144.565 80.315 146.605 80.485 ;
        RECT 144.225 76.255 144.395 80.255 ;
        RECT 146.775 76.255 146.945 80.255 ;
        RECT 144.565 76.025 146.605 76.195 ;
        RECT 147.285 75.625 147.455 80.885 ;
        RECT 148.195 82.855 158.580 83.025 ;
        RECT 148.195 79.595 148.365 82.855 ;
        RECT 149.090 82.285 157.130 82.455 ;
        RECT 148.705 80.225 148.875 82.225 ;
        RECT 157.345 80.225 157.515 82.225 ;
        RECT 149.090 79.995 157.130 80.165 ;
        RECT 157.855 79.595 158.580 82.855 ;
        RECT 148.195 79.425 158.580 79.595 ;
        RECT 148.195 76.165 148.365 79.425 ;
        RECT 149.090 78.855 157.130 79.025 ;
        RECT 148.705 76.795 148.875 78.795 ;
        RECT 157.345 76.795 157.515 78.795 ;
        RECT 149.090 76.565 157.130 76.735 ;
        RECT 157.855 76.165 158.580 79.425 ;
        RECT 148.195 75.995 158.580 76.165 ;
        RECT 153.905 75.715 158.580 75.995 ;
        RECT 143.000 75.455 147.455 75.625 ;
        RECT 143.000 70.195 143.885 75.455 ;
        RECT 144.565 74.885 146.605 75.055 ;
        RECT 144.225 70.825 144.395 74.825 ;
        RECT 146.775 70.825 146.945 74.825 ;
        RECT 144.565 70.595 146.605 70.765 ;
        RECT 147.285 70.195 147.455 75.455 ;
        RECT 143.000 70.025 147.455 70.195 ;
        RECT 143.000 64.765 143.885 70.025 ;
        RECT 144.565 69.455 146.605 69.625 ;
        RECT 144.225 65.395 144.395 69.395 ;
        RECT 146.775 65.395 146.945 69.395 ;
        RECT 144.565 65.165 146.605 65.335 ;
        RECT 147.285 64.765 147.455 70.025 ;
        RECT 143.000 64.595 147.455 64.765 ;
        RECT 148.190 75.545 158.580 75.715 ;
        RECT 148.190 70.285 148.360 75.545 ;
        RECT 149.085 74.975 153.125 75.145 ;
        RECT 148.700 70.915 148.870 74.915 ;
        RECT 153.340 70.915 153.510 74.915 ;
        RECT 153.850 74.435 158.580 75.545 ;
        RECT 149.085 70.685 153.125 70.855 ;
        RECT 153.850 70.285 154.020 74.435 ;
        RECT 148.190 70.115 154.020 70.285 ;
        RECT 148.190 64.855 148.360 70.115 ;
        RECT 149.085 69.545 153.125 69.715 ;
        RECT 148.700 65.485 148.870 69.485 ;
        RECT 153.340 65.485 153.510 69.485 ;
        RECT 149.085 65.255 153.125 65.425 ;
        RECT 153.850 64.855 154.020 70.115 ;
        RECT 154.535 74.360 156.285 74.435 ;
        RECT 154.535 67.870 154.705 74.360 ;
        RECT 155.245 73.850 155.575 74.020 ;
        RECT 155.105 68.595 155.275 73.635 ;
        RECT 155.545 68.595 155.715 73.635 ;
        RECT 155.245 68.210 155.575 68.380 ;
        RECT 156.115 67.870 156.285 74.360 ;
        RECT 154.535 67.700 156.285 67.870 ;
        RECT 148.190 64.685 154.020 64.855 ;
        RECT 143.000 64.325 144.860 64.595 ;
        RECT 143.000 64.155 147.460 64.325 ;
        RECT 143.000 62.745 144.890 64.155 ;
        RECT 145.230 63.285 145.400 63.615 ;
        RECT 145.570 63.585 146.610 63.755 ;
        RECT 145.570 63.145 146.610 63.315 ;
        RECT 146.780 63.285 146.950 63.615 ;
        RECT 147.290 62.745 147.460 64.155 ;
        RECT 143.000 62.575 147.460 62.745 ;
        RECT 148.205 64.240 154.035 64.410 ;
        RECT 148.205 62.830 148.375 64.240 ;
        RECT 148.715 63.370 148.885 63.700 ;
        RECT 149.100 63.670 153.140 63.840 ;
        RECT 149.100 63.230 153.140 63.400 ;
        RECT 153.355 63.370 153.525 63.700 ;
        RECT 153.865 62.830 154.035 64.240 ;
        RECT 148.205 62.660 154.035 62.830 ;
        RECT 143.000 62.300 144.860 62.575 ;
        RECT 157.880 62.385 158.580 74.435 ;
        RECT 143.000 62.130 147.465 62.300 ;
        RECT 143.000 60.720 143.895 62.130 ;
        RECT 144.235 61.260 144.405 61.590 ;
        RECT 144.575 61.560 146.615 61.730 ;
        RECT 144.575 61.120 146.615 61.290 ;
        RECT 146.785 61.260 146.955 61.590 ;
        RECT 147.295 60.720 147.465 62.130 ;
        RECT 131.210 60.635 141.040 60.690 ;
        RECT 143.000 60.560 147.465 60.720 ;
        RECT 148.210 62.215 158.580 62.385 ;
        RECT 148.210 60.805 148.380 62.215 ;
        RECT 148.720 61.345 148.890 61.675 ;
        RECT 149.105 61.645 157.145 61.815 ;
        RECT 149.105 61.205 157.145 61.375 ;
        RECT 157.360 61.345 157.530 61.675 ;
        RECT 157.870 60.805 158.580 62.215 ;
        RECT 148.210 60.690 158.580 60.805 ;
        RECT 148.210 60.635 158.040 60.690 ;
        RECT 75.725 60.550 79.465 60.560 ;
        RECT 92.725 60.550 96.465 60.560 ;
        RECT 109.725 60.550 113.465 60.560 ;
        RECT 126.725 60.550 130.465 60.560 ;
        RECT 143.725 60.550 147.465 60.560 ;
        RECT 22.520 59.155 58.400 59.325 ;
        RECT 22.605 58.065 23.815 59.155 ;
        RECT 23.985 58.720 29.330 59.155 ;
        RECT 22.605 57.355 23.125 57.895 ;
        RECT 23.295 57.525 23.815 58.065 ;
        RECT 22.605 56.605 23.815 57.355 ;
        RECT 25.570 57.150 25.910 57.980 ;
        RECT 27.390 57.470 27.740 58.720 ;
        RECT 30.515 58.225 30.685 58.985 ;
        RECT 30.900 58.395 31.230 59.155 ;
        RECT 30.515 58.055 31.230 58.225 ;
        RECT 31.400 58.080 31.655 58.985 ;
        RECT 30.425 57.505 30.780 57.875 ;
        RECT 31.060 57.845 31.230 58.055 ;
        RECT 31.060 57.515 31.315 57.845 ;
        RECT 31.060 57.325 31.230 57.515 ;
        RECT 31.485 57.350 31.655 58.080 ;
        RECT 31.830 58.005 32.090 59.155 ;
        RECT 32.275 58.355 32.605 59.155 ;
        RECT 32.785 58.815 34.215 58.985 ;
        RECT 32.785 58.185 33.035 58.815 ;
        RECT 32.265 58.015 33.035 58.185 ;
        RECT 30.515 57.155 31.230 57.325 ;
        RECT 23.985 56.605 29.330 57.150 ;
        RECT 30.515 56.775 30.685 57.155 ;
        RECT 30.900 56.605 31.230 56.985 ;
        RECT 31.400 56.775 31.655 57.350 ;
        RECT 31.830 56.605 32.090 57.445 ;
        RECT 32.265 57.345 32.435 58.015 ;
        RECT 32.605 57.515 33.010 57.845 ;
        RECT 33.225 57.515 33.475 58.645 ;
        RECT 33.675 57.845 33.875 58.645 ;
        RECT 34.045 58.135 34.215 58.815 ;
        RECT 34.385 58.305 34.700 59.155 ;
        RECT 34.875 58.355 35.315 58.985 ;
        RECT 34.045 57.965 34.835 58.135 ;
        RECT 33.675 57.515 33.920 57.845 ;
        RECT 34.105 57.515 34.495 57.795 ;
        RECT 34.665 57.515 34.835 57.965 ;
        RECT 35.005 57.345 35.315 58.355 ;
        RECT 35.485 57.990 35.775 59.155 ;
        RECT 36.980 58.525 37.265 58.985 ;
        RECT 37.435 58.695 37.705 59.155 ;
        RECT 36.980 58.305 37.935 58.525 ;
        RECT 36.865 57.575 37.555 58.135 ;
        RECT 37.725 57.405 37.935 58.305 ;
        RECT 32.265 56.775 32.755 57.345 ;
        RECT 32.925 57.175 34.085 57.345 ;
        RECT 32.925 56.775 33.155 57.175 ;
        RECT 33.325 56.605 33.745 57.005 ;
        RECT 33.915 56.775 34.085 57.175 ;
        RECT 34.255 56.605 34.705 57.345 ;
        RECT 34.875 56.785 35.315 57.345 ;
        RECT 35.485 56.605 35.775 57.330 ;
        RECT 36.980 57.235 37.935 57.405 ;
        RECT 38.105 58.135 38.505 58.985 ;
        RECT 38.695 58.525 38.975 58.985 ;
        RECT 39.495 58.695 39.820 59.155 ;
        RECT 38.695 58.305 39.820 58.525 ;
        RECT 38.105 57.575 39.200 58.135 ;
        RECT 39.370 57.845 39.820 58.305 ;
        RECT 39.990 58.015 40.375 58.985 ;
        RECT 36.980 56.775 37.265 57.235 ;
        RECT 37.435 56.605 37.705 57.065 ;
        RECT 38.105 56.775 38.505 57.575 ;
        RECT 39.370 57.515 39.925 57.845 ;
        RECT 39.370 57.405 39.820 57.515 ;
        RECT 38.695 57.235 39.820 57.405 ;
        RECT 40.095 57.345 40.375 58.015 ;
        RECT 41.470 58.005 41.730 59.155 ;
        RECT 41.905 58.080 42.160 58.985 ;
        RECT 42.330 58.395 42.660 59.155 ;
        RECT 42.875 58.225 43.045 58.985 ;
        RECT 43.420 58.525 43.705 58.985 ;
        RECT 43.875 58.695 44.145 59.155 ;
        RECT 43.420 58.305 44.375 58.525 ;
        RECT 38.695 56.775 38.975 57.235 ;
        RECT 39.495 56.605 39.820 57.065 ;
        RECT 39.990 56.775 40.375 57.345 ;
        RECT 41.470 56.605 41.730 57.445 ;
        RECT 41.905 57.350 42.075 58.080 ;
        RECT 42.330 58.055 43.045 58.225 ;
        RECT 42.330 57.845 42.500 58.055 ;
        RECT 42.245 57.515 42.500 57.845 ;
        RECT 41.905 56.775 42.160 57.350 ;
        RECT 42.330 57.325 42.500 57.515 ;
        RECT 42.780 57.505 43.135 57.875 ;
        RECT 43.305 57.575 43.995 58.135 ;
        RECT 44.165 57.405 44.375 58.305 ;
        RECT 42.330 57.155 43.045 57.325 ;
        RECT 42.330 56.605 42.660 56.985 ;
        RECT 42.875 56.775 43.045 57.155 ;
        RECT 43.420 57.235 44.375 57.405 ;
        RECT 44.545 58.135 44.945 58.985 ;
        RECT 45.135 58.525 45.415 58.985 ;
        RECT 45.935 58.695 46.260 59.155 ;
        RECT 45.135 58.305 46.260 58.525 ;
        RECT 44.545 57.575 45.640 58.135 ;
        RECT 45.810 57.845 46.260 58.305 ;
        RECT 46.430 58.015 46.815 58.985 ;
        RECT 47.065 58.225 47.245 58.985 ;
        RECT 47.425 58.395 47.755 59.155 ;
        RECT 47.065 58.055 47.740 58.225 ;
        RECT 47.925 58.080 48.195 58.985 ;
        RECT 43.420 56.775 43.705 57.235 ;
        RECT 43.875 56.605 44.145 57.065 ;
        RECT 44.545 56.775 44.945 57.575 ;
        RECT 45.810 57.515 46.365 57.845 ;
        RECT 45.810 57.405 46.260 57.515 ;
        RECT 45.135 57.235 46.260 57.405 ;
        RECT 46.535 57.345 46.815 58.015 ;
        RECT 47.570 57.910 47.740 58.055 ;
        RECT 47.005 57.505 47.345 57.875 ;
        RECT 47.570 57.580 47.845 57.910 ;
        RECT 45.135 56.775 45.415 57.235 ;
        RECT 45.935 56.605 46.260 57.065 ;
        RECT 46.430 56.775 46.815 57.345 ;
        RECT 47.570 57.325 47.740 57.580 ;
        RECT 47.075 57.155 47.740 57.325 ;
        RECT 48.015 57.280 48.195 58.080 ;
        RECT 48.365 57.990 48.655 59.155 ;
        RECT 49.750 58.005 50.010 59.155 ;
        RECT 50.185 58.080 50.440 58.985 ;
        RECT 50.610 58.395 50.940 59.155 ;
        RECT 51.155 58.225 51.325 58.985 ;
        RECT 47.075 56.775 47.245 57.155 ;
        RECT 47.425 56.605 47.755 56.985 ;
        RECT 47.935 56.775 48.195 57.280 ;
        RECT 48.365 56.605 48.655 57.330 ;
        RECT 49.750 56.605 50.010 57.445 ;
        RECT 50.185 57.350 50.355 58.080 ;
        RECT 50.610 58.055 51.325 58.225 ;
        RECT 51.585 58.065 52.795 59.155 ;
        RECT 50.610 57.845 50.780 58.055 ;
        RECT 50.525 57.515 50.780 57.845 ;
        RECT 50.185 56.775 50.440 57.350 ;
        RECT 50.610 57.325 50.780 57.515 ;
        RECT 51.060 57.505 51.415 57.875 ;
        RECT 51.585 57.355 52.105 57.895 ;
        RECT 52.275 57.525 52.795 58.065 ;
        RECT 52.965 58.080 53.235 58.985 ;
        RECT 53.405 58.395 53.735 59.155 ;
        RECT 53.915 58.225 54.085 58.985 ;
        RECT 50.610 57.155 51.325 57.325 ;
        RECT 50.610 56.605 50.940 56.985 ;
        RECT 51.155 56.775 51.325 57.155 ;
        RECT 51.585 56.605 52.795 57.355 ;
        RECT 52.965 57.280 53.135 58.080 ;
        RECT 53.420 58.055 54.085 58.225 ;
        RECT 54.345 58.080 54.615 58.985 ;
        RECT 54.785 58.395 55.115 59.155 ;
        RECT 55.295 58.225 55.465 58.985 ;
        RECT 53.420 57.910 53.590 58.055 ;
        RECT 53.305 57.580 53.590 57.910 ;
        RECT 53.420 57.325 53.590 57.580 ;
        RECT 53.825 57.505 54.155 57.875 ;
        RECT 52.965 56.775 53.225 57.280 ;
        RECT 53.420 57.155 54.085 57.325 ;
        RECT 53.405 56.605 53.735 56.985 ;
        RECT 53.915 56.775 54.085 57.155 ;
        RECT 54.345 57.280 54.515 58.080 ;
        RECT 54.800 58.055 55.465 58.225 ;
        RECT 55.725 58.080 55.995 58.985 ;
        RECT 56.165 58.395 56.495 59.155 ;
        RECT 56.675 58.225 56.855 58.985 ;
        RECT 54.800 57.910 54.970 58.055 ;
        RECT 54.685 57.580 54.970 57.910 ;
        RECT 54.800 57.325 54.970 57.580 ;
        RECT 55.205 57.505 55.535 57.875 ;
        RECT 54.345 56.775 54.605 57.280 ;
        RECT 54.800 57.155 55.465 57.325 ;
        RECT 54.785 56.605 55.115 56.985 ;
        RECT 55.295 56.775 55.465 57.155 ;
        RECT 55.725 57.280 55.905 58.080 ;
        RECT 56.180 58.055 56.855 58.225 ;
        RECT 57.105 58.065 58.315 59.155 ;
        RECT 89.625 58.165 90.100 58.180 ;
        RECT 106.625 58.165 107.100 58.180 ;
        RECT 123.625 58.165 124.100 58.180 ;
        RECT 140.625 58.165 141.100 58.180 ;
        RECT 157.625 58.165 158.100 58.180 ;
        RECT 89.625 58.145 90.580 58.165 ;
        RECT 106.625 58.145 107.580 58.165 ;
        RECT 123.625 58.145 124.580 58.165 ;
        RECT 140.625 58.145 141.580 58.165 ;
        RECT 157.625 58.145 158.580 58.165 ;
        RECT 56.180 57.910 56.350 58.055 ;
        RECT 56.075 57.580 56.350 57.910 ;
        RECT 56.180 57.325 56.350 57.580 ;
        RECT 56.575 57.505 56.915 57.875 ;
        RECT 57.105 57.525 57.625 58.065 ;
        RECT 57.795 57.355 58.315 57.895 ;
        RECT 55.725 56.775 55.985 57.280 ;
        RECT 56.180 57.155 56.845 57.325 ;
        RECT 56.165 56.605 56.495 56.985 ;
        RECT 56.675 56.775 56.845 57.155 ;
        RECT 57.105 56.605 58.315 57.355 ;
        RECT 75.000 57.485 75.865 58.140 ;
        RECT 80.195 57.975 90.580 58.145 ;
        RECT 75.000 57.315 79.455 57.485 ;
        RECT 22.520 56.435 58.400 56.605 ;
        RECT 22.605 55.685 23.815 56.435 ;
        RECT 22.605 55.145 23.125 55.685 ;
        RECT 23.985 55.665 27.495 56.435 ;
        RECT 28.175 55.780 28.505 56.215 ;
        RECT 28.675 55.825 28.845 56.435 ;
        RECT 28.125 55.695 28.505 55.780 ;
        RECT 29.015 55.695 29.345 56.220 ;
        RECT 29.605 55.905 29.815 56.435 ;
        RECT 30.090 55.985 30.875 56.155 ;
        RECT 31.045 55.985 31.450 56.155 ;
        RECT 23.295 54.975 23.815 55.515 ;
        RECT 23.985 55.145 25.635 55.665 ;
        RECT 28.125 55.655 28.350 55.695 ;
        RECT 25.805 54.975 27.495 55.495 ;
        RECT 22.605 53.885 23.815 54.975 ;
        RECT 23.985 53.885 27.495 54.975 ;
        RECT 28.125 55.075 28.295 55.655 ;
        RECT 29.015 55.525 29.215 55.695 ;
        RECT 30.090 55.525 30.260 55.985 ;
        RECT 28.465 55.195 29.215 55.525 ;
        RECT 29.385 55.195 30.260 55.525 ;
        RECT 28.125 55.025 28.340 55.075 ;
        RECT 28.125 54.945 28.515 55.025 ;
        RECT 28.185 54.100 28.515 54.945 ;
        RECT 29.025 54.990 29.215 55.195 ;
        RECT 28.685 53.885 28.855 54.895 ;
        RECT 29.025 54.615 29.920 54.990 ;
        RECT 29.025 54.055 29.365 54.615 ;
        RECT 29.595 53.885 29.910 54.385 ;
        RECT 30.090 54.355 30.260 55.195 ;
        RECT 30.430 55.485 30.895 55.815 ;
        RECT 31.280 55.755 31.450 55.985 ;
        RECT 31.630 55.935 32.000 56.435 ;
        RECT 32.320 55.985 32.995 56.155 ;
        RECT 33.190 55.985 33.525 56.155 ;
        RECT 30.430 54.525 30.750 55.485 ;
        RECT 31.280 55.455 32.110 55.755 ;
        RECT 30.920 54.555 31.110 55.275 ;
        RECT 31.280 54.385 31.450 55.455 ;
        RECT 31.910 55.425 32.110 55.455 ;
        RECT 31.620 55.205 31.790 55.275 ;
        RECT 32.320 55.205 32.490 55.985 ;
        RECT 33.355 55.845 33.525 55.985 ;
        RECT 33.695 55.975 33.945 56.435 ;
        RECT 31.620 55.035 32.490 55.205 ;
        RECT 32.660 55.565 33.185 55.785 ;
        RECT 33.355 55.715 33.580 55.845 ;
        RECT 31.620 54.945 32.130 55.035 ;
        RECT 30.090 54.185 30.975 54.355 ;
        RECT 31.200 54.055 31.450 54.385 ;
        RECT 31.620 53.885 31.790 54.685 ;
        RECT 31.960 54.330 32.130 54.945 ;
        RECT 32.660 54.865 32.830 55.565 ;
        RECT 32.300 54.500 32.830 54.865 ;
        RECT 33.000 54.800 33.240 55.395 ;
        RECT 33.410 54.610 33.580 55.715 ;
        RECT 33.750 54.855 34.030 55.805 ;
        RECT 33.275 54.480 33.580 54.610 ;
        RECT 31.960 54.160 33.065 54.330 ;
        RECT 33.275 54.055 33.525 54.480 ;
        RECT 33.695 53.885 33.960 54.345 ;
        RECT 34.200 54.055 34.385 56.175 ;
        RECT 34.555 56.055 34.885 56.435 ;
        RECT 35.055 55.885 35.225 56.175 ;
        RECT 34.560 55.715 35.225 55.885 ;
        RECT 35.575 55.885 35.745 56.175 ;
        RECT 35.915 56.055 36.245 56.435 ;
        RECT 35.575 55.715 36.240 55.885 ;
        RECT 34.560 54.725 34.790 55.715 ;
        RECT 34.960 54.895 35.310 55.545 ;
        RECT 35.490 54.895 35.840 55.545 ;
        RECT 36.010 54.725 36.240 55.715 ;
        RECT 34.560 54.555 35.225 54.725 ;
        RECT 34.555 53.885 34.885 54.385 ;
        RECT 35.055 54.055 35.225 54.555 ;
        RECT 35.575 54.555 36.240 54.725 ;
        RECT 35.575 54.055 35.745 54.555 ;
        RECT 35.915 53.885 36.245 54.385 ;
        RECT 36.415 54.055 36.600 56.175 ;
        RECT 36.855 55.975 37.105 56.435 ;
        RECT 37.275 55.985 37.610 56.155 ;
        RECT 37.805 55.985 38.480 56.155 ;
        RECT 37.275 55.845 37.445 55.985 ;
        RECT 36.770 54.855 37.050 55.805 ;
        RECT 37.220 55.715 37.445 55.845 ;
        RECT 37.220 54.610 37.390 55.715 ;
        RECT 37.615 55.565 38.140 55.785 ;
        RECT 37.560 54.800 37.800 55.395 ;
        RECT 37.970 54.865 38.140 55.565 ;
        RECT 38.310 55.205 38.480 55.985 ;
        RECT 38.800 55.935 39.170 56.435 ;
        RECT 39.350 55.985 39.755 56.155 ;
        RECT 39.925 55.985 40.710 56.155 ;
        RECT 39.350 55.755 39.520 55.985 ;
        RECT 38.690 55.455 39.520 55.755 ;
        RECT 39.905 55.485 40.370 55.815 ;
        RECT 38.690 55.425 38.890 55.455 ;
        RECT 39.010 55.205 39.180 55.275 ;
        RECT 38.310 55.035 39.180 55.205 ;
        RECT 38.670 54.945 39.180 55.035 ;
        RECT 37.220 54.480 37.525 54.610 ;
        RECT 37.970 54.500 38.500 54.865 ;
        RECT 36.840 53.885 37.105 54.345 ;
        RECT 37.275 54.055 37.525 54.480 ;
        RECT 38.670 54.330 38.840 54.945 ;
        RECT 37.735 54.160 38.840 54.330 ;
        RECT 39.010 53.885 39.180 54.685 ;
        RECT 39.350 54.385 39.520 55.455 ;
        RECT 39.690 54.555 39.880 55.275 ;
        RECT 40.050 54.525 40.370 55.485 ;
        RECT 40.540 55.525 40.710 55.985 ;
        RECT 40.985 55.905 41.195 56.435 ;
        RECT 41.455 55.695 41.785 56.220 ;
        RECT 41.955 55.825 42.125 56.435 ;
        RECT 42.295 55.780 42.625 56.215 ;
        RECT 42.295 55.695 42.675 55.780 ;
        RECT 41.585 55.525 41.785 55.695 ;
        RECT 42.450 55.655 42.675 55.695 ;
        RECT 40.540 55.195 41.415 55.525 ;
        RECT 41.585 55.195 42.335 55.525 ;
        RECT 39.350 54.055 39.600 54.385 ;
        RECT 40.540 54.355 40.710 55.195 ;
        RECT 41.585 54.990 41.775 55.195 ;
        RECT 42.505 55.075 42.675 55.655 ;
        RECT 42.460 55.025 42.675 55.075 ;
        RECT 40.880 54.615 41.775 54.990 ;
        RECT 42.285 54.945 42.675 55.025 ;
        RECT 42.880 55.695 43.495 56.265 ;
        RECT 43.665 55.925 43.880 56.435 ;
        RECT 44.110 55.925 44.390 56.255 ;
        RECT 44.570 55.925 44.810 56.435 ;
        RECT 39.825 54.185 40.710 54.355 ;
        RECT 40.890 53.885 41.205 54.385 ;
        RECT 41.435 54.055 41.775 54.615 ;
        RECT 41.945 53.885 42.115 54.895 ;
        RECT 42.285 54.100 42.615 54.945 ;
        RECT 42.880 54.675 43.195 55.695 ;
        RECT 43.365 55.025 43.535 55.525 ;
        RECT 43.785 55.195 44.050 55.755 ;
        RECT 44.220 55.025 44.390 55.925 ;
        RECT 45.235 55.885 45.405 56.265 ;
        RECT 45.620 56.055 45.950 56.435 ;
        RECT 44.560 55.195 44.915 55.755 ;
        RECT 45.235 55.715 45.950 55.885 ;
        RECT 45.145 55.165 45.500 55.535 ;
        RECT 45.780 55.525 45.950 55.715 ;
        RECT 46.120 55.690 46.375 56.265 ;
        RECT 45.780 55.195 46.035 55.525 ;
        RECT 43.365 54.855 44.790 55.025 ;
        RECT 45.780 54.985 45.950 55.195 ;
        RECT 42.880 54.055 43.415 54.675 ;
        RECT 43.585 53.885 43.915 54.685 ;
        RECT 44.400 54.680 44.790 54.855 ;
        RECT 45.235 54.815 45.950 54.985 ;
        RECT 46.205 54.960 46.375 55.690 ;
        RECT 46.550 55.595 46.810 56.435 ;
        RECT 47.025 55.615 47.255 56.435 ;
        RECT 47.425 55.635 47.755 56.265 ;
        RECT 47.005 55.195 47.335 55.445 ;
        RECT 47.505 55.035 47.755 55.635 ;
        RECT 47.925 55.615 48.135 56.435 ;
        RECT 48.365 55.710 48.655 56.435 ;
        RECT 48.825 55.695 49.265 56.255 ;
        RECT 49.435 55.695 49.885 56.435 ;
        RECT 50.055 55.865 50.225 56.265 ;
        RECT 50.395 56.035 50.815 56.435 ;
        RECT 50.985 55.865 51.215 56.265 ;
        RECT 50.055 55.695 51.215 55.865 ;
        RECT 51.385 55.695 51.875 56.265 ;
        RECT 45.235 54.055 45.405 54.815 ;
        RECT 45.620 53.885 45.950 54.645 ;
        RECT 46.120 54.055 46.375 54.960 ;
        RECT 46.550 53.885 46.810 55.035 ;
        RECT 47.025 53.885 47.255 55.025 ;
        RECT 47.425 54.055 47.755 55.035 ;
        RECT 47.925 53.885 48.135 55.025 ;
        RECT 48.365 53.885 48.655 55.050 ;
        RECT 48.825 54.685 49.135 55.695 ;
        RECT 49.305 55.075 49.475 55.525 ;
        RECT 49.645 55.245 50.035 55.525 ;
        RECT 50.220 55.195 50.465 55.525 ;
        RECT 49.305 54.905 50.095 55.075 ;
        RECT 48.825 54.055 49.265 54.685 ;
        RECT 49.440 53.885 49.755 54.735 ;
        RECT 49.925 54.225 50.095 54.905 ;
        RECT 50.265 54.395 50.465 55.195 ;
        RECT 50.665 54.395 50.915 55.525 ;
        RECT 51.130 55.195 51.535 55.525 ;
        RECT 51.705 55.025 51.875 55.695 ;
        RECT 52.160 55.805 52.445 56.265 ;
        RECT 52.615 55.975 52.885 56.435 ;
        RECT 52.160 55.635 53.115 55.805 ;
        RECT 51.105 54.855 51.875 55.025 ;
        RECT 52.045 54.905 52.735 55.465 ;
        RECT 51.105 54.225 51.355 54.855 ;
        RECT 52.905 54.735 53.115 55.635 ;
        RECT 49.925 54.055 51.355 54.225 ;
        RECT 51.535 53.885 51.865 54.685 ;
        RECT 52.160 54.515 53.115 54.735 ;
        RECT 53.285 55.465 53.685 56.265 ;
        RECT 53.875 55.805 54.155 56.265 ;
        RECT 54.675 55.975 55.000 56.435 ;
        RECT 53.875 55.635 55.000 55.805 ;
        RECT 55.170 55.695 55.555 56.265 ;
        RECT 54.550 55.525 55.000 55.635 ;
        RECT 53.285 54.905 54.380 55.465 ;
        RECT 54.550 55.195 55.105 55.525 ;
        RECT 52.160 54.055 52.445 54.515 ;
        RECT 52.615 53.885 52.885 54.345 ;
        RECT 53.285 54.055 53.685 54.905 ;
        RECT 54.550 54.735 55.000 55.195 ;
        RECT 55.275 55.025 55.555 55.695 ;
        RECT 53.875 54.515 55.000 54.735 ;
        RECT 53.875 54.055 54.155 54.515 ;
        RECT 54.675 53.885 55.000 54.345 ;
        RECT 55.170 54.055 55.555 55.025 ;
        RECT 55.725 55.760 55.985 56.265 ;
        RECT 56.165 56.055 56.495 56.435 ;
        RECT 56.675 55.885 56.845 56.265 ;
        RECT 55.725 54.960 55.905 55.760 ;
        RECT 56.180 55.715 56.845 55.885 ;
        RECT 56.180 55.460 56.350 55.715 ;
        RECT 57.105 55.685 58.315 56.435 ;
        RECT 56.075 55.130 56.350 55.460 ;
        RECT 56.575 55.165 56.915 55.535 ;
        RECT 56.180 54.985 56.350 55.130 ;
        RECT 55.725 54.055 55.995 54.960 ;
        RECT 56.180 54.815 56.855 54.985 ;
        RECT 56.165 53.885 56.495 54.645 ;
        RECT 56.675 54.055 56.855 54.815 ;
        RECT 57.105 54.975 57.625 55.515 ;
        RECT 57.795 55.145 58.315 55.685 ;
        RECT 57.105 53.885 58.315 54.975 ;
        RECT 22.520 53.715 58.400 53.885 ;
        RECT 22.605 52.625 23.815 53.715 ;
        RECT 24.075 53.045 24.245 53.545 ;
        RECT 24.415 53.215 24.745 53.715 ;
        RECT 24.075 52.875 24.740 53.045 ;
        RECT 22.605 51.915 23.125 52.455 ;
        RECT 23.295 52.085 23.815 52.625 ;
        RECT 23.990 52.055 24.340 52.705 ;
        RECT 22.605 51.165 23.815 51.915 ;
        RECT 24.510 51.885 24.740 52.875 ;
        RECT 24.075 51.715 24.740 51.885 ;
        RECT 24.075 51.425 24.245 51.715 ;
        RECT 24.415 51.165 24.745 51.545 ;
        RECT 24.915 51.425 25.100 53.545 ;
        RECT 25.340 53.255 25.605 53.715 ;
        RECT 25.775 53.120 26.025 53.545 ;
        RECT 26.235 53.270 27.340 53.440 ;
        RECT 25.720 52.990 26.025 53.120 ;
        RECT 25.270 51.795 25.550 52.745 ;
        RECT 25.720 51.885 25.890 52.990 ;
        RECT 26.060 52.205 26.300 52.800 ;
        RECT 26.470 52.735 27.000 53.100 ;
        RECT 26.470 52.035 26.640 52.735 ;
        RECT 27.170 52.655 27.340 53.270 ;
        RECT 27.510 52.915 27.680 53.715 ;
        RECT 27.850 53.215 28.100 53.545 ;
        RECT 28.325 53.245 29.210 53.415 ;
        RECT 27.170 52.565 27.680 52.655 ;
        RECT 25.720 51.755 25.945 51.885 ;
        RECT 26.115 51.815 26.640 52.035 ;
        RECT 26.810 52.395 27.680 52.565 ;
        RECT 25.355 51.165 25.605 51.625 ;
        RECT 25.775 51.615 25.945 51.755 ;
        RECT 26.810 51.615 26.980 52.395 ;
        RECT 27.510 52.325 27.680 52.395 ;
        RECT 27.190 52.145 27.390 52.175 ;
        RECT 27.850 52.145 28.020 53.215 ;
        RECT 28.190 52.325 28.380 53.045 ;
        RECT 27.190 51.845 28.020 52.145 ;
        RECT 28.550 52.115 28.870 53.075 ;
        RECT 25.775 51.445 26.110 51.615 ;
        RECT 26.305 51.445 26.980 51.615 ;
        RECT 27.300 51.165 27.670 51.665 ;
        RECT 27.850 51.615 28.020 51.845 ;
        RECT 28.405 51.785 28.870 52.115 ;
        RECT 29.040 52.405 29.210 53.245 ;
        RECT 29.390 53.215 29.705 53.715 ;
        RECT 29.935 52.985 30.275 53.545 ;
        RECT 29.380 52.610 30.275 52.985 ;
        RECT 30.445 52.705 30.615 53.715 ;
        RECT 30.085 52.405 30.275 52.610 ;
        RECT 30.785 52.655 31.115 53.500 ;
        RECT 30.785 52.575 31.175 52.655 ;
        RECT 30.960 52.525 31.175 52.575 ;
        RECT 29.040 52.075 29.915 52.405 ;
        RECT 30.085 52.075 30.835 52.405 ;
        RECT 29.040 51.615 29.210 52.075 ;
        RECT 30.085 51.905 30.285 52.075 ;
        RECT 31.005 51.945 31.175 52.525 ;
        RECT 30.950 51.905 31.175 51.945 ;
        RECT 27.850 51.445 28.255 51.615 ;
        RECT 28.425 51.445 29.210 51.615 ;
        RECT 29.485 51.165 29.695 51.695 ;
        RECT 29.955 51.380 30.285 51.905 ;
        RECT 30.795 51.820 31.175 51.905 ;
        RECT 31.345 52.575 31.730 53.545 ;
        RECT 31.900 53.255 32.225 53.715 ;
        RECT 32.745 53.085 33.025 53.545 ;
        RECT 31.900 52.865 33.025 53.085 ;
        RECT 31.345 51.905 31.625 52.575 ;
        RECT 31.900 52.405 32.350 52.865 ;
        RECT 33.215 52.695 33.615 53.545 ;
        RECT 34.015 53.255 34.285 53.715 ;
        RECT 34.455 53.085 34.740 53.545 ;
        RECT 31.795 52.075 32.350 52.405 ;
        RECT 32.520 52.135 33.615 52.695 ;
        RECT 31.900 51.965 32.350 52.075 ;
        RECT 30.455 51.165 30.625 51.775 ;
        RECT 30.795 51.385 31.125 51.820 ;
        RECT 31.345 51.335 31.730 51.905 ;
        RECT 31.900 51.795 33.025 51.965 ;
        RECT 31.900 51.165 32.225 51.625 ;
        RECT 32.745 51.335 33.025 51.795 ;
        RECT 33.215 51.335 33.615 52.135 ;
        RECT 33.785 52.865 34.740 53.085 ;
        RECT 33.785 51.965 33.995 52.865 ;
        RECT 34.165 52.135 34.855 52.695 ;
        RECT 35.485 52.550 35.775 53.715 ;
        RECT 35.950 52.575 36.285 53.545 ;
        RECT 36.455 52.575 36.625 53.715 ;
        RECT 36.795 53.375 38.825 53.545 ;
        RECT 33.785 51.795 34.740 51.965 ;
        RECT 35.950 51.905 36.120 52.575 ;
        RECT 36.795 52.405 36.965 53.375 ;
        RECT 36.290 52.075 36.545 52.405 ;
        RECT 36.770 52.075 36.965 52.405 ;
        RECT 37.135 53.035 38.260 53.205 ;
        RECT 36.375 51.905 36.545 52.075 ;
        RECT 37.135 51.905 37.305 53.035 ;
        RECT 34.015 51.165 34.285 51.625 ;
        RECT 34.455 51.335 34.740 51.795 ;
        RECT 35.485 51.165 35.775 51.890 ;
        RECT 35.950 51.335 36.205 51.905 ;
        RECT 36.375 51.735 37.305 51.905 ;
        RECT 37.475 52.695 38.485 52.865 ;
        RECT 37.475 51.895 37.645 52.695 ;
        RECT 37.850 52.355 38.125 52.495 ;
        RECT 37.845 52.185 38.125 52.355 ;
        RECT 37.130 51.700 37.305 51.735 ;
        RECT 36.375 51.165 36.705 51.565 ;
        RECT 37.130 51.335 37.660 51.700 ;
        RECT 37.850 51.335 38.125 52.185 ;
        RECT 38.295 51.335 38.485 52.695 ;
        RECT 38.655 52.710 38.825 53.375 ;
        RECT 38.995 52.955 39.165 53.715 ;
        RECT 39.400 52.955 39.915 53.365 ;
        RECT 38.655 52.520 39.405 52.710 ;
        RECT 39.575 52.145 39.915 52.955 ;
        RECT 40.730 52.745 41.120 52.920 ;
        RECT 41.605 52.915 41.935 53.715 ;
        RECT 42.105 52.925 42.640 53.545 ;
        RECT 40.730 52.575 42.155 52.745 ;
        RECT 38.685 51.975 39.915 52.145 ;
        RECT 38.665 51.165 39.175 51.700 ;
        RECT 39.395 51.370 39.640 51.975 ;
        RECT 40.605 51.845 40.960 52.405 ;
        RECT 41.130 51.675 41.300 52.575 ;
        RECT 41.470 51.845 41.735 52.405 ;
        RECT 41.985 52.075 42.155 52.575 ;
        RECT 42.325 51.905 42.640 52.925 ;
        RECT 42.905 52.575 43.115 53.715 ;
        RECT 43.285 52.565 43.615 53.545 ;
        RECT 43.785 52.575 44.015 53.715 ;
        RECT 44.315 53.045 44.485 53.545 ;
        RECT 44.655 53.215 44.985 53.715 ;
        RECT 44.315 52.875 44.980 53.045 ;
        RECT 40.710 51.165 40.950 51.675 ;
        RECT 41.130 51.345 41.410 51.675 ;
        RECT 41.640 51.165 41.855 51.675 ;
        RECT 42.025 51.335 42.640 51.905 ;
        RECT 42.905 51.165 43.115 51.985 ;
        RECT 43.285 51.965 43.535 52.565 ;
        RECT 43.705 52.155 44.035 52.405 ;
        RECT 44.230 52.055 44.580 52.705 ;
        RECT 43.285 51.335 43.615 51.965 ;
        RECT 43.785 51.165 44.015 51.985 ;
        RECT 44.750 51.885 44.980 52.875 ;
        RECT 44.315 51.715 44.980 51.885 ;
        RECT 44.315 51.425 44.485 51.715 ;
        RECT 44.655 51.165 44.985 51.545 ;
        RECT 45.155 51.425 45.340 53.545 ;
        RECT 45.580 53.255 45.845 53.715 ;
        RECT 46.015 53.120 46.265 53.545 ;
        RECT 46.475 53.270 47.580 53.440 ;
        RECT 45.960 52.990 46.265 53.120 ;
        RECT 45.510 51.795 45.790 52.745 ;
        RECT 45.960 51.885 46.130 52.990 ;
        RECT 46.300 52.205 46.540 52.800 ;
        RECT 46.710 52.735 47.240 53.100 ;
        RECT 46.710 52.035 46.880 52.735 ;
        RECT 47.410 52.655 47.580 53.270 ;
        RECT 47.750 52.915 47.920 53.715 ;
        RECT 48.090 53.215 48.340 53.545 ;
        RECT 48.565 53.245 49.450 53.415 ;
        RECT 47.410 52.565 47.920 52.655 ;
        RECT 45.960 51.755 46.185 51.885 ;
        RECT 46.355 51.815 46.880 52.035 ;
        RECT 47.050 52.395 47.920 52.565 ;
        RECT 45.595 51.165 45.845 51.625 ;
        RECT 46.015 51.615 46.185 51.755 ;
        RECT 47.050 51.615 47.220 52.395 ;
        RECT 47.750 52.325 47.920 52.395 ;
        RECT 47.430 52.145 47.630 52.175 ;
        RECT 48.090 52.145 48.260 53.215 ;
        RECT 48.430 52.325 48.620 53.045 ;
        RECT 47.430 51.845 48.260 52.145 ;
        RECT 48.790 52.115 49.110 53.075 ;
        RECT 46.015 51.445 46.350 51.615 ;
        RECT 46.545 51.445 47.220 51.615 ;
        RECT 47.540 51.165 47.910 51.665 ;
        RECT 48.090 51.615 48.260 51.845 ;
        RECT 48.645 51.785 49.110 52.115 ;
        RECT 49.280 52.405 49.450 53.245 ;
        RECT 49.630 53.215 49.945 53.715 ;
        RECT 50.175 52.985 50.515 53.545 ;
        RECT 49.620 52.610 50.515 52.985 ;
        RECT 50.685 52.705 50.855 53.715 ;
        RECT 50.325 52.405 50.515 52.610 ;
        RECT 51.025 52.655 51.355 53.500 ;
        RECT 52.230 52.745 52.620 52.920 ;
        RECT 53.105 52.915 53.435 53.715 ;
        RECT 53.605 52.925 54.140 53.545 ;
        RECT 51.025 52.575 51.415 52.655 ;
        RECT 52.230 52.575 53.655 52.745 ;
        RECT 51.200 52.525 51.415 52.575 ;
        RECT 49.280 52.075 50.155 52.405 ;
        RECT 50.325 52.075 51.075 52.405 ;
        RECT 49.280 51.615 49.450 52.075 ;
        RECT 50.325 51.905 50.525 52.075 ;
        RECT 51.245 51.945 51.415 52.525 ;
        RECT 51.190 51.905 51.415 51.945 ;
        RECT 48.090 51.445 48.495 51.615 ;
        RECT 48.665 51.445 49.450 51.615 ;
        RECT 49.725 51.165 49.935 51.695 ;
        RECT 50.195 51.380 50.525 51.905 ;
        RECT 51.035 51.820 51.415 51.905 ;
        RECT 52.105 51.845 52.460 52.405 ;
        RECT 50.695 51.165 50.865 51.775 ;
        RECT 51.035 51.385 51.365 51.820 ;
        RECT 52.630 51.675 52.800 52.575 ;
        RECT 52.970 51.845 53.235 52.405 ;
        RECT 53.485 52.075 53.655 52.575 ;
        RECT 53.825 51.905 54.140 52.925 ;
        RECT 54.435 52.785 54.605 53.545 ;
        RECT 54.785 52.955 55.115 53.715 ;
        RECT 54.435 52.615 55.100 52.785 ;
        RECT 55.285 52.640 55.555 53.545 ;
        RECT 54.930 52.470 55.100 52.615 ;
        RECT 54.365 52.065 54.695 52.435 ;
        RECT 54.930 52.140 55.215 52.470 ;
        RECT 52.210 51.165 52.450 51.675 ;
        RECT 52.630 51.345 52.910 51.675 ;
        RECT 53.140 51.165 53.355 51.675 ;
        RECT 53.525 51.335 54.140 51.905 ;
        RECT 54.930 51.885 55.100 52.140 ;
        RECT 54.435 51.715 55.100 51.885 ;
        RECT 55.385 51.840 55.555 52.640 ;
        RECT 54.435 51.335 54.605 51.715 ;
        RECT 54.785 51.165 55.115 51.545 ;
        RECT 55.295 51.335 55.555 51.840 ;
        RECT 55.725 52.640 55.995 53.545 ;
        RECT 56.165 52.955 56.495 53.715 ;
        RECT 56.675 52.785 56.855 53.545 ;
        RECT 55.725 51.840 55.905 52.640 ;
        RECT 56.180 52.615 56.855 52.785 ;
        RECT 57.105 52.625 58.315 53.715 ;
        RECT 56.180 52.470 56.350 52.615 ;
        RECT 56.075 52.140 56.350 52.470 ;
        RECT 56.180 51.885 56.350 52.140 ;
        RECT 56.575 52.065 56.915 52.435 ;
        RECT 57.105 52.085 57.625 52.625 ;
        RECT 57.795 51.915 58.315 52.455 ;
        RECT 55.725 51.335 55.985 51.840 ;
        RECT 56.180 51.715 56.845 51.885 ;
        RECT 56.165 51.165 56.495 51.545 ;
        RECT 56.675 51.335 56.845 51.715 ;
        RECT 57.105 51.165 58.315 51.915 ;
        RECT 75.000 52.055 75.885 57.315 ;
        RECT 76.565 56.745 78.605 56.915 ;
        RECT 76.225 52.685 76.395 56.685 ;
        RECT 78.775 52.685 78.945 56.685 ;
        RECT 76.565 52.455 78.605 52.625 ;
        RECT 79.285 52.055 79.455 57.315 ;
        RECT 80.195 54.485 80.365 57.975 ;
        RECT 80.995 57.465 88.995 57.635 ;
        RECT 80.765 55.210 80.935 57.250 ;
        RECT 89.055 55.210 89.225 57.250 ;
        RECT 80.995 54.825 88.995 54.995 ;
        RECT 89.625 54.485 90.580 57.975 ;
        RECT 80.195 54.315 90.580 54.485 ;
        RECT 89.625 54.025 90.580 54.315 ;
        RECT 75.000 51.885 79.455 52.055 ;
        RECT 22.520 50.995 58.400 51.165 ;
        RECT 22.605 50.245 23.815 50.995 ;
        RECT 22.605 49.705 23.125 50.245 ;
        RECT 23.990 50.155 24.250 50.995 ;
        RECT 24.425 50.250 24.680 50.825 ;
        RECT 24.850 50.615 25.180 50.995 ;
        RECT 25.395 50.445 25.565 50.825 ;
        RECT 24.850 50.275 25.565 50.445 ;
        RECT 23.295 49.535 23.815 50.075 ;
        RECT 22.605 48.445 23.815 49.535 ;
        RECT 23.990 48.445 24.250 49.595 ;
        RECT 24.425 49.520 24.595 50.250 ;
        RECT 24.850 50.085 25.020 50.275 ;
        RECT 25.830 50.255 26.085 50.825 ;
        RECT 26.255 50.595 26.585 50.995 ;
        RECT 27.010 50.460 27.540 50.825 ;
        RECT 27.730 50.655 28.005 50.825 ;
        RECT 27.725 50.485 28.005 50.655 ;
        RECT 27.010 50.425 27.185 50.460 ;
        RECT 26.255 50.255 27.185 50.425 ;
        RECT 24.765 49.755 25.020 50.085 ;
        RECT 24.850 49.545 25.020 49.755 ;
        RECT 25.300 49.725 25.655 50.095 ;
        RECT 25.830 49.585 26.000 50.255 ;
        RECT 26.255 50.085 26.425 50.255 ;
        RECT 26.170 49.755 26.425 50.085 ;
        RECT 26.650 49.755 26.845 50.085 ;
        RECT 24.425 48.615 24.680 49.520 ;
        RECT 24.850 49.375 25.565 49.545 ;
        RECT 24.850 48.445 25.180 49.205 ;
        RECT 25.395 48.615 25.565 49.375 ;
        RECT 25.830 48.615 26.165 49.585 ;
        RECT 26.335 48.445 26.505 49.585 ;
        RECT 26.675 48.785 26.845 49.755 ;
        RECT 27.015 49.125 27.185 50.255 ;
        RECT 27.355 49.465 27.525 50.265 ;
        RECT 27.730 49.665 28.005 50.485 ;
        RECT 28.175 49.465 28.365 50.825 ;
        RECT 28.545 50.460 29.055 50.995 ;
        RECT 29.275 50.185 29.520 50.790 ;
        RECT 29.965 50.245 31.175 50.995 ;
        RECT 31.435 50.515 31.735 50.995 ;
        RECT 31.905 50.345 32.165 50.800 ;
        RECT 32.335 50.515 32.595 50.995 ;
        RECT 32.775 50.345 33.035 50.800 ;
        RECT 33.205 50.515 33.455 50.995 ;
        RECT 33.635 50.345 33.895 50.800 ;
        RECT 34.065 50.515 34.315 50.995 ;
        RECT 34.495 50.345 34.755 50.800 ;
        RECT 34.925 50.515 35.170 50.995 ;
        RECT 35.340 50.345 35.615 50.800 ;
        RECT 35.785 50.515 36.030 50.995 ;
        RECT 36.200 50.345 36.460 50.800 ;
        RECT 36.630 50.515 36.890 50.995 ;
        RECT 37.060 50.345 37.320 50.800 ;
        RECT 37.490 50.515 37.750 50.995 ;
        RECT 37.920 50.345 38.180 50.800 ;
        RECT 38.350 50.435 38.610 50.995 ;
        RECT 28.565 50.015 29.795 50.185 ;
        RECT 27.355 49.295 28.365 49.465 ;
        RECT 28.535 49.450 29.285 49.640 ;
        RECT 27.015 48.955 28.140 49.125 ;
        RECT 28.535 48.785 28.705 49.450 ;
        RECT 29.455 49.205 29.795 50.015 ;
        RECT 29.965 49.705 30.485 50.245 ;
        RECT 31.435 50.175 38.180 50.345 ;
        RECT 30.655 49.535 31.175 50.075 ;
        RECT 26.675 48.615 28.705 48.785 ;
        RECT 28.875 48.445 29.045 49.205 ;
        RECT 29.280 48.795 29.795 49.205 ;
        RECT 29.965 48.445 31.175 49.535 ;
        RECT 31.435 49.585 32.600 50.175 ;
        RECT 38.780 50.005 39.030 50.815 ;
        RECT 39.210 50.470 39.470 50.995 ;
        RECT 39.640 50.005 39.890 50.815 ;
        RECT 40.070 50.485 40.375 50.995 ;
        RECT 32.770 49.755 39.890 50.005 ;
        RECT 40.060 49.755 40.375 50.315 ;
        RECT 40.545 50.255 40.930 50.825 ;
        RECT 41.100 50.535 41.425 50.995 ;
        RECT 41.945 50.365 42.225 50.825 ;
        RECT 31.435 49.360 38.180 49.585 ;
        RECT 31.435 48.445 31.705 49.190 ;
        RECT 31.875 48.620 32.165 49.360 ;
        RECT 32.775 49.345 38.180 49.360 ;
        RECT 32.335 48.450 32.590 49.175 ;
        RECT 32.775 48.620 33.035 49.345 ;
        RECT 33.205 48.450 33.450 49.175 ;
        RECT 33.635 48.620 33.895 49.345 ;
        RECT 34.065 48.450 34.310 49.175 ;
        RECT 34.495 48.620 34.755 49.345 ;
        RECT 34.925 48.450 35.170 49.175 ;
        RECT 35.340 48.620 35.600 49.345 ;
        RECT 35.770 48.450 36.030 49.175 ;
        RECT 36.200 48.620 36.460 49.345 ;
        RECT 36.630 48.450 36.890 49.175 ;
        RECT 37.060 48.620 37.320 49.345 ;
        RECT 37.490 48.450 37.750 49.175 ;
        RECT 37.920 48.620 38.180 49.345 ;
        RECT 38.350 48.450 38.610 49.245 ;
        RECT 38.780 48.620 39.030 49.755 ;
        RECT 32.335 48.445 38.610 48.450 ;
        RECT 39.210 48.445 39.470 49.255 ;
        RECT 39.645 48.615 39.890 49.755 ;
        RECT 40.545 49.585 40.825 50.255 ;
        RECT 41.100 50.195 42.225 50.365 ;
        RECT 41.100 50.085 41.550 50.195 ;
        RECT 40.995 49.755 41.550 50.085 ;
        RECT 42.415 50.025 42.815 50.825 ;
        RECT 43.215 50.535 43.485 50.995 ;
        RECT 43.655 50.365 43.940 50.825 ;
        RECT 40.070 48.445 40.365 49.255 ;
        RECT 40.545 48.615 40.930 49.585 ;
        RECT 41.100 49.295 41.550 49.755 ;
        RECT 41.720 49.465 42.815 50.025 ;
        RECT 41.100 49.075 42.225 49.295 ;
        RECT 41.100 48.445 41.425 48.905 ;
        RECT 41.945 48.615 42.225 49.075 ;
        RECT 42.415 48.615 42.815 49.465 ;
        RECT 42.985 50.195 43.940 50.365 ;
        RECT 44.225 50.245 45.435 50.995 ;
        RECT 45.615 50.495 45.945 50.995 ;
        RECT 46.145 50.425 46.315 50.775 ;
        RECT 46.515 50.595 46.845 50.995 ;
        RECT 47.015 50.425 47.185 50.775 ;
        RECT 47.355 50.595 47.735 50.995 ;
        RECT 42.985 49.295 43.195 50.195 ;
        RECT 43.365 49.465 44.055 50.025 ;
        RECT 44.225 49.705 44.745 50.245 ;
        RECT 44.915 49.535 45.435 50.075 ;
        RECT 45.610 49.755 45.960 50.325 ;
        RECT 46.145 50.255 47.755 50.425 ;
        RECT 47.925 50.320 48.195 50.665 ;
        RECT 47.585 50.085 47.755 50.255 ;
        RECT 42.985 49.075 43.940 49.295 ;
        RECT 43.215 48.445 43.485 48.905 ;
        RECT 43.655 48.615 43.940 49.075 ;
        RECT 44.225 48.445 45.435 49.535 ;
        RECT 45.610 49.295 45.930 49.585 ;
        RECT 46.130 49.465 46.840 50.085 ;
        RECT 47.010 49.755 47.415 50.085 ;
        RECT 47.585 49.755 47.855 50.085 ;
        RECT 47.585 49.585 47.755 49.755 ;
        RECT 48.025 49.585 48.195 50.320 ;
        RECT 48.365 50.270 48.655 50.995 ;
        RECT 48.825 50.255 49.185 50.630 ;
        RECT 49.450 50.255 49.620 50.995 ;
        RECT 49.900 50.425 50.070 50.630 ;
        RECT 49.900 50.255 50.440 50.425 ;
        RECT 47.030 49.415 47.755 49.585 ;
        RECT 47.030 49.295 47.200 49.415 ;
        RECT 45.610 49.125 47.200 49.295 ;
        RECT 45.610 48.665 47.265 48.955 ;
        RECT 47.435 48.445 47.715 49.245 ;
        RECT 47.925 48.615 48.195 49.585 ;
        RECT 48.365 48.445 48.655 49.610 ;
        RECT 48.825 49.600 49.080 50.255 ;
        RECT 49.250 49.755 49.600 50.085 ;
        RECT 49.770 49.755 50.100 50.085 ;
        RECT 48.825 48.615 49.165 49.600 ;
        RECT 49.335 49.215 49.600 49.755 ;
        RECT 50.270 49.555 50.440 50.255 ;
        RECT 49.815 49.385 50.440 49.555 ;
        RECT 50.610 49.625 50.780 50.825 ;
        RECT 51.010 50.345 51.340 50.825 ;
        RECT 51.510 50.525 51.680 50.995 ;
        RECT 51.850 50.345 52.180 50.810 ;
        RECT 51.010 50.175 52.180 50.345 ;
        RECT 52.505 50.255 52.865 50.630 ;
        RECT 53.130 50.255 53.300 50.995 ;
        RECT 53.580 50.425 53.750 50.630 ;
        RECT 53.580 50.255 54.120 50.425 ;
        RECT 50.950 49.795 51.520 50.005 ;
        RECT 51.690 49.795 52.335 50.005 ;
        RECT 50.610 49.215 51.315 49.625 ;
        RECT 52.505 49.600 52.760 50.255 ;
        RECT 52.930 49.755 53.280 50.085 ;
        RECT 53.450 49.755 53.780 50.085 ;
        RECT 49.335 49.045 51.315 49.215 ;
        RECT 49.335 48.445 49.745 48.875 ;
        RECT 50.490 48.445 50.820 48.865 ;
        RECT 50.990 48.615 51.315 49.045 ;
        RECT 51.790 48.445 52.120 49.545 ;
        RECT 52.505 48.615 52.845 49.600 ;
        RECT 53.015 49.215 53.280 49.755 ;
        RECT 53.950 49.555 54.120 50.255 ;
        RECT 53.495 49.385 54.120 49.555 ;
        RECT 54.290 49.625 54.460 50.825 ;
        RECT 54.690 50.345 55.020 50.825 ;
        RECT 55.190 50.525 55.360 50.995 ;
        RECT 55.530 50.345 55.860 50.810 ;
        RECT 54.690 50.175 55.860 50.345 ;
        RECT 57.105 50.245 58.315 50.995 ;
        RECT 54.630 49.795 55.200 50.005 ;
        RECT 55.370 49.795 56.015 50.005 ;
        RECT 54.290 49.215 54.995 49.625 ;
        RECT 53.015 49.045 54.995 49.215 ;
        RECT 53.015 48.445 53.425 48.875 ;
        RECT 54.170 48.445 54.500 48.865 ;
        RECT 54.670 48.615 54.995 49.045 ;
        RECT 55.470 48.445 55.800 49.545 ;
        RECT 57.105 49.535 57.625 50.075 ;
        RECT 57.795 49.705 58.315 50.245 ;
        RECT 57.105 48.445 58.315 49.535 ;
        RECT 22.520 48.275 58.400 48.445 ;
        RECT 22.605 47.185 23.815 48.275 ;
        RECT 22.605 46.475 23.125 47.015 ;
        RECT 23.295 46.645 23.815 47.185 ;
        RECT 23.990 47.135 24.325 48.105 ;
        RECT 24.495 47.135 24.665 48.275 ;
        RECT 24.835 47.935 26.865 48.105 ;
        RECT 22.605 45.725 23.815 46.475 ;
        RECT 23.990 46.465 24.160 47.135 ;
        RECT 24.835 46.965 25.005 47.935 ;
        RECT 24.330 46.635 24.585 46.965 ;
        RECT 24.810 46.635 25.005 46.965 ;
        RECT 25.175 47.595 26.300 47.765 ;
        RECT 24.415 46.465 24.585 46.635 ;
        RECT 25.175 46.465 25.345 47.595 ;
        RECT 23.990 45.895 24.245 46.465 ;
        RECT 24.415 46.295 25.345 46.465 ;
        RECT 25.515 47.255 26.525 47.425 ;
        RECT 25.515 46.455 25.685 47.255 ;
        RECT 25.170 46.260 25.345 46.295 ;
        RECT 24.415 45.725 24.745 46.125 ;
        RECT 25.170 45.895 25.700 46.260 ;
        RECT 25.890 46.235 26.165 47.055 ;
        RECT 25.885 46.065 26.165 46.235 ;
        RECT 25.890 45.895 26.165 46.065 ;
        RECT 26.335 45.895 26.525 47.255 ;
        RECT 26.695 47.270 26.865 47.935 ;
        RECT 27.035 47.515 27.205 48.275 ;
        RECT 27.440 47.515 27.955 47.925 ;
        RECT 26.695 47.080 27.445 47.270 ;
        RECT 27.615 46.705 27.955 47.515 ;
        RECT 28.215 47.605 28.385 48.105 ;
        RECT 28.555 47.775 28.885 48.275 ;
        RECT 28.215 47.435 28.880 47.605 ;
        RECT 26.725 46.535 27.955 46.705 ;
        RECT 28.130 46.615 28.480 47.265 ;
        RECT 26.705 45.725 27.215 46.260 ;
        RECT 27.435 45.930 27.680 46.535 ;
        RECT 28.650 46.445 28.880 47.435 ;
        RECT 28.215 46.275 28.880 46.445 ;
        RECT 28.215 45.985 28.385 46.275 ;
        RECT 28.555 45.725 28.885 46.105 ;
        RECT 29.055 45.985 29.240 48.105 ;
        RECT 29.480 47.815 29.745 48.275 ;
        RECT 29.915 47.680 30.165 48.105 ;
        RECT 30.375 47.830 31.480 48.000 ;
        RECT 29.860 47.550 30.165 47.680 ;
        RECT 29.410 46.355 29.690 47.305 ;
        RECT 29.860 46.445 30.030 47.550 ;
        RECT 30.200 46.765 30.440 47.360 ;
        RECT 30.610 47.295 31.140 47.660 ;
        RECT 30.610 46.595 30.780 47.295 ;
        RECT 31.310 47.215 31.480 47.830 ;
        RECT 31.650 47.475 31.820 48.275 ;
        RECT 31.990 47.775 32.240 48.105 ;
        RECT 32.465 47.805 33.350 47.975 ;
        RECT 31.310 47.125 31.820 47.215 ;
        RECT 29.860 46.315 30.085 46.445 ;
        RECT 30.255 46.375 30.780 46.595 ;
        RECT 30.950 46.955 31.820 47.125 ;
        RECT 29.495 45.725 29.745 46.185 ;
        RECT 29.915 46.175 30.085 46.315 ;
        RECT 30.950 46.175 31.120 46.955 ;
        RECT 31.650 46.885 31.820 46.955 ;
        RECT 31.330 46.705 31.530 46.735 ;
        RECT 31.990 46.705 32.160 47.775 ;
        RECT 32.330 46.885 32.520 47.605 ;
        RECT 31.330 46.405 32.160 46.705 ;
        RECT 32.690 46.675 33.010 47.635 ;
        RECT 29.915 46.005 30.250 46.175 ;
        RECT 30.445 46.005 31.120 46.175 ;
        RECT 31.440 45.725 31.810 46.225 ;
        RECT 31.990 46.175 32.160 46.405 ;
        RECT 32.545 46.345 33.010 46.675 ;
        RECT 33.180 46.965 33.350 47.805 ;
        RECT 33.530 47.775 33.845 48.275 ;
        RECT 34.075 47.545 34.415 48.105 ;
        RECT 33.520 47.170 34.415 47.545 ;
        RECT 34.585 47.265 34.755 48.275 ;
        RECT 34.225 46.965 34.415 47.170 ;
        RECT 34.925 47.215 35.255 48.060 ;
        RECT 34.925 47.135 35.315 47.215 ;
        RECT 35.100 47.085 35.315 47.135 ;
        RECT 35.485 47.110 35.775 48.275 ;
        RECT 36.035 47.605 36.205 48.105 ;
        RECT 36.375 47.775 36.705 48.275 ;
        RECT 36.035 47.435 36.700 47.605 ;
        RECT 33.180 46.635 34.055 46.965 ;
        RECT 34.225 46.635 34.975 46.965 ;
        RECT 33.180 46.175 33.350 46.635 ;
        RECT 34.225 46.465 34.425 46.635 ;
        RECT 35.145 46.505 35.315 47.085 ;
        RECT 35.950 46.615 36.300 47.265 ;
        RECT 35.090 46.465 35.315 46.505 ;
        RECT 31.990 46.005 32.395 46.175 ;
        RECT 32.565 46.005 33.350 46.175 ;
        RECT 33.625 45.725 33.835 46.255 ;
        RECT 34.095 45.940 34.425 46.465 ;
        RECT 34.935 46.380 35.315 46.465 ;
        RECT 34.595 45.725 34.765 46.335 ;
        RECT 34.935 45.945 35.265 46.380 ;
        RECT 35.485 45.725 35.775 46.450 ;
        RECT 36.470 46.445 36.700 47.435 ;
        RECT 36.035 46.275 36.700 46.445 ;
        RECT 36.035 45.985 36.205 46.275 ;
        RECT 36.375 45.725 36.705 46.105 ;
        RECT 36.875 45.985 37.060 48.105 ;
        RECT 37.300 47.815 37.565 48.275 ;
        RECT 37.735 47.680 37.985 48.105 ;
        RECT 38.195 47.830 39.300 48.000 ;
        RECT 37.680 47.550 37.985 47.680 ;
        RECT 37.230 46.355 37.510 47.305 ;
        RECT 37.680 46.445 37.850 47.550 ;
        RECT 38.020 46.765 38.260 47.360 ;
        RECT 38.430 47.295 38.960 47.660 ;
        RECT 38.430 46.595 38.600 47.295 ;
        RECT 39.130 47.215 39.300 47.830 ;
        RECT 39.470 47.475 39.640 48.275 ;
        RECT 39.810 47.775 40.060 48.105 ;
        RECT 40.285 47.805 41.170 47.975 ;
        RECT 39.130 47.125 39.640 47.215 ;
        RECT 37.680 46.315 37.905 46.445 ;
        RECT 38.075 46.375 38.600 46.595 ;
        RECT 38.770 46.955 39.640 47.125 ;
        RECT 37.315 45.725 37.565 46.185 ;
        RECT 37.735 46.175 37.905 46.315 ;
        RECT 38.770 46.175 38.940 46.955 ;
        RECT 39.470 46.885 39.640 46.955 ;
        RECT 39.150 46.705 39.350 46.735 ;
        RECT 39.810 46.705 39.980 47.775 ;
        RECT 40.150 46.885 40.340 47.605 ;
        RECT 39.150 46.405 39.980 46.705 ;
        RECT 40.510 46.675 40.830 47.635 ;
        RECT 37.735 46.005 38.070 46.175 ;
        RECT 38.265 46.005 38.940 46.175 ;
        RECT 39.260 45.725 39.630 46.225 ;
        RECT 39.810 46.175 39.980 46.405 ;
        RECT 40.365 46.345 40.830 46.675 ;
        RECT 41.000 46.965 41.170 47.805 ;
        RECT 41.350 47.775 41.665 48.275 ;
        RECT 41.895 47.545 42.235 48.105 ;
        RECT 41.340 47.170 42.235 47.545 ;
        RECT 42.405 47.265 42.575 48.275 ;
        RECT 42.045 46.965 42.235 47.170 ;
        RECT 42.745 47.215 43.075 48.060 ;
        RECT 43.765 47.320 44.035 48.275 ;
        RECT 44.220 47.220 44.525 48.005 ;
        RECT 44.705 47.805 45.390 48.275 ;
        RECT 44.700 47.285 45.395 47.595 ;
        RECT 42.745 47.135 43.135 47.215 ;
        RECT 42.920 47.085 43.135 47.135 ;
        RECT 41.000 46.635 41.875 46.965 ;
        RECT 42.045 46.635 42.795 46.965 ;
        RECT 41.000 46.175 41.170 46.635 ;
        RECT 42.045 46.465 42.245 46.635 ;
        RECT 42.965 46.505 43.135 47.085 ;
        RECT 42.910 46.465 43.135 46.505 ;
        RECT 39.810 46.005 40.215 46.175 ;
        RECT 40.385 46.005 41.170 46.175 ;
        RECT 41.445 45.725 41.655 46.255 ;
        RECT 41.915 45.940 42.245 46.465 ;
        RECT 42.755 46.380 43.135 46.465 ;
        RECT 44.220 46.415 44.395 47.220 ;
        RECT 45.570 47.115 45.855 48.060 ;
        RECT 46.055 47.825 46.385 48.275 ;
        RECT 46.555 47.655 46.725 48.085 ;
        RECT 44.995 46.965 45.855 47.115 ;
        RECT 44.565 46.945 45.855 46.965 ;
        RECT 46.045 47.425 46.725 47.655 ;
        RECT 47.905 47.475 48.345 48.105 ;
        RECT 44.565 46.585 45.555 46.945 ;
        RECT 46.045 46.775 46.280 47.425 ;
        RECT 42.415 45.725 42.585 46.335 ;
        RECT 42.755 45.945 43.085 46.380 ;
        RECT 43.765 45.725 44.035 46.360 ;
        RECT 44.220 45.895 44.455 46.415 ;
        RECT 45.385 46.250 45.555 46.585 ;
        RECT 45.725 46.445 46.280 46.775 ;
        RECT 46.065 46.295 46.280 46.445 ;
        RECT 46.450 46.575 46.750 47.255 ;
        RECT 46.450 46.405 46.755 46.575 ;
        RECT 47.905 46.465 48.215 47.475 ;
        RECT 48.520 47.425 48.835 48.275 ;
        RECT 49.005 47.935 50.435 48.105 ;
        RECT 49.005 47.255 49.175 47.935 ;
        RECT 48.385 47.085 49.175 47.255 ;
        RECT 48.385 46.635 48.555 47.085 ;
        RECT 49.345 46.965 49.545 47.765 ;
        RECT 48.725 46.635 49.115 46.915 ;
        RECT 49.300 46.635 49.545 46.965 ;
        RECT 49.745 46.635 49.995 47.765 ;
        RECT 50.185 47.305 50.435 47.935 ;
        RECT 50.615 47.475 50.945 48.275 ;
        RECT 51.135 47.305 51.465 48.090 ;
        RECT 50.185 47.135 50.955 47.305 ;
        RECT 51.135 47.135 51.815 47.305 ;
        RECT 51.995 47.135 52.325 48.275 ;
        RECT 50.210 46.635 50.615 46.965 ;
        RECT 50.785 46.465 50.955 47.135 ;
        RECT 51.125 46.715 51.475 46.965 ;
        RECT 51.645 46.535 51.815 47.135 ;
        RECT 52.965 47.120 53.305 48.105 ;
        RECT 53.475 47.845 53.885 48.275 ;
        RECT 54.630 47.855 54.960 48.275 ;
        RECT 55.130 47.675 55.455 48.105 ;
        RECT 53.475 47.505 55.455 47.675 ;
        RECT 51.985 46.715 52.335 46.965 ;
        RECT 44.625 45.725 45.025 46.220 ;
        RECT 45.385 46.055 45.785 46.250 ;
        RECT 45.615 45.910 45.785 46.055 ;
        RECT 46.065 45.920 46.305 46.295 ;
        RECT 46.475 45.725 46.805 46.230 ;
        RECT 47.905 45.905 48.345 46.465 ;
        RECT 48.515 45.725 48.965 46.465 ;
        RECT 49.135 46.295 50.295 46.465 ;
        RECT 49.135 45.895 49.305 46.295 ;
        RECT 49.475 45.725 49.895 46.125 ;
        RECT 50.065 45.895 50.295 46.295 ;
        RECT 50.465 45.895 50.955 46.465 ;
        RECT 51.145 45.725 51.385 46.535 ;
        RECT 51.555 45.895 51.885 46.535 ;
        RECT 52.055 45.725 52.325 46.535 ;
        RECT 52.965 46.465 53.220 47.120 ;
        RECT 53.475 46.965 53.740 47.505 ;
        RECT 53.955 47.165 54.580 47.335 ;
        RECT 53.390 46.635 53.740 46.965 ;
        RECT 53.910 46.635 54.240 46.965 ;
        RECT 54.410 46.465 54.580 47.165 ;
        RECT 52.965 46.090 53.325 46.465 ;
        RECT 53.590 45.725 53.760 46.465 ;
        RECT 54.040 46.295 54.580 46.465 ;
        RECT 54.750 47.095 55.455 47.505 ;
        RECT 55.930 47.175 56.260 48.275 ;
        RECT 57.105 47.185 58.315 48.275 ;
        RECT 54.040 46.090 54.210 46.295 ;
        RECT 54.750 45.895 54.920 47.095 ;
        RECT 55.090 46.715 55.660 46.925 ;
        RECT 55.830 46.715 56.475 46.925 ;
        RECT 57.105 46.645 57.625 47.185 ;
        RECT 55.150 46.375 56.320 46.545 ;
        RECT 57.795 46.475 58.315 47.015 ;
        RECT 55.150 45.895 55.480 46.375 ;
        RECT 55.650 45.725 55.820 46.195 ;
        RECT 55.990 45.910 56.320 46.375 ;
        RECT 57.105 45.725 58.315 46.475 ;
        RECT 75.000 46.625 75.885 51.885 ;
        RECT 76.565 51.315 78.605 51.485 ;
        RECT 76.225 47.255 76.395 51.255 ;
        RECT 78.775 47.255 78.945 51.255 ;
        RECT 76.565 47.025 78.605 47.195 ;
        RECT 79.285 46.625 79.455 51.885 ;
        RECT 80.195 53.855 90.580 54.025 ;
        RECT 80.195 50.595 80.365 53.855 ;
        RECT 81.090 53.285 89.130 53.455 ;
        RECT 80.705 51.225 80.875 53.225 ;
        RECT 89.345 51.225 89.515 53.225 ;
        RECT 81.090 50.995 89.130 51.165 ;
        RECT 89.855 50.595 90.580 53.855 ;
        RECT 80.195 50.425 90.580 50.595 ;
        RECT 80.195 47.165 80.365 50.425 ;
        RECT 81.090 49.855 89.130 50.025 ;
        RECT 80.705 47.795 80.875 49.795 ;
        RECT 89.345 47.795 89.515 49.795 ;
        RECT 81.090 47.565 89.130 47.735 ;
        RECT 89.855 47.165 90.580 50.425 ;
        RECT 80.195 46.995 90.580 47.165 ;
        RECT 85.905 46.715 90.580 46.995 ;
        RECT 75.000 46.455 79.455 46.625 ;
        RECT 22.520 45.555 58.400 45.725 ;
        RECT 22.605 44.805 23.815 45.555 ;
        RECT 24.035 44.900 24.365 45.335 ;
        RECT 24.535 44.945 24.705 45.555 ;
        RECT 23.985 44.815 24.365 44.900 ;
        RECT 24.875 44.815 25.205 45.340 ;
        RECT 25.465 45.025 25.675 45.555 ;
        RECT 25.950 45.105 26.735 45.275 ;
        RECT 26.905 45.105 27.310 45.275 ;
        RECT 22.605 44.265 23.125 44.805 ;
        RECT 23.985 44.775 24.210 44.815 ;
        RECT 23.295 44.095 23.815 44.635 ;
        RECT 22.605 43.005 23.815 44.095 ;
        RECT 23.985 44.195 24.155 44.775 ;
        RECT 24.875 44.645 25.075 44.815 ;
        RECT 25.950 44.645 26.120 45.105 ;
        RECT 24.325 44.315 25.075 44.645 ;
        RECT 25.245 44.315 26.120 44.645 ;
        RECT 23.985 44.145 24.200 44.195 ;
        RECT 23.985 44.065 24.375 44.145 ;
        RECT 24.045 43.220 24.375 44.065 ;
        RECT 24.885 44.110 25.075 44.315 ;
        RECT 24.545 43.005 24.715 44.015 ;
        RECT 24.885 43.735 25.780 44.110 ;
        RECT 24.885 43.175 25.225 43.735 ;
        RECT 25.455 43.005 25.770 43.505 ;
        RECT 25.950 43.475 26.120 44.315 ;
        RECT 26.290 44.605 26.755 44.935 ;
        RECT 27.140 44.875 27.310 45.105 ;
        RECT 27.490 45.055 27.860 45.555 ;
        RECT 28.180 45.105 28.855 45.275 ;
        RECT 29.050 45.105 29.385 45.275 ;
        RECT 26.290 43.645 26.610 44.605 ;
        RECT 27.140 44.575 27.970 44.875 ;
        RECT 26.780 43.675 26.970 44.395 ;
        RECT 27.140 43.505 27.310 44.575 ;
        RECT 27.770 44.545 27.970 44.575 ;
        RECT 27.480 44.325 27.650 44.395 ;
        RECT 28.180 44.325 28.350 45.105 ;
        RECT 29.215 44.965 29.385 45.105 ;
        RECT 29.555 45.095 29.805 45.555 ;
        RECT 27.480 44.155 28.350 44.325 ;
        RECT 28.520 44.685 29.045 44.905 ;
        RECT 29.215 44.835 29.440 44.965 ;
        RECT 27.480 44.065 27.990 44.155 ;
        RECT 25.950 43.305 26.835 43.475 ;
        RECT 27.060 43.175 27.310 43.505 ;
        RECT 27.480 43.005 27.650 43.805 ;
        RECT 27.820 43.450 27.990 44.065 ;
        RECT 28.520 43.985 28.690 44.685 ;
        RECT 28.160 43.620 28.690 43.985 ;
        RECT 28.860 43.920 29.100 44.515 ;
        RECT 29.270 43.730 29.440 44.835 ;
        RECT 29.610 43.975 29.890 44.925 ;
        RECT 29.135 43.600 29.440 43.730 ;
        RECT 27.820 43.280 28.925 43.450 ;
        RECT 29.135 43.175 29.385 43.600 ;
        RECT 29.555 43.005 29.820 43.465 ;
        RECT 30.060 43.175 30.245 45.295 ;
        RECT 30.415 45.175 30.745 45.555 ;
        RECT 30.915 45.005 31.085 45.295 ;
        RECT 30.420 44.835 31.085 45.005 ;
        RECT 30.420 43.845 30.650 44.835 ;
        RECT 31.345 44.785 33.935 45.555 ;
        RECT 34.565 45.045 34.870 45.555 ;
        RECT 30.820 44.015 31.170 44.665 ;
        RECT 31.345 44.265 32.555 44.785 ;
        RECT 32.725 44.095 33.935 44.615 ;
        RECT 34.565 44.315 34.880 44.875 ;
        RECT 35.050 44.565 35.300 45.375 ;
        RECT 35.470 45.030 35.730 45.555 ;
        RECT 35.910 44.565 36.160 45.375 ;
        RECT 36.330 44.995 36.590 45.555 ;
        RECT 36.760 44.905 37.020 45.360 ;
        RECT 37.190 45.075 37.450 45.555 ;
        RECT 37.620 44.905 37.880 45.360 ;
        RECT 38.050 45.075 38.310 45.555 ;
        RECT 38.480 44.905 38.740 45.360 ;
        RECT 38.910 45.075 39.155 45.555 ;
        RECT 39.325 44.905 39.600 45.360 ;
        RECT 39.770 45.075 40.015 45.555 ;
        RECT 40.185 44.905 40.445 45.360 ;
        RECT 40.625 45.075 40.875 45.555 ;
        RECT 41.045 44.905 41.305 45.360 ;
        RECT 41.485 45.075 41.735 45.555 ;
        RECT 41.905 44.905 42.165 45.360 ;
        RECT 42.345 45.075 42.605 45.555 ;
        RECT 42.775 44.905 43.035 45.360 ;
        RECT 43.205 45.075 43.505 45.555 ;
        RECT 36.760 44.735 43.505 44.905 ;
        RECT 35.050 44.315 42.170 44.565 ;
        RECT 30.420 43.675 31.085 43.845 ;
        RECT 30.415 43.005 30.745 43.505 ;
        RECT 30.915 43.175 31.085 43.675 ;
        RECT 31.345 43.005 33.935 44.095 ;
        RECT 34.575 43.005 34.870 43.815 ;
        RECT 35.050 43.175 35.295 44.315 ;
        RECT 35.470 43.005 35.730 43.815 ;
        RECT 35.910 43.180 36.160 44.315 ;
        RECT 42.340 44.145 43.505 44.735 ;
        RECT 36.760 43.920 43.505 44.145 ;
        RECT 43.765 44.815 44.150 45.385 ;
        RECT 44.320 45.095 44.645 45.555 ;
        RECT 45.165 44.925 45.445 45.385 ;
        RECT 43.765 44.145 44.045 44.815 ;
        RECT 44.320 44.755 45.445 44.925 ;
        RECT 44.320 44.645 44.770 44.755 ;
        RECT 44.215 44.315 44.770 44.645 ;
        RECT 45.635 44.585 46.035 45.385 ;
        RECT 46.435 45.095 46.705 45.555 ;
        RECT 46.875 44.925 47.160 45.385 ;
        RECT 36.760 43.905 42.165 43.920 ;
        RECT 36.330 43.010 36.590 43.805 ;
        RECT 36.760 43.180 37.020 43.905 ;
        RECT 37.190 43.010 37.450 43.735 ;
        RECT 37.620 43.180 37.880 43.905 ;
        RECT 38.050 43.010 38.310 43.735 ;
        RECT 38.480 43.180 38.740 43.905 ;
        RECT 38.910 43.010 39.170 43.735 ;
        RECT 39.340 43.180 39.600 43.905 ;
        RECT 39.770 43.010 40.015 43.735 ;
        RECT 40.185 43.180 40.445 43.905 ;
        RECT 40.630 43.010 40.875 43.735 ;
        RECT 41.045 43.180 41.305 43.905 ;
        RECT 41.490 43.010 41.735 43.735 ;
        RECT 41.905 43.180 42.165 43.905 ;
        RECT 42.350 43.010 42.605 43.735 ;
        RECT 42.775 43.180 43.065 43.920 ;
        RECT 36.330 43.005 42.605 43.010 ;
        RECT 43.235 43.005 43.505 43.750 ;
        RECT 43.765 43.175 44.150 44.145 ;
        RECT 44.320 43.855 44.770 44.315 ;
        RECT 44.940 44.025 46.035 44.585 ;
        RECT 44.320 43.635 45.445 43.855 ;
        RECT 44.320 43.005 44.645 43.465 ;
        RECT 45.165 43.175 45.445 43.635 ;
        RECT 45.635 43.175 46.035 44.025 ;
        RECT 46.205 44.755 47.160 44.925 ;
        RECT 48.365 44.830 48.655 45.555 ;
        RECT 48.840 44.985 49.095 45.335 ;
        RECT 49.265 45.155 49.595 45.555 ;
        RECT 49.765 44.985 49.935 45.335 ;
        RECT 50.105 45.155 50.485 45.555 ;
        RECT 48.840 44.815 50.505 44.985 ;
        RECT 50.675 44.880 50.950 45.225 ;
        RECT 46.205 43.855 46.415 44.755 ;
        RECT 50.335 44.645 50.505 44.815 ;
        RECT 46.585 44.025 47.275 44.585 ;
        RECT 48.825 44.315 49.170 44.645 ;
        RECT 49.340 44.315 50.165 44.645 ;
        RECT 50.335 44.315 50.610 44.645 ;
        RECT 46.205 43.635 47.160 43.855 ;
        RECT 46.435 43.005 46.705 43.465 ;
        RECT 46.875 43.175 47.160 43.635 ;
        RECT 48.365 43.005 48.655 44.170 ;
        RECT 48.845 43.855 49.170 44.145 ;
        RECT 49.340 44.025 49.535 44.315 ;
        RECT 50.335 44.145 50.505 44.315 ;
        RECT 50.780 44.145 50.950 44.880 ;
        RECT 51.125 44.785 53.715 45.555 ;
        RECT 51.125 44.265 52.335 44.785 ;
        RECT 54.355 44.745 54.625 45.555 ;
        RECT 54.795 44.745 55.125 45.385 ;
        RECT 55.295 44.745 55.535 45.555 ;
        RECT 55.725 44.880 55.985 45.385 ;
        RECT 56.165 45.175 56.495 45.555 ;
        RECT 56.675 45.005 56.845 45.385 ;
        RECT 49.845 43.975 50.505 44.145 ;
        RECT 49.845 43.855 50.015 43.975 ;
        RECT 48.845 43.685 50.015 43.855 ;
        RECT 48.825 43.225 50.015 43.515 ;
        RECT 50.185 43.005 50.465 43.805 ;
        RECT 50.675 43.175 50.950 44.145 ;
        RECT 52.505 44.095 53.715 44.615 ;
        RECT 54.345 44.315 54.695 44.565 ;
        RECT 54.865 44.145 55.035 44.745 ;
        RECT 55.205 44.315 55.555 44.565 ;
        RECT 51.125 43.005 53.715 44.095 ;
        RECT 54.355 43.005 54.685 44.145 ;
        RECT 54.865 43.975 55.545 44.145 ;
        RECT 55.215 43.190 55.545 43.975 ;
        RECT 55.725 44.080 55.895 44.880 ;
        RECT 56.180 44.835 56.845 45.005 ;
        RECT 56.180 44.580 56.350 44.835 ;
        RECT 57.105 44.805 58.315 45.555 ;
        RECT 56.065 44.250 56.350 44.580 ;
        RECT 56.585 44.285 56.915 44.655 ;
        RECT 56.180 44.105 56.350 44.250 ;
        RECT 55.725 43.175 55.995 44.080 ;
        RECT 56.180 43.935 56.845 44.105 ;
        RECT 56.165 43.005 56.495 43.765 ;
        RECT 56.675 43.175 56.845 43.935 ;
        RECT 57.105 44.095 57.625 44.635 ;
        RECT 57.795 44.265 58.315 44.805 ;
        RECT 57.105 43.005 58.315 44.095 ;
        RECT 22.520 42.835 58.400 43.005 ;
        RECT 22.605 41.745 23.815 42.835 ;
        RECT 23.985 41.745 25.195 42.835 ;
        RECT 25.480 42.205 25.765 42.665 ;
        RECT 25.935 42.375 26.205 42.835 ;
        RECT 25.480 41.985 26.435 42.205 ;
        RECT 22.605 41.035 23.125 41.575 ;
        RECT 23.295 41.205 23.815 41.745 ;
        RECT 23.985 41.035 24.505 41.575 ;
        RECT 24.675 41.205 25.195 41.745 ;
        RECT 25.365 41.255 26.055 41.815 ;
        RECT 26.225 41.085 26.435 41.985 ;
        RECT 22.605 40.285 23.815 41.035 ;
        RECT 23.985 40.285 25.195 41.035 ;
        RECT 25.480 40.915 26.435 41.085 ;
        RECT 26.605 41.815 27.005 42.665 ;
        RECT 27.195 42.205 27.475 42.665 ;
        RECT 27.995 42.375 28.320 42.835 ;
        RECT 27.195 41.985 28.320 42.205 ;
        RECT 26.605 41.255 27.700 41.815 ;
        RECT 27.870 41.525 28.320 41.985 ;
        RECT 28.490 41.695 28.875 42.665 ;
        RECT 25.480 40.455 25.765 40.915 ;
        RECT 25.935 40.285 26.205 40.745 ;
        RECT 26.605 40.455 27.005 41.255 ;
        RECT 27.870 41.195 28.425 41.525 ;
        RECT 27.870 41.085 28.320 41.195 ;
        RECT 27.195 40.915 28.320 41.085 ;
        RECT 28.595 41.025 28.875 41.695 ;
        RECT 27.195 40.455 27.475 40.915 ;
        RECT 27.995 40.285 28.320 40.745 ;
        RECT 28.490 40.455 28.875 41.025 ;
        RECT 29.045 41.695 29.430 42.665 ;
        RECT 29.600 42.375 29.925 42.835 ;
        RECT 30.445 42.205 30.725 42.665 ;
        RECT 29.600 41.985 30.725 42.205 ;
        RECT 29.045 41.025 29.325 41.695 ;
        RECT 29.600 41.525 30.050 41.985 ;
        RECT 30.915 41.815 31.315 42.665 ;
        RECT 31.715 42.375 31.985 42.835 ;
        RECT 32.155 42.205 32.440 42.665 ;
        RECT 29.495 41.195 30.050 41.525 ;
        RECT 30.220 41.255 31.315 41.815 ;
        RECT 29.600 41.085 30.050 41.195 ;
        RECT 29.045 40.455 29.430 41.025 ;
        RECT 29.600 40.915 30.725 41.085 ;
        RECT 29.600 40.285 29.925 40.745 ;
        RECT 30.445 40.455 30.725 40.915 ;
        RECT 30.915 40.455 31.315 41.255 ;
        RECT 31.485 41.985 32.440 42.205 ;
        RECT 31.485 41.085 31.695 41.985 ;
        RECT 31.865 41.255 32.555 41.815 ;
        RECT 32.725 41.745 35.315 42.835 ;
        RECT 31.485 40.915 32.440 41.085 ;
        RECT 31.715 40.285 31.985 40.745 ;
        RECT 32.155 40.455 32.440 40.915 ;
        RECT 32.725 41.055 33.935 41.575 ;
        RECT 34.105 41.225 35.315 41.745 ;
        RECT 35.485 41.670 35.775 42.835 ;
        RECT 35.955 41.695 36.285 42.835 ;
        RECT 36.815 41.865 37.145 42.650 ;
        RECT 36.465 41.695 37.145 41.865 ;
        RECT 37.445 41.715 37.775 42.835 ;
        RECT 35.945 41.275 36.295 41.525 ;
        RECT 36.465 41.095 36.635 41.695 ;
        RECT 36.805 41.275 37.155 41.525 ;
        RECT 37.385 41.275 37.895 41.525 ;
        RECT 38.105 41.275 38.475 42.590 ;
        RECT 38.645 41.275 38.975 42.590 ;
        RECT 39.185 41.275 39.515 42.590 ;
        RECT 39.785 41.945 40.035 42.665 ;
        RECT 40.205 42.115 40.535 42.835 ;
        RECT 39.785 41.655 40.535 41.945 ;
        RECT 40.770 41.655 41.295 42.665 ;
        RECT 40.275 41.485 40.535 41.655 ;
        RECT 39.685 41.275 40.105 41.485 ;
        RECT 40.275 41.275 40.855 41.485 ;
        RECT 40.275 41.105 40.645 41.275 ;
        RECT 32.725 40.285 35.315 41.055 ;
        RECT 35.485 40.285 35.775 41.010 ;
        RECT 35.955 40.285 36.225 41.095 ;
        RECT 36.395 40.455 36.725 41.095 ;
        RECT 36.895 40.285 37.135 41.095 ;
        RECT 37.425 40.935 39.725 41.105 ;
        RECT 37.425 40.455 37.755 40.935 ;
        RECT 37.925 40.285 38.255 40.745 ;
        RECT 38.470 40.455 38.800 40.935 ;
        RECT 39.000 40.285 39.330 40.745 ;
        RECT 39.555 40.615 39.725 40.935 ;
        RECT 39.895 40.915 40.645 41.105 ;
        RECT 41.025 41.085 41.295 41.655 ;
        RECT 39.895 40.470 40.225 40.915 ;
        RECT 40.495 40.285 40.665 40.745 ;
        RECT 40.955 40.455 41.295 41.085 ;
        RECT 41.465 41.695 41.850 42.665 ;
        RECT 42.020 42.375 42.345 42.835 ;
        RECT 42.865 42.205 43.145 42.665 ;
        RECT 42.020 41.985 43.145 42.205 ;
        RECT 41.465 41.025 41.745 41.695 ;
        RECT 42.020 41.525 42.470 41.985 ;
        RECT 43.335 41.815 43.735 42.665 ;
        RECT 44.135 42.375 44.405 42.835 ;
        RECT 44.575 42.205 44.860 42.665 ;
        RECT 41.915 41.195 42.470 41.525 ;
        RECT 42.640 41.255 43.735 41.815 ;
        RECT 42.020 41.085 42.470 41.195 ;
        RECT 41.465 40.455 41.850 41.025 ;
        RECT 42.020 40.915 43.145 41.085 ;
        RECT 42.020 40.285 42.345 40.745 ;
        RECT 42.865 40.455 43.145 40.915 ;
        RECT 43.335 40.455 43.735 41.255 ;
        RECT 43.905 41.985 44.860 42.205 ;
        RECT 43.905 41.085 44.115 41.985 ;
        RECT 44.285 41.255 44.975 41.815 ;
        RECT 45.145 41.745 46.355 42.835 ;
        RECT 43.905 40.915 44.860 41.085 ;
        RECT 44.135 40.285 44.405 40.745 ;
        RECT 44.575 40.455 44.860 40.915 ;
        RECT 45.145 41.035 45.665 41.575 ;
        RECT 45.835 41.205 46.355 41.745 ;
        RECT 46.525 41.695 46.800 42.665 ;
        RECT 47.010 42.035 47.290 42.835 ;
        RECT 47.460 42.325 49.510 42.615 ;
        RECT 47.460 41.985 49.090 42.155 ;
        RECT 47.460 41.865 47.630 41.985 ;
        RECT 46.970 41.695 47.630 41.865 ;
        RECT 45.145 40.285 46.355 41.035 ;
        RECT 46.525 40.960 46.695 41.695 ;
        RECT 46.970 41.525 47.140 41.695 ;
        RECT 46.865 41.195 47.140 41.525 ;
        RECT 47.310 41.195 47.690 41.525 ;
        RECT 47.860 41.195 48.600 41.815 ;
        RECT 48.770 41.695 49.090 41.985 ;
        RECT 49.285 41.525 49.525 42.120 ;
        RECT 49.695 41.760 50.035 42.835 ;
        RECT 50.215 41.865 50.545 42.650 ;
        RECT 50.215 41.695 50.895 41.865 ;
        RECT 51.075 41.695 51.405 42.835 ;
        RECT 51.665 41.905 51.845 42.665 ;
        RECT 52.025 42.075 52.355 42.835 ;
        RECT 51.665 41.735 52.340 41.905 ;
        RECT 52.525 41.760 52.795 42.665 ;
        RECT 48.870 41.195 49.525 41.525 ;
        RECT 46.970 41.025 47.140 41.195 ;
        RECT 46.525 40.615 46.800 40.960 ;
        RECT 46.970 40.855 48.555 41.025 ;
        RECT 46.990 40.285 47.370 40.685 ;
        RECT 47.540 40.505 47.710 40.855 ;
        RECT 47.880 40.285 48.210 40.685 ;
        RECT 48.385 40.505 48.555 40.855 ;
        RECT 48.755 40.285 49.085 40.785 ;
        RECT 49.280 40.505 49.525 41.195 ;
        RECT 49.695 40.955 50.035 41.525 ;
        RECT 50.205 41.275 50.555 41.525 ;
        RECT 50.725 41.095 50.895 41.695 ;
        RECT 52.170 41.590 52.340 41.735 ;
        RECT 51.065 41.275 51.415 41.525 ;
        RECT 51.605 41.185 51.945 41.555 ;
        RECT 52.170 41.260 52.445 41.590 ;
        RECT 49.695 40.285 50.035 40.785 ;
        RECT 50.225 40.285 50.465 41.095 ;
        RECT 50.635 40.455 50.965 41.095 ;
        RECT 51.135 40.285 51.405 41.095 ;
        RECT 52.170 41.005 52.340 41.260 ;
        RECT 51.675 40.835 52.340 41.005 ;
        RECT 52.615 40.960 52.795 41.760 ;
        RECT 53.180 41.735 53.510 42.835 ;
        RECT 53.985 42.235 54.310 42.665 ;
        RECT 54.480 42.415 54.810 42.835 ;
        RECT 55.555 42.405 55.965 42.835 ;
        RECT 53.985 42.065 55.965 42.235 ;
        RECT 53.985 41.655 54.690 42.065 ;
        RECT 52.965 41.275 53.610 41.485 ;
        RECT 53.780 41.275 54.350 41.485 ;
        RECT 51.675 40.455 51.845 40.835 ;
        RECT 52.025 40.285 52.355 40.665 ;
        RECT 52.535 40.455 52.795 40.960 ;
        RECT 53.120 40.935 54.290 41.105 ;
        RECT 53.120 40.470 53.450 40.935 ;
        RECT 53.620 40.285 53.790 40.755 ;
        RECT 53.960 40.455 54.290 40.935 ;
        RECT 54.520 40.455 54.690 41.655 ;
        RECT 54.860 41.725 55.485 41.895 ;
        RECT 54.860 41.025 55.030 41.725 ;
        RECT 55.700 41.525 55.965 42.065 ;
        RECT 56.135 41.680 56.475 42.665 ;
        RECT 55.200 41.195 55.530 41.525 ;
        RECT 55.700 41.195 56.050 41.525 ;
        RECT 56.220 41.025 56.475 41.680 ;
        RECT 57.105 41.745 58.315 42.835 ;
        RECT 57.105 41.205 57.625 41.745 ;
        RECT 57.795 41.035 58.315 41.575 ;
        RECT 54.860 40.855 55.400 41.025 ;
        RECT 55.230 40.650 55.400 40.855 ;
        RECT 55.680 40.285 55.850 41.025 ;
        RECT 56.115 40.650 56.475 41.025 ;
        RECT 57.105 40.285 58.315 41.035 ;
        RECT 75.000 41.195 75.885 46.455 ;
        RECT 76.565 45.885 78.605 46.055 ;
        RECT 76.225 41.825 76.395 45.825 ;
        RECT 78.775 41.825 78.945 45.825 ;
        RECT 76.565 41.595 78.605 41.765 ;
        RECT 79.285 41.195 79.455 46.455 ;
        RECT 75.000 41.025 79.455 41.195 ;
        RECT 22.520 40.115 58.400 40.285 ;
        RECT 22.605 39.365 23.815 40.115 ;
        RECT 22.605 38.825 23.125 39.365 ;
        RECT 23.990 39.275 24.250 40.115 ;
        RECT 24.425 39.370 24.680 39.945 ;
        RECT 24.850 39.735 25.180 40.115 ;
        RECT 25.395 39.565 25.565 39.945 ;
        RECT 24.850 39.395 25.565 39.565 ;
        RECT 23.295 38.655 23.815 39.195 ;
        RECT 22.605 37.565 23.815 38.655 ;
        RECT 23.990 37.565 24.250 38.715 ;
        RECT 24.425 38.640 24.595 39.370 ;
        RECT 24.850 39.205 25.020 39.395 ;
        RECT 26.290 39.375 26.545 39.945 ;
        RECT 26.715 39.715 27.045 40.115 ;
        RECT 27.470 39.580 28.000 39.945 ;
        RECT 28.190 39.775 28.465 39.945 ;
        RECT 28.185 39.605 28.465 39.775 ;
        RECT 27.470 39.545 27.645 39.580 ;
        RECT 26.715 39.375 27.645 39.545 ;
        RECT 24.765 38.875 25.020 39.205 ;
        RECT 24.850 38.665 25.020 38.875 ;
        RECT 25.300 38.845 25.655 39.215 ;
        RECT 26.290 38.705 26.460 39.375 ;
        RECT 26.715 39.205 26.885 39.375 ;
        RECT 26.630 38.875 26.885 39.205 ;
        RECT 27.110 38.875 27.305 39.205 ;
        RECT 24.425 37.735 24.680 38.640 ;
        RECT 24.850 38.495 25.565 38.665 ;
        RECT 24.850 37.565 25.180 38.325 ;
        RECT 25.395 37.735 25.565 38.495 ;
        RECT 26.290 37.735 26.625 38.705 ;
        RECT 26.795 37.565 26.965 38.705 ;
        RECT 27.135 37.905 27.305 38.875 ;
        RECT 27.475 38.245 27.645 39.375 ;
        RECT 27.815 38.585 27.985 39.385 ;
        RECT 28.190 38.785 28.465 39.605 ;
        RECT 28.635 38.585 28.825 39.945 ;
        RECT 29.005 39.580 29.515 40.115 ;
        RECT 29.735 39.305 29.980 39.910 ;
        RECT 30.515 39.565 30.685 39.855 ;
        RECT 30.855 39.735 31.185 40.115 ;
        RECT 30.515 39.395 31.180 39.565 ;
        RECT 29.025 39.135 30.255 39.305 ;
        RECT 27.815 38.415 28.825 38.585 ;
        RECT 28.995 38.570 29.745 38.760 ;
        RECT 27.475 38.075 28.600 38.245 ;
        RECT 28.995 37.905 29.165 38.570 ;
        RECT 29.915 38.325 30.255 39.135 ;
        RECT 30.430 38.575 30.780 39.225 ;
        RECT 30.950 38.405 31.180 39.395 ;
        RECT 27.135 37.735 29.165 37.905 ;
        RECT 29.335 37.565 29.505 38.325 ;
        RECT 29.740 37.915 30.255 38.325 ;
        RECT 30.515 38.235 31.180 38.405 ;
        RECT 30.515 37.735 30.685 38.235 ;
        RECT 30.855 37.565 31.185 38.065 ;
        RECT 31.355 37.735 31.540 39.855 ;
        RECT 31.795 39.655 32.045 40.115 ;
        RECT 32.215 39.665 32.550 39.835 ;
        RECT 32.745 39.665 33.420 39.835 ;
        RECT 32.215 39.525 32.385 39.665 ;
        RECT 31.710 38.535 31.990 39.485 ;
        RECT 32.160 39.395 32.385 39.525 ;
        RECT 32.160 38.290 32.330 39.395 ;
        RECT 32.555 39.245 33.080 39.465 ;
        RECT 32.500 38.480 32.740 39.075 ;
        RECT 32.910 38.545 33.080 39.245 ;
        RECT 33.250 38.885 33.420 39.665 ;
        RECT 33.740 39.615 34.110 40.115 ;
        RECT 34.290 39.665 34.695 39.835 ;
        RECT 34.865 39.665 35.650 39.835 ;
        RECT 34.290 39.435 34.460 39.665 ;
        RECT 33.630 39.135 34.460 39.435 ;
        RECT 34.845 39.165 35.310 39.495 ;
        RECT 33.630 39.105 33.830 39.135 ;
        RECT 33.950 38.885 34.120 38.955 ;
        RECT 33.250 38.715 34.120 38.885 ;
        RECT 33.610 38.625 34.120 38.715 ;
        RECT 32.160 38.160 32.465 38.290 ;
        RECT 32.910 38.180 33.440 38.545 ;
        RECT 31.780 37.565 32.045 38.025 ;
        RECT 32.215 37.735 32.465 38.160 ;
        RECT 33.610 38.010 33.780 38.625 ;
        RECT 32.675 37.840 33.780 38.010 ;
        RECT 33.950 37.565 34.120 38.365 ;
        RECT 34.290 38.065 34.460 39.135 ;
        RECT 34.630 38.235 34.820 38.955 ;
        RECT 34.990 38.205 35.310 39.165 ;
        RECT 35.480 39.205 35.650 39.665 ;
        RECT 35.925 39.585 36.135 40.115 ;
        RECT 36.395 39.375 36.725 39.900 ;
        RECT 36.895 39.505 37.065 40.115 ;
        RECT 37.235 39.460 37.565 39.895 ;
        RECT 37.235 39.375 37.615 39.460 ;
        RECT 36.525 39.205 36.725 39.375 ;
        RECT 37.390 39.335 37.615 39.375 ;
        RECT 35.480 38.875 36.355 39.205 ;
        RECT 36.525 38.875 37.275 39.205 ;
        RECT 34.290 37.735 34.540 38.065 ;
        RECT 35.480 38.035 35.650 38.875 ;
        RECT 36.525 38.670 36.715 38.875 ;
        RECT 37.445 38.755 37.615 39.335 ;
        RECT 37.400 38.705 37.615 38.755 ;
        RECT 35.820 38.295 36.715 38.670 ;
        RECT 37.225 38.625 37.615 38.705 ;
        RECT 37.790 39.375 38.045 39.945 ;
        RECT 38.215 39.715 38.545 40.115 ;
        RECT 38.970 39.580 39.500 39.945 ;
        RECT 38.970 39.545 39.145 39.580 ;
        RECT 38.215 39.375 39.145 39.545 ;
        RECT 37.790 38.705 37.960 39.375 ;
        RECT 38.215 39.205 38.385 39.375 ;
        RECT 38.130 38.875 38.385 39.205 ;
        RECT 38.610 38.875 38.805 39.205 ;
        RECT 34.765 37.865 35.650 38.035 ;
        RECT 35.830 37.565 36.145 38.065 ;
        RECT 36.375 37.735 36.715 38.295 ;
        RECT 36.885 37.565 37.055 38.575 ;
        RECT 37.225 37.780 37.555 38.625 ;
        RECT 37.790 37.735 38.125 38.705 ;
        RECT 38.295 37.565 38.465 38.705 ;
        RECT 38.635 37.905 38.805 38.875 ;
        RECT 38.975 38.245 39.145 39.375 ;
        RECT 39.315 38.585 39.485 39.385 ;
        RECT 39.690 39.095 39.965 39.945 ;
        RECT 39.685 38.925 39.965 39.095 ;
        RECT 39.690 38.785 39.965 38.925 ;
        RECT 40.135 38.585 40.325 39.945 ;
        RECT 40.505 39.580 41.015 40.115 ;
        RECT 41.235 39.305 41.480 39.910 ;
        RECT 41.925 39.375 42.310 39.945 ;
        RECT 42.480 39.655 42.805 40.115 ;
        RECT 43.325 39.485 43.605 39.945 ;
        RECT 40.525 39.135 41.755 39.305 ;
        RECT 39.315 38.415 40.325 38.585 ;
        RECT 40.495 38.570 41.245 38.760 ;
        RECT 38.975 38.075 40.100 38.245 ;
        RECT 40.495 37.905 40.665 38.570 ;
        RECT 41.415 38.325 41.755 39.135 ;
        RECT 38.635 37.735 40.665 37.905 ;
        RECT 40.835 37.565 41.005 38.325 ;
        RECT 41.240 37.915 41.755 38.325 ;
        RECT 41.925 38.705 42.205 39.375 ;
        RECT 42.480 39.315 43.605 39.485 ;
        RECT 42.480 39.205 42.930 39.315 ;
        RECT 42.375 38.875 42.930 39.205 ;
        RECT 43.795 39.145 44.195 39.945 ;
        RECT 44.595 39.655 44.865 40.115 ;
        RECT 45.035 39.485 45.320 39.945 ;
        RECT 41.925 37.735 42.310 38.705 ;
        RECT 42.480 38.415 42.930 38.875 ;
        RECT 43.100 38.585 44.195 39.145 ;
        RECT 42.480 38.195 43.605 38.415 ;
        RECT 42.480 37.565 42.805 38.025 ;
        RECT 43.325 37.735 43.605 38.195 ;
        RECT 43.795 37.735 44.195 38.585 ;
        RECT 44.365 39.315 45.320 39.485 ;
        RECT 45.605 39.345 48.195 40.115 ;
        RECT 48.365 39.390 48.655 40.115 ;
        RECT 49.155 39.715 49.485 40.115 ;
        RECT 49.655 39.545 49.985 39.885 ;
        RECT 51.035 39.715 51.365 40.115 ;
        RECT 49.000 39.375 51.365 39.545 ;
        RECT 51.535 39.390 51.865 39.900 ;
        RECT 44.365 38.415 44.575 39.315 ;
        RECT 44.745 38.585 45.435 39.145 ;
        RECT 45.605 38.825 46.815 39.345 ;
        RECT 46.985 38.655 48.195 39.175 ;
        RECT 44.365 38.195 45.320 38.415 ;
        RECT 44.595 37.565 44.865 38.025 ;
        RECT 45.035 37.735 45.320 38.195 ;
        RECT 45.605 37.565 48.195 38.655 ;
        RECT 48.365 37.565 48.655 38.730 ;
        RECT 49.000 38.375 49.170 39.375 ;
        RECT 51.195 39.205 51.365 39.375 ;
        RECT 49.340 38.545 49.585 39.205 ;
        RECT 49.800 38.545 50.065 39.205 ;
        RECT 50.260 38.545 50.545 39.205 ;
        RECT 50.720 38.875 51.025 39.205 ;
        RECT 51.195 38.875 51.505 39.205 ;
        RECT 50.720 38.545 50.935 38.875 ;
        RECT 49.000 38.205 49.455 38.375 ;
        RECT 49.125 37.775 49.455 38.205 ;
        RECT 49.635 38.205 50.925 38.375 ;
        RECT 49.635 37.785 49.885 38.205 ;
        RECT 50.115 37.565 50.445 38.035 ;
        RECT 50.675 37.785 50.925 38.205 ;
        RECT 51.115 37.565 51.365 38.705 ;
        RECT 51.675 38.625 51.865 39.390 ;
        RECT 53.120 39.465 53.450 39.930 ;
        RECT 53.620 39.645 53.790 40.115 ;
        RECT 53.960 39.465 54.290 39.945 ;
        RECT 53.120 39.295 54.290 39.465 ;
        RECT 52.965 38.915 53.610 39.125 ;
        RECT 53.780 38.915 54.350 39.125 ;
        RECT 54.520 38.745 54.690 39.945 ;
        RECT 55.230 39.545 55.400 39.750 ;
        RECT 51.535 37.775 51.865 38.625 ;
        RECT 53.180 37.565 53.510 38.665 ;
        RECT 53.985 38.335 54.690 38.745 ;
        RECT 54.860 39.375 55.400 39.545 ;
        RECT 55.680 39.375 55.850 40.115 ;
        RECT 56.245 39.750 56.415 39.775 ;
        RECT 56.115 39.375 56.475 39.750 ;
        RECT 54.860 38.675 55.030 39.375 ;
        RECT 55.200 38.875 55.530 39.205 ;
        RECT 55.700 38.875 56.050 39.205 ;
        RECT 54.860 38.505 55.485 38.675 ;
        RECT 55.700 38.335 55.965 38.875 ;
        RECT 56.220 38.720 56.475 39.375 ;
        RECT 57.105 39.365 58.315 40.115 ;
        RECT 53.985 38.165 55.965 38.335 ;
        RECT 53.985 37.735 54.310 38.165 ;
        RECT 54.480 37.565 54.810 37.985 ;
        RECT 55.555 37.565 55.965 37.995 ;
        RECT 56.135 37.735 56.475 38.720 ;
        RECT 57.105 38.655 57.625 39.195 ;
        RECT 57.795 38.825 58.315 39.365 ;
        RECT 57.105 37.565 58.315 38.655 ;
        RECT 22.520 37.395 58.400 37.565 ;
        RECT 22.605 36.305 23.815 37.395 ;
        RECT 24.075 36.725 24.245 37.225 ;
        RECT 24.415 36.895 24.745 37.395 ;
        RECT 24.075 36.555 24.740 36.725 ;
        RECT 22.605 35.595 23.125 36.135 ;
        RECT 23.295 35.765 23.815 36.305 ;
        RECT 23.990 35.735 24.340 36.385 ;
        RECT 22.605 34.845 23.815 35.595 ;
        RECT 24.510 35.565 24.740 36.555 ;
        RECT 24.075 35.395 24.740 35.565 ;
        RECT 24.075 35.105 24.245 35.395 ;
        RECT 24.415 34.845 24.745 35.225 ;
        RECT 24.915 35.105 25.100 37.225 ;
        RECT 25.340 36.935 25.605 37.395 ;
        RECT 25.775 36.800 26.025 37.225 ;
        RECT 26.235 36.950 27.340 37.120 ;
        RECT 25.720 36.670 26.025 36.800 ;
        RECT 25.270 35.475 25.550 36.425 ;
        RECT 25.720 35.565 25.890 36.670 ;
        RECT 26.060 35.885 26.300 36.480 ;
        RECT 26.470 36.415 27.000 36.780 ;
        RECT 26.470 35.715 26.640 36.415 ;
        RECT 27.170 36.335 27.340 36.950 ;
        RECT 27.510 36.595 27.680 37.395 ;
        RECT 27.850 36.895 28.100 37.225 ;
        RECT 28.325 36.925 29.210 37.095 ;
        RECT 27.170 36.245 27.680 36.335 ;
        RECT 25.720 35.435 25.945 35.565 ;
        RECT 26.115 35.495 26.640 35.715 ;
        RECT 26.810 36.075 27.680 36.245 ;
        RECT 25.355 34.845 25.605 35.305 ;
        RECT 25.775 35.295 25.945 35.435 ;
        RECT 26.810 35.295 26.980 36.075 ;
        RECT 27.510 36.005 27.680 36.075 ;
        RECT 27.190 35.825 27.390 35.855 ;
        RECT 27.850 35.825 28.020 36.895 ;
        RECT 28.190 36.005 28.380 36.725 ;
        RECT 27.190 35.525 28.020 35.825 ;
        RECT 28.550 35.795 28.870 36.755 ;
        RECT 25.775 35.125 26.110 35.295 ;
        RECT 26.305 35.125 26.980 35.295 ;
        RECT 27.300 34.845 27.670 35.345 ;
        RECT 27.850 35.295 28.020 35.525 ;
        RECT 28.405 35.465 28.870 35.795 ;
        RECT 29.040 36.085 29.210 36.925 ;
        RECT 29.390 36.895 29.705 37.395 ;
        RECT 29.935 36.665 30.275 37.225 ;
        RECT 29.380 36.290 30.275 36.665 ;
        RECT 30.445 36.385 30.615 37.395 ;
        RECT 30.085 36.085 30.275 36.290 ;
        RECT 30.785 36.335 31.115 37.180 ;
        RECT 30.785 36.255 31.175 36.335 ;
        RECT 31.345 36.305 34.855 37.395 ;
        RECT 30.960 36.205 31.175 36.255 ;
        RECT 29.040 35.755 29.915 36.085 ;
        RECT 30.085 35.755 30.835 36.085 ;
        RECT 29.040 35.295 29.210 35.755 ;
        RECT 30.085 35.585 30.285 35.755 ;
        RECT 31.005 35.625 31.175 36.205 ;
        RECT 30.950 35.585 31.175 35.625 ;
        RECT 27.850 35.125 28.255 35.295 ;
        RECT 28.425 35.125 29.210 35.295 ;
        RECT 29.485 34.845 29.695 35.375 ;
        RECT 29.955 35.060 30.285 35.585 ;
        RECT 30.795 35.500 31.175 35.585 ;
        RECT 31.345 35.615 32.995 36.135 ;
        RECT 33.165 35.785 34.855 36.305 ;
        RECT 35.485 36.230 35.775 37.395 ;
        RECT 36.035 36.725 36.205 37.225 ;
        RECT 36.375 36.895 36.705 37.395 ;
        RECT 36.035 36.555 36.700 36.725 ;
        RECT 35.950 35.735 36.300 36.385 ;
        RECT 30.455 34.845 30.625 35.455 ;
        RECT 30.795 35.065 31.125 35.500 ;
        RECT 31.345 34.845 34.855 35.615 ;
        RECT 35.485 34.845 35.775 35.570 ;
        RECT 36.470 35.565 36.700 36.555 ;
        RECT 36.035 35.395 36.700 35.565 ;
        RECT 36.035 35.105 36.205 35.395 ;
        RECT 36.375 34.845 36.705 35.225 ;
        RECT 36.875 35.105 37.060 37.225 ;
        RECT 37.300 36.935 37.565 37.395 ;
        RECT 37.735 36.800 37.985 37.225 ;
        RECT 38.195 36.950 39.300 37.120 ;
        RECT 37.680 36.670 37.985 36.800 ;
        RECT 37.230 35.475 37.510 36.425 ;
        RECT 37.680 35.565 37.850 36.670 ;
        RECT 38.020 35.885 38.260 36.480 ;
        RECT 38.430 36.415 38.960 36.780 ;
        RECT 38.430 35.715 38.600 36.415 ;
        RECT 39.130 36.335 39.300 36.950 ;
        RECT 39.470 36.595 39.640 37.395 ;
        RECT 39.810 36.895 40.060 37.225 ;
        RECT 40.285 36.925 41.170 37.095 ;
        RECT 39.130 36.245 39.640 36.335 ;
        RECT 37.680 35.435 37.905 35.565 ;
        RECT 38.075 35.495 38.600 35.715 ;
        RECT 38.770 36.075 39.640 36.245 ;
        RECT 37.315 34.845 37.565 35.305 ;
        RECT 37.735 35.295 37.905 35.435 ;
        RECT 38.770 35.295 38.940 36.075 ;
        RECT 39.470 36.005 39.640 36.075 ;
        RECT 39.150 35.825 39.350 35.855 ;
        RECT 39.810 35.825 39.980 36.895 ;
        RECT 40.150 36.005 40.340 36.725 ;
        RECT 39.150 35.525 39.980 35.825 ;
        RECT 40.510 35.795 40.830 36.755 ;
        RECT 37.735 35.125 38.070 35.295 ;
        RECT 38.265 35.125 38.940 35.295 ;
        RECT 39.260 34.845 39.630 35.345 ;
        RECT 39.810 35.295 39.980 35.525 ;
        RECT 40.365 35.465 40.830 35.795 ;
        RECT 41.000 36.085 41.170 36.925 ;
        RECT 41.350 36.895 41.665 37.395 ;
        RECT 41.895 36.665 42.235 37.225 ;
        RECT 41.340 36.290 42.235 36.665 ;
        RECT 42.405 36.385 42.575 37.395 ;
        RECT 42.045 36.085 42.235 36.290 ;
        RECT 42.745 36.335 43.075 37.180 ;
        RECT 43.395 36.775 43.565 37.205 ;
        RECT 43.735 36.945 44.065 37.395 ;
        RECT 43.395 36.545 44.075 36.775 ;
        RECT 42.745 36.255 43.135 36.335 ;
        RECT 42.920 36.205 43.135 36.255 ;
        RECT 43.365 36.205 43.670 36.375 ;
        RECT 41.000 35.755 41.875 36.085 ;
        RECT 42.045 35.755 42.795 36.085 ;
        RECT 41.000 35.295 41.170 35.755 ;
        RECT 42.045 35.585 42.245 35.755 ;
        RECT 42.965 35.625 43.135 36.205 ;
        RECT 42.910 35.585 43.135 35.625 ;
        RECT 39.810 35.125 40.215 35.295 ;
        RECT 40.385 35.125 41.170 35.295 ;
        RECT 41.445 34.845 41.655 35.375 ;
        RECT 41.915 35.060 42.245 35.585 ;
        RECT 42.755 35.500 43.135 35.585 ;
        RECT 43.370 35.525 43.670 36.205 ;
        RECT 43.840 35.895 44.075 36.545 ;
        RECT 44.265 36.235 44.550 37.180 ;
        RECT 44.730 36.925 45.415 37.395 ;
        RECT 44.725 36.405 45.420 36.715 ;
        RECT 45.595 36.340 45.900 37.125 ;
        RECT 46.085 36.440 46.355 37.395 ;
        RECT 44.265 36.085 45.125 36.235 ;
        RECT 44.265 36.065 45.555 36.085 ;
        RECT 43.840 35.565 44.395 35.895 ;
        RECT 44.565 35.705 45.555 36.065 ;
        RECT 42.415 34.845 42.585 35.455 ;
        RECT 42.755 35.065 43.085 35.500 ;
        RECT 43.840 35.415 44.055 35.565 ;
        RECT 43.315 34.845 43.645 35.350 ;
        RECT 43.815 35.040 44.055 35.415 ;
        RECT 44.565 35.370 44.735 35.705 ;
        RECT 45.725 35.535 45.900 36.340 ;
        RECT 46.525 36.305 49.115 37.395 ;
        RECT 49.860 36.765 50.145 37.225 ;
        RECT 50.315 36.935 50.585 37.395 ;
        RECT 49.860 36.545 50.815 36.765 ;
        RECT 44.335 35.175 44.735 35.370 ;
        RECT 44.335 35.030 44.505 35.175 ;
        RECT 45.095 34.845 45.495 35.340 ;
        RECT 45.665 35.015 45.900 35.535 ;
        RECT 46.525 35.615 47.735 36.135 ;
        RECT 47.905 35.785 49.115 36.305 ;
        RECT 49.745 35.815 50.435 36.375 ;
        RECT 50.605 35.645 50.815 36.545 ;
        RECT 46.085 34.845 46.355 35.480 ;
        RECT 46.525 34.845 49.115 35.615 ;
        RECT 49.860 35.475 50.815 35.645 ;
        RECT 50.985 36.375 51.385 37.225 ;
        RECT 51.575 36.765 51.855 37.225 ;
        RECT 52.375 36.935 52.700 37.395 ;
        RECT 51.575 36.545 52.700 36.765 ;
        RECT 50.985 35.815 52.080 36.375 ;
        RECT 52.250 36.085 52.700 36.545 ;
        RECT 52.870 36.255 53.255 37.225 ;
        RECT 49.860 35.015 50.145 35.475 ;
        RECT 50.315 34.845 50.585 35.305 ;
        RECT 50.985 35.015 51.385 35.815 ;
        RECT 52.250 35.755 52.805 36.085 ;
        RECT 52.250 35.645 52.700 35.755 ;
        RECT 51.575 35.475 52.700 35.645 ;
        RECT 52.975 35.585 53.255 36.255 ;
        RECT 51.575 35.015 51.855 35.475 ;
        RECT 52.375 34.845 52.700 35.305 ;
        RECT 52.870 35.015 53.255 35.585 ;
        RECT 53.425 36.595 53.865 37.225 ;
        RECT 53.425 35.585 53.735 36.595 ;
        RECT 54.040 36.545 54.355 37.395 ;
        RECT 54.525 37.055 55.955 37.225 ;
        RECT 54.525 36.375 54.695 37.055 ;
        RECT 53.905 36.205 54.695 36.375 ;
        RECT 53.905 35.755 54.075 36.205 ;
        RECT 54.865 36.085 55.065 36.885 ;
        RECT 54.245 35.755 54.635 36.035 ;
        RECT 54.820 35.755 55.065 36.085 ;
        RECT 55.265 35.755 55.515 36.885 ;
        RECT 55.705 36.425 55.955 37.055 ;
        RECT 56.135 36.595 56.465 37.395 ;
        RECT 55.705 36.255 56.475 36.425 ;
        RECT 55.730 35.755 56.135 36.085 ;
        RECT 56.305 35.585 56.475 36.255 ;
        RECT 57.105 36.305 58.315 37.395 ;
        RECT 57.105 35.765 57.625 36.305 ;
        RECT 57.795 35.595 58.315 36.135 ;
        RECT 53.425 35.025 53.865 35.585 ;
        RECT 54.035 34.845 54.485 35.585 ;
        RECT 54.655 35.415 55.815 35.585 ;
        RECT 54.655 35.015 54.825 35.415 ;
        RECT 54.995 34.845 55.415 35.245 ;
        RECT 55.585 35.015 55.815 35.415 ;
        RECT 55.985 35.015 56.475 35.585 ;
        RECT 57.105 34.845 58.315 35.595 ;
        RECT 75.000 35.765 75.885 41.025 ;
        RECT 76.565 40.455 78.605 40.625 ;
        RECT 76.225 36.395 76.395 40.395 ;
        RECT 78.775 36.395 78.945 40.395 ;
        RECT 76.565 36.165 78.605 36.335 ;
        RECT 79.285 35.765 79.455 41.025 ;
        RECT 75.000 35.595 79.455 35.765 ;
        RECT 80.190 46.545 90.580 46.715 ;
        RECT 80.190 41.285 80.360 46.545 ;
        RECT 81.085 45.975 85.125 46.145 ;
        RECT 80.700 41.915 80.870 45.915 ;
        RECT 85.340 41.915 85.510 45.915 ;
        RECT 85.850 45.435 90.580 46.545 ;
        RECT 81.085 41.685 85.125 41.855 ;
        RECT 85.850 41.285 86.020 45.435 ;
        RECT 80.190 41.115 86.020 41.285 ;
        RECT 80.190 35.855 80.360 41.115 ;
        RECT 81.085 40.545 85.125 40.715 ;
        RECT 80.700 36.485 80.870 40.485 ;
        RECT 85.340 36.485 85.510 40.485 ;
        RECT 81.085 36.255 85.125 36.425 ;
        RECT 85.850 35.855 86.020 41.115 ;
        RECT 86.535 45.360 88.285 45.435 ;
        RECT 86.535 38.870 86.705 45.360 ;
        RECT 87.245 44.850 87.575 45.020 ;
        RECT 87.105 39.595 87.275 44.635 ;
        RECT 87.545 39.595 87.715 44.635 ;
        RECT 87.245 39.210 87.575 39.380 ;
        RECT 88.115 38.870 88.285 45.360 ;
        RECT 86.535 38.700 88.285 38.870 ;
        RECT 80.190 35.685 86.020 35.855 ;
        RECT 75.000 35.325 76.860 35.595 ;
        RECT 75.000 35.155 79.460 35.325 ;
        RECT 22.520 34.675 58.400 34.845 ;
        RECT 22.605 33.925 23.815 34.675 ;
        RECT 22.605 33.385 23.125 33.925 ;
        RECT 23.990 33.835 24.250 34.675 ;
        RECT 24.425 33.930 24.680 34.505 ;
        RECT 24.850 34.295 25.180 34.675 ;
        RECT 25.395 34.125 25.565 34.505 ;
        RECT 24.850 33.955 25.565 34.125 ;
        RECT 26.860 34.045 27.145 34.505 ;
        RECT 27.315 34.215 27.585 34.675 ;
        RECT 23.295 33.215 23.815 33.755 ;
        RECT 22.605 32.125 23.815 33.215 ;
        RECT 23.990 32.125 24.250 33.275 ;
        RECT 24.425 33.200 24.595 33.930 ;
        RECT 24.850 33.765 25.020 33.955 ;
        RECT 26.860 33.875 27.815 34.045 ;
        RECT 24.765 33.435 25.020 33.765 ;
        RECT 24.850 33.225 25.020 33.435 ;
        RECT 25.300 33.405 25.655 33.775 ;
        RECT 24.425 32.295 24.680 33.200 ;
        RECT 24.850 33.055 25.565 33.225 ;
        RECT 26.745 33.145 27.435 33.705 ;
        RECT 24.850 32.125 25.180 32.885 ;
        RECT 25.395 32.295 25.565 33.055 ;
        RECT 27.605 32.975 27.815 33.875 ;
        RECT 26.860 32.755 27.815 32.975 ;
        RECT 27.985 33.705 28.385 34.505 ;
        RECT 28.575 34.045 28.855 34.505 ;
        RECT 29.375 34.215 29.700 34.675 ;
        RECT 28.575 33.875 29.700 34.045 ;
        RECT 29.870 33.935 30.255 34.505 ;
        RECT 29.250 33.765 29.700 33.875 ;
        RECT 27.985 33.145 29.080 33.705 ;
        RECT 29.250 33.435 29.805 33.765 ;
        RECT 26.860 32.295 27.145 32.755 ;
        RECT 27.315 32.125 27.585 32.585 ;
        RECT 27.985 32.295 28.385 33.145 ;
        RECT 29.250 32.975 29.700 33.435 ;
        RECT 29.975 33.265 30.255 33.935 ;
        RECT 31.460 34.045 31.745 34.505 ;
        RECT 31.915 34.215 32.185 34.675 ;
        RECT 31.460 33.875 32.415 34.045 ;
        RECT 28.575 32.755 29.700 32.975 ;
        RECT 28.575 32.295 28.855 32.755 ;
        RECT 29.375 32.125 29.700 32.585 ;
        RECT 29.870 32.295 30.255 33.265 ;
        RECT 31.345 33.145 32.035 33.705 ;
        RECT 32.205 32.975 32.415 33.875 ;
        RECT 31.460 32.755 32.415 32.975 ;
        RECT 32.585 33.705 32.985 34.505 ;
        RECT 33.175 34.045 33.455 34.505 ;
        RECT 33.975 34.215 34.300 34.675 ;
        RECT 33.175 33.875 34.300 34.045 ;
        RECT 34.470 33.935 34.855 34.505 ;
        RECT 33.850 33.765 34.300 33.875 ;
        RECT 32.585 33.145 33.680 33.705 ;
        RECT 33.850 33.435 34.405 33.765 ;
        RECT 31.460 32.295 31.745 32.755 ;
        RECT 31.915 32.125 32.185 32.585 ;
        RECT 32.585 32.295 32.985 33.145 ;
        RECT 33.850 32.975 34.300 33.435 ;
        RECT 34.575 33.265 34.855 33.935 ;
        RECT 35.300 33.865 35.545 34.470 ;
        RECT 35.765 34.140 36.275 34.675 ;
        RECT 33.175 32.755 34.300 32.975 ;
        RECT 33.175 32.295 33.455 32.755 ;
        RECT 33.975 32.125 34.300 32.585 ;
        RECT 34.470 32.295 34.855 33.265 ;
        RECT 35.025 33.695 36.255 33.865 ;
        RECT 35.025 32.885 35.365 33.695 ;
        RECT 35.535 33.130 36.285 33.320 ;
        RECT 35.025 32.475 35.540 32.885 ;
        RECT 35.775 32.125 35.945 32.885 ;
        RECT 36.115 32.465 36.285 33.130 ;
        RECT 36.455 33.145 36.645 34.505 ;
        RECT 36.815 33.655 37.090 34.505 ;
        RECT 37.280 34.140 37.810 34.505 ;
        RECT 38.235 34.275 38.565 34.675 ;
        RECT 37.635 34.105 37.810 34.140 ;
        RECT 36.815 33.485 37.095 33.655 ;
        RECT 36.815 33.345 37.090 33.485 ;
        RECT 37.295 33.145 37.465 33.945 ;
        RECT 36.455 32.975 37.465 33.145 ;
        RECT 37.635 33.935 38.565 34.105 ;
        RECT 38.735 33.935 38.990 34.505 ;
        RECT 37.635 32.805 37.805 33.935 ;
        RECT 38.395 33.765 38.565 33.935 ;
        RECT 36.680 32.635 37.805 32.805 ;
        RECT 37.975 33.435 38.170 33.765 ;
        RECT 38.395 33.435 38.650 33.765 ;
        RECT 37.975 32.465 38.145 33.435 ;
        RECT 38.820 33.265 38.990 33.935 ;
        RECT 39.165 33.905 40.835 34.675 ;
        RECT 41.095 34.125 41.265 34.415 ;
        RECT 41.435 34.295 41.765 34.675 ;
        RECT 41.095 33.955 41.760 34.125 ;
        RECT 39.165 33.385 39.915 33.905 ;
        RECT 36.115 32.295 38.145 32.465 ;
        RECT 38.315 32.125 38.485 33.265 ;
        RECT 38.655 32.295 38.990 33.265 ;
        RECT 40.085 33.215 40.835 33.735 ;
        RECT 39.165 32.125 40.835 33.215 ;
        RECT 41.010 33.135 41.360 33.785 ;
        RECT 41.530 32.965 41.760 33.955 ;
        RECT 41.095 32.795 41.760 32.965 ;
        RECT 41.095 32.295 41.265 32.795 ;
        RECT 41.435 32.125 41.765 32.625 ;
        RECT 41.935 32.295 42.120 34.415 ;
        RECT 42.375 34.215 42.625 34.675 ;
        RECT 42.795 34.225 43.130 34.395 ;
        RECT 43.325 34.225 44.000 34.395 ;
        RECT 42.795 34.085 42.965 34.225 ;
        RECT 42.290 33.095 42.570 34.045 ;
        RECT 42.740 33.955 42.965 34.085 ;
        RECT 42.740 32.850 42.910 33.955 ;
        RECT 43.135 33.805 43.660 34.025 ;
        RECT 43.080 33.040 43.320 33.635 ;
        RECT 43.490 33.105 43.660 33.805 ;
        RECT 43.830 33.445 44.000 34.225 ;
        RECT 44.320 34.175 44.690 34.675 ;
        RECT 44.870 34.225 45.275 34.395 ;
        RECT 45.445 34.225 46.230 34.395 ;
        RECT 44.870 33.995 45.040 34.225 ;
        RECT 44.210 33.695 45.040 33.995 ;
        RECT 45.425 33.725 45.890 34.055 ;
        RECT 44.210 33.665 44.410 33.695 ;
        RECT 44.530 33.445 44.700 33.515 ;
        RECT 43.830 33.275 44.700 33.445 ;
        RECT 44.190 33.185 44.700 33.275 ;
        RECT 42.740 32.720 43.045 32.850 ;
        RECT 43.490 32.740 44.020 33.105 ;
        RECT 42.360 32.125 42.625 32.585 ;
        RECT 42.795 32.295 43.045 32.720 ;
        RECT 44.190 32.570 44.360 33.185 ;
        RECT 43.255 32.400 44.360 32.570 ;
        RECT 44.530 32.125 44.700 32.925 ;
        RECT 44.870 32.625 45.040 33.695 ;
        RECT 45.210 32.795 45.400 33.515 ;
        RECT 45.570 32.765 45.890 33.725 ;
        RECT 46.060 33.765 46.230 34.225 ;
        RECT 46.505 34.145 46.715 34.675 ;
        RECT 46.975 33.935 47.305 34.460 ;
        RECT 47.475 34.065 47.645 34.675 ;
        RECT 47.815 34.020 48.145 34.455 ;
        RECT 47.815 33.935 48.195 34.020 ;
        RECT 48.365 33.950 48.655 34.675 ;
        RECT 47.105 33.765 47.305 33.935 ;
        RECT 47.970 33.895 48.195 33.935 ;
        RECT 46.060 33.435 46.935 33.765 ;
        RECT 47.105 33.435 47.855 33.765 ;
        RECT 44.870 32.295 45.120 32.625 ;
        RECT 46.060 32.595 46.230 33.435 ;
        RECT 47.105 33.230 47.295 33.435 ;
        RECT 48.025 33.315 48.195 33.895 ;
        RECT 47.980 33.265 48.195 33.315 ;
        RECT 48.830 33.935 49.085 34.505 ;
        RECT 49.255 34.275 49.585 34.675 ;
        RECT 50.010 34.140 50.540 34.505 ;
        RECT 50.730 34.335 51.005 34.505 ;
        RECT 50.725 34.165 51.005 34.335 ;
        RECT 50.010 34.105 50.185 34.140 ;
        RECT 49.255 33.935 50.185 34.105 ;
        RECT 46.400 32.855 47.295 33.230 ;
        RECT 47.805 33.185 48.195 33.265 ;
        RECT 45.345 32.425 46.230 32.595 ;
        RECT 46.410 32.125 46.725 32.625 ;
        RECT 46.955 32.295 47.295 32.855 ;
        RECT 47.465 32.125 47.635 33.135 ;
        RECT 47.805 32.340 48.135 33.185 ;
        RECT 48.365 32.125 48.655 33.290 ;
        RECT 48.830 33.265 49.000 33.935 ;
        RECT 49.255 33.765 49.425 33.935 ;
        RECT 49.170 33.435 49.425 33.765 ;
        RECT 49.650 33.435 49.845 33.765 ;
        RECT 48.830 32.295 49.165 33.265 ;
        RECT 49.335 32.125 49.505 33.265 ;
        RECT 49.675 32.465 49.845 33.435 ;
        RECT 50.015 32.805 50.185 33.935 ;
        RECT 50.355 33.145 50.525 33.945 ;
        RECT 50.730 33.345 51.005 34.165 ;
        RECT 51.175 33.145 51.365 34.505 ;
        RECT 51.545 34.140 52.055 34.675 ;
        RECT 52.275 33.865 52.520 34.470 ;
        RECT 53.055 34.125 53.225 34.505 ;
        RECT 53.405 34.295 53.735 34.675 ;
        RECT 53.055 33.955 53.720 34.125 ;
        RECT 53.915 34.000 54.175 34.505 ;
        RECT 51.565 33.695 52.795 33.865 ;
        RECT 50.355 32.975 51.365 33.145 ;
        RECT 51.535 33.130 52.285 33.320 ;
        RECT 50.015 32.635 51.140 32.805 ;
        RECT 51.535 32.465 51.705 33.130 ;
        RECT 52.455 32.885 52.795 33.695 ;
        RECT 52.985 33.405 53.315 33.775 ;
        RECT 53.550 33.700 53.720 33.955 ;
        RECT 53.550 33.370 53.835 33.700 ;
        RECT 53.550 33.225 53.720 33.370 ;
        RECT 49.675 32.295 51.705 32.465 ;
        RECT 51.875 32.125 52.045 32.885 ;
        RECT 52.280 32.475 52.795 32.885 ;
        RECT 53.055 33.055 53.720 33.225 ;
        RECT 54.005 33.200 54.175 34.000 ;
        RECT 53.055 32.295 53.225 33.055 ;
        RECT 53.405 32.125 53.735 32.885 ;
        RECT 53.905 32.295 54.175 33.200 ;
        RECT 54.345 34.000 54.615 34.345 ;
        RECT 54.805 34.275 55.185 34.675 ;
        RECT 55.355 34.105 55.525 34.455 ;
        RECT 55.695 34.275 56.025 34.675 ;
        RECT 56.225 34.105 56.395 34.455 ;
        RECT 56.595 34.175 56.925 34.675 ;
        RECT 54.345 33.265 54.515 34.000 ;
        RECT 54.785 33.935 56.395 34.105 ;
        RECT 54.785 33.765 54.955 33.935 ;
        RECT 54.685 33.435 54.955 33.765 ;
        RECT 55.125 33.435 55.530 33.765 ;
        RECT 54.785 33.265 54.955 33.435 ;
        RECT 54.345 32.295 54.615 33.265 ;
        RECT 54.785 33.095 55.510 33.265 ;
        RECT 55.700 33.145 56.410 33.765 ;
        RECT 56.580 33.435 56.930 34.005 ;
        RECT 57.105 33.925 58.315 34.675 ;
        RECT 55.340 32.975 55.510 33.095 ;
        RECT 56.610 32.975 56.930 33.265 ;
        RECT 54.825 32.125 55.105 32.925 ;
        RECT 55.340 32.805 56.930 32.975 ;
        RECT 57.105 33.215 57.625 33.755 ;
        RECT 57.795 33.385 58.315 33.925 ;
        RECT 75.000 33.745 76.890 35.155 ;
        RECT 77.230 34.285 77.400 34.615 ;
        RECT 77.570 34.585 78.610 34.755 ;
        RECT 77.570 34.145 78.610 34.315 ;
        RECT 78.780 34.285 78.950 34.615 ;
        RECT 79.290 33.745 79.460 35.155 ;
        RECT 75.000 33.575 79.460 33.745 ;
        RECT 80.205 35.240 86.035 35.410 ;
        RECT 80.205 33.830 80.375 35.240 ;
        RECT 80.715 34.370 80.885 34.700 ;
        RECT 81.100 34.670 85.140 34.840 ;
        RECT 81.100 34.230 85.140 34.400 ;
        RECT 85.355 34.370 85.525 34.700 ;
        RECT 85.865 33.830 86.035 35.240 ;
        RECT 80.205 33.660 86.035 33.830 ;
        RECT 75.000 33.300 76.860 33.575 ;
        RECT 89.880 33.385 90.580 45.435 ;
        RECT 55.275 32.345 56.930 32.635 ;
        RECT 57.105 32.125 58.315 33.215 ;
        RECT 75.000 33.130 79.465 33.300 ;
        RECT 22.520 31.955 58.400 32.125 ;
        RECT 22.605 30.865 23.815 31.955 ;
        RECT 24.045 30.895 24.375 31.740 ;
        RECT 24.545 30.945 24.715 31.955 ;
        RECT 24.885 31.225 25.225 31.785 ;
        RECT 25.455 31.455 25.770 31.955 ;
        RECT 25.950 31.485 26.835 31.655 ;
        RECT 22.605 30.155 23.125 30.695 ;
        RECT 23.295 30.325 23.815 30.865 ;
        RECT 23.985 30.815 24.375 30.895 ;
        RECT 24.885 30.850 25.780 31.225 ;
        RECT 23.985 30.765 24.200 30.815 ;
        RECT 23.985 30.185 24.155 30.765 ;
        RECT 24.885 30.645 25.075 30.850 ;
        RECT 25.950 30.645 26.120 31.485 ;
        RECT 27.060 31.455 27.310 31.785 ;
        RECT 24.325 30.315 25.075 30.645 ;
        RECT 25.245 30.315 26.120 30.645 ;
        RECT 22.605 29.405 23.815 30.155 ;
        RECT 23.985 30.145 24.210 30.185 ;
        RECT 24.875 30.145 25.075 30.315 ;
        RECT 23.985 30.060 24.365 30.145 ;
        RECT 24.035 29.625 24.365 30.060 ;
        RECT 24.535 29.405 24.705 30.015 ;
        RECT 24.875 29.620 25.205 30.145 ;
        RECT 25.465 29.405 25.675 29.935 ;
        RECT 25.950 29.855 26.120 30.315 ;
        RECT 26.290 30.355 26.610 31.315 ;
        RECT 26.780 30.565 26.970 31.285 ;
        RECT 27.140 30.385 27.310 31.455 ;
        RECT 27.480 31.155 27.650 31.955 ;
        RECT 27.820 31.510 28.925 31.680 ;
        RECT 27.820 30.895 27.990 31.510 ;
        RECT 29.135 31.360 29.385 31.785 ;
        RECT 29.555 31.495 29.820 31.955 ;
        RECT 28.160 30.975 28.690 31.340 ;
        RECT 29.135 31.230 29.440 31.360 ;
        RECT 27.480 30.805 27.990 30.895 ;
        RECT 27.480 30.635 28.350 30.805 ;
        RECT 27.480 30.565 27.650 30.635 ;
        RECT 27.770 30.385 27.970 30.415 ;
        RECT 26.290 30.025 26.755 30.355 ;
        RECT 27.140 30.085 27.970 30.385 ;
        RECT 27.140 29.855 27.310 30.085 ;
        RECT 25.950 29.685 26.735 29.855 ;
        RECT 26.905 29.685 27.310 29.855 ;
        RECT 27.490 29.405 27.860 29.905 ;
        RECT 28.180 29.855 28.350 30.635 ;
        RECT 28.520 30.275 28.690 30.975 ;
        RECT 28.860 30.445 29.100 31.040 ;
        RECT 28.520 30.055 29.045 30.275 ;
        RECT 29.270 30.125 29.440 31.230 ;
        RECT 29.215 29.995 29.440 30.125 ;
        RECT 29.610 30.035 29.890 30.985 ;
        RECT 29.215 29.855 29.385 29.995 ;
        RECT 28.180 29.685 28.855 29.855 ;
        RECT 29.050 29.685 29.385 29.855 ;
        RECT 29.555 29.405 29.805 29.865 ;
        RECT 30.060 29.665 30.245 31.785 ;
        RECT 30.415 31.455 30.745 31.955 ;
        RECT 30.915 31.285 31.085 31.785 ;
        RECT 30.420 31.115 31.085 31.285 ;
        RECT 30.420 30.125 30.650 31.115 ;
        RECT 30.820 30.295 31.170 30.945 ;
        RECT 31.345 30.865 34.855 31.955 ;
        RECT 31.345 30.175 32.995 30.695 ;
        RECT 33.165 30.345 34.855 30.865 ;
        RECT 35.485 30.790 35.775 31.955 ;
        RECT 35.955 31.145 36.250 31.955 ;
        RECT 36.430 30.645 36.675 31.785 ;
        RECT 36.850 31.145 37.110 31.955 ;
        RECT 37.710 31.950 43.985 31.955 ;
        RECT 37.290 30.645 37.540 31.780 ;
        RECT 37.710 31.155 37.970 31.950 ;
        RECT 38.140 31.055 38.400 31.780 ;
        RECT 38.570 31.225 38.830 31.950 ;
        RECT 39.000 31.055 39.260 31.780 ;
        RECT 39.430 31.225 39.690 31.950 ;
        RECT 39.860 31.055 40.120 31.780 ;
        RECT 40.290 31.225 40.550 31.950 ;
        RECT 40.720 31.055 40.980 31.780 ;
        RECT 41.150 31.225 41.395 31.950 ;
        RECT 41.565 31.055 41.825 31.780 ;
        RECT 42.010 31.225 42.255 31.950 ;
        RECT 42.425 31.055 42.685 31.780 ;
        RECT 42.870 31.225 43.115 31.950 ;
        RECT 43.285 31.055 43.545 31.780 ;
        RECT 43.730 31.225 43.985 31.950 ;
        RECT 38.140 31.040 43.545 31.055 ;
        RECT 44.155 31.040 44.445 31.780 ;
        RECT 44.615 31.210 44.885 31.955 ;
        RECT 38.140 30.815 44.885 31.040 ;
        RECT 45.145 30.865 46.355 31.955 ;
        RECT 30.420 29.955 31.085 30.125 ;
        RECT 30.415 29.405 30.745 29.785 ;
        RECT 30.915 29.665 31.085 29.955 ;
        RECT 31.345 29.405 34.855 30.175 ;
        RECT 35.485 29.405 35.775 30.130 ;
        RECT 35.945 30.085 36.260 30.645 ;
        RECT 36.430 30.395 43.550 30.645 ;
        RECT 35.945 29.405 36.250 29.915 ;
        RECT 36.430 29.585 36.680 30.395 ;
        RECT 36.850 29.405 37.110 29.930 ;
        RECT 37.290 29.585 37.540 30.395 ;
        RECT 43.720 30.225 44.885 30.815 ;
        RECT 38.140 30.055 44.885 30.225 ;
        RECT 45.145 30.155 45.665 30.695 ;
        RECT 45.835 30.325 46.355 30.865 ;
        RECT 46.615 31.025 46.785 31.785 ;
        RECT 46.965 31.195 47.295 31.955 ;
        RECT 46.615 30.855 47.280 31.025 ;
        RECT 47.465 30.880 47.735 31.785 ;
        RECT 47.110 30.710 47.280 30.855 ;
        RECT 46.545 30.305 46.875 30.675 ;
        RECT 47.110 30.380 47.395 30.710 ;
        RECT 37.710 29.405 37.970 29.965 ;
        RECT 38.140 29.600 38.400 30.055 ;
        RECT 38.570 29.405 38.830 29.885 ;
        RECT 39.000 29.600 39.260 30.055 ;
        RECT 39.430 29.405 39.690 29.885 ;
        RECT 39.860 29.600 40.120 30.055 ;
        RECT 40.290 29.405 40.535 29.885 ;
        RECT 40.705 29.600 40.980 30.055 ;
        RECT 41.150 29.405 41.395 29.885 ;
        RECT 41.565 29.600 41.825 30.055 ;
        RECT 42.005 29.405 42.255 29.885 ;
        RECT 42.425 29.600 42.685 30.055 ;
        RECT 42.865 29.405 43.115 29.885 ;
        RECT 43.285 29.600 43.545 30.055 ;
        RECT 43.725 29.405 43.985 29.885 ;
        RECT 44.155 29.600 44.415 30.055 ;
        RECT 44.585 29.405 44.885 29.885 ;
        RECT 45.145 29.405 46.355 30.155 ;
        RECT 47.110 30.125 47.280 30.380 ;
        RECT 46.615 29.955 47.280 30.125 ;
        RECT 47.565 30.080 47.735 30.880 ;
        RECT 47.995 31.025 48.165 31.785 ;
        RECT 48.345 31.195 48.675 31.955 ;
        RECT 47.995 30.855 48.660 31.025 ;
        RECT 48.845 30.880 49.115 31.785 ;
        RECT 48.490 30.710 48.660 30.855 ;
        RECT 47.925 30.305 48.255 30.675 ;
        RECT 48.490 30.380 48.775 30.710 ;
        RECT 48.490 30.125 48.660 30.380 ;
        RECT 46.615 29.575 46.785 29.955 ;
        RECT 46.965 29.405 47.295 29.785 ;
        RECT 47.475 29.575 47.735 30.080 ;
        RECT 47.995 29.955 48.660 30.125 ;
        RECT 48.945 30.080 49.115 30.880 ;
        RECT 49.375 31.025 49.545 31.785 ;
        RECT 49.725 31.195 50.055 31.955 ;
        RECT 49.375 30.855 50.040 31.025 ;
        RECT 50.225 30.880 50.495 31.785 ;
        RECT 49.870 30.710 50.040 30.855 ;
        RECT 49.305 30.305 49.635 30.675 ;
        RECT 49.870 30.380 50.155 30.710 ;
        RECT 49.870 30.125 50.040 30.380 ;
        RECT 47.995 29.575 48.165 29.955 ;
        RECT 48.345 29.405 48.675 29.785 ;
        RECT 48.855 29.575 49.115 30.080 ;
        RECT 49.375 29.955 50.040 30.125 ;
        RECT 50.325 30.080 50.495 30.880 ;
        RECT 50.755 31.025 50.925 31.785 ;
        RECT 51.105 31.195 51.435 31.955 ;
        RECT 50.755 30.855 51.420 31.025 ;
        RECT 51.605 30.880 51.875 31.785 ;
        RECT 51.250 30.710 51.420 30.855 ;
        RECT 50.685 30.305 51.015 30.675 ;
        RECT 51.250 30.380 51.535 30.710 ;
        RECT 51.250 30.125 51.420 30.380 ;
        RECT 49.375 29.575 49.545 29.955 ;
        RECT 49.725 29.405 50.055 29.785 ;
        RECT 50.235 29.575 50.495 30.080 ;
        RECT 50.755 29.955 51.420 30.125 ;
        RECT 51.705 30.080 51.875 30.880 ;
        RECT 52.055 30.815 52.385 31.955 ;
        RECT 52.915 30.985 53.245 31.770 ;
        RECT 52.565 30.815 53.245 30.985 ;
        RECT 52.045 30.395 52.395 30.645 ;
        RECT 52.565 30.215 52.735 30.815 ;
        RECT 53.425 30.800 53.765 31.785 ;
        RECT 53.935 31.525 54.345 31.955 ;
        RECT 55.090 31.535 55.420 31.955 ;
        RECT 55.590 31.355 55.915 31.785 ;
        RECT 53.935 31.185 55.915 31.355 ;
        RECT 52.905 30.395 53.255 30.645 ;
        RECT 50.755 29.575 50.925 29.955 ;
        RECT 51.105 29.405 51.435 29.785 ;
        RECT 51.615 29.575 51.875 30.080 ;
        RECT 52.055 29.405 52.325 30.215 ;
        RECT 52.495 29.575 52.825 30.215 ;
        RECT 52.995 29.405 53.235 30.215 ;
        RECT 53.425 30.145 53.680 30.800 ;
        RECT 53.935 30.645 54.200 31.185 ;
        RECT 54.415 30.845 55.040 31.015 ;
        RECT 53.850 30.315 54.200 30.645 ;
        RECT 54.370 30.315 54.700 30.645 ;
        RECT 54.870 30.145 55.040 30.845 ;
        RECT 53.425 29.770 53.785 30.145 ;
        RECT 54.050 29.405 54.220 30.145 ;
        RECT 54.500 29.975 55.040 30.145 ;
        RECT 55.210 30.775 55.915 31.185 ;
        RECT 56.390 30.855 56.720 31.955 ;
        RECT 57.105 30.865 58.315 31.955 ;
        RECT 75.000 31.720 75.895 33.130 ;
        RECT 76.235 32.260 76.405 32.590 ;
        RECT 76.575 32.560 78.615 32.730 ;
        RECT 76.575 32.120 78.615 32.290 ;
        RECT 78.785 32.260 78.955 32.590 ;
        RECT 79.295 31.720 79.465 33.130 ;
        RECT 75.000 31.560 79.465 31.720 ;
        RECT 80.210 33.215 90.580 33.385 ;
        RECT 80.210 31.805 80.380 33.215 ;
        RECT 80.720 32.345 80.890 32.675 ;
        RECT 81.105 32.645 89.145 32.815 ;
        RECT 81.105 32.205 89.145 32.375 ;
        RECT 89.360 32.345 89.530 32.675 ;
        RECT 89.870 31.805 90.580 33.215 ;
        RECT 80.210 31.690 90.580 31.805 ;
        RECT 92.000 57.485 92.865 58.140 ;
        RECT 97.195 57.975 107.580 58.145 ;
        RECT 92.000 57.315 96.455 57.485 ;
        RECT 92.000 52.055 92.885 57.315 ;
        RECT 93.565 56.745 95.605 56.915 ;
        RECT 93.225 52.685 93.395 56.685 ;
        RECT 95.775 52.685 95.945 56.685 ;
        RECT 93.565 52.455 95.605 52.625 ;
        RECT 96.285 52.055 96.455 57.315 ;
        RECT 97.195 54.485 97.365 57.975 ;
        RECT 97.995 57.465 105.995 57.635 ;
        RECT 97.765 55.210 97.935 57.250 ;
        RECT 106.055 55.210 106.225 57.250 ;
        RECT 97.995 54.825 105.995 54.995 ;
        RECT 106.625 54.485 107.580 57.975 ;
        RECT 97.195 54.315 107.580 54.485 ;
        RECT 106.625 54.025 107.580 54.315 ;
        RECT 92.000 51.885 96.455 52.055 ;
        RECT 92.000 46.625 92.885 51.885 ;
        RECT 93.565 51.315 95.605 51.485 ;
        RECT 93.225 47.255 93.395 51.255 ;
        RECT 95.775 47.255 95.945 51.255 ;
        RECT 93.565 47.025 95.605 47.195 ;
        RECT 96.285 46.625 96.455 51.885 ;
        RECT 97.195 53.855 107.580 54.025 ;
        RECT 97.195 50.595 97.365 53.855 ;
        RECT 98.090 53.285 106.130 53.455 ;
        RECT 97.705 51.225 97.875 53.225 ;
        RECT 106.345 51.225 106.515 53.225 ;
        RECT 98.090 50.995 106.130 51.165 ;
        RECT 106.855 50.595 107.580 53.855 ;
        RECT 97.195 50.425 107.580 50.595 ;
        RECT 97.195 47.165 97.365 50.425 ;
        RECT 98.090 49.855 106.130 50.025 ;
        RECT 97.705 47.795 97.875 49.795 ;
        RECT 106.345 47.795 106.515 49.795 ;
        RECT 98.090 47.565 106.130 47.735 ;
        RECT 106.855 47.165 107.580 50.425 ;
        RECT 97.195 46.995 107.580 47.165 ;
        RECT 102.905 46.715 107.580 46.995 ;
        RECT 92.000 46.455 96.455 46.625 ;
        RECT 92.000 41.195 92.885 46.455 ;
        RECT 93.565 45.885 95.605 46.055 ;
        RECT 93.225 41.825 93.395 45.825 ;
        RECT 95.775 41.825 95.945 45.825 ;
        RECT 93.565 41.595 95.605 41.765 ;
        RECT 96.285 41.195 96.455 46.455 ;
        RECT 92.000 41.025 96.455 41.195 ;
        RECT 92.000 35.765 92.885 41.025 ;
        RECT 93.565 40.455 95.605 40.625 ;
        RECT 93.225 36.395 93.395 40.395 ;
        RECT 95.775 36.395 95.945 40.395 ;
        RECT 93.565 36.165 95.605 36.335 ;
        RECT 96.285 35.765 96.455 41.025 ;
        RECT 92.000 35.595 96.455 35.765 ;
        RECT 97.190 46.545 107.580 46.715 ;
        RECT 97.190 41.285 97.360 46.545 ;
        RECT 98.085 45.975 102.125 46.145 ;
        RECT 97.700 41.915 97.870 45.915 ;
        RECT 102.340 41.915 102.510 45.915 ;
        RECT 102.850 45.435 107.580 46.545 ;
        RECT 98.085 41.685 102.125 41.855 ;
        RECT 102.850 41.285 103.020 45.435 ;
        RECT 97.190 41.115 103.020 41.285 ;
        RECT 97.190 35.855 97.360 41.115 ;
        RECT 98.085 40.545 102.125 40.715 ;
        RECT 97.700 36.485 97.870 40.485 ;
        RECT 102.340 36.485 102.510 40.485 ;
        RECT 98.085 36.255 102.125 36.425 ;
        RECT 102.850 35.855 103.020 41.115 ;
        RECT 103.535 45.360 105.285 45.435 ;
        RECT 103.535 38.870 103.705 45.360 ;
        RECT 104.245 44.850 104.575 45.020 ;
        RECT 104.105 39.595 104.275 44.635 ;
        RECT 104.545 39.595 104.715 44.635 ;
        RECT 104.245 39.210 104.575 39.380 ;
        RECT 105.115 38.870 105.285 45.360 ;
        RECT 103.535 38.700 105.285 38.870 ;
        RECT 97.190 35.685 103.020 35.855 ;
        RECT 92.000 35.325 93.860 35.595 ;
        RECT 92.000 35.155 96.460 35.325 ;
        RECT 92.000 33.745 93.890 35.155 ;
        RECT 94.230 34.285 94.400 34.615 ;
        RECT 94.570 34.585 95.610 34.755 ;
        RECT 94.570 34.145 95.610 34.315 ;
        RECT 95.780 34.285 95.950 34.615 ;
        RECT 96.290 33.745 96.460 35.155 ;
        RECT 92.000 33.575 96.460 33.745 ;
        RECT 97.205 35.240 103.035 35.410 ;
        RECT 97.205 33.830 97.375 35.240 ;
        RECT 97.715 34.370 97.885 34.700 ;
        RECT 98.100 34.670 102.140 34.840 ;
        RECT 98.100 34.230 102.140 34.400 ;
        RECT 102.355 34.370 102.525 34.700 ;
        RECT 102.865 33.830 103.035 35.240 ;
        RECT 97.205 33.660 103.035 33.830 ;
        RECT 92.000 33.300 93.860 33.575 ;
        RECT 106.880 33.385 107.580 45.435 ;
        RECT 92.000 33.130 96.465 33.300 ;
        RECT 92.000 31.720 92.895 33.130 ;
        RECT 93.235 32.260 93.405 32.590 ;
        RECT 93.575 32.560 95.615 32.730 ;
        RECT 93.575 32.120 95.615 32.290 ;
        RECT 95.785 32.260 95.955 32.590 ;
        RECT 96.295 31.720 96.465 33.130 ;
        RECT 80.210 31.635 90.040 31.690 ;
        RECT 92.000 31.560 96.465 31.720 ;
        RECT 97.210 33.215 107.580 33.385 ;
        RECT 97.210 31.805 97.380 33.215 ;
        RECT 97.720 32.345 97.890 32.675 ;
        RECT 98.105 32.645 106.145 32.815 ;
        RECT 98.105 32.205 106.145 32.375 ;
        RECT 106.360 32.345 106.530 32.675 ;
        RECT 106.870 31.805 107.580 33.215 ;
        RECT 97.210 31.690 107.580 31.805 ;
        RECT 109.000 57.485 109.865 58.140 ;
        RECT 114.195 57.975 124.580 58.145 ;
        RECT 109.000 57.315 113.455 57.485 ;
        RECT 109.000 52.055 109.885 57.315 ;
        RECT 110.565 56.745 112.605 56.915 ;
        RECT 110.225 52.685 110.395 56.685 ;
        RECT 112.775 52.685 112.945 56.685 ;
        RECT 110.565 52.455 112.605 52.625 ;
        RECT 113.285 52.055 113.455 57.315 ;
        RECT 114.195 54.485 114.365 57.975 ;
        RECT 114.995 57.465 122.995 57.635 ;
        RECT 114.765 55.210 114.935 57.250 ;
        RECT 123.055 55.210 123.225 57.250 ;
        RECT 114.995 54.825 122.995 54.995 ;
        RECT 123.625 54.485 124.580 57.975 ;
        RECT 114.195 54.315 124.580 54.485 ;
        RECT 123.625 54.025 124.580 54.315 ;
        RECT 109.000 51.885 113.455 52.055 ;
        RECT 109.000 46.625 109.885 51.885 ;
        RECT 110.565 51.315 112.605 51.485 ;
        RECT 110.225 47.255 110.395 51.255 ;
        RECT 112.775 47.255 112.945 51.255 ;
        RECT 110.565 47.025 112.605 47.195 ;
        RECT 113.285 46.625 113.455 51.885 ;
        RECT 114.195 53.855 124.580 54.025 ;
        RECT 114.195 50.595 114.365 53.855 ;
        RECT 115.090 53.285 123.130 53.455 ;
        RECT 114.705 51.225 114.875 53.225 ;
        RECT 123.345 51.225 123.515 53.225 ;
        RECT 115.090 50.995 123.130 51.165 ;
        RECT 123.855 50.595 124.580 53.855 ;
        RECT 114.195 50.425 124.580 50.595 ;
        RECT 114.195 47.165 114.365 50.425 ;
        RECT 115.090 49.855 123.130 50.025 ;
        RECT 114.705 47.795 114.875 49.795 ;
        RECT 123.345 47.795 123.515 49.795 ;
        RECT 115.090 47.565 123.130 47.735 ;
        RECT 123.855 47.165 124.580 50.425 ;
        RECT 114.195 46.995 124.580 47.165 ;
        RECT 119.905 46.715 124.580 46.995 ;
        RECT 109.000 46.455 113.455 46.625 ;
        RECT 109.000 41.195 109.885 46.455 ;
        RECT 110.565 45.885 112.605 46.055 ;
        RECT 110.225 41.825 110.395 45.825 ;
        RECT 112.775 41.825 112.945 45.825 ;
        RECT 110.565 41.595 112.605 41.765 ;
        RECT 113.285 41.195 113.455 46.455 ;
        RECT 109.000 41.025 113.455 41.195 ;
        RECT 109.000 35.765 109.885 41.025 ;
        RECT 110.565 40.455 112.605 40.625 ;
        RECT 110.225 36.395 110.395 40.395 ;
        RECT 112.775 36.395 112.945 40.395 ;
        RECT 110.565 36.165 112.605 36.335 ;
        RECT 113.285 35.765 113.455 41.025 ;
        RECT 109.000 35.595 113.455 35.765 ;
        RECT 114.190 46.545 124.580 46.715 ;
        RECT 114.190 41.285 114.360 46.545 ;
        RECT 115.085 45.975 119.125 46.145 ;
        RECT 114.700 41.915 114.870 45.915 ;
        RECT 119.340 41.915 119.510 45.915 ;
        RECT 119.850 45.435 124.580 46.545 ;
        RECT 115.085 41.685 119.125 41.855 ;
        RECT 119.850 41.285 120.020 45.435 ;
        RECT 114.190 41.115 120.020 41.285 ;
        RECT 114.190 35.855 114.360 41.115 ;
        RECT 115.085 40.545 119.125 40.715 ;
        RECT 114.700 36.485 114.870 40.485 ;
        RECT 119.340 36.485 119.510 40.485 ;
        RECT 115.085 36.255 119.125 36.425 ;
        RECT 119.850 35.855 120.020 41.115 ;
        RECT 120.535 45.360 122.285 45.435 ;
        RECT 120.535 38.870 120.705 45.360 ;
        RECT 121.245 44.850 121.575 45.020 ;
        RECT 121.105 39.595 121.275 44.635 ;
        RECT 121.545 39.595 121.715 44.635 ;
        RECT 121.245 39.210 121.575 39.380 ;
        RECT 122.115 38.870 122.285 45.360 ;
        RECT 120.535 38.700 122.285 38.870 ;
        RECT 114.190 35.685 120.020 35.855 ;
        RECT 109.000 35.325 110.860 35.595 ;
        RECT 109.000 35.155 113.460 35.325 ;
        RECT 109.000 33.745 110.890 35.155 ;
        RECT 111.230 34.285 111.400 34.615 ;
        RECT 111.570 34.585 112.610 34.755 ;
        RECT 111.570 34.145 112.610 34.315 ;
        RECT 112.780 34.285 112.950 34.615 ;
        RECT 113.290 33.745 113.460 35.155 ;
        RECT 109.000 33.575 113.460 33.745 ;
        RECT 114.205 35.240 120.035 35.410 ;
        RECT 114.205 33.830 114.375 35.240 ;
        RECT 114.715 34.370 114.885 34.700 ;
        RECT 115.100 34.670 119.140 34.840 ;
        RECT 115.100 34.230 119.140 34.400 ;
        RECT 119.355 34.370 119.525 34.700 ;
        RECT 119.865 33.830 120.035 35.240 ;
        RECT 114.205 33.660 120.035 33.830 ;
        RECT 109.000 33.300 110.860 33.575 ;
        RECT 123.880 33.385 124.580 45.435 ;
        RECT 109.000 33.130 113.465 33.300 ;
        RECT 109.000 31.720 109.895 33.130 ;
        RECT 110.235 32.260 110.405 32.590 ;
        RECT 110.575 32.560 112.615 32.730 ;
        RECT 110.575 32.120 112.615 32.290 ;
        RECT 112.785 32.260 112.955 32.590 ;
        RECT 113.295 31.720 113.465 33.130 ;
        RECT 97.210 31.635 107.040 31.690 ;
        RECT 109.000 31.560 113.465 31.720 ;
        RECT 114.210 33.215 124.580 33.385 ;
        RECT 114.210 31.805 114.380 33.215 ;
        RECT 114.720 32.345 114.890 32.675 ;
        RECT 115.105 32.645 123.145 32.815 ;
        RECT 115.105 32.205 123.145 32.375 ;
        RECT 123.360 32.345 123.530 32.675 ;
        RECT 123.870 31.805 124.580 33.215 ;
        RECT 114.210 31.690 124.580 31.805 ;
        RECT 126.000 57.485 126.865 58.140 ;
        RECT 131.195 57.975 141.580 58.145 ;
        RECT 126.000 57.315 130.455 57.485 ;
        RECT 126.000 52.055 126.885 57.315 ;
        RECT 127.565 56.745 129.605 56.915 ;
        RECT 127.225 52.685 127.395 56.685 ;
        RECT 129.775 52.685 129.945 56.685 ;
        RECT 127.565 52.455 129.605 52.625 ;
        RECT 130.285 52.055 130.455 57.315 ;
        RECT 131.195 54.485 131.365 57.975 ;
        RECT 131.995 57.465 139.995 57.635 ;
        RECT 131.765 55.210 131.935 57.250 ;
        RECT 140.055 55.210 140.225 57.250 ;
        RECT 131.995 54.825 139.995 54.995 ;
        RECT 140.625 54.485 141.580 57.975 ;
        RECT 131.195 54.315 141.580 54.485 ;
        RECT 140.625 54.025 141.580 54.315 ;
        RECT 126.000 51.885 130.455 52.055 ;
        RECT 126.000 46.625 126.885 51.885 ;
        RECT 127.565 51.315 129.605 51.485 ;
        RECT 127.225 47.255 127.395 51.255 ;
        RECT 129.775 47.255 129.945 51.255 ;
        RECT 127.565 47.025 129.605 47.195 ;
        RECT 130.285 46.625 130.455 51.885 ;
        RECT 131.195 53.855 141.580 54.025 ;
        RECT 131.195 50.595 131.365 53.855 ;
        RECT 132.090 53.285 140.130 53.455 ;
        RECT 131.705 51.225 131.875 53.225 ;
        RECT 140.345 51.225 140.515 53.225 ;
        RECT 132.090 50.995 140.130 51.165 ;
        RECT 140.855 50.595 141.580 53.855 ;
        RECT 131.195 50.425 141.580 50.595 ;
        RECT 131.195 47.165 131.365 50.425 ;
        RECT 132.090 49.855 140.130 50.025 ;
        RECT 131.705 47.795 131.875 49.795 ;
        RECT 140.345 47.795 140.515 49.795 ;
        RECT 132.090 47.565 140.130 47.735 ;
        RECT 140.855 47.165 141.580 50.425 ;
        RECT 131.195 46.995 141.580 47.165 ;
        RECT 136.905 46.715 141.580 46.995 ;
        RECT 126.000 46.455 130.455 46.625 ;
        RECT 126.000 41.195 126.885 46.455 ;
        RECT 127.565 45.885 129.605 46.055 ;
        RECT 127.225 41.825 127.395 45.825 ;
        RECT 129.775 41.825 129.945 45.825 ;
        RECT 127.565 41.595 129.605 41.765 ;
        RECT 130.285 41.195 130.455 46.455 ;
        RECT 126.000 41.025 130.455 41.195 ;
        RECT 126.000 35.765 126.885 41.025 ;
        RECT 127.565 40.455 129.605 40.625 ;
        RECT 127.225 36.395 127.395 40.395 ;
        RECT 129.775 36.395 129.945 40.395 ;
        RECT 127.565 36.165 129.605 36.335 ;
        RECT 130.285 35.765 130.455 41.025 ;
        RECT 126.000 35.595 130.455 35.765 ;
        RECT 131.190 46.545 141.580 46.715 ;
        RECT 131.190 41.285 131.360 46.545 ;
        RECT 132.085 45.975 136.125 46.145 ;
        RECT 131.700 41.915 131.870 45.915 ;
        RECT 136.340 41.915 136.510 45.915 ;
        RECT 136.850 45.435 141.580 46.545 ;
        RECT 132.085 41.685 136.125 41.855 ;
        RECT 136.850 41.285 137.020 45.435 ;
        RECT 131.190 41.115 137.020 41.285 ;
        RECT 131.190 35.855 131.360 41.115 ;
        RECT 132.085 40.545 136.125 40.715 ;
        RECT 131.700 36.485 131.870 40.485 ;
        RECT 136.340 36.485 136.510 40.485 ;
        RECT 132.085 36.255 136.125 36.425 ;
        RECT 136.850 35.855 137.020 41.115 ;
        RECT 137.535 45.360 139.285 45.435 ;
        RECT 137.535 38.870 137.705 45.360 ;
        RECT 138.245 44.850 138.575 45.020 ;
        RECT 138.105 39.595 138.275 44.635 ;
        RECT 138.545 39.595 138.715 44.635 ;
        RECT 138.245 39.210 138.575 39.380 ;
        RECT 139.115 38.870 139.285 45.360 ;
        RECT 137.535 38.700 139.285 38.870 ;
        RECT 131.190 35.685 137.020 35.855 ;
        RECT 126.000 35.325 127.860 35.595 ;
        RECT 126.000 35.155 130.460 35.325 ;
        RECT 126.000 33.745 127.890 35.155 ;
        RECT 128.230 34.285 128.400 34.615 ;
        RECT 128.570 34.585 129.610 34.755 ;
        RECT 128.570 34.145 129.610 34.315 ;
        RECT 129.780 34.285 129.950 34.615 ;
        RECT 130.290 33.745 130.460 35.155 ;
        RECT 126.000 33.575 130.460 33.745 ;
        RECT 131.205 35.240 137.035 35.410 ;
        RECT 131.205 33.830 131.375 35.240 ;
        RECT 131.715 34.370 131.885 34.700 ;
        RECT 132.100 34.670 136.140 34.840 ;
        RECT 132.100 34.230 136.140 34.400 ;
        RECT 136.355 34.370 136.525 34.700 ;
        RECT 136.865 33.830 137.035 35.240 ;
        RECT 131.205 33.660 137.035 33.830 ;
        RECT 126.000 33.300 127.860 33.575 ;
        RECT 140.880 33.385 141.580 45.435 ;
        RECT 126.000 33.130 130.465 33.300 ;
        RECT 126.000 31.720 126.895 33.130 ;
        RECT 127.235 32.260 127.405 32.590 ;
        RECT 127.575 32.560 129.615 32.730 ;
        RECT 127.575 32.120 129.615 32.290 ;
        RECT 129.785 32.260 129.955 32.590 ;
        RECT 130.295 31.720 130.465 33.130 ;
        RECT 114.210 31.635 124.040 31.690 ;
        RECT 126.000 31.560 130.465 31.720 ;
        RECT 131.210 33.215 141.580 33.385 ;
        RECT 131.210 31.805 131.380 33.215 ;
        RECT 131.720 32.345 131.890 32.675 ;
        RECT 132.105 32.645 140.145 32.815 ;
        RECT 132.105 32.205 140.145 32.375 ;
        RECT 140.360 32.345 140.530 32.675 ;
        RECT 140.870 31.805 141.580 33.215 ;
        RECT 131.210 31.690 141.580 31.805 ;
        RECT 143.000 57.485 143.865 58.140 ;
        RECT 148.195 57.975 158.580 58.145 ;
        RECT 143.000 57.315 147.455 57.485 ;
        RECT 143.000 52.055 143.885 57.315 ;
        RECT 144.565 56.745 146.605 56.915 ;
        RECT 144.225 52.685 144.395 56.685 ;
        RECT 146.775 52.685 146.945 56.685 ;
        RECT 144.565 52.455 146.605 52.625 ;
        RECT 147.285 52.055 147.455 57.315 ;
        RECT 148.195 54.485 148.365 57.975 ;
        RECT 148.995 57.465 156.995 57.635 ;
        RECT 148.765 55.210 148.935 57.250 ;
        RECT 157.055 55.210 157.225 57.250 ;
        RECT 148.995 54.825 156.995 54.995 ;
        RECT 157.625 54.485 158.580 57.975 ;
        RECT 148.195 54.315 158.580 54.485 ;
        RECT 157.625 54.025 158.580 54.315 ;
        RECT 143.000 51.885 147.455 52.055 ;
        RECT 143.000 46.625 143.885 51.885 ;
        RECT 144.565 51.315 146.605 51.485 ;
        RECT 144.225 47.255 144.395 51.255 ;
        RECT 146.775 47.255 146.945 51.255 ;
        RECT 144.565 47.025 146.605 47.195 ;
        RECT 147.285 46.625 147.455 51.885 ;
        RECT 148.195 53.855 158.580 54.025 ;
        RECT 148.195 50.595 148.365 53.855 ;
        RECT 149.090 53.285 157.130 53.455 ;
        RECT 148.705 51.225 148.875 53.225 ;
        RECT 157.345 51.225 157.515 53.225 ;
        RECT 149.090 50.995 157.130 51.165 ;
        RECT 157.855 50.595 158.580 53.855 ;
        RECT 148.195 50.425 158.580 50.595 ;
        RECT 148.195 47.165 148.365 50.425 ;
        RECT 149.090 49.855 157.130 50.025 ;
        RECT 148.705 47.795 148.875 49.795 ;
        RECT 157.345 47.795 157.515 49.795 ;
        RECT 149.090 47.565 157.130 47.735 ;
        RECT 157.855 47.165 158.580 50.425 ;
        RECT 148.195 46.995 158.580 47.165 ;
        RECT 153.905 46.715 158.580 46.995 ;
        RECT 143.000 46.455 147.455 46.625 ;
        RECT 143.000 41.195 143.885 46.455 ;
        RECT 144.565 45.885 146.605 46.055 ;
        RECT 144.225 41.825 144.395 45.825 ;
        RECT 146.775 41.825 146.945 45.825 ;
        RECT 144.565 41.595 146.605 41.765 ;
        RECT 147.285 41.195 147.455 46.455 ;
        RECT 143.000 41.025 147.455 41.195 ;
        RECT 143.000 35.765 143.885 41.025 ;
        RECT 144.565 40.455 146.605 40.625 ;
        RECT 144.225 36.395 144.395 40.395 ;
        RECT 146.775 36.395 146.945 40.395 ;
        RECT 144.565 36.165 146.605 36.335 ;
        RECT 147.285 35.765 147.455 41.025 ;
        RECT 143.000 35.595 147.455 35.765 ;
        RECT 148.190 46.545 158.580 46.715 ;
        RECT 148.190 41.285 148.360 46.545 ;
        RECT 149.085 45.975 153.125 46.145 ;
        RECT 148.700 41.915 148.870 45.915 ;
        RECT 153.340 41.915 153.510 45.915 ;
        RECT 153.850 45.435 158.580 46.545 ;
        RECT 149.085 41.685 153.125 41.855 ;
        RECT 153.850 41.285 154.020 45.435 ;
        RECT 148.190 41.115 154.020 41.285 ;
        RECT 148.190 35.855 148.360 41.115 ;
        RECT 149.085 40.545 153.125 40.715 ;
        RECT 148.700 36.485 148.870 40.485 ;
        RECT 153.340 36.485 153.510 40.485 ;
        RECT 149.085 36.255 153.125 36.425 ;
        RECT 153.850 35.855 154.020 41.115 ;
        RECT 154.535 45.360 156.285 45.435 ;
        RECT 154.535 38.870 154.705 45.360 ;
        RECT 155.245 44.850 155.575 45.020 ;
        RECT 155.105 39.595 155.275 44.635 ;
        RECT 155.545 39.595 155.715 44.635 ;
        RECT 155.245 39.210 155.575 39.380 ;
        RECT 156.115 38.870 156.285 45.360 ;
        RECT 154.535 38.700 156.285 38.870 ;
        RECT 148.190 35.685 154.020 35.855 ;
        RECT 143.000 35.325 144.860 35.595 ;
        RECT 143.000 35.155 147.460 35.325 ;
        RECT 143.000 33.745 144.890 35.155 ;
        RECT 145.230 34.285 145.400 34.615 ;
        RECT 145.570 34.585 146.610 34.755 ;
        RECT 145.570 34.145 146.610 34.315 ;
        RECT 146.780 34.285 146.950 34.615 ;
        RECT 147.290 33.745 147.460 35.155 ;
        RECT 143.000 33.575 147.460 33.745 ;
        RECT 148.205 35.240 154.035 35.410 ;
        RECT 148.205 33.830 148.375 35.240 ;
        RECT 148.715 34.370 148.885 34.700 ;
        RECT 149.100 34.670 153.140 34.840 ;
        RECT 149.100 34.230 153.140 34.400 ;
        RECT 153.355 34.370 153.525 34.700 ;
        RECT 153.865 33.830 154.035 35.240 ;
        RECT 148.205 33.660 154.035 33.830 ;
        RECT 143.000 33.300 144.860 33.575 ;
        RECT 157.880 33.385 158.580 45.435 ;
        RECT 143.000 33.130 147.465 33.300 ;
        RECT 143.000 31.720 143.895 33.130 ;
        RECT 144.235 32.260 144.405 32.590 ;
        RECT 144.575 32.560 146.615 32.730 ;
        RECT 144.575 32.120 146.615 32.290 ;
        RECT 146.785 32.260 146.955 32.590 ;
        RECT 147.295 31.720 147.465 33.130 ;
        RECT 131.210 31.635 141.040 31.690 ;
        RECT 143.000 31.560 147.465 31.720 ;
        RECT 148.210 33.215 158.580 33.385 ;
        RECT 148.210 31.805 148.380 33.215 ;
        RECT 148.720 32.345 148.890 32.675 ;
        RECT 149.105 32.645 157.145 32.815 ;
        RECT 149.105 32.205 157.145 32.375 ;
        RECT 157.360 32.345 157.530 32.675 ;
        RECT 157.870 31.805 158.580 33.215 ;
        RECT 148.210 31.690 158.580 31.805 ;
        RECT 148.210 31.635 158.040 31.690 ;
        RECT 75.725 31.550 79.465 31.560 ;
        RECT 92.725 31.550 96.465 31.560 ;
        RECT 109.725 31.550 113.465 31.560 ;
        RECT 126.725 31.550 130.465 31.560 ;
        RECT 143.725 31.550 147.465 31.560 ;
        RECT 54.500 29.770 54.670 29.975 ;
        RECT 55.210 29.575 55.380 30.775 ;
        RECT 55.550 30.395 56.120 30.605 ;
        RECT 56.290 30.395 56.935 30.605 ;
        RECT 57.105 30.325 57.625 30.865 ;
        RECT 55.610 30.055 56.780 30.225 ;
        RECT 57.795 30.155 58.315 30.695 ;
        RECT 55.610 29.575 55.940 30.055 ;
        RECT 56.110 29.405 56.280 29.875 ;
        RECT 56.450 29.590 56.780 30.055 ;
        RECT 57.105 29.405 58.315 30.155 ;
        RECT 22.520 29.235 58.400 29.405 ;
        RECT 22.605 28.485 23.815 29.235 ;
        RECT 22.605 27.945 23.125 28.485 ;
        RECT 23.990 28.395 24.250 29.235 ;
        RECT 24.425 28.490 24.680 29.065 ;
        RECT 24.850 28.855 25.180 29.235 ;
        RECT 25.395 28.685 25.565 29.065 ;
        RECT 24.850 28.515 25.565 28.685 ;
        RECT 23.295 27.775 23.815 28.315 ;
        RECT 22.605 26.685 23.815 27.775 ;
        RECT 23.990 26.685 24.250 27.835 ;
        RECT 24.425 27.760 24.595 28.490 ;
        RECT 24.850 28.325 25.020 28.515 ;
        RECT 26.750 28.495 27.005 29.065 ;
        RECT 27.175 28.835 27.505 29.235 ;
        RECT 27.930 28.700 28.460 29.065 ;
        RECT 28.650 28.895 28.925 29.065 ;
        RECT 28.645 28.725 28.925 28.895 ;
        RECT 27.930 28.665 28.105 28.700 ;
        RECT 27.175 28.495 28.105 28.665 ;
        RECT 24.765 27.995 25.020 28.325 ;
        RECT 24.850 27.785 25.020 27.995 ;
        RECT 25.300 27.965 25.655 28.335 ;
        RECT 26.750 27.825 26.920 28.495 ;
        RECT 27.175 28.325 27.345 28.495 ;
        RECT 27.090 27.995 27.345 28.325 ;
        RECT 27.570 27.995 27.765 28.325 ;
        RECT 24.425 26.855 24.680 27.760 ;
        RECT 24.850 27.615 25.565 27.785 ;
        RECT 24.850 26.685 25.180 27.445 ;
        RECT 25.395 26.855 25.565 27.615 ;
        RECT 26.750 26.855 27.085 27.825 ;
        RECT 27.255 26.685 27.425 27.825 ;
        RECT 27.595 27.025 27.765 27.995 ;
        RECT 27.935 27.365 28.105 28.495 ;
        RECT 28.275 27.705 28.445 28.505 ;
        RECT 28.650 27.905 28.925 28.725 ;
        RECT 29.095 27.705 29.285 29.065 ;
        RECT 29.465 28.700 29.975 29.235 ;
        RECT 30.195 28.425 30.440 29.030 ;
        RECT 30.885 28.465 34.395 29.235 ;
        RECT 34.565 28.485 35.775 29.235 ;
        RECT 35.995 28.580 36.325 29.015 ;
        RECT 36.495 28.625 36.665 29.235 ;
        RECT 35.945 28.495 36.325 28.580 ;
        RECT 36.835 28.495 37.165 29.020 ;
        RECT 37.425 28.705 37.635 29.235 ;
        RECT 37.910 28.785 38.695 28.955 ;
        RECT 38.865 28.785 39.270 28.955 ;
        RECT 29.485 28.255 30.715 28.425 ;
        RECT 28.275 27.535 29.285 27.705 ;
        RECT 29.455 27.690 30.205 27.880 ;
        RECT 27.935 27.195 29.060 27.365 ;
        RECT 29.455 27.025 29.625 27.690 ;
        RECT 30.375 27.445 30.715 28.255 ;
        RECT 30.885 27.945 32.535 28.465 ;
        RECT 32.705 27.775 34.395 28.295 ;
        RECT 34.565 27.945 35.085 28.485 ;
        RECT 35.945 28.455 36.170 28.495 ;
        RECT 35.255 27.775 35.775 28.315 ;
        RECT 27.595 26.855 29.625 27.025 ;
        RECT 29.795 26.685 29.965 27.445 ;
        RECT 30.200 27.035 30.715 27.445 ;
        RECT 30.885 26.685 34.395 27.775 ;
        RECT 34.565 26.685 35.775 27.775 ;
        RECT 35.945 27.875 36.115 28.455 ;
        RECT 36.835 28.325 37.035 28.495 ;
        RECT 37.910 28.325 38.080 28.785 ;
        RECT 36.285 27.995 37.035 28.325 ;
        RECT 37.205 27.995 38.080 28.325 ;
        RECT 35.945 27.825 36.160 27.875 ;
        RECT 35.945 27.745 36.335 27.825 ;
        RECT 36.005 26.900 36.335 27.745 ;
        RECT 36.845 27.790 37.035 27.995 ;
        RECT 36.505 26.685 36.675 27.695 ;
        RECT 36.845 27.415 37.740 27.790 ;
        RECT 36.845 26.855 37.185 27.415 ;
        RECT 37.415 26.685 37.730 27.185 ;
        RECT 37.910 27.155 38.080 27.995 ;
        RECT 38.250 28.285 38.715 28.615 ;
        RECT 39.100 28.555 39.270 28.785 ;
        RECT 39.450 28.735 39.820 29.235 ;
        RECT 40.140 28.785 40.815 28.955 ;
        RECT 41.010 28.785 41.345 28.955 ;
        RECT 38.250 27.325 38.570 28.285 ;
        RECT 39.100 28.255 39.930 28.555 ;
        RECT 38.740 27.355 38.930 28.075 ;
        RECT 39.100 27.185 39.270 28.255 ;
        RECT 39.730 28.225 39.930 28.255 ;
        RECT 39.440 28.005 39.610 28.075 ;
        RECT 40.140 28.005 40.310 28.785 ;
        RECT 41.175 28.645 41.345 28.785 ;
        RECT 41.515 28.775 41.765 29.235 ;
        RECT 39.440 27.835 40.310 28.005 ;
        RECT 40.480 28.365 41.005 28.585 ;
        RECT 41.175 28.515 41.400 28.645 ;
        RECT 39.440 27.745 39.950 27.835 ;
        RECT 37.910 26.985 38.795 27.155 ;
        RECT 39.020 26.855 39.270 27.185 ;
        RECT 39.440 26.685 39.610 27.485 ;
        RECT 39.780 27.130 39.950 27.745 ;
        RECT 40.480 27.665 40.650 28.365 ;
        RECT 40.120 27.300 40.650 27.665 ;
        RECT 40.820 27.600 41.060 28.195 ;
        RECT 41.230 27.410 41.400 28.515 ;
        RECT 41.570 27.655 41.850 28.605 ;
        RECT 41.095 27.280 41.400 27.410 ;
        RECT 39.780 26.960 40.885 27.130 ;
        RECT 41.095 26.855 41.345 27.280 ;
        RECT 41.515 26.685 41.780 27.145 ;
        RECT 42.020 26.855 42.205 28.975 ;
        RECT 42.375 28.855 42.705 29.235 ;
        RECT 42.875 28.685 43.045 28.975 ;
        RECT 42.380 28.515 43.045 28.685 ;
        RECT 42.380 27.525 42.610 28.515 ;
        RECT 43.310 28.495 43.565 29.065 ;
        RECT 43.735 28.835 44.065 29.235 ;
        RECT 44.490 28.700 45.020 29.065 ;
        RECT 44.490 28.665 44.665 28.700 ;
        RECT 43.735 28.495 44.665 28.665 ;
        RECT 42.780 27.695 43.130 28.345 ;
        RECT 43.310 27.825 43.480 28.495 ;
        RECT 43.735 28.325 43.905 28.495 ;
        RECT 43.650 27.995 43.905 28.325 ;
        RECT 44.130 27.995 44.325 28.325 ;
        RECT 42.380 27.355 43.045 27.525 ;
        RECT 42.375 26.685 42.705 27.185 ;
        RECT 42.875 26.855 43.045 27.355 ;
        RECT 43.310 26.855 43.645 27.825 ;
        RECT 43.815 26.685 43.985 27.825 ;
        RECT 44.155 27.025 44.325 27.995 ;
        RECT 44.495 27.365 44.665 28.495 ;
        RECT 44.835 27.705 45.005 28.505 ;
        RECT 45.210 28.215 45.485 29.065 ;
        RECT 45.205 28.045 45.485 28.215 ;
        RECT 45.210 27.905 45.485 28.045 ;
        RECT 45.655 27.705 45.845 29.065 ;
        RECT 46.025 28.700 46.535 29.235 ;
        RECT 46.755 28.425 47.000 29.030 ;
        RECT 48.365 28.510 48.655 29.235 ;
        RECT 48.825 28.495 49.210 29.065 ;
        RECT 49.380 28.775 49.705 29.235 ;
        RECT 50.225 28.605 50.505 29.065 ;
        RECT 46.045 28.255 47.275 28.425 ;
        RECT 44.835 27.535 45.845 27.705 ;
        RECT 46.015 27.690 46.765 27.880 ;
        RECT 44.495 27.195 45.620 27.365 ;
        RECT 46.015 27.025 46.185 27.690 ;
        RECT 46.935 27.445 47.275 28.255 ;
        RECT 44.155 26.855 46.185 27.025 ;
        RECT 46.355 26.685 46.525 27.445 ;
        RECT 46.760 27.035 47.275 27.445 ;
        RECT 48.365 26.685 48.655 27.850 ;
        RECT 48.825 27.825 49.105 28.495 ;
        RECT 49.380 28.435 50.505 28.605 ;
        RECT 49.380 28.325 49.830 28.435 ;
        RECT 49.275 27.995 49.830 28.325 ;
        RECT 50.695 28.265 51.095 29.065 ;
        RECT 51.495 28.775 51.765 29.235 ;
        RECT 51.935 28.605 52.220 29.065 ;
        RECT 48.825 26.855 49.210 27.825 ;
        RECT 49.380 27.535 49.830 27.995 ;
        RECT 50.000 27.705 51.095 28.265 ;
        RECT 49.380 27.315 50.505 27.535 ;
        RECT 49.380 26.685 49.705 27.145 ;
        RECT 50.225 26.855 50.505 27.315 ;
        RECT 50.695 26.855 51.095 27.705 ;
        RECT 51.265 28.435 52.220 28.605 ;
        RECT 53.425 28.605 53.765 29.065 ;
        RECT 53.935 28.775 54.105 29.235 ;
        RECT 54.735 28.800 55.095 29.065 ;
        RECT 54.740 28.795 55.095 28.800 ;
        RECT 54.745 28.785 55.095 28.795 ;
        RECT 54.750 28.780 55.095 28.785 ;
        RECT 54.755 28.770 55.095 28.780 ;
        RECT 55.335 28.775 55.505 29.235 ;
        RECT 54.760 28.765 55.095 28.770 ;
        RECT 54.770 28.755 55.095 28.765 ;
        RECT 54.780 28.745 55.095 28.755 ;
        RECT 54.275 28.605 54.605 28.685 ;
        RECT 51.265 27.535 51.475 28.435 ;
        RECT 53.425 28.415 54.605 28.605 ;
        RECT 54.795 28.605 55.095 28.745 ;
        RECT 54.795 28.415 55.505 28.605 ;
        RECT 51.645 27.705 52.335 28.265 ;
        RECT 53.425 28.045 53.755 28.245 ;
        RECT 54.065 28.225 54.395 28.245 ;
        RECT 53.945 28.045 54.395 28.225 ;
        RECT 53.425 27.705 53.655 28.045 ;
        RECT 51.265 27.315 52.220 27.535 ;
        RECT 51.495 26.685 51.765 27.145 ;
        RECT 51.935 26.855 52.220 27.315 ;
        RECT 53.435 26.685 53.765 27.405 ;
        RECT 53.945 26.930 54.160 28.045 ;
        RECT 54.565 28.015 55.035 28.245 ;
        RECT 55.220 27.845 55.505 28.415 ;
        RECT 55.675 28.290 56.015 29.065 ;
        RECT 57.105 28.485 58.315 29.235 ;
        RECT 89.625 29.165 90.100 29.180 ;
        RECT 106.625 29.165 107.100 29.180 ;
        RECT 123.625 29.165 124.100 29.180 ;
        RECT 140.625 29.165 141.100 29.180 ;
        RECT 157.625 29.165 158.100 29.180 ;
        RECT 89.625 29.145 90.580 29.165 ;
        RECT 106.625 29.145 107.580 29.165 ;
        RECT 123.625 29.145 124.580 29.165 ;
        RECT 140.625 29.145 141.580 29.165 ;
        RECT 157.625 29.145 158.580 29.165 ;
        RECT 54.355 27.630 55.505 27.845 ;
        RECT 54.355 26.855 54.685 27.630 ;
        RECT 54.855 26.685 55.565 27.460 ;
        RECT 55.735 26.855 56.015 28.290 ;
        RECT 57.105 27.775 57.625 28.315 ;
        RECT 57.795 27.945 58.315 28.485 ;
        RECT 75.000 28.485 75.865 29.140 ;
        RECT 80.195 28.975 90.580 29.145 ;
        RECT 75.000 28.315 79.455 28.485 ;
        RECT 57.105 26.685 58.315 27.775 ;
        RECT 22.520 26.515 58.400 26.685 ;
        RECT 22.605 25.425 23.815 26.515 ;
        RECT 23.985 26.080 29.330 26.515 ;
        RECT 22.605 24.715 23.125 25.255 ;
        RECT 23.295 24.885 23.815 25.425 ;
        RECT 22.605 23.965 23.815 24.715 ;
        RECT 25.570 24.510 25.910 25.340 ;
        RECT 27.390 24.830 27.740 26.080 ;
        RECT 29.505 25.425 33.015 26.515 ;
        RECT 29.505 24.735 31.155 25.255 ;
        RECT 31.325 24.905 33.015 25.425 ;
        RECT 33.735 25.585 33.905 26.345 ;
        RECT 34.120 25.755 34.450 26.515 ;
        RECT 33.735 25.415 34.450 25.585 ;
        RECT 34.620 25.440 34.875 26.345 ;
        RECT 33.645 24.865 34.000 25.235 ;
        RECT 34.280 25.205 34.450 25.415 ;
        RECT 34.280 24.875 34.535 25.205 ;
        RECT 23.985 23.965 29.330 24.510 ;
        RECT 29.505 23.965 33.015 24.735 ;
        RECT 34.280 24.685 34.450 24.875 ;
        RECT 34.705 24.710 34.875 25.440 ;
        RECT 35.050 25.365 35.310 26.515 ;
        RECT 35.485 25.350 35.775 26.515 ;
        RECT 36.410 25.365 36.670 26.515 ;
        RECT 36.845 25.440 37.100 26.345 ;
        RECT 37.270 25.755 37.600 26.515 ;
        RECT 37.815 25.585 37.985 26.345 ;
        RECT 38.335 25.845 38.505 26.345 ;
        RECT 38.675 26.015 39.005 26.515 ;
        RECT 38.335 25.675 39.000 25.845 ;
        RECT 33.735 24.515 34.450 24.685 ;
        RECT 33.735 24.135 33.905 24.515 ;
        RECT 34.120 23.965 34.450 24.345 ;
        RECT 34.620 24.135 34.875 24.710 ;
        RECT 35.050 23.965 35.310 24.805 ;
        RECT 35.485 23.965 35.775 24.690 ;
        RECT 36.410 23.965 36.670 24.805 ;
        RECT 36.845 24.710 37.015 25.440 ;
        RECT 37.270 25.415 37.985 25.585 ;
        RECT 37.270 25.205 37.440 25.415 ;
        RECT 37.185 24.875 37.440 25.205 ;
        RECT 36.845 24.135 37.100 24.710 ;
        RECT 37.270 24.685 37.440 24.875 ;
        RECT 37.720 24.865 38.075 25.235 ;
        RECT 38.250 24.855 38.600 25.505 ;
        RECT 38.770 24.685 39.000 25.675 ;
        RECT 37.270 24.515 37.985 24.685 ;
        RECT 37.270 23.965 37.600 24.345 ;
        RECT 37.815 24.135 37.985 24.515 ;
        RECT 38.335 24.515 39.000 24.685 ;
        RECT 38.335 24.225 38.505 24.515 ;
        RECT 38.675 23.965 39.005 24.345 ;
        RECT 39.175 24.225 39.360 26.345 ;
        RECT 39.600 26.055 39.865 26.515 ;
        RECT 40.035 25.920 40.285 26.345 ;
        RECT 40.495 26.070 41.600 26.240 ;
        RECT 39.980 25.790 40.285 25.920 ;
        RECT 39.530 24.595 39.810 25.545 ;
        RECT 39.980 24.685 40.150 25.790 ;
        RECT 40.320 25.005 40.560 25.600 ;
        RECT 40.730 25.535 41.260 25.900 ;
        RECT 40.730 24.835 40.900 25.535 ;
        RECT 41.430 25.455 41.600 26.070 ;
        RECT 41.770 25.715 41.940 26.515 ;
        RECT 42.110 26.015 42.360 26.345 ;
        RECT 42.585 26.045 43.470 26.215 ;
        RECT 41.430 25.365 41.940 25.455 ;
        RECT 39.980 24.555 40.205 24.685 ;
        RECT 40.375 24.615 40.900 24.835 ;
        RECT 41.070 25.195 41.940 25.365 ;
        RECT 39.615 23.965 39.865 24.425 ;
        RECT 40.035 24.415 40.205 24.555 ;
        RECT 41.070 24.415 41.240 25.195 ;
        RECT 41.770 25.125 41.940 25.195 ;
        RECT 41.450 24.945 41.650 24.975 ;
        RECT 42.110 24.945 42.280 26.015 ;
        RECT 42.450 25.125 42.640 25.845 ;
        RECT 41.450 24.645 42.280 24.945 ;
        RECT 42.810 24.915 43.130 25.875 ;
        RECT 40.035 24.245 40.370 24.415 ;
        RECT 40.565 24.245 41.240 24.415 ;
        RECT 41.560 23.965 41.930 24.465 ;
        RECT 42.110 24.415 42.280 24.645 ;
        RECT 42.665 24.585 43.130 24.915 ;
        RECT 43.300 25.205 43.470 26.045 ;
        RECT 43.650 26.015 43.965 26.515 ;
        RECT 44.195 25.785 44.535 26.345 ;
        RECT 43.640 25.410 44.535 25.785 ;
        RECT 44.705 25.505 44.875 26.515 ;
        RECT 44.345 25.205 44.535 25.410 ;
        RECT 45.045 25.455 45.375 26.300 ;
        RECT 45.045 25.375 45.435 25.455 ;
        RECT 45.220 25.325 45.435 25.375 ;
        RECT 45.610 25.365 45.870 26.515 ;
        RECT 46.045 25.440 46.300 26.345 ;
        RECT 46.470 25.755 46.800 26.515 ;
        RECT 47.015 25.585 47.185 26.345 ;
        RECT 43.300 24.875 44.175 25.205 ;
        RECT 44.345 24.875 45.095 25.205 ;
        RECT 43.300 24.415 43.470 24.875 ;
        RECT 44.345 24.705 44.545 24.875 ;
        RECT 45.265 24.745 45.435 25.325 ;
        RECT 45.210 24.705 45.435 24.745 ;
        RECT 42.110 24.245 42.515 24.415 ;
        RECT 42.685 24.245 43.470 24.415 ;
        RECT 43.745 23.965 43.955 24.495 ;
        RECT 44.215 24.180 44.545 24.705 ;
        RECT 45.055 24.620 45.435 24.705 ;
        RECT 44.715 23.965 44.885 24.575 ;
        RECT 45.055 24.185 45.385 24.620 ;
        RECT 45.610 23.965 45.870 24.805 ;
        RECT 46.045 24.710 46.215 25.440 ;
        RECT 46.470 25.415 47.185 25.585 ;
        RECT 46.470 25.205 46.640 25.415 ;
        RECT 48.365 25.350 48.655 26.515 ;
        RECT 49.835 25.585 50.005 26.345 ;
        RECT 50.220 25.755 50.550 26.515 ;
        RECT 49.835 25.415 50.550 25.585 ;
        RECT 50.720 25.440 50.975 26.345 ;
        RECT 46.385 24.875 46.640 25.205 ;
        RECT 46.045 24.135 46.300 24.710 ;
        RECT 46.470 24.685 46.640 24.875 ;
        RECT 46.920 24.865 47.275 25.235 ;
        RECT 49.745 24.865 50.100 25.235 ;
        RECT 50.380 25.205 50.550 25.415 ;
        RECT 50.380 24.875 50.635 25.205 ;
        RECT 46.470 24.515 47.185 24.685 ;
        RECT 46.470 23.965 46.800 24.345 ;
        RECT 47.015 24.135 47.185 24.515 ;
        RECT 48.365 23.965 48.655 24.690 ;
        RECT 50.380 24.685 50.550 24.875 ;
        RECT 50.805 24.710 50.975 25.440 ;
        RECT 51.150 25.365 51.410 26.515 ;
        RECT 51.585 25.440 51.855 26.345 ;
        RECT 52.025 25.755 52.355 26.515 ;
        RECT 52.535 25.585 52.715 26.345 ;
        RECT 53.975 25.895 54.145 26.325 ;
        RECT 54.315 26.065 54.645 26.515 ;
        RECT 53.975 25.665 54.650 25.895 ;
        RECT 49.835 24.515 50.550 24.685 ;
        RECT 49.835 24.135 50.005 24.515 ;
        RECT 50.220 23.965 50.550 24.345 ;
        RECT 50.720 24.135 50.975 24.710 ;
        RECT 51.150 23.965 51.410 24.805 ;
        RECT 51.585 24.640 51.765 25.440 ;
        RECT 52.040 25.415 52.715 25.585 ;
        RECT 52.040 25.270 52.210 25.415 ;
        RECT 51.935 24.940 52.210 25.270 ;
        RECT 52.040 24.685 52.210 24.940 ;
        RECT 52.435 24.865 52.775 25.235 ;
        RECT 51.585 24.135 51.845 24.640 ;
        RECT 52.040 24.515 52.705 24.685 ;
        RECT 53.945 24.645 54.245 25.495 ;
        RECT 54.415 25.015 54.650 25.665 ;
        RECT 54.820 25.355 55.105 26.300 ;
        RECT 55.285 26.045 55.970 26.515 ;
        RECT 55.280 25.525 55.975 25.835 ;
        RECT 56.150 25.460 56.455 26.245 ;
        RECT 54.820 25.205 55.680 25.355 ;
        RECT 54.820 25.185 56.105 25.205 ;
        RECT 54.415 24.685 54.950 25.015 ;
        RECT 55.120 24.825 56.105 25.185 ;
        RECT 54.415 24.535 54.635 24.685 ;
        RECT 52.025 23.965 52.355 24.345 ;
        RECT 52.535 24.135 52.705 24.515 ;
        RECT 53.890 23.965 54.225 24.470 ;
        RECT 54.395 24.160 54.635 24.535 ;
        RECT 55.120 24.490 55.290 24.825 ;
        RECT 56.280 24.655 56.455 25.460 ;
        RECT 57.105 25.425 58.315 26.515 ;
        RECT 57.105 24.885 57.625 25.425 ;
        RECT 57.795 24.715 58.315 25.255 ;
        RECT 54.915 24.295 55.290 24.490 ;
        RECT 54.915 24.150 55.085 24.295 ;
        RECT 55.650 23.965 56.045 24.460 ;
        RECT 56.215 24.135 56.455 24.655 ;
        RECT 57.105 23.965 58.315 24.715 ;
        RECT 22.520 23.795 58.400 23.965 ;
        RECT 75.000 23.055 75.885 28.315 ;
        RECT 76.565 27.745 78.605 27.915 ;
        RECT 76.225 23.685 76.395 27.685 ;
        RECT 78.775 23.685 78.945 27.685 ;
        RECT 76.565 23.455 78.605 23.625 ;
        RECT 79.285 23.055 79.455 28.315 ;
        RECT 80.195 25.485 80.365 28.975 ;
        RECT 80.995 28.465 88.995 28.635 ;
        RECT 80.765 26.210 80.935 28.250 ;
        RECT 89.055 26.210 89.225 28.250 ;
        RECT 80.995 25.825 88.995 25.995 ;
        RECT 89.625 25.485 90.580 28.975 ;
        RECT 80.195 25.315 90.580 25.485 ;
        RECT 89.625 25.025 90.580 25.315 ;
        RECT 75.000 22.885 79.455 23.055 ;
        RECT 75.000 17.625 75.885 22.885 ;
        RECT 76.565 22.315 78.605 22.485 ;
        RECT 76.225 18.255 76.395 22.255 ;
        RECT 78.775 18.255 78.945 22.255 ;
        RECT 76.565 18.025 78.605 18.195 ;
        RECT 79.285 17.625 79.455 22.885 ;
        RECT 80.195 24.855 90.580 25.025 ;
        RECT 80.195 21.595 80.365 24.855 ;
        RECT 81.090 24.285 89.130 24.455 ;
        RECT 80.705 22.225 80.875 24.225 ;
        RECT 89.345 22.225 89.515 24.225 ;
        RECT 81.090 21.995 89.130 22.165 ;
        RECT 89.855 21.595 90.580 24.855 ;
        RECT 80.195 21.425 90.580 21.595 ;
        RECT 80.195 18.165 80.365 21.425 ;
        RECT 81.090 20.855 89.130 21.025 ;
        RECT 80.705 18.795 80.875 20.795 ;
        RECT 89.345 18.795 89.515 20.795 ;
        RECT 81.090 18.565 89.130 18.735 ;
        RECT 89.855 18.165 90.580 21.425 ;
        RECT 80.195 17.995 90.580 18.165 ;
        RECT 85.905 17.715 90.580 17.995 ;
        RECT 75.000 17.455 79.455 17.625 ;
        RECT 75.000 12.195 75.885 17.455 ;
        RECT 76.565 16.885 78.605 17.055 ;
        RECT 76.225 12.825 76.395 16.825 ;
        RECT 78.775 12.825 78.945 16.825 ;
        RECT 76.565 12.595 78.605 12.765 ;
        RECT 79.285 12.195 79.455 17.455 ;
        RECT 75.000 12.025 79.455 12.195 ;
        RECT 75.000 6.765 75.885 12.025 ;
        RECT 76.565 11.455 78.605 11.625 ;
        RECT 76.225 7.395 76.395 11.395 ;
        RECT 78.775 7.395 78.945 11.395 ;
        RECT 76.565 7.165 78.605 7.335 ;
        RECT 79.285 6.765 79.455 12.025 ;
        RECT 75.000 6.595 79.455 6.765 ;
        RECT 80.190 17.545 90.580 17.715 ;
        RECT 80.190 12.285 80.360 17.545 ;
        RECT 81.085 16.975 85.125 17.145 ;
        RECT 80.700 12.915 80.870 16.915 ;
        RECT 85.340 12.915 85.510 16.915 ;
        RECT 85.850 16.435 90.580 17.545 ;
        RECT 81.085 12.685 85.125 12.855 ;
        RECT 85.850 12.285 86.020 16.435 ;
        RECT 80.190 12.115 86.020 12.285 ;
        RECT 80.190 6.855 80.360 12.115 ;
        RECT 81.085 11.545 85.125 11.715 ;
        RECT 80.700 7.485 80.870 11.485 ;
        RECT 85.340 7.485 85.510 11.485 ;
        RECT 81.085 7.255 85.125 7.425 ;
        RECT 85.850 6.855 86.020 12.115 ;
        RECT 86.535 16.360 88.285 16.435 ;
        RECT 86.535 9.870 86.705 16.360 ;
        RECT 87.245 15.850 87.575 16.020 ;
        RECT 87.105 10.595 87.275 15.635 ;
        RECT 87.545 10.595 87.715 15.635 ;
        RECT 87.245 10.210 87.575 10.380 ;
        RECT 88.115 9.870 88.285 16.360 ;
        RECT 86.535 9.700 88.285 9.870 ;
        RECT 80.190 6.685 86.020 6.855 ;
        RECT 75.000 6.325 76.860 6.595 ;
        RECT 75.000 6.155 79.460 6.325 ;
        RECT 75.000 4.745 76.890 6.155 ;
        RECT 77.230 5.285 77.400 5.615 ;
        RECT 77.570 5.585 78.610 5.755 ;
        RECT 77.570 5.145 78.610 5.315 ;
        RECT 78.780 5.285 78.950 5.615 ;
        RECT 79.290 4.745 79.460 6.155 ;
        RECT 75.000 4.575 79.460 4.745 ;
        RECT 80.205 6.240 86.035 6.410 ;
        RECT 80.205 4.830 80.375 6.240 ;
        RECT 80.715 5.370 80.885 5.700 ;
        RECT 81.100 5.670 85.140 5.840 ;
        RECT 81.100 5.230 85.140 5.400 ;
        RECT 85.355 5.370 85.525 5.700 ;
        RECT 85.865 4.830 86.035 6.240 ;
        RECT 80.205 4.660 86.035 4.830 ;
        RECT 75.000 4.300 76.860 4.575 ;
        RECT 89.880 4.385 90.580 16.435 ;
        RECT 75.000 4.130 79.465 4.300 ;
        RECT 75.000 2.720 75.895 4.130 ;
        RECT 76.235 3.260 76.405 3.590 ;
        RECT 76.575 3.560 78.615 3.730 ;
        RECT 76.575 3.120 78.615 3.290 ;
        RECT 78.785 3.260 78.955 3.590 ;
        RECT 79.295 2.720 79.465 4.130 ;
        RECT 75.000 2.560 79.465 2.720 ;
        RECT 80.210 4.215 90.580 4.385 ;
        RECT 80.210 2.805 80.380 4.215 ;
        RECT 80.720 3.345 80.890 3.675 ;
        RECT 81.105 3.645 89.145 3.815 ;
        RECT 81.105 3.205 89.145 3.375 ;
        RECT 89.360 3.345 89.530 3.675 ;
        RECT 89.870 2.805 90.580 4.215 ;
        RECT 80.210 2.690 90.580 2.805 ;
        RECT 92.000 28.485 92.865 29.140 ;
        RECT 97.195 28.975 107.580 29.145 ;
        RECT 92.000 28.315 96.455 28.485 ;
        RECT 92.000 23.055 92.885 28.315 ;
        RECT 93.565 27.745 95.605 27.915 ;
        RECT 93.225 23.685 93.395 27.685 ;
        RECT 95.775 23.685 95.945 27.685 ;
        RECT 93.565 23.455 95.605 23.625 ;
        RECT 96.285 23.055 96.455 28.315 ;
        RECT 97.195 25.485 97.365 28.975 ;
        RECT 97.995 28.465 105.995 28.635 ;
        RECT 97.765 26.210 97.935 28.250 ;
        RECT 106.055 26.210 106.225 28.250 ;
        RECT 97.995 25.825 105.995 25.995 ;
        RECT 106.625 25.485 107.580 28.975 ;
        RECT 97.195 25.315 107.580 25.485 ;
        RECT 106.625 25.025 107.580 25.315 ;
        RECT 92.000 22.885 96.455 23.055 ;
        RECT 92.000 17.625 92.885 22.885 ;
        RECT 93.565 22.315 95.605 22.485 ;
        RECT 93.225 18.255 93.395 22.255 ;
        RECT 95.775 18.255 95.945 22.255 ;
        RECT 93.565 18.025 95.605 18.195 ;
        RECT 96.285 17.625 96.455 22.885 ;
        RECT 97.195 24.855 107.580 25.025 ;
        RECT 97.195 21.595 97.365 24.855 ;
        RECT 98.090 24.285 106.130 24.455 ;
        RECT 97.705 22.225 97.875 24.225 ;
        RECT 106.345 22.225 106.515 24.225 ;
        RECT 98.090 21.995 106.130 22.165 ;
        RECT 106.855 21.595 107.580 24.855 ;
        RECT 97.195 21.425 107.580 21.595 ;
        RECT 97.195 18.165 97.365 21.425 ;
        RECT 98.090 20.855 106.130 21.025 ;
        RECT 97.705 18.795 97.875 20.795 ;
        RECT 106.345 18.795 106.515 20.795 ;
        RECT 98.090 18.565 106.130 18.735 ;
        RECT 106.855 18.165 107.580 21.425 ;
        RECT 97.195 17.995 107.580 18.165 ;
        RECT 102.905 17.715 107.580 17.995 ;
        RECT 92.000 17.455 96.455 17.625 ;
        RECT 92.000 12.195 92.885 17.455 ;
        RECT 93.565 16.885 95.605 17.055 ;
        RECT 93.225 12.825 93.395 16.825 ;
        RECT 95.775 12.825 95.945 16.825 ;
        RECT 93.565 12.595 95.605 12.765 ;
        RECT 96.285 12.195 96.455 17.455 ;
        RECT 92.000 12.025 96.455 12.195 ;
        RECT 92.000 6.765 92.885 12.025 ;
        RECT 93.565 11.455 95.605 11.625 ;
        RECT 93.225 7.395 93.395 11.395 ;
        RECT 95.775 7.395 95.945 11.395 ;
        RECT 93.565 7.165 95.605 7.335 ;
        RECT 96.285 6.765 96.455 12.025 ;
        RECT 92.000 6.595 96.455 6.765 ;
        RECT 97.190 17.545 107.580 17.715 ;
        RECT 97.190 12.285 97.360 17.545 ;
        RECT 98.085 16.975 102.125 17.145 ;
        RECT 97.700 12.915 97.870 16.915 ;
        RECT 102.340 12.915 102.510 16.915 ;
        RECT 102.850 16.435 107.580 17.545 ;
        RECT 98.085 12.685 102.125 12.855 ;
        RECT 102.850 12.285 103.020 16.435 ;
        RECT 97.190 12.115 103.020 12.285 ;
        RECT 97.190 6.855 97.360 12.115 ;
        RECT 98.085 11.545 102.125 11.715 ;
        RECT 97.700 7.485 97.870 11.485 ;
        RECT 102.340 7.485 102.510 11.485 ;
        RECT 98.085 7.255 102.125 7.425 ;
        RECT 102.850 6.855 103.020 12.115 ;
        RECT 103.535 16.360 105.285 16.435 ;
        RECT 103.535 9.870 103.705 16.360 ;
        RECT 104.245 15.850 104.575 16.020 ;
        RECT 104.105 10.595 104.275 15.635 ;
        RECT 104.545 10.595 104.715 15.635 ;
        RECT 104.245 10.210 104.575 10.380 ;
        RECT 105.115 9.870 105.285 16.360 ;
        RECT 103.535 9.700 105.285 9.870 ;
        RECT 97.190 6.685 103.020 6.855 ;
        RECT 92.000 6.325 93.860 6.595 ;
        RECT 92.000 6.155 96.460 6.325 ;
        RECT 92.000 4.745 93.890 6.155 ;
        RECT 94.230 5.285 94.400 5.615 ;
        RECT 94.570 5.585 95.610 5.755 ;
        RECT 94.570 5.145 95.610 5.315 ;
        RECT 95.780 5.285 95.950 5.615 ;
        RECT 96.290 4.745 96.460 6.155 ;
        RECT 92.000 4.575 96.460 4.745 ;
        RECT 97.205 6.240 103.035 6.410 ;
        RECT 97.205 4.830 97.375 6.240 ;
        RECT 97.715 5.370 97.885 5.700 ;
        RECT 98.100 5.670 102.140 5.840 ;
        RECT 98.100 5.230 102.140 5.400 ;
        RECT 102.355 5.370 102.525 5.700 ;
        RECT 102.865 4.830 103.035 6.240 ;
        RECT 97.205 4.660 103.035 4.830 ;
        RECT 92.000 4.300 93.860 4.575 ;
        RECT 106.880 4.385 107.580 16.435 ;
        RECT 92.000 4.130 96.465 4.300 ;
        RECT 92.000 2.720 92.895 4.130 ;
        RECT 93.235 3.260 93.405 3.590 ;
        RECT 93.575 3.560 95.615 3.730 ;
        RECT 93.575 3.120 95.615 3.290 ;
        RECT 95.785 3.260 95.955 3.590 ;
        RECT 96.295 2.720 96.465 4.130 ;
        RECT 80.210 2.635 90.040 2.690 ;
        RECT 92.000 2.560 96.465 2.720 ;
        RECT 97.210 4.215 107.580 4.385 ;
        RECT 97.210 2.805 97.380 4.215 ;
        RECT 97.720 3.345 97.890 3.675 ;
        RECT 98.105 3.645 106.145 3.815 ;
        RECT 98.105 3.205 106.145 3.375 ;
        RECT 106.360 3.345 106.530 3.675 ;
        RECT 106.870 2.805 107.580 4.215 ;
        RECT 97.210 2.690 107.580 2.805 ;
        RECT 109.000 28.485 109.865 29.140 ;
        RECT 114.195 28.975 124.580 29.145 ;
        RECT 109.000 28.315 113.455 28.485 ;
        RECT 109.000 23.055 109.885 28.315 ;
        RECT 110.565 27.745 112.605 27.915 ;
        RECT 110.225 23.685 110.395 27.685 ;
        RECT 112.775 23.685 112.945 27.685 ;
        RECT 110.565 23.455 112.605 23.625 ;
        RECT 113.285 23.055 113.455 28.315 ;
        RECT 114.195 25.485 114.365 28.975 ;
        RECT 114.995 28.465 122.995 28.635 ;
        RECT 114.765 26.210 114.935 28.250 ;
        RECT 123.055 26.210 123.225 28.250 ;
        RECT 114.995 25.825 122.995 25.995 ;
        RECT 123.625 25.485 124.580 28.975 ;
        RECT 114.195 25.315 124.580 25.485 ;
        RECT 123.625 25.025 124.580 25.315 ;
        RECT 109.000 22.885 113.455 23.055 ;
        RECT 109.000 17.625 109.885 22.885 ;
        RECT 110.565 22.315 112.605 22.485 ;
        RECT 110.225 18.255 110.395 22.255 ;
        RECT 112.775 18.255 112.945 22.255 ;
        RECT 110.565 18.025 112.605 18.195 ;
        RECT 113.285 17.625 113.455 22.885 ;
        RECT 114.195 24.855 124.580 25.025 ;
        RECT 114.195 21.595 114.365 24.855 ;
        RECT 115.090 24.285 123.130 24.455 ;
        RECT 114.705 22.225 114.875 24.225 ;
        RECT 123.345 22.225 123.515 24.225 ;
        RECT 115.090 21.995 123.130 22.165 ;
        RECT 123.855 21.595 124.580 24.855 ;
        RECT 114.195 21.425 124.580 21.595 ;
        RECT 114.195 18.165 114.365 21.425 ;
        RECT 115.090 20.855 123.130 21.025 ;
        RECT 114.705 18.795 114.875 20.795 ;
        RECT 123.345 18.795 123.515 20.795 ;
        RECT 115.090 18.565 123.130 18.735 ;
        RECT 123.855 18.165 124.580 21.425 ;
        RECT 114.195 17.995 124.580 18.165 ;
        RECT 119.905 17.715 124.580 17.995 ;
        RECT 109.000 17.455 113.455 17.625 ;
        RECT 109.000 12.195 109.885 17.455 ;
        RECT 110.565 16.885 112.605 17.055 ;
        RECT 110.225 12.825 110.395 16.825 ;
        RECT 112.775 12.825 112.945 16.825 ;
        RECT 110.565 12.595 112.605 12.765 ;
        RECT 113.285 12.195 113.455 17.455 ;
        RECT 109.000 12.025 113.455 12.195 ;
        RECT 109.000 6.765 109.885 12.025 ;
        RECT 110.565 11.455 112.605 11.625 ;
        RECT 110.225 7.395 110.395 11.395 ;
        RECT 112.775 7.395 112.945 11.395 ;
        RECT 110.565 7.165 112.605 7.335 ;
        RECT 113.285 6.765 113.455 12.025 ;
        RECT 109.000 6.595 113.455 6.765 ;
        RECT 114.190 17.545 124.580 17.715 ;
        RECT 114.190 12.285 114.360 17.545 ;
        RECT 115.085 16.975 119.125 17.145 ;
        RECT 114.700 12.915 114.870 16.915 ;
        RECT 119.340 12.915 119.510 16.915 ;
        RECT 119.850 16.435 124.580 17.545 ;
        RECT 115.085 12.685 119.125 12.855 ;
        RECT 119.850 12.285 120.020 16.435 ;
        RECT 114.190 12.115 120.020 12.285 ;
        RECT 114.190 6.855 114.360 12.115 ;
        RECT 115.085 11.545 119.125 11.715 ;
        RECT 114.700 7.485 114.870 11.485 ;
        RECT 119.340 7.485 119.510 11.485 ;
        RECT 115.085 7.255 119.125 7.425 ;
        RECT 119.850 6.855 120.020 12.115 ;
        RECT 120.535 16.360 122.285 16.435 ;
        RECT 120.535 9.870 120.705 16.360 ;
        RECT 121.245 15.850 121.575 16.020 ;
        RECT 121.105 10.595 121.275 15.635 ;
        RECT 121.545 10.595 121.715 15.635 ;
        RECT 121.245 10.210 121.575 10.380 ;
        RECT 122.115 9.870 122.285 16.360 ;
        RECT 120.535 9.700 122.285 9.870 ;
        RECT 114.190 6.685 120.020 6.855 ;
        RECT 109.000 6.325 110.860 6.595 ;
        RECT 109.000 6.155 113.460 6.325 ;
        RECT 109.000 4.745 110.890 6.155 ;
        RECT 111.230 5.285 111.400 5.615 ;
        RECT 111.570 5.585 112.610 5.755 ;
        RECT 111.570 5.145 112.610 5.315 ;
        RECT 112.780 5.285 112.950 5.615 ;
        RECT 113.290 4.745 113.460 6.155 ;
        RECT 109.000 4.575 113.460 4.745 ;
        RECT 114.205 6.240 120.035 6.410 ;
        RECT 114.205 4.830 114.375 6.240 ;
        RECT 114.715 5.370 114.885 5.700 ;
        RECT 115.100 5.670 119.140 5.840 ;
        RECT 115.100 5.230 119.140 5.400 ;
        RECT 119.355 5.370 119.525 5.700 ;
        RECT 119.865 4.830 120.035 6.240 ;
        RECT 114.205 4.660 120.035 4.830 ;
        RECT 109.000 4.300 110.860 4.575 ;
        RECT 123.880 4.385 124.580 16.435 ;
        RECT 109.000 4.130 113.465 4.300 ;
        RECT 109.000 2.720 109.895 4.130 ;
        RECT 110.235 3.260 110.405 3.590 ;
        RECT 110.575 3.560 112.615 3.730 ;
        RECT 110.575 3.120 112.615 3.290 ;
        RECT 112.785 3.260 112.955 3.590 ;
        RECT 113.295 2.720 113.465 4.130 ;
        RECT 97.210 2.635 107.040 2.690 ;
        RECT 109.000 2.560 113.465 2.720 ;
        RECT 114.210 4.215 124.580 4.385 ;
        RECT 114.210 2.805 114.380 4.215 ;
        RECT 114.720 3.345 114.890 3.675 ;
        RECT 115.105 3.645 123.145 3.815 ;
        RECT 115.105 3.205 123.145 3.375 ;
        RECT 123.360 3.345 123.530 3.675 ;
        RECT 123.870 2.805 124.580 4.215 ;
        RECT 114.210 2.690 124.580 2.805 ;
        RECT 126.000 28.485 126.865 29.140 ;
        RECT 131.195 28.975 141.580 29.145 ;
        RECT 126.000 28.315 130.455 28.485 ;
        RECT 126.000 23.055 126.885 28.315 ;
        RECT 127.565 27.745 129.605 27.915 ;
        RECT 127.225 23.685 127.395 27.685 ;
        RECT 129.775 23.685 129.945 27.685 ;
        RECT 127.565 23.455 129.605 23.625 ;
        RECT 130.285 23.055 130.455 28.315 ;
        RECT 131.195 25.485 131.365 28.975 ;
        RECT 131.995 28.465 139.995 28.635 ;
        RECT 131.765 26.210 131.935 28.250 ;
        RECT 140.055 26.210 140.225 28.250 ;
        RECT 131.995 25.825 139.995 25.995 ;
        RECT 140.625 25.485 141.580 28.975 ;
        RECT 131.195 25.315 141.580 25.485 ;
        RECT 140.625 25.025 141.580 25.315 ;
        RECT 126.000 22.885 130.455 23.055 ;
        RECT 126.000 17.625 126.885 22.885 ;
        RECT 127.565 22.315 129.605 22.485 ;
        RECT 127.225 18.255 127.395 22.255 ;
        RECT 129.775 18.255 129.945 22.255 ;
        RECT 127.565 18.025 129.605 18.195 ;
        RECT 130.285 17.625 130.455 22.885 ;
        RECT 131.195 24.855 141.580 25.025 ;
        RECT 131.195 21.595 131.365 24.855 ;
        RECT 132.090 24.285 140.130 24.455 ;
        RECT 131.705 22.225 131.875 24.225 ;
        RECT 140.345 22.225 140.515 24.225 ;
        RECT 132.090 21.995 140.130 22.165 ;
        RECT 140.855 21.595 141.580 24.855 ;
        RECT 131.195 21.425 141.580 21.595 ;
        RECT 131.195 18.165 131.365 21.425 ;
        RECT 132.090 20.855 140.130 21.025 ;
        RECT 131.705 18.795 131.875 20.795 ;
        RECT 140.345 18.795 140.515 20.795 ;
        RECT 132.090 18.565 140.130 18.735 ;
        RECT 140.855 18.165 141.580 21.425 ;
        RECT 131.195 17.995 141.580 18.165 ;
        RECT 136.905 17.715 141.580 17.995 ;
        RECT 126.000 17.455 130.455 17.625 ;
        RECT 126.000 12.195 126.885 17.455 ;
        RECT 127.565 16.885 129.605 17.055 ;
        RECT 127.225 12.825 127.395 16.825 ;
        RECT 129.775 12.825 129.945 16.825 ;
        RECT 127.565 12.595 129.605 12.765 ;
        RECT 130.285 12.195 130.455 17.455 ;
        RECT 126.000 12.025 130.455 12.195 ;
        RECT 126.000 6.765 126.885 12.025 ;
        RECT 127.565 11.455 129.605 11.625 ;
        RECT 127.225 7.395 127.395 11.395 ;
        RECT 129.775 7.395 129.945 11.395 ;
        RECT 127.565 7.165 129.605 7.335 ;
        RECT 130.285 6.765 130.455 12.025 ;
        RECT 126.000 6.595 130.455 6.765 ;
        RECT 131.190 17.545 141.580 17.715 ;
        RECT 131.190 12.285 131.360 17.545 ;
        RECT 132.085 16.975 136.125 17.145 ;
        RECT 131.700 12.915 131.870 16.915 ;
        RECT 136.340 12.915 136.510 16.915 ;
        RECT 136.850 16.435 141.580 17.545 ;
        RECT 132.085 12.685 136.125 12.855 ;
        RECT 136.850 12.285 137.020 16.435 ;
        RECT 131.190 12.115 137.020 12.285 ;
        RECT 131.190 6.855 131.360 12.115 ;
        RECT 132.085 11.545 136.125 11.715 ;
        RECT 131.700 7.485 131.870 11.485 ;
        RECT 136.340 7.485 136.510 11.485 ;
        RECT 132.085 7.255 136.125 7.425 ;
        RECT 136.850 6.855 137.020 12.115 ;
        RECT 137.535 16.360 139.285 16.435 ;
        RECT 137.535 9.870 137.705 16.360 ;
        RECT 138.245 15.850 138.575 16.020 ;
        RECT 138.105 10.595 138.275 15.635 ;
        RECT 138.545 10.595 138.715 15.635 ;
        RECT 138.245 10.210 138.575 10.380 ;
        RECT 139.115 9.870 139.285 16.360 ;
        RECT 137.535 9.700 139.285 9.870 ;
        RECT 131.190 6.685 137.020 6.855 ;
        RECT 126.000 6.325 127.860 6.595 ;
        RECT 126.000 6.155 130.460 6.325 ;
        RECT 126.000 4.745 127.890 6.155 ;
        RECT 128.230 5.285 128.400 5.615 ;
        RECT 128.570 5.585 129.610 5.755 ;
        RECT 128.570 5.145 129.610 5.315 ;
        RECT 129.780 5.285 129.950 5.615 ;
        RECT 130.290 4.745 130.460 6.155 ;
        RECT 126.000 4.575 130.460 4.745 ;
        RECT 131.205 6.240 137.035 6.410 ;
        RECT 131.205 4.830 131.375 6.240 ;
        RECT 131.715 5.370 131.885 5.700 ;
        RECT 132.100 5.670 136.140 5.840 ;
        RECT 132.100 5.230 136.140 5.400 ;
        RECT 136.355 5.370 136.525 5.700 ;
        RECT 136.865 4.830 137.035 6.240 ;
        RECT 131.205 4.660 137.035 4.830 ;
        RECT 126.000 4.300 127.860 4.575 ;
        RECT 140.880 4.385 141.580 16.435 ;
        RECT 126.000 4.130 130.465 4.300 ;
        RECT 126.000 2.720 126.895 4.130 ;
        RECT 127.235 3.260 127.405 3.590 ;
        RECT 127.575 3.560 129.615 3.730 ;
        RECT 127.575 3.120 129.615 3.290 ;
        RECT 129.785 3.260 129.955 3.590 ;
        RECT 130.295 2.720 130.465 4.130 ;
        RECT 114.210 2.635 124.040 2.690 ;
        RECT 126.000 2.560 130.465 2.720 ;
        RECT 131.210 4.215 141.580 4.385 ;
        RECT 131.210 2.805 131.380 4.215 ;
        RECT 131.720 3.345 131.890 3.675 ;
        RECT 132.105 3.645 140.145 3.815 ;
        RECT 132.105 3.205 140.145 3.375 ;
        RECT 140.360 3.345 140.530 3.675 ;
        RECT 140.870 2.805 141.580 4.215 ;
        RECT 131.210 2.690 141.580 2.805 ;
        RECT 143.000 28.485 143.865 29.140 ;
        RECT 148.195 28.975 158.580 29.145 ;
        RECT 143.000 28.315 147.455 28.485 ;
        RECT 143.000 23.055 143.885 28.315 ;
        RECT 144.565 27.745 146.605 27.915 ;
        RECT 144.225 23.685 144.395 27.685 ;
        RECT 146.775 23.685 146.945 27.685 ;
        RECT 144.565 23.455 146.605 23.625 ;
        RECT 147.285 23.055 147.455 28.315 ;
        RECT 148.195 25.485 148.365 28.975 ;
        RECT 148.995 28.465 156.995 28.635 ;
        RECT 148.765 26.210 148.935 28.250 ;
        RECT 157.055 26.210 157.225 28.250 ;
        RECT 148.995 25.825 156.995 25.995 ;
        RECT 157.625 25.485 158.580 28.975 ;
        RECT 148.195 25.315 158.580 25.485 ;
        RECT 157.625 25.025 158.580 25.315 ;
        RECT 143.000 22.885 147.455 23.055 ;
        RECT 143.000 17.625 143.885 22.885 ;
        RECT 144.565 22.315 146.605 22.485 ;
        RECT 144.225 18.255 144.395 22.255 ;
        RECT 146.775 18.255 146.945 22.255 ;
        RECT 144.565 18.025 146.605 18.195 ;
        RECT 147.285 17.625 147.455 22.885 ;
        RECT 148.195 24.855 158.580 25.025 ;
        RECT 148.195 21.595 148.365 24.855 ;
        RECT 149.090 24.285 157.130 24.455 ;
        RECT 148.705 22.225 148.875 24.225 ;
        RECT 157.345 22.225 157.515 24.225 ;
        RECT 149.090 21.995 157.130 22.165 ;
        RECT 157.855 21.595 158.580 24.855 ;
        RECT 148.195 21.425 158.580 21.595 ;
        RECT 148.195 18.165 148.365 21.425 ;
        RECT 149.090 20.855 157.130 21.025 ;
        RECT 148.705 18.795 148.875 20.795 ;
        RECT 157.345 18.795 157.515 20.795 ;
        RECT 149.090 18.565 157.130 18.735 ;
        RECT 157.855 18.165 158.580 21.425 ;
        RECT 148.195 17.995 158.580 18.165 ;
        RECT 153.905 17.715 158.580 17.995 ;
        RECT 143.000 17.455 147.455 17.625 ;
        RECT 143.000 12.195 143.885 17.455 ;
        RECT 144.565 16.885 146.605 17.055 ;
        RECT 144.225 12.825 144.395 16.825 ;
        RECT 146.775 12.825 146.945 16.825 ;
        RECT 144.565 12.595 146.605 12.765 ;
        RECT 147.285 12.195 147.455 17.455 ;
        RECT 143.000 12.025 147.455 12.195 ;
        RECT 143.000 6.765 143.885 12.025 ;
        RECT 144.565 11.455 146.605 11.625 ;
        RECT 144.225 7.395 144.395 11.395 ;
        RECT 146.775 7.395 146.945 11.395 ;
        RECT 144.565 7.165 146.605 7.335 ;
        RECT 147.285 6.765 147.455 12.025 ;
        RECT 143.000 6.595 147.455 6.765 ;
        RECT 148.190 17.545 158.580 17.715 ;
        RECT 148.190 12.285 148.360 17.545 ;
        RECT 149.085 16.975 153.125 17.145 ;
        RECT 148.700 12.915 148.870 16.915 ;
        RECT 153.340 12.915 153.510 16.915 ;
        RECT 153.850 16.435 158.580 17.545 ;
        RECT 149.085 12.685 153.125 12.855 ;
        RECT 153.850 12.285 154.020 16.435 ;
        RECT 148.190 12.115 154.020 12.285 ;
        RECT 148.190 6.855 148.360 12.115 ;
        RECT 149.085 11.545 153.125 11.715 ;
        RECT 148.700 7.485 148.870 11.485 ;
        RECT 153.340 7.485 153.510 11.485 ;
        RECT 149.085 7.255 153.125 7.425 ;
        RECT 153.850 6.855 154.020 12.115 ;
        RECT 154.535 16.360 156.285 16.435 ;
        RECT 154.535 9.870 154.705 16.360 ;
        RECT 155.245 15.850 155.575 16.020 ;
        RECT 155.105 10.595 155.275 15.635 ;
        RECT 155.545 10.595 155.715 15.635 ;
        RECT 155.245 10.210 155.575 10.380 ;
        RECT 156.115 9.870 156.285 16.360 ;
        RECT 154.535 9.700 156.285 9.870 ;
        RECT 148.190 6.685 154.020 6.855 ;
        RECT 143.000 6.325 144.860 6.595 ;
        RECT 143.000 6.155 147.460 6.325 ;
        RECT 143.000 4.745 144.890 6.155 ;
        RECT 145.230 5.285 145.400 5.615 ;
        RECT 145.570 5.585 146.610 5.755 ;
        RECT 145.570 5.145 146.610 5.315 ;
        RECT 146.780 5.285 146.950 5.615 ;
        RECT 147.290 4.745 147.460 6.155 ;
        RECT 143.000 4.575 147.460 4.745 ;
        RECT 148.205 6.240 154.035 6.410 ;
        RECT 148.205 4.830 148.375 6.240 ;
        RECT 148.715 5.370 148.885 5.700 ;
        RECT 149.100 5.670 153.140 5.840 ;
        RECT 149.100 5.230 153.140 5.400 ;
        RECT 153.355 5.370 153.525 5.700 ;
        RECT 153.865 4.830 154.035 6.240 ;
        RECT 148.205 4.660 154.035 4.830 ;
        RECT 143.000 4.300 144.860 4.575 ;
        RECT 157.880 4.385 158.580 16.435 ;
        RECT 143.000 4.130 147.465 4.300 ;
        RECT 143.000 2.720 143.895 4.130 ;
        RECT 144.235 3.260 144.405 3.590 ;
        RECT 144.575 3.560 146.615 3.730 ;
        RECT 144.575 3.120 146.615 3.290 ;
        RECT 146.785 3.260 146.955 3.590 ;
        RECT 147.295 2.720 147.465 4.130 ;
        RECT 131.210 2.635 141.040 2.690 ;
        RECT 143.000 2.560 147.465 2.720 ;
        RECT 148.210 4.215 158.580 4.385 ;
        RECT 148.210 2.805 148.380 4.215 ;
        RECT 148.720 3.345 148.890 3.675 ;
        RECT 149.105 3.645 157.145 3.815 ;
        RECT 149.105 3.205 157.145 3.375 ;
        RECT 157.360 3.345 157.530 3.675 ;
        RECT 157.870 2.805 158.580 4.215 ;
        RECT 148.210 2.690 158.580 2.805 ;
        RECT 148.210 2.635 158.040 2.690 ;
        RECT 75.725 2.550 79.465 2.560 ;
        RECT 92.725 2.550 96.465 2.560 ;
        RECT 109.725 2.550 113.465 2.560 ;
        RECT 126.725 2.550 130.465 2.560 ;
        RECT 143.725 2.550 147.465 2.560 ;
      LAYER met1 ;
        RECT 74.630 130.980 87.440 131.000 ;
        RECT 74.610 130.170 87.450 130.980 ;
        RECT 74.630 130.110 87.440 130.170 ;
        RECT 75.630 129.750 76.070 130.110 ;
        RECT 77.210 130.000 78.370 130.110 ;
        RECT 77.210 129.750 77.650 130.000 ;
        RECT 78.800 129.750 79.240 130.110 ;
        RECT 80.390 129.750 80.830 130.110 ;
        RECT 74.770 129.700 75.000 129.730 ;
        RECT 75.160 129.700 75.390 129.750 ;
        RECT 74.770 123.810 75.390 129.700 ;
        RECT 74.770 123.530 75.010 123.810 ;
        RECT 75.160 123.750 75.390 123.810 ;
        RECT 75.600 123.810 76.070 129.750 ;
        RECT 76.740 129.680 76.970 129.750 ;
        RECT 76.440 123.830 76.970 129.680 ;
        RECT 76.440 123.810 76.600 123.830 ;
        RECT 75.600 123.750 75.830 123.810 ;
        RECT 76.450 123.570 76.600 123.810 ;
        RECT 76.740 123.750 76.970 123.830 ;
        RECT 77.180 123.830 77.650 129.750 ;
        RECT 78.320 129.680 78.550 129.750 ;
        RECT 77.950 125.090 78.560 129.680 ;
        RECT 77.180 123.750 77.410 123.830 ;
        RECT 77.930 123.800 78.560 125.090 ;
        RECT 78.760 123.840 79.240 129.750 ;
        RECT 79.900 129.700 80.130 129.750 ;
        RECT 74.770 121.100 75.150 123.530 ;
        RECT 75.350 123.520 75.640 123.545 ;
        RECT 75.340 122.790 75.660 123.520 ;
        RECT 75.290 121.790 76.290 122.790 ;
        RECT 75.340 121.100 75.660 121.790 ;
        RECT 74.770 120.790 75.010 121.100 ;
        RECT 75.360 121.060 75.660 121.100 ;
        RECT 75.360 121.050 75.650 121.060 ;
        RECT 76.450 121.040 76.650 123.570 ;
        RECT 76.930 123.540 77.220 123.545 ;
        RECT 76.920 122.840 77.260 123.540 ;
        RECT 76.790 121.840 77.790 122.840 ;
        RECT 76.920 121.070 77.260 121.840 ;
        RECT 76.940 121.050 77.230 121.070 ;
        RECT 75.170 120.790 75.400 120.890 ;
        RECT 74.770 120.780 75.400 120.790 ;
        RECT 74.740 118.980 75.400 120.780 ;
        RECT 74.770 118.960 75.000 118.980 ;
        RECT 75.170 118.890 75.400 118.980 ;
        RECT 75.610 120.820 75.840 120.890 ;
        RECT 75.610 119.010 76.170 120.820 ;
        RECT 76.450 120.780 76.600 121.040 ;
        RECT 76.750 120.780 76.980 120.890 ;
        RECT 76.450 120.770 76.980 120.780 ;
        RECT 75.610 118.890 75.840 119.010 ;
        RECT 76.000 118.690 76.170 119.010 ;
        RECT 76.410 118.970 76.980 120.770 ;
        RECT 76.460 118.960 76.980 118.970 ;
        RECT 76.750 118.890 76.980 118.960 ;
        RECT 77.190 120.840 77.420 120.890 ;
        RECT 77.190 120.810 77.700 120.840 ;
        RECT 77.190 119.000 77.730 120.810 ;
        RECT 77.930 120.790 78.120 123.800 ;
        RECT 78.320 123.750 78.550 123.800 ;
        RECT 78.760 123.750 78.990 123.840 ;
        RECT 79.510 123.800 80.130 129.700 ;
        RECT 78.480 122.840 78.840 123.550 ;
        RECT 78.300 121.840 79.300 122.840 ;
        RECT 78.480 121.050 78.840 121.840 ;
        RECT 78.330 120.790 78.560 120.890 ;
        RECT 77.930 120.120 78.560 120.790 ;
        RECT 77.190 118.890 77.420 119.000 ;
        RECT 77.560 118.770 77.730 119.000 ;
        RECT 77.950 118.920 78.560 120.120 ;
        RECT 78.330 118.890 78.560 118.920 ;
        RECT 78.770 120.840 79.000 120.890 ;
        RECT 78.770 118.960 79.310 120.840 ;
        RECT 79.530 120.820 79.700 123.800 ;
        RECT 79.900 123.750 80.130 123.800 ;
        RECT 80.340 123.830 80.830 129.750 ;
        RECT 81.480 129.670 81.710 129.750 ;
        RECT 80.340 123.750 80.570 123.830 ;
        RECT 81.070 123.790 81.710 129.670 ;
        RECT 80.090 123.540 80.380 123.545 ;
        RECT 80.080 122.870 80.420 123.540 ;
        RECT 79.910 121.870 80.910 122.870 ;
        RECT 80.080 121.060 80.420 121.870 ;
        RECT 80.100 121.050 80.390 121.060 ;
        RECT 79.910 120.820 80.140 120.890 ;
        RECT 79.530 120.780 80.140 120.820 ;
        RECT 79.510 118.980 80.140 120.780 ;
        RECT 79.540 118.960 80.140 118.980 ;
        RECT 78.770 118.890 79.000 118.960 ;
        RECT 74.640 118.550 75.640 118.560 ;
        RECT 75.920 118.550 76.170 118.690 ;
        RECT 77.550 118.550 77.730 118.770 ;
        RECT 79.140 118.720 79.310 118.960 ;
        RECT 79.910 118.890 80.140 118.960 ;
        RECT 80.350 120.820 80.580 120.890 ;
        RECT 80.350 118.940 80.890 120.820 ;
        RECT 81.080 120.810 81.270 123.790 ;
        RECT 81.480 123.750 81.710 123.790 ;
        RECT 81.910 123.780 82.350 130.110 ;
        RECT 83.530 129.750 83.970 130.110 ;
        RECT 85.120 129.750 85.560 130.110 ;
        RECT 86.700 129.750 87.140 130.110 ;
        RECT 83.060 129.730 83.290 129.750 ;
        RECT 82.610 123.800 83.290 129.730 ;
        RECT 81.920 123.750 82.150 123.780 ;
        RECT 81.670 123.540 81.960 123.545 ;
        RECT 81.650 122.840 82.010 123.540 ;
        RECT 81.460 121.840 82.460 122.840 ;
        RECT 81.650 121.050 82.010 121.840 ;
        RECT 81.490 120.810 81.720 120.890 ;
        RECT 81.080 118.960 81.720 120.810 ;
        RECT 80.350 118.890 80.580 118.940 ;
        RECT 79.130 118.550 79.310 118.720 ;
        RECT 80.720 118.550 80.890 118.940 ;
        RECT 81.490 118.890 81.720 118.960 ;
        RECT 81.930 120.840 82.160 120.890 ;
        RECT 82.620 120.850 82.880 123.800 ;
        RECT 83.060 123.750 83.290 123.800 ;
        RECT 83.500 123.810 83.970 129.750 ;
        RECT 84.640 129.710 84.870 129.750 ;
        RECT 83.500 123.750 83.730 123.810 ;
        RECT 84.190 123.800 84.870 129.710 ;
        RECT 83.250 123.540 83.540 123.545 ;
        RECT 83.220 122.870 83.560 123.540 ;
        RECT 83.080 121.870 84.080 122.870 ;
        RECT 83.220 121.050 83.560 121.870 ;
        RECT 83.070 120.850 83.300 120.890 ;
        RECT 81.930 118.960 82.470 120.840 ;
        RECT 81.930 118.890 82.160 118.960 ;
        RECT 82.300 118.550 82.470 118.960 ;
        RECT 82.620 118.930 83.300 120.850 ;
        RECT 83.070 118.890 83.300 118.930 ;
        RECT 83.510 120.830 83.740 120.890 ;
        RECT 83.510 118.950 84.060 120.830 ;
        RECT 84.240 120.810 84.500 123.800 ;
        RECT 84.640 123.750 84.870 123.800 ;
        RECT 85.080 123.790 85.560 129.750 ;
        RECT 86.220 129.710 86.450 129.750 ;
        RECT 85.790 123.820 86.450 129.710 ;
        RECT 85.790 123.800 86.050 123.820 ;
        RECT 85.080 123.750 85.310 123.790 ;
        RECT 85.800 123.590 86.050 123.800 ;
        RECT 86.220 123.750 86.450 123.820 ;
        RECT 86.660 123.840 87.140 129.750 ;
        RECT 142.375 126.805 146.455 127.305 ;
        RECT 86.660 123.750 86.890 123.840 ;
        RECT 84.830 123.540 85.120 123.545 ;
        RECT 84.820 122.840 85.150 123.540 ;
        RECT 84.650 121.840 85.650 122.840 ;
        RECT 84.820 121.050 85.150 121.840 ;
        RECT 85.800 121.490 86.100 123.590 ;
        RECT 86.410 123.540 86.700 123.545 ;
        RECT 86.390 122.860 86.750 123.540 ;
        RECT 86.310 121.860 87.310 122.860 ;
        RECT 85.880 121.040 86.100 121.490 ;
        RECT 86.390 121.050 86.750 121.860 ;
        RECT 84.650 120.810 84.880 120.890 ;
        RECT 84.220 118.960 84.880 120.810 ;
        RECT 83.510 118.890 83.740 118.950 ;
        RECT 83.900 118.550 84.060 118.950 ;
        RECT 84.650 118.890 84.880 118.960 ;
        RECT 85.090 120.830 85.320 120.890 ;
        RECT 85.090 118.940 85.640 120.830 ;
        RECT 85.880 120.800 86.060 121.040 ;
        RECT 86.230 120.800 86.460 120.890 ;
        RECT 85.880 120.650 86.460 120.800 ;
        RECT 85.850 118.980 86.460 120.650 ;
        RECT 85.860 118.950 86.460 118.980 ;
        RECT 85.090 118.890 85.320 118.940 ;
        RECT 85.470 118.550 85.640 118.940 ;
        RECT 86.230 118.890 86.460 118.950 ;
        RECT 86.670 120.830 86.900 120.890 ;
        RECT 86.670 118.980 87.360 120.830 ;
        RECT 86.670 118.890 86.900 118.980 ;
        RECT 87.050 118.730 87.360 118.980 ;
        RECT 87.030 118.690 87.360 118.730 ;
        RECT 87.030 118.550 87.520 118.690 ;
        RECT 74.640 118.520 87.520 118.550 ;
        RECT 74.620 117.530 87.520 118.520 ;
        RECT 142.375 118.010 142.875 126.805 ;
        RECT 145.850 118.830 146.850 119.150 ;
        RECT 147.350 118.880 148.350 119.200 ;
        RECT 148.860 118.880 149.860 119.200 ;
        RECT 150.470 118.910 151.470 119.230 ;
        RECT 152.020 118.880 153.020 119.200 ;
        RECT 153.640 118.910 154.640 119.230 ;
        RECT 155.210 118.880 156.210 119.200 ;
        RECT 156.870 118.900 157.870 119.220 ;
        RECT 74.640 117.490 87.520 117.530 ;
        RECT 75.180 114.810 75.790 117.150 ;
        RECT 76.620 116.960 77.280 117.280 ;
        RECT 76.670 114.840 77.280 116.960 ;
        RECT 77.120 114.810 77.280 114.840 ;
        RECT 78.140 114.800 78.690 117.150 ;
        RECT 79.650 114.780 80.200 117.130 ;
        RECT 81.110 114.810 81.660 117.160 ;
        RECT 82.590 114.840 83.140 117.190 ;
        RECT 84.040 114.830 84.590 117.180 ;
        RECT 85.540 114.840 86.090 117.190 ;
        RECT 86.960 117.050 87.520 117.490 ;
        RECT 121.890 117.510 142.875 118.010 ;
        RECT 86.960 114.890 87.530 117.050 ;
        RECT 121.890 117.010 122.390 117.510 ;
        RECT 121.335 116.975 123.200 117.010 ;
        RECT 121.210 116.915 123.200 116.975 ;
        RECT 121.210 116.435 123.250 116.915 ;
        RECT 127.870 116.905 128.315 116.920 ;
        RECT 124.830 116.845 128.315 116.905 ;
        RECT 121.215 116.360 123.250 116.435 ;
        RECT 124.695 116.490 128.315 116.845 ;
        RECT 86.960 114.880 87.520 114.890 ;
        RECT 74.620 113.630 75.010 113.640 ;
        RECT 74.620 111.470 75.640 113.630 ;
        RECT 74.620 107.650 75.010 111.470 ;
        RECT 76.100 111.230 77.100 113.630 ;
        RECT 77.590 111.500 78.590 113.650 ;
        RECT 75.850 111.000 77.100 111.230 ;
        RECT 75.290 110.840 77.100 111.000 ;
        RECT 77.360 110.860 78.590 111.500 ;
        RECT 79.070 111.490 80.070 113.640 ;
        RECT 80.530 111.490 81.530 113.630 ;
        RECT 75.290 110.540 76.570 110.840 ;
        RECT 75.290 108.660 76.290 110.540 ;
        RECT 77.360 110.390 78.040 110.860 ;
        RECT 78.850 110.850 80.070 111.490 ;
        RECT 78.850 110.390 79.530 110.850 ;
        RECT 80.340 110.840 81.530 111.490 ;
        RECT 82.030 111.460 83.030 113.650 ;
        RECT 84.970 113.630 87.280 113.640 ;
        RECT 81.790 110.860 83.030 111.460 ;
        RECT 83.540 111.450 84.540 113.630 ;
        RECT 84.970 111.460 87.450 113.630 ;
        RECT 121.215 113.355 123.385 116.360 ;
        RECT 123.955 115.890 124.300 116.150 ;
        RECT 123.975 115.860 124.265 115.890 ;
        RECT 123.785 115.625 124.015 115.655 ;
        RECT 80.340 110.390 81.020 110.840 ;
        RECT 81.790 110.390 82.470 110.860 ;
        RECT 76.740 109.920 78.040 110.390 ;
        RECT 76.740 108.750 77.780 109.920 ;
        RECT 78.250 109.910 79.530 110.390 ;
        RECT 79.720 109.910 81.020 110.390 ;
        RECT 78.250 108.750 79.290 109.910 ;
        RECT 79.720 108.750 80.760 109.910 ;
        RECT 81.210 109.880 82.470 110.390 ;
        RECT 83.290 110.840 84.540 111.450 ;
        RECT 84.800 110.850 87.450 111.460 ;
        RECT 83.290 110.380 83.970 110.840 ;
        RECT 84.800 110.390 85.480 110.850 ;
        RECT 86.450 110.840 87.450 110.850 ;
        RECT 118.590 112.160 123.385 113.355 ;
        RECT 75.290 108.210 76.520 108.660 ;
        RECT 76.740 108.210 78.070 108.750 ;
        RECT 78.250 108.210 79.560 108.750 ;
        RECT 79.720 108.210 81.050 108.750 ;
        RECT 81.210 108.740 82.250 109.880 ;
        RECT 82.690 109.870 83.970 110.380 ;
        RECT 84.170 109.880 85.480 110.390 ;
        RECT 82.690 108.740 83.730 109.870 ;
        RECT 81.210 108.210 82.480 108.740 ;
        RECT 75.840 107.650 76.520 108.210 ;
        RECT 77.390 107.660 78.070 108.210 ;
        RECT 78.880 107.670 79.560 108.210 ;
        RECT 80.370 107.670 81.050 108.210 ;
        RECT 81.800 107.670 82.480 108.210 ;
        RECT 82.690 108.200 83.990 108.740 ;
        RECT 84.170 108.210 85.210 109.880 ;
        RECT 83.310 107.670 83.990 108.200 ;
        RECT 74.620 105.500 75.640 107.650 ;
        RECT 75.840 107.080 77.150 107.650 ;
        RECT 77.390 107.170 78.600 107.660 ;
        RECT 78.880 107.170 80.110 107.670 ;
        RECT 80.370 107.170 81.580 107.670 ;
        RECT 76.110 105.490 77.150 107.080 ;
        RECT 77.560 105.480 78.600 107.170 ;
        RECT 79.070 105.490 80.110 107.170 ;
        RECT 80.540 105.490 81.580 107.170 ;
        RECT 81.800 107.160 83.070 107.670 ;
        RECT 83.310 107.160 84.540 107.670 ;
        RECT 82.030 105.490 83.070 107.160 ;
        RECT 83.500 105.490 84.540 107.160 ;
        RECT 118.590 99.125 119.785 112.160 ;
        RECT 121.215 110.435 123.385 112.160 ;
        RECT 121.230 109.585 121.535 110.435 ;
        RECT 121.925 109.885 122.270 110.145 ;
        RECT 121.955 109.865 122.245 109.885 ;
        RECT 121.765 109.585 121.995 109.660 ;
        RECT 121.230 108.725 121.995 109.585 ;
        RECT 121.250 105.720 121.995 108.725 ;
        RECT 121.765 105.660 121.995 105.720 ;
        RECT 122.205 109.550 122.435 109.660 ;
        RECT 122.205 105.925 123.120 109.550 ;
        RECT 122.205 105.755 123.180 105.925 ;
        RECT 122.205 105.660 122.435 105.755 ;
        RECT 122.890 105.465 123.180 105.755 ;
        RECT 123.600 105.720 124.015 115.625 ;
        RECT 123.785 105.655 124.015 105.720 ;
        RECT 124.225 115.595 124.455 115.655 ;
        RECT 124.695 115.595 125.140 116.490 ;
        RECT 125.535 115.890 125.880 116.150 ;
        RECT 125.555 115.860 125.845 115.890 ;
        RECT 127.115 115.880 127.460 116.140 ;
        RECT 127.135 115.860 127.425 115.880 ;
        RECT 125.365 115.595 125.595 115.655 ;
        RECT 124.225 105.745 125.595 115.595 ;
        RECT 124.225 105.655 124.455 105.745 ;
        RECT 125.365 105.655 125.595 105.745 ;
        RECT 125.805 115.595 126.035 115.655 ;
        RECT 126.390 115.595 126.650 115.625 ;
        RECT 126.945 115.595 127.175 115.655 ;
        RECT 125.805 105.745 127.175 115.595 ;
        RECT 125.805 105.655 126.035 105.745 ;
        RECT 126.945 105.655 127.175 105.745 ;
        RECT 127.385 115.605 127.615 115.655 ;
        RECT 127.870 115.605 128.315 116.490 ;
        RECT 128.690 115.895 129.035 116.155 ;
        RECT 134.470 116.040 134.970 117.510 ;
        RECT 128.715 115.860 129.005 115.895 ;
        RECT 128.525 115.605 128.755 115.655 ;
        RECT 127.385 105.755 128.755 115.605 ;
        RECT 127.385 105.655 127.615 105.755 ;
        RECT 128.525 105.655 128.755 105.755 ;
        RECT 128.965 115.625 129.195 115.655 ;
        RECT 128.965 115.305 129.410 115.625 ;
        RECT 128.965 105.720 129.400 115.305 ;
        RECT 143.840 114.000 146.560 114.800 ;
        RECT 128.965 105.655 129.195 105.720 ;
        RECT 121.955 105.435 122.245 105.455 ;
        RECT 121.600 104.945 122.600 105.435 ;
        RECT 122.890 105.140 129.040 105.465 ;
        RECT 121.600 103.945 122.640 104.945 ;
        RECT 121.600 103.400 122.600 103.945 ;
        RECT 121.950 103.375 122.240 103.400 ;
        RECT 121.760 103.135 121.990 103.215 ;
        RECT 121.260 102.525 121.990 103.135 ;
        RECT 121.250 102.290 121.990 102.525 ;
        RECT 121.250 101.520 121.505 102.290 ;
        RECT 121.750 102.270 121.990 102.290 ;
        RECT 121.760 102.215 121.990 102.270 ;
        RECT 122.200 103.165 122.430 103.215 ;
        RECT 122.890 103.165 123.180 105.140 ;
        RECT 129.995 104.705 130.995 105.705 ;
        RECT 145.180 105.345 145.570 107.855 ;
        RECT 142.885 104.955 145.570 105.345 ;
        RECT 124.385 104.250 124.615 104.540 ;
        RECT 127.865 104.515 128.245 104.590 ;
        RECT 130.355 104.515 130.580 104.705 ;
        RECT 127.865 104.290 130.580 104.515 ;
        RECT 124.405 103.675 124.590 104.250 ;
        RECT 127.865 104.230 128.245 104.290 ;
        RECT 134.320 104.210 134.580 104.530 ;
        RECT 129.955 103.955 130.985 104.130 ;
        RECT 123.950 103.375 129.050 103.675 ;
        RECT 123.975 103.370 124.265 103.375 ;
        RECT 125.555 103.370 125.845 103.375 ;
        RECT 127.135 103.370 127.425 103.375 ;
        RECT 128.715 103.370 129.005 103.375 ;
        RECT 129.245 103.345 130.985 103.955 ;
        RECT 122.200 102.300 123.240 103.165 ;
        RECT 123.785 103.120 124.015 103.210 ;
        RECT 122.200 102.215 122.430 102.300 ;
        RECT 121.950 102.025 122.240 102.055 ;
        RECT 121.905 101.765 122.250 102.025 ;
        RECT 121.240 101.485 121.505 101.520 ;
        RECT 106.520 97.930 119.785 99.125 ;
        RECT 69.130 90.285 70.440 90.340 ;
        RECT 106.520 90.285 107.715 97.930 ;
        RECT 121.220 97.455 123.370 101.485 ;
        RECT 123.620 98.285 124.015 103.120 ;
        RECT 123.785 98.210 124.015 98.285 ;
        RECT 124.225 103.145 124.455 103.210 ;
        RECT 125.365 103.145 125.595 103.210 ;
        RECT 124.225 98.305 125.595 103.145 ;
        RECT 124.225 98.210 124.455 98.305 ;
        RECT 123.975 98.020 124.265 98.050 ;
        RECT 123.950 97.760 124.295 98.020 ;
        RECT 124.725 97.495 125.085 98.305 ;
        RECT 125.365 98.210 125.595 98.305 ;
        RECT 125.805 103.170 126.035 103.210 ;
        RECT 126.945 103.170 127.175 103.210 ;
        RECT 125.805 98.330 127.175 103.170 ;
        RECT 125.805 98.210 126.035 98.330 ;
        RECT 126.345 98.325 126.605 98.330 ;
        RECT 126.945 98.210 127.175 98.330 ;
        RECT 127.385 103.125 127.615 103.210 ;
        RECT 128.525 103.125 128.755 103.210 ;
        RECT 127.385 98.285 128.755 103.125 ;
        RECT 127.385 98.210 127.615 98.285 ;
        RECT 125.555 98.025 125.845 98.050 ;
        RECT 127.135 98.025 127.425 98.050 ;
        RECT 125.530 97.765 125.875 98.025 ;
        RECT 127.115 97.765 127.460 98.025 ;
        RECT 127.850 97.495 128.210 98.285 ;
        RECT 128.525 98.210 128.755 98.285 ;
        RECT 128.965 103.170 129.195 103.210 ;
        RECT 129.350 103.170 130.985 103.345 ;
        RECT 142.760 103.300 143.080 103.560 ;
        RECT 128.965 103.040 130.985 103.170 ;
        RECT 128.965 102.580 130.285 103.040 ;
        RECT 128.965 98.310 129.400 102.580 ;
        RECT 128.965 98.210 129.195 98.310 ;
        RECT 128.715 98.025 129.005 98.050 ;
        RECT 128.700 97.765 129.045 98.025 ;
        RECT 121.220 97.410 123.400 97.455 ;
        RECT 121.220 97.335 123.420 97.410 ;
        RECT 121.230 97.010 123.420 97.335 ;
        RECT 124.725 97.135 128.210 97.495 ;
        RECT 124.725 97.105 128.155 97.135 ;
        RECT 121.230 97.000 123.400 97.010 ;
        RECT 121.325 96.580 122.590 97.000 ;
        RECT 134.110 96.580 135.310 98.080 ;
        RECT 121.325 96.430 135.310 96.580 ;
        RECT 69.130 89.090 107.715 90.285 ;
        RECT 108.905 96.380 135.310 96.430 ;
        RECT 143.870 96.380 144.670 99.580 ;
        RECT 150.420 98.840 150.770 99.665 ;
        RECT 150.075 98.560 150.770 98.840 ;
        RECT 150.030 98.280 150.770 98.560 ;
        RECT 150.075 98.060 150.770 98.280 ;
        RECT 150.420 97.535 150.770 98.060 ;
        RECT 151.950 97.550 153.705 99.665 ;
        RECT 154.900 97.550 156.655 99.665 ;
        RECT 157.880 99.645 158.130 99.650 ;
        RECT 157.865 98.690 158.750 99.645 ;
        RECT 151.960 97.545 152.210 97.550 ;
        RECT 153.440 97.545 153.690 97.550 ;
        RECT 154.920 97.545 155.170 97.550 ;
        RECT 156.400 97.545 156.650 97.550 ;
        RECT 157.865 97.535 158.860 98.690 ;
        RECT 150.480 96.930 150.730 96.955 ;
        RECT 151.960 96.930 152.210 96.955 ;
        RECT 153.440 96.945 153.690 96.955 ;
        RECT 154.920 96.945 155.170 96.955 ;
        RECT 156.400 96.945 156.650 96.955 ;
        RECT 157.880 96.945 158.130 96.955 ;
        RECT 108.905 95.580 144.670 96.380 ;
        RECT 108.905 95.380 135.310 95.580 ;
        RECT 108.905 95.165 122.590 95.380 ;
        RECT 125.745 95.225 130.890 95.380 ;
        RECT 69.130 89.040 70.440 89.090 ;
        RECT 75.005 87.935 92.760 88.225 ;
        RECT 108.905 88.065 110.170 95.165 ;
        RECT 97.775 87.935 110.170 88.065 ;
        RECT 75.005 87.855 110.170 87.935 ;
        RECT 124.530 94.670 130.890 95.225 ;
        RECT 124.530 94.235 130.780 94.670 ;
        RECT 124.530 90.950 126.210 94.235 ;
        RECT 126.800 93.600 127.050 93.660 ;
        RECT 128.280 93.600 128.530 93.660 ;
        RECT 129.760 93.600 130.010 93.660 ;
        RECT 131.240 93.600 131.490 93.660 ;
        RECT 132.720 93.600 132.970 93.660 ;
        RECT 134.200 93.600 134.450 93.660 ;
        RECT 135.680 93.600 135.930 93.660 ;
        RECT 137.160 93.600 137.410 93.660 ;
        RECT 138.640 93.600 138.890 93.660 ;
        RECT 140.120 93.600 140.370 93.660 ;
        RECT 141.600 93.600 141.850 93.660 ;
        RECT 143.080 93.600 143.330 93.660 ;
        RECT 144.560 93.600 144.810 93.660 ;
        RECT 146.040 93.600 146.290 93.660 ;
        RECT 147.520 93.600 147.770 93.660 ;
        RECT 149.000 93.600 149.250 93.660 ;
        RECT 126.800 91.600 128.600 93.600 ;
        RECT 129.700 91.600 131.500 93.600 ;
        RECT 132.700 91.600 134.500 93.600 ;
        RECT 135.680 91.600 137.500 93.600 ;
        RECT 138.600 91.600 140.400 93.600 ;
        RECT 141.600 91.600 143.400 93.600 ;
        RECT 144.500 91.600 146.300 93.600 ;
        RECT 147.500 91.600 149.300 93.600 ;
        RECT 126.800 91.555 127.050 91.600 ;
        RECT 128.280 91.555 128.530 91.600 ;
        RECT 129.760 91.555 130.010 91.600 ;
        RECT 131.240 91.555 131.490 91.600 ;
        RECT 132.720 91.555 132.970 91.600 ;
        RECT 134.200 91.555 134.450 91.600 ;
        RECT 135.680 91.555 135.930 91.600 ;
        RECT 137.160 91.555 137.410 91.600 ;
        RECT 138.640 91.555 138.890 91.600 ;
        RECT 140.120 91.555 140.370 91.600 ;
        RECT 141.600 91.555 141.850 91.600 ;
        RECT 143.080 91.555 143.330 91.600 ;
        RECT 144.560 91.555 144.810 91.600 ;
        RECT 146.040 91.555 146.290 91.600 ;
        RECT 147.520 91.555 147.770 91.600 ;
        RECT 149.000 91.555 149.250 91.600 ;
        RECT 126.800 90.950 127.050 90.965 ;
        RECT 124.530 88.860 127.050 90.950 ;
        RECT 128.280 90.800 128.530 90.965 ;
        RECT 129.760 90.800 130.010 90.965 ;
        RECT 131.240 90.800 131.490 90.965 ;
        RECT 132.720 90.800 132.970 90.965 ;
        RECT 134.200 90.900 134.450 90.965 ;
        RECT 135.680 90.900 135.930 90.965 ;
        RECT 128.200 88.860 130.010 90.800 ;
        RECT 124.530 87.885 127.010 88.860 ;
        RECT 128.200 88.800 130.000 88.860 ;
        RECT 131.200 88.800 133.000 90.800 ;
        RECT 134.200 88.900 136.000 90.900 ;
        RECT 137.160 90.800 137.410 90.965 ;
        RECT 138.640 90.800 138.890 90.965 ;
        RECT 140.120 90.800 140.370 90.965 ;
        RECT 141.600 90.800 141.850 90.965 ;
        RECT 143.080 90.900 143.330 90.965 ;
        RECT 144.560 90.900 144.810 90.965 ;
        RECT 146.040 90.900 146.290 90.965 ;
        RECT 147.520 90.900 147.770 90.965 ;
        RECT 134.200 88.860 134.450 88.900 ;
        RECT 135.680 88.860 135.930 88.900 ;
        RECT 137.100 88.800 138.900 90.800 ;
        RECT 140.100 88.800 141.900 90.800 ;
        RECT 143.000 88.900 144.810 90.900 ;
        RECT 146.000 88.900 147.800 90.900 ;
        RECT 149.000 90.800 149.250 90.965 ;
        RECT 149.760 90.800 150.040 95.950 ;
        RECT 150.435 94.850 152.210 96.930 ;
        RECT 153.410 94.850 155.170 96.945 ;
        RECT 150.435 94.815 152.190 94.850 ;
        RECT 153.410 94.830 155.165 94.850 ;
        RECT 156.380 94.830 158.135 96.945 ;
        RECT 150.480 93.600 150.730 93.660 ;
        RECT 151.960 93.600 152.210 93.660 ;
        RECT 150.400 91.600 152.210 93.600 ;
        RECT 153.400 91.700 155.200 93.700 ;
        RECT 156.400 93.600 156.650 93.660 ;
        RECT 157.880 93.600 158.130 93.660 ;
        RECT 150.480 91.555 150.730 91.600 ;
        RECT 151.960 91.555 152.210 91.600 ;
        RECT 153.440 91.555 153.690 91.700 ;
        RECT 154.920 91.555 155.170 91.700 ;
        RECT 156.400 91.600 158.200 93.600 ;
        RECT 156.400 91.555 156.650 91.600 ;
        RECT 157.880 91.555 158.130 91.600 ;
        RECT 150.480 90.800 150.730 90.965 ;
        RECT 151.960 90.800 152.210 90.965 ;
        RECT 153.440 90.800 153.690 90.965 ;
        RECT 154.920 90.800 155.170 90.965 ;
        RECT 156.400 90.800 156.650 90.965 ;
        RECT 157.880 90.900 158.130 90.965 ;
        RECT 158.520 90.900 158.860 97.535 ;
        RECT 143.080 88.860 143.330 88.900 ;
        RECT 144.560 88.860 144.810 88.900 ;
        RECT 146.040 88.860 146.290 88.900 ;
        RECT 147.520 88.860 147.770 88.900 ;
        RECT 149.000 88.800 150.800 90.800 ;
        RECT 151.900 88.800 153.700 90.800 ;
        RECT 154.900 88.800 156.700 90.800 ;
        RECT 157.880 88.860 158.860 90.900 ;
        RECT 157.900 88.775 158.860 88.860 ;
        RECT 157.900 88.725 158.600 88.775 ;
        RECT 124.530 87.875 144.875 87.885 ;
        RECT 114.255 87.855 144.875 87.875 ;
        RECT 75.005 87.470 144.875 87.855 ;
        RECT 75.005 87.140 81.375 87.470 ;
        RECT 92.005 87.320 144.875 87.470 ;
        RECT 92.005 87.310 123.720 87.320 ;
        RECT 75.000 87.025 81.375 87.140 ;
        RECT 75.000 86.665 81.445 87.025 ;
        RECT 75.000 86.530 88.975 86.665 ;
        RECT 75.000 86.085 75.875 86.530 ;
        RECT 81.015 86.435 88.975 86.530 ;
        RECT 75.000 85.860 75.885 86.085 ;
        RECT 76.595 86.000 77.815 86.085 ;
        RECT 76.595 85.945 77.830 86.000 ;
        RECT 75.000 81.185 75.875 85.860 ;
        RECT 76.585 85.715 78.585 85.945 ;
        RECT 76.195 84.465 76.425 85.665 ;
        RECT 76.970 84.465 78.135 85.715 ;
        RECT 78.745 84.465 78.975 85.665 ;
        RECT 76.195 83.675 78.975 84.465 ;
        RECT 80.735 85.510 80.965 86.230 ;
        RECT 80.735 85.485 81.100 85.510 ;
        RECT 81.260 85.485 81.580 85.540 ;
        RECT 80.735 85.335 81.580 85.485 ;
        RECT 80.735 85.305 81.100 85.335 ;
        RECT 80.735 84.230 80.965 85.305 ;
        RECT 81.260 85.280 81.580 85.335 ;
        RECT 83.865 84.055 85.680 86.435 ;
        RECT 89.025 86.195 89.255 86.230 ;
        RECT 89.880 86.195 90.580 87.165 ;
        RECT 92.005 87.140 98.530 87.310 ;
        RECT 108.835 87.290 123.720 87.310 ;
        RECT 124.740 87.290 140.700 87.320 ;
        RECT 89.025 84.285 90.580 86.195 ;
        RECT 89.025 84.230 89.255 84.285 ;
        RECT 81.265 84.025 88.895 84.055 ;
        RECT 81.015 83.795 88.975 84.025 ;
        RECT 76.195 81.705 76.425 83.675 ;
        RECT 78.745 83.005 78.975 83.675 ;
        RECT 78.745 82.725 81.610 83.005 ;
        RECT 78.745 82.635 89.030 82.725 ;
        RECT 78.745 81.705 78.975 82.635 ;
        RECT 81.170 82.485 89.030 82.635 ;
        RECT 81.110 82.255 89.110 82.485 ;
        RECT 80.675 81.765 80.905 82.205 ;
        RECT 89.315 82.195 89.545 82.205 ;
        RECT 81.395 81.765 82.395 81.835 ;
        RECT 89.315 81.765 89.550 82.195 ;
        RECT 76.585 81.425 78.585 81.655 ;
        RECT 76.675 81.185 78.500 81.425 ;
        RECT 75.000 80.695 78.500 81.185 ;
        RECT 75.000 75.860 75.875 80.695 ;
        RECT 76.675 80.515 78.500 80.695 ;
        RECT 80.675 80.875 89.550 81.765 ;
        RECT 76.585 80.285 78.585 80.515 ;
        RECT 80.675 80.245 80.905 80.875 ;
        RECT 81.395 80.820 82.395 80.875 ;
        RECT 89.315 80.310 89.550 80.875 ;
        RECT 89.315 80.245 89.545 80.310 ;
        RECT 76.195 78.800 76.425 80.235 ;
        RECT 78.745 78.800 78.975 80.235 ;
        RECT 81.110 79.965 89.110 80.195 ;
        RECT 81.180 79.840 89.010 79.965 ;
        RECT 81.200 79.055 89.000 79.840 ;
        RECT 81.110 78.825 89.110 79.055 ;
        RECT 76.195 77.460 78.975 78.800 ;
        RECT 80.675 78.750 80.905 78.775 ;
        RECT 76.195 76.275 76.425 77.460 ;
        RECT 76.770 76.225 78.365 77.460 ;
        RECT 78.745 76.570 78.975 77.460 ;
        RECT 80.670 78.305 80.905 78.750 ;
        RECT 89.315 78.750 89.545 78.775 ;
        RECT 80.670 78.295 81.085 78.305 ;
        RECT 81.225 78.295 82.225 78.365 ;
        RECT 80.670 78.290 82.225 78.295 ;
        RECT 82.635 78.290 84.255 78.295 ;
        RECT 89.315 78.290 89.550 78.750 ;
        RECT 80.670 77.400 89.550 78.290 ;
        RECT 80.670 77.385 82.225 77.400 ;
        RECT 82.635 77.395 84.255 77.400 ;
        RECT 80.670 77.295 81.085 77.385 ;
        RECT 81.225 77.335 82.225 77.385 ;
        RECT 80.670 76.865 80.905 77.295 ;
        RECT 80.675 76.815 80.905 76.865 ;
        RECT 89.315 76.865 89.550 77.400 ;
        RECT 89.315 76.815 89.545 76.865 ;
        RECT 81.110 76.570 89.110 76.765 ;
        RECT 78.745 76.535 89.110 76.570 ;
        RECT 78.745 76.390 89.030 76.535 ;
        RECT 78.745 76.375 81.245 76.390 ;
        RECT 78.745 76.275 78.975 76.375 ;
        RECT 76.585 75.995 78.585 76.225 ;
        RECT 89.880 76.115 90.580 84.285 ;
        RECT 84.955 75.985 85.230 76.055 ;
        RECT 79.260 75.860 85.230 75.985 ;
        RECT 75.000 75.845 76.405 75.860 ;
        RECT 78.750 75.845 85.230 75.860 ;
        RECT 75.000 75.795 85.230 75.845 ;
        RECT 75.000 75.670 79.450 75.795 ;
        RECT 84.955 75.720 85.230 75.795 ;
        RECT 75.000 70.390 75.875 75.670 ;
        RECT 77.825 75.365 81.610 75.370 ;
        RECT 77.825 75.300 85.060 75.365 ;
        RECT 76.645 75.175 85.060 75.300 ;
        RECT 76.645 75.085 85.105 75.175 ;
        RECT 76.585 75.075 85.105 75.085 ;
        RECT 76.585 74.855 78.585 75.075 ;
        RECT 81.105 74.945 85.105 75.075 ;
        RECT 76.195 73.425 76.425 74.805 ;
        RECT 78.745 73.425 78.975 74.805 ;
        RECT 76.195 72.470 78.975 73.425 ;
        RECT 76.195 70.845 76.425 72.470 ;
        RECT 78.745 70.845 78.975 72.470 ;
        RECT 80.670 73.640 80.900 74.895 ;
        RECT 82.340 73.640 83.725 74.945 ;
        RECT 85.310 73.640 85.540 74.895 ;
        RECT 85.905 74.435 90.580 76.115 ;
        RECT 87.265 74.095 87.540 74.125 ;
        RECT 87.250 73.840 87.580 74.095 ;
        RECT 87.265 73.820 87.555 73.840 ;
        RECT 87.265 73.790 87.540 73.820 ;
        RECT 80.670 73.570 85.540 73.640 ;
        RECT 87.075 73.570 87.305 73.615 ;
        RECT 80.670 72.295 85.545 73.570 ;
        RECT 80.670 70.935 80.900 72.295 ;
        RECT 85.310 70.935 85.545 72.295 ;
        RECT 76.585 70.565 78.585 70.795 ;
        RECT 76.650 70.390 78.520 70.565 ;
        RECT 75.000 69.835 78.520 70.390 ;
        RECT 75.000 64.730 75.875 69.835 ;
        RECT 76.650 69.655 78.520 69.835 ;
        RECT 76.585 69.425 78.585 69.655 ;
        RECT 80.710 69.465 80.870 70.935 ;
        RECT 85.340 70.925 85.545 70.935 ;
        RECT 81.105 70.655 85.105 70.885 ;
        RECT 81.185 70.410 85.010 70.655 ;
        RECT 87.065 70.410 87.305 73.570 ;
        RECT 81.185 69.920 87.305 70.410 ;
        RECT 81.185 69.745 85.010 69.920 ;
        RECT 81.105 69.515 85.105 69.745 ;
        RECT 76.195 67.980 76.425 69.375 ;
        RECT 78.745 67.980 78.975 69.375 ;
        RECT 76.195 67.025 78.975 67.980 ;
        RECT 76.195 65.415 76.425 67.025 ;
        RECT 78.745 65.415 78.975 67.025 ;
        RECT 80.670 68.090 80.900 69.465 ;
        RECT 85.310 69.350 85.540 69.465 ;
        RECT 85.310 68.715 85.545 69.350 ;
        RECT 87.065 68.715 87.305 69.920 ;
        RECT 85.310 68.090 85.540 68.715 ;
        RECT 87.075 68.615 87.305 68.715 ;
        RECT 87.515 73.600 87.745 73.615 ;
        RECT 88.165 73.600 88.645 74.435 ;
        RECT 87.515 68.675 88.655 73.600 ;
        RECT 87.515 68.615 87.745 68.675 ;
        RECT 87.265 68.405 87.555 68.410 ;
        RECT 87.250 68.150 87.580 68.405 ;
        RECT 80.670 66.745 85.540 68.090 ;
        RECT 80.670 65.505 80.900 66.745 ;
        RECT 85.310 65.505 85.540 66.745 ;
        RECT 76.585 65.340 78.585 65.365 ;
        RECT 81.105 65.340 85.105 65.455 ;
        RECT 76.585 65.265 78.590 65.340 ;
        RECT 79.125 65.265 85.105 65.340 ;
        RECT 76.585 65.225 85.105 65.265 ;
        RECT 76.585 65.135 85.040 65.225 ;
        RECT 76.640 65.000 85.040 65.135 ;
        RECT 75.000 64.290 76.860 64.730 ;
        RECT 75.000 64.280 77.850 64.290 ;
        RECT 75.000 63.935 78.520 64.280 ;
        RECT 75.000 62.310 76.860 63.935 ;
        RECT 77.660 63.785 78.520 63.935 ;
        RECT 77.155 63.595 77.405 63.610 ;
        RECT 77.155 63.305 77.430 63.595 ;
        RECT 77.590 63.555 78.590 63.785 ;
        RECT 79.010 63.690 79.280 65.000 ;
        RECT 89.880 64.570 90.580 74.435 ;
        RECT 84.300 64.235 90.580 64.570 ;
        RECT 81.185 64.095 90.580 64.235 ;
        RECT 81.185 63.870 85.045 64.095 ;
        RECT 77.155 63.275 77.405 63.305 ;
        RECT 77.590 63.115 78.590 63.345 ;
        RECT 78.735 63.270 80.925 63.690 ;
        RECT 81.120 63.640 85.120 63.870 ;
        RECT 85.355 63.680 85.605 63.700 ;
        RECT 81.120 63.200 85.120 63.430 ;
        RECT 85.325 63.390 85.605 63.680 ;
        RECT 85.355 63.365 85.605 63.390 ;
        RECT 77.660 62.975 78.545 63.115 ;
        RECT 81.170 63.035 85.095 63.200 ;
        RECT 78.730 62.975 85.095 63.035 ;
        RECT 77.660 62.920 85.095 62.975 ;
        RECT 77.660 62.850 81.540 62.920 ;
        RECT 78.215 62.735 81.540 62.850 ;
        RECT 89.880 62.770 90.580 64.095 ;
        RECT 75.000 62.265 77.385 62.310 ;
        RECT 42.055 61.285 42.315 61.605 ;
        RECT 42.115 60.640 42.255 61.285 ;
        RECT 49.120 60.640 49.380 60.730 ;
        RECT 42.115 60.500 49.380 60.640 ;
        RECT 75.000 60.535 75.875 62.265 ;
        RECT 76.240 61.990 77.385 62.265 ;
        RECT 79.570 62.105 79.975 62.735 ;
        RECT 88.575 62.235 90.580 62.770 ;
        RECT 76.240 61.925 78.490 61.990 ;
        RECT 76.680 61.760 78.490 61.925 ;
        RECT 76.165 61.570 76.415 61.595 ;
        RECT 76.165 61.280 76.435 61.570 ;
        RECT 76.595 61.530 78.595 61.760 ;
        RECT 79.555 61.740 79.980 62.105 ;
        RECT 81.220 62.090 90.580 62.235 ;
        RECT 81.220 61.845 89.075 62.090 ;
        RECT 76.165 61.260 76.415 61.280 ;
        RECT 76.595 61.090 78.595 61.320 ;
        RECT 78.745 61.230 80.935 61.740 ;
        RECT 81.125 61.615 89.125 61.845 ;
        RECT 89.355 61.655 89.605 61.670 ;
        RECT 78.745 61.225 79.445 61.230 ;
        RECT 80.445 61.225 80.935 61.230 ;
        RECT 81.125 61.175 89.125 61.405 ;
        RECT 89.330 61.365 89.605 61.655 ;
        RECT 89.355 61.335 89.605 61.365 ;
        RECT 76.665 60.925 78.530 61.090 ;
        RECT 79.415 60.925 80.415 61.000 ;
        RECT 81.200 60.925 89.050 61.175 ;
        RECT 76.665 60.630 89.050 60.925 ;
        RECT 89.880 60.690 90.580 62.090 ;
        RECT 92.000 86.665 98.530 87.140 ;
        RECT 92.000 86.530 105.975 86.665 ;
        RECT 92.000 86.085 92.875 86.530 ;
        RECT 98.015 86.435 105.975 86.530 ;
        RECT 92.000 85.860 92.885 86.085 ;
        RECT 93.595 86.000 94.815 86.085 ;
        RECT 93.595 85.945 94.830 86.000 ;
        RECT 92.000 81.185 92.875 85.860 ;
        RECT 93.585 85.715 95.585 85.945 ;
        RECT 93.195 84.465 93.425 85.665 ;
        RECT 93.970 84.465 95.135 85.715 ;
        RECT 95.745 84.465 95.975 85.665 ;
        RECT 93.195 83.675 95.975 84.465 ;
        RECT 97.735 85.510 97.965 86.230 ;
        RECT 97.735 85.485 98.100 85.510 ;
        RECT 98.260 85.485 98.580 85.540 ;
        RECT 97.735 85.335 98.580 85.485 ;
        RECT 97.735 85.305 98.100 85.335 ;
        RECT 97.735 84.230 97.965 85.305 ;
        RECT 98.260 85.280 98.580 85.335 ;
        RECT 100.865 84.055 102.680 86.435 ;
        RECT 106.025 86.195 106.255 86.230 ;
        RECT 106.880 86.195 107.580 87.165 ;
        RECT 108.835 87.120 123.530 87.290 ;
        RECT 108.835 86.920 115.590 87.120 ;
        RECT 108.835 86.665 115.445 86.920 ;
        RECT 108.835 86.530 122.975 86.665 ;
        RECT 108.835 86.425 109.875 86.530 ;
        RECT 115.015 86.435 122.975 86.530 ;
        RECT 106.025 84.285 107.580 86.195 ;
        RECT 106.025 84.230 106.255 84.285 ;
        RECT 98.265 84.025 105.895 84.055 ;
        RECT 98.015 83.795 105.975 84.025 ;
        RECT 93.195 81.705 93.425 83.675 ;
        RECT 95.745 83.005 95.975 83.675 ;
        RECT 95.745 82.725 98.610 83.005 ;
        RECT 95.745 82.635 106.030 82.725 ;
        RECT 95.745 81.705 95.975 82.635 ;
        RECT 98.170 82.485 106.030 82.635 ;
        RECT 98.110 82.255 106.110 82.485 ;
        RECT 97.675 81.765 97.905 82.205 ;
        RECT 106.315 82.195 106.545 82.205 ;
        RECT 98.395 81.765 99.395 81.835 ;
        RECT 106.315 81.765 106.550 82.195 ;
        RECT 93.585 81.425 95.585 81.655 ;
        RECT 93.675 81.185 95.500 81.425 ;
        RECT 92.000 80.695 95.500 81.185 ;
        RECT 92.000 75.860 92.875 80.695 ;
        RECT 93.675 80.515 95.500 80.695 ;
        RECT 97.675 80.875 106.550 81.765 ;
        RECT 93.585 80.285 95.585 80.515 ;
        RECT 97.675 80.245 97.905 80.875 ;
        RECT 98.395 80.820 99.395 80.875 ;
        RECT 106.315 80.310 106.550 80.875 ;
        RECT 106.315 80.245 106.545 80.310 ;
        RECT 93.195 78.800 93.425 80.235 ;
        RECT 95.745 78.800 95.975 80.235 ;
        RECT 98.110 79.965 106.110 80.195 ;
        RECT 98.180 79.840 106.010 79.965 ;
        RECT 98.200 79.055 106.000 79.840 ;
        RECT 98.110 78.825 106.110 79.055 ;
        RECT 93.195 77.460 95.975 78.800 ;
        RECT 97.675 78.750 97.905 78.775 ;
        RECT 93.195 76.275 93.425 77.460 ;
        RECT 93.770 76.225 95.365 77.460 ;
        RECT 95.745 76.570 95.975 77.460 ;
        RECT 97.670 78.305 97.905 78.750 ;
        RECT 106.315 78.750 106.545 78.775 ;
        RECT 97.670 78.295 98.085 78.305 ;
        RECT 98.225 78.295 99.225 78.365 ;
        RECT 97.670 78.290 99.225 78.295 ;
        RECT 99.635 78.290 101.255 78.295 ;
        RECT 106.315 78.290 106.550 78.750 ;
        RECT 97.670 77.400 106.550 78.290 ;
        RECT 97.670 77.385 99.225 77.400 ;
        RECT 99.635 77.395 101.255 77.400 ;
        RECT 97.670 77.295 98.085 77.385 ;
        RECT 98.225 77.335 99.225 77.385 ;
        RECT 97.670 76.865 97.905 77.295 ;
        RECT 97.675 76.815 97.905 76.865 ;
        RECT 106.315 76.865 106.550 77.400 ;
        RECT 106.315 76.815 106.545 76.865 ;
        RECT 98.110 76.570 106.110 76.765 ;
        RECT 95.745 76.535 106.110 76.570 ;
        RECT 95.745 76.390 106.030 76.535 ;
        RECT 95.745 76.375 98.245 76.390 ;
        RECT 95.745 76.275 95.975 76.375 ;
        RECT 93.585 75.995 95.585 76.225 ;
        RECT 106.880 76.115 107.580 84.285 ;
        RECT 101.955 75.985 102.230 76.055 ;
        RECT 96.260 75.860 102.230 75.985 ;
        RECT 92.000 75.845 93.405 75.860 ;
        RECT 95.750 75.845 102.230 75.860 ;
        RECT 92.000 75.795 102.230 75.845 ;
        RECT 92.000 75.670 96.450 75.795 ;
        RECT 101.955 75.720 102.230 75.795 ;
        RECT 92.000 70.390 92.875 75.670 ;
        RECT 94.825 75.365 98.610 75.370 ;
        RECT 94.825 75.300 102.060 75.365 ;
        RECT 93.645 75.175 102.060 75.300 ;
        RECT 93.645 75.085 102.105 75.175 ;
        RECT 93.585 75.075 102.105 75.085 ;
        RECT 93.585 74.855 95.585 75.075 ;
        RECT 98.105 74.945 102.105 75.075 ;
        RECT 93.195 73.425 93.425 74.805 ;
        RECT 95.745 73.425 95.975 74.805 ;
        RECT 93.195 72.470 95.975 73.425 ;
        RECT 93.195 70.845 93.425 72.470 ;
        RECT 95.745 70.845 95.975 72.470 ;
        RECT 97.670 73.640 97.900 74.895 ;
        RECT 99.340 73.640 100.725 74.945 ;
        RECT 102.310 73.640 102.540 74.895 ;
        RECT 102.905 74.435 107.580 76.115 ;
        RECT 104.265 74.095 104.540 74.125 ;
        RECT 104.250 73.840 104.580 74.095 ;
        RECT 104.265 73.820 104.555 73.840 ;
        RECT 104.265 73.790 104.540 73.820 ;
        RECT 97.670 73.570 102.540 73.640 ;
        RECT 104.075 73.570 104.305 73.615 ;
        RECT 97.670 72.295 102.545 73.570 ;
        RECT 97.670 70.935 97.900 72.295 ;
        RECT 102.310 70.935 102.545 72.295 ;
        RECT 93.585 70.565 95.585 70.795 ;
        RECT 93.650 70.390 95.520 70.565 ;
        RECT 92.000 69.835 95.520 70.390 ;
        RECT 92.000 64.730 92.875 69.835 ;
        RECT 93.650 69.655 95.520 69.835 ;
        RECT 93.585 69.425 95.585 69.655 ;
        RECT 97.710 69.465 97.870 70.935 ;
        RECT 102.340 70.925 102.545 70.935 ;
        RECT 98.105 70.655 102.105 70.885 ;
        RECT 98.185 70.410 102.010 70.655 ;
        RECT 104.065 70.410 104.305 73.570 ;
        RECT 98.185 69.920 104.305 70.410 ;
        RECT 98.185 69.745 102.010 69.920 ;
        RECT 98.105 69.515 102.105 69.745 ;
        RECT 93.195 67.980 93.425 69.375 ;
        RECT 95.745 67.980 95.975 69.375 ;
        RECT 93.195 67.025 95.975 67.980 ;
        RECT 93.195 65.415 93.425 67.025 ;
        RECT 95.745 65.415 95.975 67.025 ;
        RECT 97.670 68.090 97.900 69.465 ;
        RECT 102.310 69.350 102.540 69.465 ;
        RECT 102.310 68.715 102.545 69.350 ;
        RECT 104.065 68.715 104.305 69.920 ;
        RECT 102.310 68.090 102.540 68.715 ;
        RECT 104.075 68.615 104.305 68.715 ;
        RECT 104.515 73.600 104.745 73.615 ;
        RECT 105.165 73.600 105.645 74.435 ;
        RECT 104.515 68.675 105.655 73.600 ;
        RECT 104.515 68.615 104.745 68.675 ;
        RECT 104.265 68.405 104.555 68.410 ;
        RECT 104.250 68.150 104.580 68.405 ;
        RECT 97.670 66.745 102.540 68.090 ;
        RECT 97.670 65.505 97.900 66.745 ;
        RECT 102.310 65.505 102.540 66.745 ;
        RECT 93.585 65.340 95.585 65.365 ;
        RECT 98.105 65.340 102.105 65.455 ;
        RECT 93.585 65.265 95.590 65.340 ;
        RECT 96.125 65.265 102.105 65.340 ;
        RECT 93.585 65.225 102.105 65.265 ;
        RECT 93.585 65.135 102.040 65.225 ;
        RECT 93.640 65.000 102.040 65.135 ;
        RECT 92.000 64.290 93.860 64.730 ;
        RECT 92.000 64.280 94.850 64.290 ;
        RECT 92.000 63.935 95.520 64.280 ;
        RECT 92.000 62.310 93.860 63.935 ;
        RECT 94.660 63.785 95.520 63.935 ;
        RECT 94.155 63.595 94.405 63.610 ;
        RECT 94.155 63.305 94.430 63.595 ;
        RECT 94.590 63.555 95.590 63.785 ;
        RECT 96.010 63.690 96.280 65.000 ;
        RECT 106.880 64.570 107.580 74.435 ;
        RECT 101.300 64.235 107.580 64.570 ;
        RECT 98.185 64.095 107.580 64.235 ;
        RECT 98.185 63.870 102.045 64.095 ;
        RECT 94.155 63.275 94.405 63.305 ;
        RECT 94.590 63.115 95.590 63.345 ;
        RECT 95.735 63.270 97.925 63.690 ;
        RECT 98.120 63.640 102.120 63.870 ;
        RECT 102.355 63.680 102.605 63.700 ;
        RECT 98.120 63.200 102.120 63.430 ;
        RECT 102.325 63.390 102.605 63.680 ;
        RECT 102.355 63.365 102.605 63.390 ;
        RECT 94.660 62.975 95.545 63.115 ;
        RECT 98.170 63.035 102.095 63.200 ;
        RECT 95.730 62.975 102.095 63.035 ;
        RECT 94.660 62.920 102.095 62.975 ;
        RECT 94.660 62.850 98.540 62.920 ;
        RECT 95.215 62.735 98.540 62.850 ;
        RECT 106.880 62.770 107.580 64.095 ;
        RECT 92.000 62.265 94.385 62.310 ;
        RECT 76.665 60.560 81.730 60.630 ;
        RECT 78.205 60.555 81.730 60.560 ;
        RECT 49.120 60.410 49.380 60.500 ;
        RECT 46.080 60.235 46.400 60.240 ;
        RECT 79.415 60.235 80.415 60.555 ;
        RECT 92.000 60.535 92.875 62.265 ;
        RECT 93.240 61.990 94.385 62.265 ;
        RECT 96.570 62.105 96.975 62.735 ;
        RECT 105.575 62.235 107.580 62.770 ;
        RECT 93.240 61.925 95.490 61.990 ;
        RECT 93.680 61.760 95.490 61.925 ;
        RECT 93.165 61.570 93.415 61.595 ;
        RECT 93.165 61.280 93.435 61.570 ;
        RECT 93.595 61.530 95.595 61.760 ;
        RECT 96.555 61.740 96.980 62.105 ;
        RECT 98.220 62.090 107.580 62.235 ;
        RECT 98.220 61.845 106.075 62.090 ;
        RECT 93.165 61.260 93.415 61.280 ;
        RECT 93.595 61.090 95.595 61.320 ;
        RECT 95.745 61.230 97.935 61.740 ;
        RECT 98.125 61.615 106.125 61.845 ;
        RECT 106.355 61.655 106.605 61.670 ;
        RECT 95.745 61.225 96.445 61.230 ;
        RECT 97.445 61.225 97.935 61.230 ;
        RECT 98.125 61.175 106.125 61.405 ;
        RECT 106.330 61.365 106.605 61.655 ;
        RECT 106.355 61.335 106.605 61.365 ;
        RECT 93.665 60.925 95.530 61.090 ;
        RECT 96.415 60.925 97.415 61.000 ;
        RECT 98.200 60.925 106.050 61.175 ;
        RECT 93.665 60.630 106.050 60.925 ;
        RECT 106.880 60.690 107.580 62.090 ;
        RECT 109.000 86.085 109.875 86.425 ;
        RECT 109.000 85.860 109.885 86.085 ;
        RECT 110.595 86.000 111.815 86.085 ;
        RECT 110.595 85.945 111.830 86.000 ;
        RECT 109.000 81.185 109.875 85.860 ;
        RECT 110.585 85.715 112.585 85.945 ;
        RECT 110.195 84.465 110.425 85.665 ;
        RECT 110.970 84.465 112.135 85.715 ;
        RECT 112.745 84.465 112.975 85.665 ;
        RECT 110.195 83.675 112.975 84.465 ;
        RECT 114.735 85.510 114.965 86.230 ;
        RECT 114.735 85.485 115.100 85.510 ;
        RECT 115.260 85.485 115.580 85.540 ;
        RECT 114.735 85.335 115.580 85.485 ;
        RECT 114.735 85.305 115.100 85.335 ;
        RECT 114.735 84.230 114.965 85.305 ;
        RECT 115.260 85.280 115.580 85.335 ;
        RECT 117.865 84.055 119.680 86.435 ;
        RECT 123.025 86.195 123.255 86.230 ;
        RECT 123.880 86.195 124.580 87.165 ;
        RECT 124.790 87.130 140.470 87.290 ;
        RECT 124.790 87.120 132.605 87.130 ;
        RECT 123.025 84.285 124.580 86.195 ;
        RECT 123.025 84.230 123.255 84.285 ;
        RECT 115.265 84.025 122.895 84.055 ;
        RECT 115.015 83.795 122.975 84.025 ;
        RECT 110.195 81.705 110.425 83.675 ;
        RECT 112.745 83.005 112.975 83.675 ;
        RECT 112.745 82.725 115.610 83.005 ;
        RECT 112.745 82.635 123.030 82.725 ;
        RECT 112.745 81.705 112.975 82.635 ;
        RECT 115.170 82.485 123.030 82.635 ;
        RECT 115.110 82.255 123.110 82.485 ;
        RECT 114.675 81.765 114.905 82.205 ;
        RECT 123.315 82.195 123.545 82.205 ;
        RECT 115.395 81.765 116.395 81.835 ;
        RECT 123.315 81.765 123.550 82.195 ;
        RECT 110.585 81.425 112.585 81.655 ;
        RECT 110.675 81.185 112.500 81.425 ;
        RECT 109.000 80.695 112.500 81.185 ;
        RECT 109.000 75.860 109.875 80.695 ;
        RECT 110.675 80.515 112.500 80.695 ;
        RECT 114.675 80.875 123.550 81.765 ;
        RECT 110.585 80.285 112.585 80.515 ;
        RECT 114.675 80.245 114.905 80.875 ;
        RECT 115.395 80.820 116.395 80.875 ;
        RECT 123.315 80.310 123.550 80.875 ;
        RECT 123.315 80.245 123.545 80.310 ;
        RECT 110.195 78.800 110.425 80.235 ;
        RECT 112.745 78.800 112.975 80.235 ;
        RECT 115.110 79.965 123.110 80.195 ;
        RECT 115.180 79.840 123.010 79.965 ;
        RECT 115.200 79.055 123.000 79.840 ;
        RECT 115.110 78.825 123.110 79.055 ;
        RECT 110.195 77.460 112.975 78.800 ;
        RECT 114.675 78.750 114.905 78.775 ;
        RECT 110.195 76.275 110.425 77.460 ;
        RECT 110.770 76.225 112.365 77.460 ;
        RECT 112.745 76.570 112.975 77.460 ;
        RECT 114.670 78.305 114.905 78.750 ;
        RECT 123.315 78.750 123.545 78.775 ;
        RECT 114.670 78.295 115.085 78.305 ;
        RECT 115.225 78.295 116.225 78.365 ;
        RECT 114.670 78.290 116.225 78.295 ;
        RECT 116.635 78.290 118.255 78.295 ;
        RECT 123.315 78.290 123.550 78.750 ;
        RECT 114.670 77.400 123.550 78.290 ;
        RECT 114.670 77.385 116.225 77.400 ;
        RECT 116.635 77.395 118.255 77.400 ;
        RECT 114.670 77.295 115.085 77.385 ;
        RECT 115.225 77.335 116.225 77.385 ;
        RECT 114.670 76.865 114.905 77.295 ;
        RECT 114.675 76.815 114.905 76.865 ;
        RECT 123.315 76.865 123.550 77.400 ;
        RECT 123.315 76.815 123.545 76.865 ;
        RECT 115.110 76.570 123.110 76.765 ;
        RECT 112.745 76.535 123.110 76.570 ;
        RECT 112.745 76.390 123.030 76.535 ;
        RECT 112.745 76.375 115.245 76.390 ;
        RECT 112.745 76.275 112.975 76.375 ;
        RECT 110.585 75.995 112.585 76.225 ;
        RECT 123.880 76.115 124.580 84.285 ;
        RECT 118.955 75.985 119.230 76.055 ;
        RECT 113.260 75.860 119.230 75.985 ;
        RECT 109.000 75.845 110.405 75.860 ;
        RECT 112.750 75.845 119.230 75.860 ;
        RECT 109.000 75.795 119.230 75.845 ;
        RECT 109.000 75.670 113.450 75.795 ;
        RECT 118.955 75.720 119.230 75.795 ;
        RECT 109.000 70.390 109.875 75.670 ;
        RECT 111.825 75.365 115.610 75.370 ;
        RECT 111.825 75.300 119.060 75.365 ;
        RECT 110.645 75.175 119.060 75.300 ;
        RECT 110.645 75.085 119.105 75.175 ;
        RECT 110.585 75.075 119.105 75.085 ;
        RECT 110.585 74.855 112.585 75.075 ;
        RECT 115.105 74.945 119.105 75.075 ;
        RECT 110.195 73.425 110.425 74.805 ;
        RECT 112.745 73.425 112.975 74.805 ;
        RECT 110.195 72.470 112.975 73.425 ;
        RECT 110.195 70.845 110.425 72.470 ;
        RECT 112.745 70.845 112.975 72.470 ;
        RECT 114.670 73.640 114.900 74.895 ;
        RECT 116.340 73.640 117.725 74.945 ;
        RECT 119.310 73.640 119.540 74.895 ;
        RECT 119.905 74.435 124.580 76.115 ;
        RECT 121.265 74.095 121.540 74.125 ;
        RECT 121.250 73.840 121.580 74.095 ;
        RECT 121.265 73.820 121.555 73.840 ;
        RECT 121.265 73.790 121.540 73.820 ;
        RECT 114.670 73.570 119.540 73.640 ;
        RECT 121.075 73.570 121.305 73.615 ;
        RECT 114.670 72.295 119.545 73.570 ;
        RECT 114.670 70.935 114.900 72.295 ;
        RECT 119.310 70.935 119.545 72.295 ;
        RECT 110.585 70.565 112.585 70.795 ;
        RECT 110.650 70.390 112.520 70.565 ;
        RECT 109.000 69.835 112.520 70.390 ;
        RECT 109.000 64.730 109.875 69.835 ;
        RECT 110.650 69.655 112.520 69.835 ;
        RECT 110.585 69.425 112.585 69.655 ;
        RECT 114.710 69.465 114.870 70.935 ;
        RECT 119.340 70.925 119.545 70.935 ;
        RECT 115.105 70.655 119.105 70.885 ;
        RECT 115.185 70.410 119.010 70.655 ;
        RECT 121.065 70.410 121.305 73.570 ;
        RECT 115.185 69.920 121.305 70.410 ;
        RECT 115.185 69.745 119.010 69.920 ;
        RECT 115.105 69.515 119.105 69.745 ;
        RECT 110.195 67.980 110.425 69.375 ;
        RECT 112.745 67.980 112.975 69.375 ;
        RECT 110.195 67.025 112.975 67.980 ;
        RECT 110.195 65.415 110.425 67.025 ;
        RECT 112.745 65.415 112.975 67.025 ;
        RECT 114.670 68.090 114.900 69.465 ;
        RECT 119.310 69.350 119.540 69.465 ;
        RECT 119.310 68.715 119.545 69.350 ;
        RECT 121.065 68.715 121.305 69.920 ;
        RECT 119.310 68.090 119.540 68.715 ;
        RECT 121.075 68.615 121.305 68.715 ;
        RECT 121.515 73.600 121.745 73.615 ;
        RECT 122.165 73.600 122.645 74.435 ;
        RECT 121.515 68.675 122.655 73.600 ;
        RECT 121.515 68.615 121.745 68.675 ;
        RECT 121.265 68.405 121.555 68.410 ;
        RECT 121.250 68.150 121.580 68.405 ;
        RECT 114.670 66.745 119.540 68.090 ;
        RECT 114.670 65.505 114.900 66.745 ;
        RECT 119.310 65.505 119.540 66.745 ;
        RECT 110.585 65.340 112.585 65.365 ;
        RECT 115.105 65.340 119.105 65.455 ;
        RECT 110.585 65.265 112.590 65.340 ;
        RECT 113.125 65.265 119.105 65.340 ;
        RECT 110.585 65.225 119.105 65.265 ;
        RECT 110.585 65.135 119.040 65.225 ;
        RECT 110.640 65.000 119.040 65.135 ;
        RECT 109.000 64.290 110.860 64.730 ;
        RECT 109.000 64.280 111.850 64.290 ;
        RECT 109.000 63.935 112.520 64.280 ;
        RECT 109.000 62.310 110.860 63.935 ;
        RECT 111.660 63.785 112.520 63.935 ;
        RECT 111.155 63.595 111.405 63.610 ;
        RECT 111.155 63.305 111.430 63.595 ;
        RECT 111.590 63.555 112.590 63.785 ;
        RECT 113.010 63.690 113.280 65.000 ;
        RECT 123.880 64.570 124.580 74.435 ;
        RECT 118.300 64.235 124.580 64.570 ;
        RECT 115.185 64.095 124.580 64.235 ;
        RECT 115.185 63.870 119.045 64.095 ;
        RECT 111.155 63.275 111.405 63.305 ;
        RECT 111.590 63.115 112.590 63.345 ;
        RECT 112.735 63.270 114.925 63.690 ;
        RECT 115.120 63.640 119.120 63.870 ;
        RECT 119.355 63.680 119.605 63.700 ;
        RECT 115.120 63.200 119.120 63.430 ;
        RECT 119.325 63.390 119.605 63.680 ;
        RECT 119.355 63.365 119.605 63.390 ;
        RECT 111.660 62.975 112.545 63.115 ;
        RECT 115.170 63.035 119.095 63.200 ;
        RECT 112.730 62.975 119.095 63.035 ;
        RECT 111.660 62.920 119.095 62.975 ;
        RECT 111.660 62.850 115.540 62.920 ;
        RECT 112.215 62.735 115.540 62.850 ;
        RECT 123.880 62.770 124.580 64.095 ;
        RECT 109.000 62.265 111.385 62.310 ;
        RECT 93.665 60.560 98.730 60.630 ;
        RECT 95.205 60.555 98.730 60.560 ;
        RECT 46.080 60.000 80.415 60.235 ;
        RECT 96.415 60.000 97.415 60.555 ;
        RECT 109.000 60.535 109.875 62.265 ;
        RECT 110.240 61.990 111.385 62.265 ;
        RECT 113.570 62.105 113.975 62.735 ;
        RECT 122.575 62.235 124.580 62.770 ;
        RECT 110.240 61.925 112.490 61.990 ;
        RECT 110.680 61.760 112.490 61.925 ;
        RECT 110.165 61.570 110.415 61.595 ;
        RECT 110.165 61.280 110.435 61.570 ;
        RECT 110.595 61.530 112.595 61.760 ;
        RECT 113.555 61.740 113.980 62.105 ;
        RECT 115.220 62.090 124.580 62.235 ;
        RECT 115.220 61.845 123.075 62.090 ;
        RECT 110.165 61.260 110.415 61.280 ;
        RECT 110.595 61.090 112.595 61.320 ;
        RECT 112.745 61.230 114.935 61.740 ;
        RECT 115.125 61.615 123.125 61.845 ;
        RECT 123.355 61.655 123.605 61.670 ;
        RECT 112.745 61.225 113.445 61.230 ;
        RECT 114.445 61.225 114.935 61.230 ;
        RECT 115.125 61.175 123.125 61.405 ;
        RECT 123.330 61.365 123.605 61.655 ;
        RECT 123.355 61.335 123.605 61.365 ;
        RECT 110.665 60.925 112.530 61.090 ;
        RECT 113.415 60.925 114.415 61.000 ;
        RECT 115.200 60.925 123.050 61.175 ;
        RECT 110.665 60.630 123.050 60.925 ;
        RECT 123.880 60.690 124.580 62.090 ;
        RECT 126.000 86.860 132.605 87.120 ;
        RECT 126.000 86.665 132.800 86.860 ;
        RECT 126.000 86.530 139.975 86.665 ;
        RECT 126.000 86.425 127.010 86.530 ;
        RECT 132.015 86.435 139.975 86.530 ;
        RECT 126.000 86.085 126.875 86.425 ;
        RECT 126.000 85.860 126.885 86.085 ;
        RECT 127.595 86.000 128.815 86.085 ;
        RECT 127.595 85.945 128.830 86.000 ;
        RECT 126.000 81.185 126.875 85.860 ;
        RECT 127.585 85.715 129.585 85.945 ;
        RECT 127.195 84.465 127.425 85.665 ;
        RECT 127.970 84.465 129.135 85.715 ;
        RECT 129.745 84.465 129.975 85.665 ;
        RECT 127.195 83.675 129.975 84.465 ;
        RECT 131.735 85.510 131.965 86.230 ;
        RECT 131.735 85.485 132.100 85.510 ;
        RECT 132.260 85.485 132.580 85.540 ;
        RECT 131.735 85.335 132.580 85.485 ;
        RECT 131.735 85.305 132.100 85.335 ;
        RECT 131.735 84.230 131.965 85.305 ;
        RECT 132.260 85.280 132.580 85.335 ;
        RECT 134.865 84.055 136.680 86.435 ;
        RECT 140.025 86.195 140.255 86.230 ;
        RECT 140.880 86.195 141.580 87.165 ;
        RECT 141.760 87.130 144.875 87.320 ;
        RECT 157.900 87.165 158.600 87.285 ;
        RECT 140.025 84.285 141.580 86.195 ;
        RECT 140.025 84.230 140.255 84.285 ;
        RECT 132.265 84.025 139.895 84.055 ;
        RECT 132.015 83.795 139.975 84.025 ;
        RECT 127.195 81.705 127.425 83.675 ;
        RECT 129.745 83.005 129.975 83.675 ;
        RECT 129.745 82.725 132.610 83.005 ;
        RECT 129.745 82.635 140.030 82.725 ;
        RECT 129.745 81.705 129.975 82.635 ;
        RECT 132.170 82.485 140.030 82.635 ;
        RECT 132.110 82.255 140.110 82.485 ;
        RECT 131.675 81.765 131.905 82.205 ;
        RECT 140.315 82.195 140.545 82.205 ;
        RECT 132.395 81.765 133.395 81.835 ;
        RECT 140.315 81.765 140.550 82.195 ;
        RECT 127.585 81.425 129.585 81.655 ;
        RECT 127.675 81.185 129.500 81.425 ;
        RECT 126.000 80.695 129.500 81.185 ;
        RECT 126.000 75.860 126.875 80.695 ;
        RECT 127.675 80.515 129.500 80.695 ;
        RECT 131.675 80.875 140.550 81.765 ;
        RECT 127.585 80.285 129.585 80.515 ;
        RECT 131.675 80.245 131.905 80.875 ;
        RECT 132.395 80.820 133.395 80.875 ;
        RECT 140.315 80.310 140.550 80.875 ;
        RECT 140.315 80.245 140.545 80.310 ;
        RECT 127.195 78.800 127.425 80.235 ;
        RECT 129.745 78.800 129.975 80.235 ;
        RECT 132.110 79.965 140.110 80.195 ;
        RECT 132.180 79.840 140.010 79.965 ;
        RECT 132.200 79.055 140.000 79.840 ;
        RECT 132.110 78.825 140.110 79.055 ;
        RECT 127.195 77.460 129.975 78.800 ;
        RECT 131.675 78.750 131.905 78.775 ;
        RECT 127.195 76.275 127.425 77.460 ;
        RECT 127.770 76.225 129.365 77.460 ;
        RECT 129.745 76.570 129.975 77.460 ;
        RECT 131.670 78.305 131.905 78.750 ;
        RECT 140.315 78.750 140.545 78.775 ;
        RECT 131.670 78.295 132.085 78.305 ;
        RECT 132.225 78.295 133.225 78.365 ;
        RECT 131.670 78.290 133.225 78.295 ;
        RECT 133.635 78.290 135.255 78.295 ;
        RECT 140.315 78.290 140.550 78.750 ;
        RECT 131.670 77.400 140.550 78.290 ;
        RECT 131.670 77.385 133.225 77.400 ;
        RECT 133.635 77.395 135.255 77.400 ;
        RECT 131.670 77.295 132.085 77.385 ;
        RECT 132.225 77.335 133.225 77.385 ;
        RECT 131.670 76.865 131.905 77.295 ;
        RECT 131.675 76.815 131.905 76.865 ;
        RECT 140.315 76.865 140.550 77.400 ;
        RECT 140.315 76.815 140.545 76.865 ;
        RECT 132.110 76.570 140.110 76.765 ;
        RECT 129.745 76.535 140.110 76.570 ;
        RECT 129.745 76.390 140.030 76.535 ;
        RECT 129.745 76.375 132.245 76.390 ;
        RECT 129.745 76.275 129.975 76.375 ;
        RECT 127.585 75.995 129.585 76.225 ;
        RECT 140.880 76.115 141.580 84.285 ;
        RECT 135.955 75.985 136.230 76.055 ;
        RECT 130.260 75.860 136.230 75.985 ;
        RECT 126.000 75.845 127.405 75.860 ;
        RECT 129.750 75.845 136.230 75.860 ;
        RECT 126.000 75.795 136.230 75.845 ;
        RECT 126.000 75.670 130.450 75.795 ;
        RECT 135.955 75.720 136.230 75.795 ;
        RECT 126.000 70.390 126.875 75.670 ;
        RECT 128.825 75.365 132.610 75.370 ;
        RECT 128.825 75.300 136.060 75.365 ;
        RECT 127.645 75.175 136.060 75.300 ;
        RECT 127.645 75.085 136.105 75.175 ;
        RECT 127.585 75.075 136.105 75.085 ;
        RECT 127.585 74.855 129.585 75.075 ;
        RECT 132.105 74.945 136.105 75.075 ;
        RECT 127.195 73.425 127.425 74.805 ;
        RECT 129.745 73.425 129.975 74.805 ;
        RECT 127.195 72.470 129.975 73.425 ;
        RECT 127.195 70.845 127.425 72.470 ;
        RECT 129.745 70.845 129.975 72.470 ;
        RECT 131.670 73.640 131.900 74.895 ;
        RECT 133.340 73.640 134.725 74.945 ;
        RECT 136.310 73.640 136.540 74.895 ;
        RECT 136.905 74.435 141.580 76.115 ;
        RECT 138.265 74.095 138.540 74.125 ;
        RECT 138.250 73.840 138.580 74.095 ;
        RECT 138.265 73.820 138.555 73.840 ;
        RECT 138.265 73.790 138.540 73.820 ;
        RECT 131.670 73.570 136.540 73.640 ;
        RECT 138.075 73.570 138.305 73.615 ;
        RECT 131.670 72.295 136.545 73.570 ;
        RECT 131.670 70.935 131.900 72.295 ;
        RECT 136.310 70.935 136.545 72.295 ;
        RECT 127.585 70.565 129.585 70.795 ;
        RECT 127.650 70.390 129.520 70.565 ;
        RECT 126.000 69.835 129.520 70.390 ;
        RECT 126.000 64.730 126.875 69.835 ;
        RECT 127.650 69.655 129.520 69.835 ;
        RECT 127.585 69.425 129.585 69.655 ;
        RECT 131.710 69.465 131.870 70.935 ;
        RECT 136.340 70.925 136.545 70.935 ;
        RECT 132.105 70.655 136.105 70.885 ;
        RECT 132.185 70.410 136.010 70.655 ;
        RECT 138.065 70.410 138.305 73.570 ;
        RECT 132.185 69.920 138.305 70.410 ;
        RECT 132.185 69.745 136.010 69.920 ;
        RECT 132.105 69.515 136.105 69.745 ;
        RECT 127.195 67.980 127.425 69.375 ;
        RECT 129.745 67.980 129.975 69.375 ;
        RECT 127.195 67.025 129.975 67.980 ;
        RECT 127.195 65.415 127.425 67.025 ;
        RECT 129.745 65.415 129.975 67.025 ;
        RECT 131.670 68.090 131.900 69.465 ;
        RECT 136.310 69.350 136.540 69.465 ;
        RECT 136.310 68.715 136.545 69.350 ;
        RECT 138.065 68.715 138.305 69.920 ;
        RECT 136.310 68.090 136.540 68.715 ;
        RECT 138.075 68.615 138.305 68.715 ;
        RECT 138.515 73.600 138.745 73.615 ;
        RECT 139.165 73.600 139.645 74.435 ;
        RECT 138.515 68.675 139.655 73.600 ;
        RECT 138.515 68.615 138.745 68.675 ;
        RECT 138.265 68.405 138.555 68.410 ;
        RECT 138.250 68.150 138.580 68.405 ;
        RECT 131.670 66.745 136.540 68.090 ;
        RECT 131.670 65.505 131.900 66.745 ;
        RECT 136.310 65.505 136.540 66.745 ;
        RECT 127.585 65.340 129.585 65.365 ;
        RECT 132.105 65.340 136.105 65.455 ;
        RECT 127.585 65.265 129.590 65.340 ;
        RECT 130.125 65.265 136.105 65.340 ;
        RECT 127.585 65.225 136.105 65.265 ;
        RECT 127.585 65.135 136.040 65.225 ;
        RECT 127.640 65.000 136.040 65.135 ;
        RECT 126.000 64.290 127.860 64.730 ;
        RECT 126.000 64.280 128.850 64.290 ;
        RECT 126.000 63.935 129.520 64.280 ;
        RECT 126.000 62.310 127.860 63.935 ;
        RECT 128.660 63.785 129.520 63.935 ;
        RECT 128.155 63.595 128.405 63.610 ;
        RECT 128.155 63.305 128.430 63.595 ;
        RECT 128.590 63.555 129.590 63.785 ;
        RECT 130.010 63.690 130.280 65.000 ;
        RECT 140.880 64.570 141.580 74.435 ;
        RECT 135.300 64.235 141.580 64.570 ;
        RECT 132.185 64.095 141.580 64.235 ;
        RECT 132.185 63.870 136.045 64.095 ;
        RECT 128.155 63.275 128.405 63.305 ;
        RECT 128.590 63.115 129.590 63.345 ;
        RECT 129.735 63.270 131.925 63.690 ;
        RECT 132.120 63.640 136.120 63.870 ;
        RECT 136.355 63.680 136.605 63.700 ;
        RECT 132.120 63.200 136.120 63.430 ;
        RECT 136.325 63.390 136.605 63.680 ;
        RECT 136.355 63.365 136.605 63.390 ;
        RECT 128.660 62.975 129.545 63.115 ;
        RECT 132.170 63.035 136.095 63.200 ;
        RECT 129.730 62.975 136.095 63.035 ;
        RECT 128.660 62.920 136.095 62.975 ;
        RECT 128.660 62.850 132.540 62.920 ;
        RECT 129.215 62.735 132.540 62.850 ;
        RECT 140.880 62.770 141.580 64.095 ;
        RECT 126.000 62.265 128.385 62.310 ;
        RECT 110.665 60.560 115.730 60.630 ;
        RECT 112.205 60.555 115.730 60.560 ;
        RECT 113.415 60.000 114.415 60.555 ;
        RECT 126.000 60.535 126.875 62.265 ;
        RECT 127.240 61.990 128.385 62.265 ;
        RECT 130.570 62.105 130.975 62.735 ;
        RECT 139.575 62.235 141.580 62.770 ;
        RECT 127.240 61.925 129.490 61.990 ;
        RECT 127.680 61.760 129.490 61.925 ;
        RECT 127.165 61.570 127.415 61.595 ;
        RECT 127.165 61.280 127.435 61.570 ;
        RECT 127.595 61.530 129.595 61.760 ;
        RECT 130.555 61.740 130.980 62.105 ;
        RECT 132.220 62.090 141.580 62.235 ;
        RECT 132.220 61.845 140.075 62.090 ;
        RECT 127.165 61.260 127.415 61.280 ;
        RECT 127.595 61.090 129.595 61.320 ;
        RECT 129.745 61.230 131.935 61.740 ;
        RECT 132.125 61.615 140.125 61.845 ;
        RECT 140.355 61.655 140.605 61.670 ;
        RECT 129.745 61.225 130.445 61.230 ;
        RECT 131.445 61.225 131.935 61.230 ;
        RECT 132.125 61.175 140.125 61.405 ;
        RECT 140.330 61.365 140.605 61.655 ;
        RECT 140.355 61.335 140.605 61.365 ;
        RECT 127.665 60.925 129.530 61.090 ;
        RECT 130.415 60.925 131.415 61.000 ;
        RECT 132.200 60.925 140.050 61.175 ;
        RECT 127.665 60.630 140.050 60.925 ;
        RECT 140.880 60.690 141.580 62.090 ;
        RECT 143.000 87.025 144.875 87.130 ;
        RECT 143.000 86.665 149.445 87.025 ;
        RECT 157.880 86.800 158.600 87.165 ;
        RECT 143.000 86.530 156.975 86.665 ;
        RECT 143.000 86.085 143.875 86.530 ;
        RECT 144.120 86.400 144.875 86.530 ;
        RECT 149.015 86.435 156.975 86.530 ;
        RECT 143.000 85.860 143.885 86.085 ;
        RECT 144.595 86.000 145.815 86.085 ;
        RECT 144.595 85.945 145.830 86.000 ;
        RECT 143.000 81.185 143.875 85.860 ;
        RECT 144.585 85.715 146.585 85.945 ;
        RECT 144.195 84.465 144.425 85.665 ;
        RECT 144.970 84.465 146.135 85.715 ;
        RECT 146.745 84.465 146.975 85.665 ;
        RECT 144.195 83.675 146.975 84.465 ;
        RECT 148.735 85.510 148.965 86.230 ;
        RECT 148.735 85.485 149.100 85.510 ;
        RECT 149.260 85.485 149.580 85.540 ;
        RECT 148.735 85.335 149.580 85.485 ;
        RECT 148.735 85.305 149.100 85.335 ;
        RECT 148.735 84.230 148.965 85.305 ;
        RECT 149.260 85.280 149.580 85.335 ;
        RECT 151.865 84.055 153.680 86.435 ;
        RECT 157.025 86.195 157.255 86.230 ;
        RECT 157.880 86.195 158.580 86.800 ;
        RECT 157.025 84.285 158.580 86.195 ;
        RECT 157.025 84.230 157.255 84.285 ;
        RECT 149.265 84.025 156.895 84.055 ;
        RECT 149.015 83.795 156.975 84.025 ;
        RECT 144.195 81.705 144.425 83.675 ;
        RECT 146.745 83.005 146.975 83.675 ;
        RECT 146.745 82.725 149.610 83.005 ;
        RECT 146.745 82.635 157.030 82.725 ;
        RECT 146.745 81.705 146.975 82.635 ;
        RECT 149.170 82.485 157.030 82.635 ;
        RECT 149.110 82.255 157.110 82.485 ;
        RECT 148.675 81.765 148.905 82.205 ;
        RECT 157.315 82.195 157.545 82.205 ;
        RECT 149.395 81.765 150.395 81.835 ;
        RECT 157.315 81.765 157.550 82.195 ;
        RECT 144.585 81.425 146.585 81.655 ;
        RECT 144.675 81.185 146.500 81.425 ;
        RECT 143.000 80.695 146.500 81.185 ;
        RECT 143.000 75.860 143.875 80.695 ;
        RECT 144.675 80.515 146.500 80.695 ;
        RECT 148.675 80.875 157.550 81.765 ;
        RECT 144.585 80.285 146.585 80.515 ;
        RECT 148.675 80.245 148.905 80.875 ;
        RECT 149.395 80.820 150.395 80.875 ;
        RECT 157.315 80.310 157.550 80.875 ;
        RECT 157.315 80.245 157.545 80.310 ;
        RECT 144.195 78.800 144.425 80.235 ;
        RECT 146.745 78.800 146.975 80.235 ;
        RECT 149.110 79.965 157.110 80.195 ;
        RECT 149.180 79.840 157.010 79.965 ;
        RECT 149.200 79.055 157.000 79.840 ;
        RECT 149.110 78.825 157.110 79.055 ;
        RECT 144.195 77.460 146.975 78.800 ;
        RECT 148.675 78.750 148.905 78.775 ;
        RECT 144.195 76.275 144.425 77.460 ;
        RECT 144.770 76.225 146.365 77.460 ;
        RECT 146.745 76.570 146.975 77.460 ;
        RECT 148.670 78.305 148.905 78.750 ;
        RECT 157.315 78.750 157.545 78.775 ;
        RECT 148.670 78.295 149.085 78.305 ;
        RECT 149.225 78.295 150.225 78.365 ;
        RECT 148.670 78.290 150.225 78.295 ;
        RECT 150.635 78.290 152.255 78.295 ;
        RECT 157.315 78.290 157.550 78.750 ;
        RECT 148.670 77.400 157.550 78.290 ;
        RECT 148.670 77.385 150.225 77.400 ;
        RECT 150.635 77.395 152.255 77.400 ;
        RECT 148.670 77.295 149.085 77.385 ;
        RECT 149.225 77.335 150.225 77.385 ;
        RECT 148.670 76.865 148.905 77.295 ;
        RECT 148.675 76.815 148.905 76.865 ;
        RECT 157.315 76.865 157.550 77.400 ;
        RECT 157.315 76.815 157.545 76.865 ;
        RECT 149.110 76.570 157.110 76.765 ;
        RECT 146.745 76.535 157.110 76.570 ;
        RECT 146.745 76.390 157.030 76.535 ;
        RECT 146.745 76.375 149.245 76.390 ;
        RECT 146.745 76.275 146.975 76.375 ;
        RECT 144.585 75.995 146.585 76.225 ;
        RECT 157.880 76.115 158.580 84.285 ;
        RECT 152.955 75.985 153.230 76.055 ;
        RECT 147.260 75.860 153.230 75.985 ;
        RECT 143.000 75.845 144.405 75.860 ;
        RECT 146.750 75.845 153.230 75.860 ;
        RECT 143.000 75.795 153.230 75.845 ;
        RECT 143.000 75.670 147.450 75.795 ;
        RECT 152.955 75.720 153.230 75.795 ;
        RECT 143.000 70.390 143.875 75.670 ;
        RECT 145.825 75.365 149.610 75.370 ;
        RECT 145.825 75.300 153.060 75.365 ;
        RECT 144.645 75.175 153.060 75.300 ;
        RECT 144.645 75.085 153.105 75.175 ;
        RECT 144.585 75.075 153.105 75.085 ;
        RECT 144.585 74.855 146.585 75.075 ;
        RECT 149.105 74.945 153.105 75.075 ;
        RECT 144.195 73.425 144.425 74.805 ;
        RECT 146.745 73.425 146.975 74.805 ;
        RECT 144.195 72.470 146.975 73.425 ;
        RECT 144.195 70.845 144.425 72.470 ;
        RECT 146.745 70.845 146.975 72.470 ;
        RECT 148.670 73.640 148.900 74.895 ;
        RECT 150.340 73.640 151.725 74.945 ;
        RECT 153.310 73.640 153.540 74.895 ;
        RECT 153.905 74.435 158.580 76.115 ;
        RECT 155.265 74.095 155.540 74.125 ;
        RECT 155.250 73.840 155.580 74.095 ;
        RECT 155.265 73.820 155.555 73.840 ;
        RECT 155.265 73.790 155.540 73.820 ;
        RECT 148.670 73.570 153.540 73.640 ;
        RECT 155.075 73.570 155.305 73.615 ;
        RECT 148.670 72.295 153.545 73.570 ;
        RECT 148.670 70.935 148.900 72.295 ;
        RECT 153.310 70.935 153.545 72.295 ;
        RECT 144.585 70.565 146.585 70.795 ;
        RECT 144.650 70.390 146.520 70.565 ;
        RECT 143.000 69.835 146.520 70.390 ;
        RECT 143.000 64.730 143.875 69.835 ;
        RECT 144.650 69.655 146.520 69.835 ;
        RECT 144.585 69.425 146.585 69.655 ;
        RECT 148.710 69.465 148.870 70.935 ;
        RECT 153.340 70.925 153.545 70.935 ;
        RECT 149.105 70.655 153.105 70.885 ;
        RECT 149.185 70.410 153.010 70.655 ;
        RECT 155.065 70.410 155.305 73.570 ;
        RECT 149.185 69.920 155.305 70.410 ;
        RECT 149.185 69.745 153.010 69.920 ;
        RECT 149.105 69.515 153.105 69.745 ;
        RECT 144.195 67.980 144.425 69.375 ;
        RECT 146.745 67.980 146.975 69.375 ;
        RECT 144.195 67.025 146.975 67.980 ;
        RECT 144.195 65.415 144.425 67.025 ;
        RECT 146.745 65.415 146.975 67.025 ;
        RECT 148.670 68.090 148.900 69.465 ;
        RECT 153.310 69.350 153.540 69.465 ;
        RECT 153.310 68.715 153.545 69.350 ;
        RECT 155.065 68.715 155.305 69.920 ;
        RECT 153.310 68.090 153.540 68.715 ;
        RECT 155.075 68.615 155.305 68.715 ;
        RECT 155.515 73.600 155.745 73.615 ;
        RECT 156.165 73.600 156.645 74.435 ;
        RECT 155.515 68.675 156.655 73.600 ;
        RECT 155.515 68.615 155.745 68.675 ;
        RECT 155.265 68.405 155.555 68.410 ;
        RECT 155.250 68.150 155.580 68.405 ;
        RECT 148.670 66.745 153.540 68.090 ;
        RECT 148.670 65.505 148.900 66.745 ;
        RECT 153.310 65.505 153.540 66.745 ;
        RECT 144.585 65.340 146.585 65.365 ;
        RECT 149.105 65.340 153.105 65.455 ;
        RECT 144.585 65.265 146.590 65.340 ;
        RECT 147.125 65.265 153.105 65.340 ;
        RECT 144.585 65.225 153.105 65.265 ;
        RECT 144.585 65.135 153.040 65.225 ;
        RECT 144.640 65.000 153.040 65.135 ;
        RECT 143.000 64.290 144.860 64.730 ;
        RECT 143.000 64.280 145.850 64.290 ;
        RECT 143.000 63.935 146.520 64.280 ;
        RECT 143.000 62.310 144.860 63.935 ;
        RECT 145.660 63.785 146.520 63.935 ;
        RECT 145.155 63.595 145.405 63.610 ;
        RECT 145.155 63.305 145.430 63.595 ;
        RECT 145.590 63.555 146.590 63.785 ;
        RECT 147.010 63.690 147.280 65.000 ;
        RECT 157.880 64.570 158.580 74.435 ;
        RECT 152.300 64.235 158.580 64.570 ;
        RECT 149.185 64.095 158.580 64.235 ;
        RECT 149.185 63.870 153.045 64.095 ;
        RECT 145.155 63.275 145.405 63.305 ;
        RECT 145.590 63.115 146.590 63.345 ;
        RECT 146.735 63.270 148.925 63.690 ;
        RECT 149.120 63.640 153.120 63.870 ;
        RECT 153.355 63.680 153.605 63.700 ;
        RECT 149.120 63.200 153.120 63.430 ;
        RECT 153.325 63.390 153.605 63.680 ;
        RECT 153.355 63.365 153.605 63.390 ;
        RECT 145.660 62.975 146.545 63.115 ;
        RECT 149.170 63.035 153.095 63.200 ;
        RECT 146.730 62.975 153.095 63.035 ;
        RECT 145.660 62.920 153.095 62.975 ;
        RECT 145.660 62.850 149.540 62.920 ;
        RECT 146.215 62.735 149.540 62.850 ;
        RECT 157.880 62.770 158.580 64.095 ;
        RECT 143.000 62.265 145.385 62.310 ;
        RECT 127.665 60.560 132.730 60.630 ;
        RECT 129.205 60.555 132.730 60.560 ;
        RECT 130.415 60.000 131.415 60.555 ;
        RECT 143.000 60.535 143.875 62.265 ;
        RECT 144.240 61.990 145.385 62.265 ;
        RECT 147.570 62.105 147.975 62.735 ;
        RECT 156.575 62.235 158.580 62.770 ;
        RECT 144.240 61.925 146.490 61.990 ;
        RECT 144.680 61.760 146.490 61.925 ;
        RECT 144.165 61.570 144.415 61.595 ;
        RECT 144.165 61.280 144.435 61.570 ;
        RECT 144.595 61.530 146.595 61.760 ;
        RECT 147.555 61.740 147.980 62.105 ;
        RECT 149.220 62.090 158.580 62.235 ;
        RECT 149.220 61.845 157.075 62.090 ;
        RECT 144.165 61.260 144.415 61.280 ;
        RECT 144.595 61.090 146.595 61.320 ;
        RECT 146.745 61.230 148.935 61.740 ;
        RECT 149.125 61.615 157.125 61.845 ;
        RECT 157.355 61.655 157.605 61.670 ;
        RECT 146.745 61.225 147.445 61.230 ;
        RECT 148.445 61.225 148.935 61.230 ;
        RECT 149.125 61.175 157.125 61.405 ;
        RECT 157.330 61.365 157.605 61.655 ;
        RECT 157.355 61.335 157.605 61.365 ;
        RECT 144.665 60.925 146.530 61.090 ;
        RECT 147.415 60.925 148.415 61.000 ;
        RECT 149.200 60.925 157.050 61.175 ;
        RECT 144.665 60.630 157.050 60.925 ;
        RECT 157.880 60.690 158.580 62.090 ;
        RECT 144.665 60.560 149.730 60.630 ;
        RECT 146.205 60.555 149.730 60.560 ;
        RECT 147.415 60.000 148.415 60.555 ;
        RECT 46.080 59.985 80.040 60.000 ;
        RECT 46.080 59.980 46.400 59.985 ;
        RECT 60.715 59.625 61.035 59.655 ;
        RECT 96.815 59.625 97.020 60.000 ;
        RECT 22.520 59.000 58.400 59.480 ;
        RECT 60.095 59.235 60.355 59.470 ;
        RECT 60.715 59.420 97.020 59.625 ;
        RECT 60.715 59.395 61.035 59.420 ;
        RECT 113.845 59.235 113.990 60.000 ;
        RECT 60.095 59.150 113.990 59.235 ;
        RECT 60.150 59.090 113.990 59.150 ;
        RECT 59.330 58.900 59.650 58.930 ;
        RECT 130.815 58.900 131.015 60.000 ;
        RECT 31.345 58.800 31.635 58.845 ;
        RECT 36.390 58.800 36.710 58.860 ;
        RECT 31.345 58.660 36.710 58.800 ;
        RECT 31.345 58.615 31.635 58.660 ;
        RECT 36.390 58.600 36.710 58.660 ;
        RECT 41.925 58.800 42.215 58.845 ;
        RECT 42.830 58.800 43.150 58.860 ;
        RECT 41.925 58.660 43.150 58.800 ;
        RECT 41.925 58.615 42.215 58.660 ;
        RECT 42.830 58.600 43.150 58.660 ;
        RECT 49.270 58.800 49.590 58.860 ;
        RECT 50.205 58.800 50.495 58.845 ;
        RECT 49.270 58.660 50.495 58.800 ;
        RECT 59.330 58.700 131.015 58.900 ;
        RECT 59.330 58.670 59.650 58.700 ;
        RECT 49.270 58.600 49.590 58.660 ;
        RECT 50.205 58.615 50.495 58.660 ;
        RECT 58.665 58.530 58.985 58.565 ;
        RECT 147.820 58.530 148.015 60.000 ;
        RECT 33.645 58.460 33.935 58.505 ;
        RECT 40.990 58.460 41.310 58.520 ;
        RECT 47.890 58.460 48.210 58.520 ;
        RECT 33.645 58.320 41.310 58.460 ;
        RECT 33.645 58.275 33.935 58.320 ;
        RECT 40.990 58.260 41.310 58.320 ;
        RECT 42.460 58.320 48.210 58.460 ;
        RECT 36.865 58.120 37.155 58.165 ;
        RECT 30.500 57.980 37.155 58.120 ;
        RECT 28.110 57.780 28.430 57.840 ;
        RECT 30.500 57.825 30.640 57.980 ;
        RECT 36.865 57.935 37.155 57.980 ;
        RECT 30.425 57.780 30.715 57.825 ;
        RECT 28.110 57.640 30.715 57.780 ;
        RECT 28.110 57.580 28.430 57.640 ;
        RECT 30.425 57.595 30.715 57.640 ;
        RECT 32.710 57.580 33.030 57.840 ;
        RECT 33.170 57.580 33.490 57.840 ;
        RECT 34.105 57.780 34.395 57.825 ;
        RECT 42.460 57.780 42.600 58.320 ;
        RECT 47.890 58.260 48.210 58.320 ;
        RECT 58.665 58.335 148.015 58.530 ;
        RECT 58.665 58.305 58.985 58.335 ;
        RECT 75.000 58.025 75.875 58.140 ;
        RECT 34.105 57.640 42.600 57.780 ;
        RECT 42.845 57.780 43.135 57.825 ;
        RECT 43.290 57.780 43.610 57.840 ;
        RECT 42.845 57.640 43.610 57.780 ;
        RECT 34.105 57.595 34.395 57.640 ;
        RECT 42.845 57.595 43.135 57.640 ;
        RECT 43.290 57.580 43.610 57.640 ;
        RECT 46.050 57.780 46.370 57.840 ;
        RECT 46.985 57.780 47.275 57.825 ;
        RECT 46.050 57.640 47.275 57.780 ;
        RECT 46.050 57.580 46.370 57.640 ;
        RECT 46.985 57.595 47.275 57.640 ;
        RECT 51.110 57.580 51.430 57.840 ;
        RECT 53.870 57.580 54.190 57.840 ;
        RECT 55.250 57.580 55.570 57.840 ;
        RECT 56.630 57.580 56.950 57.840 ;
        RECT 75.000 57.665 81.445 58.025 ;
        RECT 75.000 57.530 88.975 57.665 ;
        RECT 35.010 56.900 35.330 57.160 ;
        RECT 40.070 56.900 40.390 57.160 ;
        RECT 43.750 57.100 44.070 57.160 ;
        RECT 46.525 57.100 46.815 57.145 ;
        RECT 43.750 56.960 46.815 57.100 ;
        RECT 43.750 56.900 44.070 56.960 ;
        RECT 46.525 56.915 46.815 56.960 ;
        RECT 49.730 57.100 50.050 57.160 ;
        RECT 52.965 57.100 53.255 57.145 ;
        RECT 49.730 56.960 53.255 57.100 ;
        RECT 49.730 56.900 50.050 56.960 ;
        RECT 52.965 56.915 53.255 56.960 ;
        RECT 53.410 57.100 53.730 57.160 ;
        RECT 54.345 57.100 54.635 57.145 ;
        RECT 53.410 56.960 54.635 57.100 ;
        RECT 53.410 56.900 53.730 56.960 ;
        RECT 54.345 56.915 54.635 56.960 ;
        RECT 55.725 57.100 56.015 57.145 ;
        RECT 56.170 57.100 56.490 57.160 ;
        RECT 55.725 56.960 56.490 57.100 ;
        RECT 55.725 56.915 56.015 56.960 ;
        RECT 56.170 56.900 56.490 56.960 ;
        RECT 75.000 57.085 75.875 57.530 ;
        RECT 81.015 57.435 88.975 57.530 ;
        RECT 75.000 56.860 75.885 57.085 ;
        RECT 76.595 57.000 77.815 57.085 ;
        RECT 76.595 56.945 77.830 57.000 ;
        RECT 22.520 56.280 58.400 56.760 ;
        RECT 28.110 55.880 28.430 56.140 ;
        RECT 32.710 56.080 33.030 56.140 ;
        RECT 42.385 56.080 42.675 56.125 ;
        RECT 43.290 56.080 43.610 56.140 ;
        RECT 32.710 55.940 38.000 56.080 ;
        RECT 32.710 55.880 33.030 55.940 ;
        RECT 35.010 55.740 35.330 55.800 ;
        RECT 36.710 55.740 37.000 55.785 ;
        RECT 35.010 55.600 37.000 55.740 ;
        RECT 37.860 55.740 38.000 55.940 ;
        RECT 42.385 55.940 43.610 56.080 ;
        RECT 42.385 55.895 42.675 55.940 ;
        RECT 43.290 55.880 43.610 55.940 ;
        RECT 42.845 55.740 43.135 55.785 ;
        RECT 37.860 55.600 43.135 55.740 ;
        RECT 35.010 55.540 35.330 55.600 ;
        RECT 36.710 55.555 37.000 55.600 ;
        RECT 42.845 55.555 43.135 55.600 ;
        RECT 43.750 55.540 44.070 55.800 ;
        RECT 33.745 55.400 34.035 55.445 ;
        RECT 35.930 55.400 36.250 55.460 ;
        RECT 33.745 55.260 36.250 55.400 ;
        RECT 33.745 55.215 34.035 55.260 ;
        RECT 35.930 55.200 36.250 55.260 ;
        RECT 44.670 55.200 44.990 55.460 ;
        RECT 45.145 55.215 45.435 55.445 ;
        RECT 46.050 55.400 46.370 55.460 ;
        RECT 46.985 55.400 47.275 55.445 ;
        RECT 46.050 55.260 47.275 55.400 ;
        RECT 30.435 55.060 30.725 55.105 ;
        RECT 32.955 55.060 33.245 55.105 ;
        RECT 34.145 55.060 34.435 55.105 ;
        RECT 30.435 54.920 34.435 55.060 ;
        RECT 30.435 54.875 30.725 54.920 ;
        RECT 32.955 54.875 33.245 54.920 ;
        RECT 34.145 54.875 34.435 54.920 ;
        RECT 35.025 55.060 35.315 55.105 ;
        RECT 35.485 55.060 35.775 55.105 ;
        RECT 35.025 54.920 35.775 55.060 ;
        RECT 35.025 54.875 35.315 54.920 ;
        RECT 35.485 54.875 35.775 54.920 ;
        RECT 36.365 55.060 36.655 55.105 ;
        RECT 37.555 55.060 37.845 55.105 ;
        RECT 40.075 55.060 40.365 55.105 ;
        RECT 36.365 54.920 40.365 55.060 ;
        RECT 36.365 54.875 36.655 54.920 ;
        RECT 37.555 54.875 37.845 54.920 ;
        RECT 40.075 54.875 40.365 54.920 ;
        RECT 41.450 55.060 41.770 55.120 ;
        RECT 45.220 55.060 45.360 55.215 ;
        RECT 46.050 55.200 46.370 55.260 ;
        RECT 46.985 55.215 47.275 55.260 ;
        RECT 47.890 55.400 48.210 55.460 ;
        RECT 49.745 55.400 50.035 55.445 ;
        RECT 47.890 55.260 50.035 55.400 ;
        RECT 47.890 55.200 48.210 55.260 ;
        RECT 49.745 55.215 50.035 55.260 ;
        RECT 50.650 55.200 50.970 55.460 ;
        RECT 51.125 55.400 51.415 55.445 ;
        RECT 53.870 55.400 54.190 55.460 ;
        RECT 51.125 55.260 54.190 55.400 ;
        RECT 51.125 55.215 51.415 55.260 ;
        RECT 53.870 55.200 54.190 55.260 ;
        RECT 56.630 55.200 56.950 55.460 ;
        RECT 41.450 54.920 45.360 55.060 ;
        RECT 45.590 55.060 45.910 55.120 ;
        RECT 47.980 55.060 48.120 55.200 ;
        RECT 45.590 54.920 48.120 55.060 ;
        RECT 30.870 54.720 31.160 54.765 ;
        RECT 32.440 54.720 32.730 54.765 ;
        RECT 34.540 54.720 34.830 54.765 ;
        RECT 30.870 54.580 34.830 54.720 ;
        RECT 30.870 54.535 31.160 54.580 ;
        RECT 32.440 54.535 32.730 54.580 ;
        RECT 34.540 54.535 34.830 54.580 ;
        RECT 33.630 54.380 33.950 54.440 ;
        RECT 35.560 54.380 35.700 54.875 ;
        RECT 41.450 54.860 41.770 54.920 ;
        RECT 45.590 54.860 45.910 54.920 ;
        RECT 52.045 54.875 52.335 55.105 ;
        RECT 35.970 54.720 36.260 54.765 ;
        RECT 38.070 54.720 38.360 54.765 ;
        RECT 39.640 54.720 39.930 54.765 ;
        RECT 35.970 54.580 39.930 54.720 ;
        RECT 35.970 54.535 36.260 54.580 ;
        RECT 38.070 54.535 38.360 54.580 ;
        RECT 39.640 54.535 39.930 54.580 ;
        RECT 40.530 54.720 40.850 54.780 ;
        RECT 46.065 54.720 46.355 54.765 ;
        RECT 40.530 54.580 46.355 54.720 ;
        RECT 40.530 54.520 40.850 54.580 ;
        RECT 46.065 54.535 46.355 54.580 ;
        RECT 47.445 54.720 47.735 54.765 ;
        RECT 50.205 54.720 50.495 54.765 ;
        RECT 47.445 54.580 50.495 54.720 ;
        RECT 47.445 54.535 47.735 54.580 ;
        RECT 50.205 54.535 50.495 54.580 ;
        RECT 51.110 54.720 51.430 54.780 ;
        RECT 52.120 54.720 52.260 54.875 ;
        RECT 51.110 54.580 52.260 54.720 ;
        RECT 54.330 54.720 54.650 54.780 ;
        RECT 55.725 54.720 56.015 54.765 ;
        RECT 54.330 54.580 56.015 54.720 ;
        RECT 51.110 54.520 51.430 54.580 ;
        RECT 54.330 54.520 54.650 54.580 ;
        RECT 55.725 54.535 56.015 54.580 ;
        RECT 44.210 54.380 44.530 54.440 ;
        RECT 33.630 54.240 44.530 54.380 ;
        RECT 33.630 54.180 33.950 54.240 ;
        RECT 44.210 54.180 44.530 54.240 ;
        RECT 46.970 54.380 47.290 54.440 ;
        RECT 48.825 54.380 49.115 54.425 ;
        RECT 46.970 54.240 49.115 54.380 ;
        RECT 46.970 54.180 47.290 54.240 ;
        RECT 48.825 54.195 49.115 54.240 ;
        RECT 52.950 54.380 53.270 54.440 ;
        RECT 55.265 54.380 55.555 54.425 ;
        RECT 52.950 54.240 55.555 54.380 ;
        RECT 52.950 54.180 53.270 54.240 ;
        RECT 55.265 54.195 55.555 54.240 ;
        RECT 22.520 53.560 58.400 54.040 ;
        RECT 35.930 53.160 36.250 53.420 ;
        RECT 40.990 53.360 41.310 53.420 ;
        RECT 43.305 53.360 43.595 53.405 ;
        RECT 46.050 53.360 46.370 53.420 ;
        RECT 40.990 53.220 43.595 53.360 ;
        RECT 40.990 53.160 41.310 53.220 ;
        RECT 43.305 53.175 43.595 53.220 ;
        RECT 44.300 53.220 49.500 53.360 ;
        RECT 24.470 53.020 24.760 53.065 ;
        RECT 26.570 53.020 26.860 53.065 ;
        RECT 28.140 53.020 28.430 53.065 ;
        RECT 44.300 53.020 44.440 53.220 ;
        RECT 46.050 53.160 46.370 53.220 ;
        RECT 24.470 52.880 28.430 53.020 ;
        RECT 24.470 52.835 24.760 52.880 ;
        RECT 26.570 52.835 26.860 52.880 ;
        RECT 28.140 52.835 28.430 52.880 ;
        RECT 39.240 52.880 44.440 53.020 ;
        RECT 44.710 53.020 45.000 53.065 ;
        RECT 46.810 53.020 47.100 53.065 ;
        RECT 48.380 53.020 48.670 53.065 ;
        RECT 44.710 52.880 48.670 53.020 ;
        RECT 39.240 52.725 39.380 52.880 ;
        RECT 44.710 52.835 45.000 52.880 ;
        RECT 46.810 52.835 47.100 52.880 ;
        RECT 48.380 52.835 48.670 52.880 ;
        RECT 24.865 52.680 25.155 52.725 ;
        RECT 26.055 52.680 26.345 52.725 ;
        RECT 28.575 52.680 28.865 52.725 ;
        RECT 24.865 52.540 28.865 52.680 ;
        RECT 24.865 52.495 25.155 52.540 ;
        RECT 26.055 52.495 26.345 52.540 ;
        RECT 28.575 52.495 28.865 52.540 ;
        RECT 39.165 52.495 39.455 52.725 ;
        RECT 44.210 52.480 44.530 52.740 ;
        RECT 45.105 52.680 45.395 52.725 ;
        RECT 46.295 52.680 46.585 52.725 ;
        RECT 48.815 52.680 49.105 52.725 ;
        RECT 45.105 52.540 49.105 52.680 ;
        RECT 45.105 52.495 45.395 52.540 ;
        RECT 46.295 52.495 46.585 52.540 ;
        RECT 48.815 52.495 49.105 52.540 ;
        RECT 23.985 52.340 24.275 52.385 ;
        RECT 33.630 52.340 33.950 52.400 ;
        RECT 23.985 52.200 33.950 52.340 ;
        RECT 23.985 52.155 24.275 52.200 ;
        RECT 33.630 52.140 33.950 52.200 ;
        RECT 34.105 52.155 34.395 52.385 ;
        RECT 37.785 52.340 38.075 52.385 ;
        RECT 40.070 52.340 40.390 52.400 ;
        RECT 37.785 52.200 40.390 52.340 ;
        RECT 37.785 52.155 38.075 52.200 ;
        RECT 25.320 52.000 25.610 52.045 ;
        RECT 25.810 52.000 26.130 52.060 ;
        RECT 34.180 52.000 34.320 52.155 ;
        RECT 40.070 52.140 40.390 52.200 ;
        RECT 40.530 52.140 40.850 52.400 ;
        RECT 41.450 52.340 41.770 52.400 ;
        RECT 43.290 52.340 43.610 52.400 ;
        RECT 41.450 52.200 43.610 52.340 ;
        RECT 41.450 52.140 41.770 52.200 ;
        RECT 43.290 52.140 43.610 52.200 ;
        RECT 43.750 52.340 44.070 52.400 ;
        RECT 44.670 52.340 44.990 52.400 ;
        RECT 43.750 52.200 44.990 52.340 ;
        RECT 43.750 52.140 44.070 52.200 ;
        RECT 44.670 52.140 44.990 52.200 ;
        RECT 45.560 52.340 45.850 52.385 ;
        RECT 46.970 52.340 47.290 52.400 ;
        RECT 45.560 52.200 47.290 52.340 ;
        RECT 49.360 52.340 49.500 53.220 ;
        RECT 51.110 53.160 51.430 53.420 ;
        RECT 53.870 53.160 54.190 53.420 ;
        RECT 52.045 52.340 52.335 52.385 ;
        RECT 49.360 52.200 52.335 52.340 ;
        RECT 45.560 52.155 45.850 52.200 ;
        RECT 46.970 52.140 47.290 52.200 ;
        RECT 52.045 52.155 52.335 52.200 ;
        RECT 52.950 52.140 53.270 52.400 ;
        RECT 54.330 52.140 54.650 52.400 ;
        RECT 56.630 52.140 56.950 52.400 ;
        RECT 75.000 52.185 75.875 56.860 ;
        RECT 76.585 56.715 78.585 56.945 ;
        RECT 76.195 55.465 76.425 56.665 ;
        RECT 76.970 55.465 78.135 56.715 ;
        RECT 78.745 55.465 78.975 56.665 ;
        RECT 76.195 54.675 78.975 55.465 ;
        RECT 80.735 56.510 80.965 57.230 ;
        RECT 80.735 56.485 81.100 56.510 ;
        RECT 81.260 56.485 81.580 56.540 ;
        RECT 80.735 56.335 81.580 56.485 ;
        RECT 80.735 56.305 81.100 56.335 ;
        RECT 80.735 55.230 80.965 56.305 ;
        RECT 81.260 56.280 81.580 56.335 ;
        RECT 83.865 55.055 85.680 57.435 ;
        RECT 89.025 57.195 89.255 57.230 ;
        RECT 89.880 57.195 90.580 58.165 ;
        RECT 89.025 55.285 90.580 57.195 ;
        RECT 89.025 55.230 89.255 55.285 ;
        RECT 81.265 55.025 88.895 55.055 ;
        RECT 81.015 54.795 88.975 55.025 ;
        RECT 76.195 52.705 76.425 54.675 ;
        RECT 78.745 54.005 78.975 54.675 ;
        RECT 78.745 53.725 81.610 54.005 ;
        RECT 78.745 53.635 89.030 53.725 ;
        RECT 78.745 52.705 78.975 53.635 ;
        RECT 81.170 53.485 89.030 53.635 ;
        RECT 81.110 53.255 89.110 53.485 ;
        RECT 80.675 52.765 80.905 53.205 ;
        RECT 89.315 53.195 89.545 53.205 ;
        RECT 81.395 52.765 82.395 52.835 ;
        RECT 89.315 52.765 89.550 53.195 ;
        RECT 76.585 52.425 78.585 52.655 ;
        RECT 76.675 52.185 78.500 52.425 ;
        RECT 25.320 51.860 26.130 52.000 ;
        RECT 25.320 51.815 25.610 51.860 ;
        RECT 25.810 51.800 26.130 51.860 ;
        RECT 30.960 51.860 34.320 52.000 ;
        RECT 38.245 52.000 38.535 52.045 ;
        RECT 46.050 52.000 46.370 52.060 ;
        RECT 38.245 51.860 46.370 52.000 ;
        RECT 30.960 51.720 31.100 51.860 ;
        RECT 38.245 51.815 38.535 51.860 ;
        RECT 46.050 51.800 46.370 51.860 ;
        RECT 30.870 51.460 31.190 51.720 ;
        RECT 31.330 51.460 31.650 51.720 ;
        RECT 40.070 51.660 40.390 51.720 ;
        RECT 42.385 51.660 42.675 51.705 ;
        RECT 40.070 51.520 42.675 51.660 ;
        RECT 40.070 51.460 40.390 51.520 ;
        RECT 42.385 51.475 42.675 51.520 ;
        RECT 55.250 51.460 55.570 51.720 ;
        RECT 55.710 51.460 56.030 51.720 ;
        RECT 75.000 51.695 78.500 52.185 ;
        RECT 22.520 50.840 58.400 51.320 ;
        RECT 23.510 50.640 23.830 50.700 ;
        RECT 24.445 50.640 24.735 50.685 ;
        RECT 23.510 50.500 24.735 50.640 ;
        RECT 23.510 50.440 23.830 50.500 ;
        RECT 24.445 50.455 24.735 50.500 ;
        RECT 25.810 50.440 26.130 50.700 ;
        RECT 27.665 50.640 27.955 50.685 ;
        RECT 31.330 50.640 31.650 50.700 ;
        RECT 27.665 50.500 31.650 50.640 ;
        RECT 27.665 50.455 27.955 50.500 ;
        RECT 31.330 50.440 31.650 50.500 ;
        RECT 33.630 50.640 33.950 50.700 ;
        RECT 35.930 50.640 36.250 50.700 ;
        RECT 33.630 50.500 36.250 50.640 ;
        RECT 33.630 50.440 33.950 50.500 ;
        RECT 35.930 50.440 36.250 50.500 ;
        RECT 36.850 50.640 37.170 50.700 ;
        RECT 40.530 50.640 40.850 50.700 ;
        RECT 53.410 50.640 53.730 50.700 ;
        RECT 36.850 50.500 40.850 50.640 ;
        RECT 36.850 50.440 37.170 50.500 ;
        RECT 40.530 50.440 40.850 50.500 ;
        RECT 47.060 50.500 53.730 50.640 ;
        RECT 45.590 50.100 45.910 50.360 ;
        RECT 25.365 49.960 25.655 50.005 ;
        RECT 30.870 49.960 31.190 50.020 ;
        RECT 25.365 49.820 31.190 49.960 ;
        RECT 25.365 49.775 25.655 49.820 ;
        RECT 30.870 49.760 31.190 49.820 ;
        RECT 40.085 49.960 40.375 50.005 ;
        RECT 40.530 49.960 40.850 50.020 ;
        RECT 47.060 50.005 47.200 50.500 ;
        RECT 53.410 50.440 53.730 50.500 ;
        RECT 55.710 50.440 56.030 50.700 ;
        RECT 48.825 50.300 49.115 50.345 ;
        RECT 50.190 50.300 50.510 50.360 ;
        RECT 48.825 50.160 50.510 50.300 ;
        RECT 48.825 50.115 49.115 50.160 ;
        RECT 50.190 50.100 50.510 50.160 ;
        RECT 50.650 50.300 50.970 50.360 ;
        RECT 55.800 50.300 55.940 50.440 ;
        RECT 50.650 50.160 55.940 50.300 ;
        RECT 50.650 50.100 50.970 50.160 ;
        RECT 40.085 49.820 40.850 49.960 ;
        RECT 40.085 49.775 40.375 49.820 ;
        RECT 40.530 49.760 40.850 49.820 ;
        RECT 46.985 49.775 47.275 50.005 ;
        RECT 49.730 49.760 50.050 50.020 ;
        RECT 52.120 50.005 52.260 50.160 ;
        RECT 51.125 49.775 51.415 50.005 ;
        RECT 52.045 49.775 52.335 50.005 ;
        RECT 28.125 49.435 28.415 49.665 ;
        RECT 29.045 49.620 29.335 49.665 ;
        RECT 29.490 49.620 29.810 49.680 ;
        RECT 29.045 49.480 29.810 49.620 ;
        RECT 29.045 49.435 29.335 49.480 ;
        RECT 26.270 49.280 26.590 49.340 ;
        RECT 28.200 49.280 28.340 49.435 ;
        RECT 29.490 49.420 29.810 49.480 ;
        RECT 43.765 49.620 44.055 49.665 ;
        RECT 44.210 49.620 44.530 49.680 ;
        RECT 43.765 49.480 44.530 49.620 ;
        RECT 43.765 49.435 44.055 49.480 ;
        RECT 44.210 49.420 44.530 49.480 ;
        RECT 46.525 49.620 46.815 49.665 ;
        RECT 49.820 49.620 49.960 49.760 ;
        RECT 46.525 49.480 49.960 49.620 ;
        RECT 51.200 49.620 51.340 49.775 ;
        RECT 53.410 49.760 53.730 50.020 ;
        RECT 54.790 49.760 55.110 50.020 ;
        RECT 55.725 49.960 56.015 50.005 ;
        RECT 56.170 49.960 56.490 50.020 ;
        RECT 55.725 49.820 56.490 49.960 ;
        RECT 55.725 49.775 56.015 49.820 ;
        RECT 56.170 49.760 56.490 49.820 ;
        RECT 52.505 49.620 52.795 49.665 ;
        RECT 51.200 49.480 52.795 49.620 ;
        RECT 46.525 49.435 46.815 49.480 ;
        RECT 52.505 49.435 52.795 49.480 ;
        RECT 46.050 49.280 46.370 49.340 ;
        RECT 50.650 49.280 50.970 49.340 ;
        RECT 26.270 49.140 46.370 49.280 ;
        RECT 26.270 49.080 26.590 49.140 ;
        RECT 46.050 49.080 46.370 49.140 ;
        RECT 47.060 49.140 50.970 49.280 ;
        RECT 40.545 48.940 40.835 48.985 ;
        RECT 40.990 48.940 41.310 49.000 ;
        RECT 47.060 48.985 47.200 49.140 ;
        RECT 50.650 49.080 50.970 49.140 ;
        RECT 40.545 48.800 41.310 48.940 ;
        RECT 40.545 48.755 40.835 48.800 ;
        RECT 40.990 48.740 41.310 48.800 ;
        RECT 46.985 48.755 47.275 48.985 ;
        RECT 47.890 48.740 48.210 49.000 ;
        RECT 22.520 48.120 58.400 48.600 ;
        RECT 36.850 47.920 37.170 47.980 ;
        RECT 28.200 47.780 37.170 47.920 ;
        RECT 26.270 47.040 26.590 47.300 ;
        RECT 27.205 47.240 27.495 47.285 ;
        RECT 28.200 47.240 28.340 47.780 ;
        RECT 36.850 47.720 37.170 47.780 ;
        RECT 42.845 47.920 43.135 47.965 ;
        RECT 43.290 47.920 43.610 47.980 ;
        RECT 42.845 47.780 43.610 47.920 ;
        RECT 42.845 47.735 43.135 47.780 ;
        RECT 43.290 47.720 43.610 47.780 ;
        RECT 52.965 47.920 53.255 47.965 ;
        RECT 54.790 47.920 55.110 47.980 ;
        RECT 52.965 47.780 55.110 47.920 ;
        RECT 52.965 47.735 53.255 47.780 ;
        RECT 54.790 47.720 55.110 47.780 ;
        RECT 28.610 47.580 28.900 47.625 ;
        RECT 30.710 47.580 31.000 47.625 ;
        RECT 32.280 47.580 32.570 47.625 ;
        RECT 28.610 47.440 32.570 47.580 ;
        RECT 28.610 47.395 28.900 47.440 ;
        RECT 30.710 47.395 31.000 47.440 ;
        RECT 32.280 47.395 32.570 47.440 ;
        RECT 35.025 47.395 35.315 47.625 ;
        RECT 36.430 47.580 36.720 47.625 ;
        RECT 38.530 47.580 38.820 47.625 ;
        RECT 40.100 47.580 40.390 47.625 ;
        RECT 36.430 47.440 40.390 47.580 ;
        RECT 36.430 47.395 36.720 47.440 ;
        RECT 38.530 47.395 38.820 47.440 ;
        RECT 40.100 47.395 40.390 47.440 ;
        RECT 27.205 47.100 28.340 47.240 ;
        RECT 29.005 47.240 29.295 47.285 ;
        RECT 30.195 47.240 30.485 47.285 ;
        RECT 32.715 47.240 33.005 47.285 ;
        RECT 29.005 47.100 33.005 47.240 ;
        RECT 27.205 47.055 27.495 47.100 ;
        RECT 29.005 47.055 29.295 47.100 ;
        RECT 30.195 47.055 30.485 47.100 ;
        RECT 32.715 47.055 33.005 47.100 ;
        RECT 28.125 46.900 28.415 46.945 ;
        RECT 30.870 46.900 31.190 46.960 ;
        RECT 33.630 46.900 33.950 46.960 ;
        RECT 28.125 46.760 33.950 46.900 ;
        RECT 35.100 46.900 35.240 47.395 ;
        RECT 44.670 47.380 44.990 47.640 ;
        RECT 51.570 47.580 51.890 47.640 ;
        RECT 56.170 47.580 56.490 47.640 ;
        RECT 49.360 47.440 56.490 47.580 ;
        RECT 35.930 47.040 36.250 47.300 ;
        RECT 49.360 47.285 49.500 47.440 ;
        RECT 51.570 47.380 51.890 47.440 ;
        RECT 56.170 47.380 56.490 47.440 ;
        RECT 36.825 47.240 37.115 47.285 ;
        RECT 38.015 47.240 38.305 47.285 ;
        RECT 40.535 47.240 40.825 47.285 ;
        RECT 36.825 47.100 40.825 47.240 ;
        RECT 36.825 47.055 37.115 47.100 ;
        RECT 38.015 47.055 38.305 47.100 ;
        RECT 40.535 47.055 40.825 47.100 ;
        RECT 49.285 47.055 49.575 47.285 ;
        RECT 49.745 47.240 50.035 47.285 ;
        RECT 52.490 47.240 52.810 47.300 ;
        RECT 49.745 47.100 52.810 47.240 ;
        RECT 49.745 47.055 50.035 47.100 ;
        RECT 52.490 47.040 52.810 47.100 ;
        RECT 44.210 46.900 44.530 46.960 ;
        RECT 35.100 46.760 45.360 46.900 ;
        RECT 28.125 46.715 28.415 46.760 ;
        RECT 30.870 46.700 31.190 46.760 ;
        RECT 33.630 46.700 33.950 46.760 ;
        RECT 44.210 46.700 44.530 46.760 ;
        RECT 45.220 46.620 45.360 46.760 ;
        RECT 48.825 46.715 49.115 46.945 ;
        RECT 50.205 46.715 50.495 46.945 ;
        RECT 50.650 46.900 50.970 46.960 ;
        RECT 51.125 46.900 51.415 46.945 ;
        RECT 50.650 46.760 51.415 46.900 ;
        RECT 29.490 46.605 29.810 46.620 ;
        RECT 29.460 46.560 29.810 46.605 ;
        RECT 37.280 46.560 37.570 46.605 ;
        RECT 43.750 46.560 44.070 46.620 ;
        RECT 29.055 46.420 37.080 46.560 ;
        RECT 29.460 46.375 29.810 46.420 ;
        RECT 29.490 46.360 29.810 46.375 ;
        RECT 23.970 46.020 24.290 46.280 ;
        RECT 25.825 46.220 26.115 46.265 ;
        RECT 28.570 46.220 28.890 46.280 ;
        RECT 25.825 46.080 28.890 46.220 ;
        RECT 36.940 46.220 37.080 46.420 ;
        RECT 37.280 46.420 44.070 46.560 ;
        RECT 37.280 46.375 37.570 46.420 ;
        RECT 43.750 46.360 44.070 46.420 ;
        RECT 45.130 46.560 45.450 46.620 ;
        RECT 46.525 46.560 46.815 46.605 ;
        RECT 45.130 46.420 46.815 46.560 ;
        RECT 48.900 46.560 49.040 46.715 ;
        RECT 50.280 46.560 50.420 46.715 ;
        RECT 50.650 46.700 50.970 46.760 ;
        RECT 51.125 46.715 51.415 46.760 ;
        RECT 52.045 46.900 52.335 46.945 ;
        RECT 53.410 46.900 53.730 46.960 ;
        RECT 52.045 46.760 53.730 46.900 ;
        RECT 52.045 46.715 52.335 46.760 ;
        RECT 53.410 46.700 53.730 46.760 ;
        RECT 53.870 46.700 54.190 46.960 ;
        RECT 55.250 46.700 55.570 46.960 ;
        RECT 55.710 46.900 56.030 46.960 ;
        RECT 56.185 46.900 56.475 46.945 ;
        RECT 55.710 46.760 56.475 46.900 ;
        RECT 55.710 46.700 56.030 46.760 ;
        RECT 56.185 46.715 56.475 46.760 ;
        RECT 75.000 46.860 75.875 51.695 ;
        RECT 76.675 51.515 78.500 51.695 ;
        RECT 80.675 51.875 89.550 52.765 ;
        RECT 76.585 51.285 78.585 51.515 ;
        RECT 80.675 51.245 80.905 51.875 ;
        RECT 81.395 51.820 82.395 51.875 ;
        RECT 89.315 51.310 89.550 51.875 ;
        RECT 89.315 51.245 89.545 51.310 ;
        RECT 76.195 49.800 76.425 51.235 ;
        RECT 78.745 49.800 78.975 51.235 ;
        RECT 81.110 50.965 89.110 51.195 ;
        RECT 81.180 50.840 89.010 50.965 ;
        RECT 81.200 50.055 89.000 50.840 ;
        RECT 81.110 49.825 89.110 50.055 ;
        RECT 76.195 48.460 78.975 49.800 ;
        RECT 80.675 49.750 80.905 49.775 ;
        RECT 76.195 47.275 76.425 48.460 ;
        RECT 76.770 47.225 78.365 48.460 ;
        RECT 78.745 47.570 78.975 48.460 ;
        RECT 80.670 49.305 80.905 49.750 ;
        RECT 89.315 49.750 89.545 49.775 ;
        RECT 80.670 49.295 81.085 49.305 ;
        RECT 81.225 49.295 82.225 49.365 ;
        RECT 80.670 49.290 82.225 49.295 ;
        RECT 82.635 49.290 84.255 49.295 ;
        RECT 89.315 49.290 89.550 49.750 ;
        RECT 80.670 48.400 89.550 49.290 ;
        RECT 80.670 48.385 82.225 48.400 ;
        RECT 82.635 48.395 84.255 48.400 ;
        RECT 80.670 48.295 81.085 48.385 ;
        RECT 81.225 48.335 82.225 48.385 ;
        RECT 80.670 47.865 80.905 48.295 ;
        RECT 80.675 47.815 80.905 47.865 ;
        RECT 89.315 47.865 89.550 48.400 ;
        RECT 89.315 47.815 89.545 47.865 ;
        RECT 81.110 47.570 89.110 47.765 ;
        RECT 78.745 47.535 89.110 47.570 ;
        RECT 78.745 47.390 89.030 47.535 ;
        RECT 78.745 47.375 81.245 47.390 ;
        RECT 78.745 47.275 78.975 47.375 ;
        RECT 76.585 46.995 78.585 47.225 ;
        RECT 89.880 47.115 90.580 55.285 ;
        RECT 84.955 46.985 85.230 47.055 ;
        RECT 79.260 46.860 85.230 46.985 ;
        RECT 75.000 46.845 76.405 46.860 ;
        RECT 78.750 46.845 85.230 46.860 ;
        RECT 75.000 46.795 85.230 46.845 ;
        RECT 51.585 46.560 51.875 46.605 ;
        RECT 48.900 46.420 49.500 46.560 ;
        RECT 50.280 46.420 51.875 46.560 ;
        RECT 45.130 46.360 45.450 46.420 ;
        RECT 46.525 46.375 46.815 46.420 ;
        RECT 43.290 46.220 43.610 46.280 ;
        RECT 44.225 46.220 44.515 46.265 ;
        RECT 36.940 46.080 44.515 46.220 ;
        RECT 25.825 46.035 26.115 46.080 ;
        RECT 28.570 46.020 28.890 46.080 ;
        RECT 43.290 46.020 43.610 46.080 ;
        RECT 44.225 46.035 44.515 46.080 ;
        RECT 47.905 46.220 48.195 46.265 ;
        RECT 48.810 46.220 49.130 46.280 ;
        RECT 47.905 46.080 49.130 46.220 ;
        RECT 49.360 46.220 49.500 46.420 ;
        RECT 51.585 46.375 51.875 46.420 ;
        RECT 53.960 46.220 54.100 46.700 ;
        RECT 49.360 46.080 54.100 46.220 ;
        RECT 75.000 46.670 79.450 46.795 ;
        RECT 84.955 46.720 85.230 46.795 ;
        RECT 47.905 46.035 48.195 46.080 ;
        RECT 48.810 46.020 49.130 46.080 ;
        RECT 22.520 45.400 58.400 45.880 ;
        RECT 43.750 45.000 44.070 45.260 ;
        RECT 46.050 45.200 46.370 45.260 ;
        RECT 50.665 45.200 50.955 45.245 ;
        RECT 46.050 45.060 50.955 45.200 ;
        RECT 46.050 45.000 46.370 45.060 ;
        RECT 50.665 45.015 50.955 45.060 ;
        RECT 55.725 45.015 56.015 45.245 ;
        RECT 23.970 44.860 24.290 44.920 ;
        RECT 29.550 44.860 29.840 44.905 ;
        RECT 23.970 44.720 29.840 44.860 ;
        RECT 23.970 44.660 24.290 44.720 ;
        RECT 29.550 44.675 29.840 44.720 ;
        RECT 34.550 44.660 34.870 44.920 ;
        RECT 55.800 44.860 55.940 45.015 ;
        RECT 54.420 44.720 55.940 44.860 ;
        RECT 54.420 44.580 54.560 44.720 ;
        RECT 30.870 44.320 31.190 44.580 ;
        RECT 48.810 44.320 49.130 44.580 ;
        RECT 49.730 44.320 50.050 44.580 ;
        RECT 54.330 44.320 54.650 44.580 ;
        RECT 55.265 44.520 55.555 44.565 ;
        RECT 55.710 44.520 56.030 44.580 ;
        RECT 55.265 44.380 56.030 44.520 ;
        RECT 55.265 44.335 55.555 44.380 ;
        RECT 55.710 44.320 56.030 44.380 ;
        RECT 56.630 44.320 56.950 44.580 ;
        RECT 26.295 44.180 26.585 44.225 ;
        RECT 28.815 44.180 29.105 44.225 ;
        RECT 30.005 44.180 30.295 44.225 ;
        RECT 26.295 44.040 30.295 44.180 ;
        RECT 26.295 43.995 26.585 44.040 ;
        RECT 28.815 43.995 29.105 44.040 ;
        RECT 30.005 43.995 30.295 44.040 ;
        RECT 40.990 44.180 41.310 44.240 ;
        RECT 46.525 44.180 46.815 44.225 ;
        RECT 40.990 44.040 46.815 44.180 ;
        RECT 40.990 43.980 41.310 44.040 ;
        RECT 46.525 43.995 46.815 44.040 ;
        RECT 26.730 43.840 27.020 43.885 ;
        RECT 28.300 43.840 28.590 43.885 ;
        RECT 30.400 43.840 30.690 43.885 ;
        RECT 26.730 43.700 30.690 43.840 ;
        RECT 26.730 43.655 27.020 43.700 ;
        RECT 28.300 43.655 28.590 43.700 ;
        RECT 30.400 43.655 30.690 43.700 ;
        RECT 23.970 43.300 24.290 43.560 ;
        RECT 40.530 43.500 40.850 43.560 ;
        RECT 41.005 43.500 41.295 43.545 ;
        RECT 40.530 43.360 41.295 43.500 ;
        RECT 40.530 43.300 40.850 43.360 ;
        RECT 41.005 43.315 41.295 43.360 ;
        RECT 45.590 43.500 45.910 43.560 ;
        RECT 48.825 43.500 49.115 43.545 ;
        RECT 45.590 43.360 49.115 43.500 ;
        RECT 45.590 43.300 45.910 43.360 ;
        RECT 48.825 43.315 49.115 43.360 ;
        RECT 52.030 43.500 52.350 43.560 ;
        RECT 55.265 43.500 55.555 43.545 ;
        RECT 52.030 43.360 55.555 43.500 ;
        RECT 52.030 43.300 52.350 43.360 ;
        RECT 55.265 43.315 55.555 43.360 ;
        RECT 22.520 42.680 58.400 43.160 ;
        RECT 28.570 42.280 28.890 42.540 ;
        RECT 36.850 42.280 37.170 42.540 ;
        RECT 37.310 42.480 37.630 42.540 ;
        RECT 39.165 42.480 39.455 42.525 ;
        RECT 37.310 42.340 39.455 42.480 ;
        RECT 37.310 42.280 37.630 42.340 ;
        RECT 39.165 42.295 39.455 42.340 ;
        RECT 47.890 42.280 48.210 42.540 ;
        RECT 55.250 42.480 55.570 42.540 ;
        RECT 56.185 42.480 56.475 42.525 ;
        RECT 55.250 42.340 56.475 42.480 ;
        RECT 55.250 42.280 55.570 42.340 ;
        RECT 56.185 42.295 56.475 42.340 ;
        RECT 38.245 42.140 38.535 42.185 ;
        RECT 41.450 42.140 41.770 42.200 ;
        RECT 45.590 42.140 45.910 42.200 ;
        RECT 38.245 42.000 41.770 42.140 ;
        RECT 38.245 41.955 38.535 42.000 ;
        RECT 23.970 41.800 24.290 41.860 ;
        RECT 25.365 41.800 25.655 41.845 ;
        RECT 38.320 41.800 38.460 41.955 ;
        RECT 41.450 41.940 41.770 42.000 ;
        RECT 44.300 42.000 45.910 42.140 ;
        RECT 23.970 41.660 25.655 41.800 ;
        RECT 23.970 41.600 24.290 41.660 ;
        RECT 25.365 41.615 25.655 41.660 ;
        RECT 36.940 41.660 38.460 41.800 ;
        RECT 38.705 41.800 38.995 41.845 ;
        RECT 44.300 41.800 44.440 42.000 ;
        RECT 45.590 41.940 45.910 42.000 ;
        RECT 53.870 41.940 54.190 42.200 ;
        RECT 38.705 41.660 44.440 41.800 ;
        RECT 31.790 41.260 32.110 41.520 ;
        RECT 36.940 41.505 37.080 41.660 ;
        RECT 38.705 41.615 38.995 41.660 ;
        RECT 44.670 41.600 44.990 41.860 ;
        RECT 53.960 41.800 54.100 41.940 ;
        RECT 47.520 41.660 54.100 41.800 ;
        RECT 35.945 41.275 36.235 41.505 ;
        RECT 36.865 41.275 37.155 41.505 ;
        RECT 36.020 41.120 36.160 41.275 ;
        RECT 37.310 41.260 37.630 41.520 ;
        RECT 39.625 41.460 39.915 41.505 ;
        RECT 40.070 41.460 40.390 41.520 ;
        RECT 39.625 41.320 40.390 41.460 ;
        RECT 39.625 41.275 39.915 41.320 ;
        RECT 40.070 41.260 40.390 41.320 ;
        RECT 40.990 41.260 41.310 41.520 ;
        RECT 47.520 41.505 47.660 41.660 ;
        RECT 47.445 41.275 47.735 41.505 ;
        RECT 48.365 41.460 48.655 41.505 ;
        RECT 50.205 41.460 50.495 41.505 ;
        RECT 50.650 41.460 50.970 41.520 ;
        RECT 51.200 41.505 51.340 41.660 ;
        RECT 48.365 41.320 50.970 41.460 ;
        RECT 48.365 41.275 48.655 41.320 ;
        RECT 50.205 41.275 50.495 41.320 ;
        RECT 50.650 41.260 50.970 41.320 ;
        RECT 51.125 41.275 51.415 41.505 ;
        RECT 51.570 41.260 51.890 41.520 ;
        RECT 52.965 41.275 53.255 41.505 ;
        RECT 41.465 41.120 41.755 41.165 ;
        RECT 36.020 40.980 41.755 41.120 ;
        RECT 41.465 40.935 41.755 40.980 ;
        RECT 49.745 41.120 50.035 41.165 ;
        RECT 52.030 41.120 52.350 41.180 ;
        RECT 53.040 41.120 53.180 41.275 ;
        RECT 53.870 41.260 54.190 41.520 ;
        RECT 54.330 41.460 54.650 41.520 ;
        RECT 55.265 41.460 55.555 41.505 ;
        RECT 54.330 41.320 55.555 41.460 ;
        RECT 54.330 41.260 54.650 41.320 ;
        RECT 55.265 41.275 55.555 41.320 ;
        RECT 75.000 41.390 75.875 46.670 ;
        RECT 77.825 46.365 81.610 46.370 ;
        RECT 77.825 46.300 85.060 46.365 ;
        RECT 76.645 46.175 85.060 46.300 ;
        RECT 76.645 46.085 85.105 46.175 ;
        RECT 76.585 46.075 85.105 46.085 ;
        RECT 76.585 45.855 78.585 46.075 ;
        RECT 81.105 45.945 85.105 46.075 ;
        RECT 76.195 44.425 76.425 45.805 ;
        RECT 78.745 44.425 78.975 45.805 ;
        RECT 76.195 43.470 78.975 44.425 ;
        RECT 76.195 41.845 76.425 43.470 ;
        RECT 78.745 41.845 78.975 43.470 ;
        RECT 80.670 44.640 80.900 45.895 ;
        RECT 82.340 44.640 83.725 45.945 ;
        RECT 85.310 44.640 85.540 45.895 ;
        RECT 85.905 45.435 90.580 47.115 ;
        RECT 87.265 45.095 87.540 45.125 ;
        RECT 87.250 44.840 87.580 45.095 ;
        RECT 87.265 44.820 87.555 44.840 ;
        RECT 87.265 44.790 87.540 44.820 ;
        RECT 80.670 44.570 85.540 44.640 ;
        RECT 87.075 44.570 87.305 44.615 ;
        RECT 80.670 43.295 85.545 44.570 ;
        RECT 80.670 41.935 80.900 43.295 ;
        RECT 85.310 41.935 85.545 43.295 ;
        RECT 76.585 41.565 78.585 41.795 ;
        RECT 76.650 41.390 78.520 41.565 ;
        RECT 54.790 41.120 55.110 41.180 ;
        RECT 49.745 40.980 52.350 41.120 ;
        RECT 49.745 40.935 50.035 40.980 ;
        RECT 52.030 40.920 52.350 40.980 ;
        RECT 52.580 40.980 55.110 41.120 ;
        RECT 29.030 40.580 29.350 40.840 ;
        RECT 46.525 40.780 46.815 40.825 ;
        RECT 47.430 40.780 47.750 40.840 ;
        RECT 46.525 40.640 47.750 40.780 ;
        RECT 46.525 40.595 46.815 40.640 ;
        RECT 47.430 40.580 47.750 40.640 ;
        RECT 50.190 40.780 50.510 40.840 ;
        RECT 52.580 40.825 52.720 40.980 ;
        RECT 54.790 40.920 55.110 40.980 ;
        RECT 75.000 40.835 78.520 41.390 ;
        RECT 50.665 40.780 50.955 40.825 ;
        RECT 50.190 40.640 50.955 40.780 ;
        RECT 50.190 40.580 50.510 40.640 ;
        RECT 50.665 40.595 50.955 40.640 ;
        RECT 52.505 40.595 52.795 40.825 ;
        RECT 22.520 39.960 58.400 40.440 ;
        RECT 23.510 39.760 23.830 39.820 ;
        RECT 24.445 39.760 24.735 39.805 ;
        RECT 23.510 39.620 24.735 39.760 ;
        RECT 23.510 39.560 23.830 39.620 ;
        RECT 24.445 39.575 24.735 39.620 ;
        RECT 28.125 39.760 28.415 39.805 ;
        RECT 29.030 39.760 29.350 39.820 ;
        RECT 28.125 39.620 29.350 39.760 ;
        RECT 28.125 39.575 28.415 39.620 ;
        RECT 29.030 39.560 29.350 39.620 ;
        RECT 37.310 39.760 37.630 39.820 ;
        RECT 44.210 39.760 44.530 39.820 ;
        RECT 37.310 39.620 44.530 39.760 ;
        RECT 37.310 39.560 37.630 39.620 ;
        RECT 44.210 39.560 44.530 39.620 ;
        RECT 53.870 39.760 54.190 39.820 ;
        RECT 56.185 39.760 56.475 39.805 ;
        RECT 53.870 39.620 56.475 39.760 ;
        RECT 53.870 39.560 54.190 39.620 ;
        RECT 56.185 39.575 56.475 39.620 ;
        RECT 31.760 39.420 32.050 39.465 ;
        RECT 35.470 39.420 35.790 39.480 ;
        RECT 36.850 39.420 37.170 39.480 ;
        RECT 52.030 39.420 52.350 39.480 ;
        RECT 31.760 39.280 37.170 39.420 ;
        RECT 31.760 39.235 32.050 39.280 ;
        RECT 35.470 39.220 35.790 39.280 ;
        RECT 36.850 39.220 37.170 39.280 ;
        RECT 49.820 39.280 52.350 39.420 ;
        RECT 23.970 39.080 24.290 39.140 ;
        RECT 25.365 39.080 25.655 39.125 ;
        RECT 23.970 38.940 25.655 39.080 ;
        RECT 23.970 38.880 24.290 38.940 ;
        RECT 25.365 38.895 25.655 38.940 ;
        RECT 39.625 39.080 39.915 39.125 ;
        RECT 41.925 39.080 42.215 39.125 ;
        RECT 39.625 38.940 42.215 39.080 ;
        RECT 39.625 38.895 39.915 38.940 ;
        RECT 41.925 38.895 42.215 38.940 ;
        RECT 47.890 39.080 48.210 39.140 ;
        RECT 49.820 39.125 49.960 39.280 ;
        RECT 52.030 39.220 52.350 39.280 ;
        RECT 49.285 39.080 49.575 39.125 ;
        RECT 47.890 38.940 49.575 39.080 ;
        RECT 47.890 38.880 48.210 38.940 ;
        RECT 49.285 38.895 49.575 38.940 ;
        RECT 49.745 38.895 50.035 39.125 ;
        RECT 50.190 38.880 50.510 39.140 ;
        RECT 52.965 39.080 53.255 39.125 ;
        RECT 53.410 39.080 53.730 39.140 ;
        RECT 52.965 38.940 53.730 39.080 ;
        RECT 52.965 38.895 53.255 38.940 ;
        RECT 53.410 38.880 53.730 38.940 ;
        RECT 53.870 38.880 54.190 39.140 ;
        RECT 55.265 39.080 55.555 39.125 ;
        RECT 55.710 39.080 56.030 39.140 ;
        RECT 55.265 38.940 56.030 39.080 ;
        RECT 55.265 38.895 55.555 38.940 ;
        RECT 55.710 38.880 56.030 38.940 ;
        RECT 28.585 38.740 28.875 38.785 ;
        RECT 29.030 38.740 29.350 38.800 ;
        RECT 28.585 38.600 29.350 38.740 ;
        RECT 28.585 38.555 28.875 38.600 ;
        RECT 29.030 38.540 29.350 38.600 ;
        RECT 29.490 38.540 29.810 38.800 ;
        RECT 30.425 38.555 30.715 38.785 ;
        RECT 31.305 38.740 31.595 38.785 ;
        RECT 32.495 38.740 32.785 38.785 ;
        RECT 35.015 38.740 35.305 38.785 ;
        RECT 31.305 38.600 35.305 38.740 ;
        RECT 31.305 38.555 31.595 38.600 ;
        RECT 32.495 38.555 32.785 38.600 ;
        RECT 35.015 38.555 35.305 38.600 ;
        RECT 40.085 38.555 40.375 38.785 ;
        RECT 41.005 38.740 41.295 38.785 ;
        RECT 43.290 38.740 43.610 38.800 ;
        RECT 41.005 38.600 43.610 38.740 ;
        RECT 41.005 38.555 41.295 38.600 ;
        RECT 23.970 38.400 24.290 38.460 ;
        RECT 30.500 38.400 30.640 38.555 ;
        RECT 23.970 38.260 30.640 38.400 ;
        RECT 30.910 38.400 31.200 38.445 ;
        RECT 33.010 38.400 33.300 38.445 ;
        RECT 34.580 38.400 34.870 38.445 ;
        RECT 30.910 38.260 34.870 38.400 ;
        RECT 23.970 38.200 24.290 38.260 ;
        RECT 30.910 38.215 31.200 38.260 ;
        RECT 33.010 38.215 33.300 38.260 ;
        RECT 34.580 38.215 34.870 38.260 ;
        RECT 36.850 38.400 37.170 38.460 ;
        RECT 37.785 38.400 38.075 38.445 ;
        RECT 36.850 38.260 38.075 38.400 ;
        RECT 40.160 38.400 40.300 38.555 ;
        RECT 43.290 38.540 43.610 38.600 ;
        RECT 43.750 38.740 44.070 38.800 ;
        RECT 44.685 38.740 44.975 38.785 ;
        RECT 43.750 38.600 44.975 38.740 ;
        RECT 43.750 38.540 44.070 38.600 ;
        RECT 44.685 38.555 44.975 38.600 ;
        RECT 50.665 38.740 50.955 38.785 ;
        RECT 54.330 38.740 54.650 38.800 ;
        RECT 50.665 38.600 54.650 38.740 ;
        RECT 50.665 38.555 50.955 38.600 ;
        RECT 54.330 38.540 54.650 38.600 ;
        RECT 45.590 38.400 45.910 38.460 ;
        RECT 51.585 38.400 51.875 38.445 ;
        RECT 40.160 38.260 51.875 38.400 ;
        RECT 36.850 38.200 37.170 38.260 ;
        RECT 37.785 38.215 38.075 38.260 ;
        RECT 45.590 38.200 45.910 38.260 ;
        RECT 51.585 38.215 51.875 38.260 ;
        RECT 26.270 37.860 26.590 38.120 ;
        RECT 22.520 37.240 58.400 37.720 ;
        RECT 30.885 37.040 31.175 37.085 ;
        RECT 31.790 37.040 32.110 37.100 ;
        RECT 30.885 36.900 32.110 37.040 ;
        RECT 30.885 36.855 31.175 36.900 ;
        RECT 31.790 36.840 32.110 36.900 ;
        RECT 45.605 37.040 45.895 37.085 ;
        RECT 46.510 37.040 46.830 37.100 ;
        RECT 45.605 36.900 46.830 37.040 ;
        RECT 45.605 36.855 45.895 36.900 ;
        RECT 46.510 36.840 46.830 36.900 ;
        RECT 52.490 37.040 52.810 37.100 ;
        RECT 53.425 37.040 53.715 37.085 ;
        RECT 52.490 36.900 53.715 37.040 ;
        RECT 52.490 36.840 52.810 36.900 ;
        RECT 53.425 36.855 53.715 36.900 ;
        RECT 24.470 36.700 24.760 36.745 ;
        RECT 26.570 36.700 26.860 36.745 ;
        RECT 28.140 36.700 28.430 36.745 ;
        RECT 24.470 36.560 28.430 36.700 ;
        RECT 24.470 36.515 24.760 36.560 ;
        RECT 26.570 36.515 26.860 36.560 ;
        RECT 28.140 36.515 28.430 36.560 ;
        RECT 36.430 36.700 36.720 36.745 ;
        RECT 38.530 36.700 38.820 36.745 ;
        RECT 40.100 36.700 40.390 36.745 ;
        RECT 36.430 36.560 40.390 36.700 ;
        RECT 36.430 36.515 36.720 36.560 ;
        RECT 38.530 36.515 38.820 36.560 ;
        RECT 40.100 36.515 40.390 36.560 ;
        RECT 45.130 36.500 45.450 36.760 ;
        RECT 23.970 36.160 24.290 36.420 ;
        RECT 24.865 36.360 25.155 36.405 ;
        RECT 26.055 36.360 26.345 36.405 ;
        RECT 28.575 36.360 28.865 36.405 ;
        RECT 24.865 36.220 28.865 36.360 ;
        RECT 24.865 36.175 25.155 36.220 ;
        RECT 26.055 36.175 26.345 36.220 ;
        RECT 28.575 36.175 28.865 36.220 ;
        RECT 36.825 36.360 37.115 36.405 ;
        RECT 38.015 36.360 38.305 36.405 ;
        RECT 40.535 36.360 40.825 36.405 ;
        RECT 36.825 36.220 40.825 36.360 ;
        RECT 36.825 36.175 37.115 36.220 ;
        RECT 38.015 36.175 38.305 36.220 ;
        RECT 40.535 36.175 40.825 36.220 ;
        RECT 43.305 36.360 43.595 36.405 ;
        RECT 44.210 36.360 44.530 36.420 ;
        RECT 43.305 36.220 44.530 36.360 ;
        RECT 43.305 36.175 43.595 36.220 ;
        RECT 44.210 36.160 44.530 36.220 ;
        RECT 52.030 36.360 52.350 36.420 ;
        RECT 52.030 36.220 55.940 36.360 ;
        RECT 52.030 36.160 52.350 36.220 ;
        RECT 24.060 36.020 24.200 36.160 ;
        RECT 30.870 36.020 31.190 36.080 ;
        RECT 35.945 36.020 36.235 36.065 ;
        RECT 24.060 35.880 36.235 36.020 ;
        RECT 30.870 35.820 31.190 35.880 ;
        RECT 35.945 35.835 36.235 35.880 ;
        RECT 37.280 35.835 37.570 36.065 ;
        RECT 25.320 35.680 25.610 35.725 ;
        RECT 26.270 35.680 26.590 35.740 ;
        RECT 25.320 35.540 26.590 35.680 ;
        RECT 25.320 35.495 25.610 35.540 ;
        RECT 26.270 35.480 26.590 35.540 ;
        RECT 36.020 35.340 36.160 35.835 ;
        RECT 36.850 35.680 37.170 35.740 ;
        RECT 37.400 35.680 37.540 35.835 ;
        RECT 49.730 35.820 50.050 36.080 ;
        RECT 52.490 36.020 52.810 36.080 ;
        RECT 54.345 36.020 54.635 36.065 ;
        RECT 52.490 35.880 54.635 36.020 ;
        RECT 52.490 35.820 52.810 35.880 ;
        RECT 54.345 35.835 54.635 35.880 ;
        RECT 54.790 35.820 55.110 36.080 ;
        RECT 55.250 35.820 55.570 36.080 ;
        RECT 55.800 36.065 55.940 36.220 ;
        RECT 55.725 35.835 56.015 36.065 ;
        RECT 36.850 35.540 37.540 35.680 ;
        RECT 75.000 35.730 75.875 40.835 ;
        RECT 76.650 40.655 78.520 40.835 ;
        RECT 76.585 40.425 78.585 40.655 ;
        RECT 80.710 40.465 80.870 41.935 ;
        RECT 85.340 41.925 85.545 41.935 ;
        RECT 81.105 41.655 85.105 41.885 ;
        RECT 81.185 41.410 85.010 41.655 ;
        RECT 87.065 41.410 87.305 44.570 ;
        RECT 81.185 40.920 87.305 41.410 ;
        RECT 81.185 40.745 85.010 40.920 ;
        RECT 81.105 40.515 85.105 40.745 ;
        RECT 76.195 38.980 76.425 40.375 ;
        RECT 78.745 38.980 78.975 40.375 ;
        RECT 76.195 38.025 78.975 38.980 ;
        RECT 76.195 36.415 76.425 38.025 ;
        RECT 78.745 36.415 78.975 38.025 ;
        RECT 80.670 39.090 80.900 40.465 ;
        RECT 85.310 40.350 85.540 40.465 ;
        RECT 85.310 39.715 85.545 40.350 ;
        RECT 87.065 39.715 87.305 40.920 ;
        RECT 85.310 39.090 85.540 39.715 ;
        RECT 87.075 39.615 87.305 39.715 ;
        RECT 87.515 44.600 87.745 44.615 ;
        RECT 88.165 44.600 88.645 45.435 ;
        RECT 87.515 39.675 88.655 44.600 ;
        RECT 87.515 39.615 87.745 39.675 ;
        RECT 87.265 39.405 87.555 39.410 ;
        RECT 87.250 39.150 87.580 39.405 ;
        RECT 80.670 37.745 85.540 39.090 ;
        RECT 80.670 36.505 80.900 37.745 ;
        RECT 85.310 36.505 85.540 37.745 ;
        RECT 76.585 36.340 78.585 36.365 ;
        RECT 81.105 36.340 85.105 36.455 ;
        RECT 76.585 36.265 78.590 36.340 ;
        RECT 79.125 36.265 85.105 36.340 ;
        RECT 76.585 36.225 85.105 36.265 ;
        RECT 76.585 36.135 85.040 36.225 ;
        RECT 76.640 36.000 85.040 36.135 ;
        RECT 36.850 35.480 37.170 35.540 ;
        RECT 40.990 35.340 41.310 35.400 ;
        RECT 36.020 35.200 41.310 35.340 ;
        RECT 40.990 35.140 41.310 35.200 ;
        RECT 42.845 35.340 43.135 35.385 ;
        RECT 43.750 35.340 44.070 35.400 ;
        RECT 42.845 35.200 44.070 35.340 ;
        RECT 42.845 35.155 43.135 35.200 ;
        RECT 43.750 35.140 44.070 35.200 ;
        RECT 50.650 35.340 50.970 35.400 ;
        RECT 52.965 35.340 53.255 35.385 ;
        RECT 50.650 35.200 53.255 35.340 ;
        RECT 50.650 35.140 50.970 35.200 ;
        RECT 52.965 35.155 53.255 35.200 ;
        RECT 75.000 35.290 76.860 35.730 ;
        RECT 75.000 35.280 77.850 35.290 ;
        RECT 22.520 34.520 58.400 35.000 ;
        RECT 75.000 34.935 78.520 35.280 ;
        RECT 50.650 34.120 50.970 34.380 ;
        RECT 54.330 34.120 54.650 34.380 ;
        RECT 45.590 33.980 45.910 34.040 ;
        RECT 40.620 33.840 45.910 33.980 ;
        RECT 25.365 33.640 25.655 33.685 ;
        RECT 31.790 33.640 32.110 33.700 ;
        RECT 25.365 33.500 32.110 33.640 ;
        RECT 25.365 33.455 25.655 33.500 ;
        RECT 31.790 33.440 32.110 33.500 ;
        RECT 34.565 33.640 34.855 33.685 ;
        RECT 36.865 33.640 37.155 33.685 ;
        RECT 34.565 33.500 37.155 33.640 ;
        RECT 34.565 33.455 34.855 33.500 ;
        RECT 36.865 33.455 37.155 33.500 ;
        RECT 23.970 33.300 24.290 33.360 ;
        RECT 26.745 33.300 27.035 33.345 ;
        RECT 23.970 33.160 27.035 33.300 ;
        RECT 23.970 33.100 24.290 33.160 ;
        RECT 26.745 33.115 27.035 33.160 ;
        RECT 31.330 33.100 31.650 33.360 ;
        RECT 35.470 33.100 35.790 33.360 ;
        RECT 36.405 33.300 36.695 33.345 ;
        RECT 40.620 33.300 40.760 33.840 ;
        RECT 45.590 33.780 45.910 33.840 ;
        RECT 54.790 33.980 55.110 34.040 ;
        RECT 56.645 33.980 56.935 34.025 ;
        RECT 54.790 33.840 56.935 33.980 ;
        RECT 54.790 33.780 55.110 33.840 ;
        RECT 56.645 33.795 56.935 33.840 ;
        RECT 40.990 33.440 41.310 33.700 ;
        RECT 42.340 33.640 42.630 33.685 ;
        RECT 46.510 33.640 46.830 33.700 ;
        RECT 42.340 33.500 46.280 33.640 ;
        RECT 42.340 33.455 42.630 33.500 ;
        RECT 36.405 33.160 40.760 33.300 ;
        RECT 41.885 33.300 42.175 33.345 ;
        RECT 43.075 33.300 43.365 33.345 ;
        RECT 45.595 33.300 45.885 33.345 ;
        RECT 41.885 33.160 45.885 33.300 ;
        RECT 36.405 33.115 36.695 33.160 ;
        RECT 41.885 33.115 42.175 33.160 ;
        RECT 43.075 33.115 43.365 33.160 ;
        RECT 45.595 33.115 45.885 33.160 ;
        RECT 23.510 32.960 23.830 33.020 ;
        RECT 24.445 32.960 24.735 33.005 ;
        RECT 23.510 32.820 24.735 32.960 ;
        RECT 23.510 32.760 23.830 32.820 ;
        RECT 24.445 32.775 24.735 32.820 ;
        RECT 29.030 32.960 29.350 33.020 ;
        RECT 41.490 32.960 41.780 33.005 ;
        RECT 43.590 32.960 43.880 33.005 ;
        RECT 45.160 32.960 45.450 33.005 ;
        RECT 29.030 32.820 41.220 32.960 ;
        RECT 29.030 32.760 29.350 32.820 ;
        RECT 28.570 32.620 28.890 32.680 ;
        RECT 29.965 32.620 30.255 32.665 ;
        RECT 28.570 32.480 30.255 32.620 ;
        RECT 28.570 32.420 28.890 32.480 ;
        RECT 29.965 32.435 30.255 32.480 ;
        RECT 38.705 32.620 38.995 32.665 ;
        RECT 40.070 32.620 40.390 32.680 ;
        RECT 38.705 32.480 40.390 32.620 ;
        RECT 41.080 32.620 41.220 32.820 ;
        RECT 41.490 32.820 45.450 32.960 ;
        RECT 46.140 32.960 46.280 33.500 ;
        RECT 46.510 33.500 51.800 33.640 ;
        RECT 46.510 33.440 46.830 33.500 ;
        RECT 47.430 33.300 47.750 33.360 ;
        RECT 51.660 33.345 51.800 33.500 ;
        RECT 52.950 33.440 53.270 33.700 ;
        RECT 54.330 33.640 54.650 33.700 ;
        RECT 55.265 33.640 55.555 33.685 ;
        RECT 54.330 33.500 55.555 33.640 ;
        RECT 54.330 33.440 54.650 33.500 ;
        RECT 55.265 33.455 55.555 33.500 ;
        RECT 51.125 33.300 51.415 33.345 ;
        RECT 47.430 33.160 51.415 33.300 ;
        RECT 47.430 33.100 47.750 33.160 ;
        RECT 51.125 33.115 51.415 33.160 ;
        RECT 51.585 33.115 51.875 33.345 ;
        RECT 52.490 33.300 52.810 33.360 ;
        RECT 55.710 33.300 56.030 33.360 ;
        RECT 52.490 33.160 56.030 33.300 ;
        RECT 52.490 33.100 52.810 33.160 ;
        RECT 55.710 33.100 56.030 33.160 ;
        RECT 75.000 33.310 76.860 34.935 ;
        RECT 77.660 34.785 78.520 34.935 ;
        RECT 77.155 34.595 77.405 34.610 ;
        RECT 77.155 34.305 77.430 34.595 ;
        RECT 77.590 34.555 78.590 34.785 ;
        RECT 79.010 34.690 79.280 36.000 ;
        RECT 89.880 35.570 90.580 45.435 ;
        RECT 84.300 35.235 90.580 35.570 ;
        RECT 81.185 35.095 90.580 35.235 ;
        RECT 81.185 34.870 85.045 35.095 ;
        RECT 77.155 34.275 77.405 34.305 ;
        RECT 77.590 34.115 78.590 34.345 ;
        RECT 78.735 34.270 80.925 34.690 ;
        RECT 81.120 34.640 85.120 34.870 ;
        RECT 85.355 34.680 85.605 34.700 ;
        RECT 81.120 34.200 85.120 34.430 ;
        RECT 85.325 34.390 85.605 34.680 ;
        RECT 85.355 34.365 85.605 34.390 ;
        RECT 77.660 33.975 78.545 34.115 ;
        RECT 81.170 34.035 85.095 34.200 ;
        RECT 78.730 33.975 85.095 34.035 ;
        RECT 77.660 33.920 85.095 33.975 ;
        RECT 77.660 33.850 81.540 33.920 ;
        RECT 78.215 33.735 81.540 33.850 ;
        RECT 89.880 33.770 90.580 35.095 ;
        RECT 75.000 33.265 77.385 33.310 ;
        RECT 48.825 32.960 49.115 33.005 ;
        RECT 46.140 32.820 49.115 32.960 ;
        RECT 41.490 32.775 41.780 32.820 ;
        RECT 43.590 32.775 43.880 32.820 ;
        RECT 45.160 32.775 45.450 32.820 ;
        RECT 48.825 32.775 49.115 32.820 ;
        RECT 53.885 32.960 54.175 33.005 ;
        RECT 56.630 32.960 56.950 33.020 ;
        RECT 53.885 32.820 56.950 32.960 ;
        RECT 53.885 32.775 54.175 32.820 ;
        RECT 56.630 32.760 56.950 32.820 ;
        RECT 47.430 32.620 47.750 32.680 ;
        RECT 41.080 32.480 47.750 32.620 ;
        RECT 38.705 32.435 38.995 32.480 ;
        RECT 40.070 32.420 40.390 32.480 ;
        RECT 47.430 32.420 47.750 32.480 ;
        RECT 47.905 32.620 48.195 32.665 ;
        RECT 49.730 32.620 50.050 32.680 ;
        RECT 47.905 32.480 50.050 32.620 ;
        RECT 47.905 32.435 48.195 32.480 ;
        RECT 49.730 32.420 50.050 32.480 ;
        RECT 53.410 32.620 53.730 32.680 ;
        RECT 55.265 32.620 55.555 32.665 ;
        RECT 53.410 32.480 55.555 32.620 ;
        RECT 53.410 32.420 53.730 32.480 ;
        RECT 55.265 32.435 55.555 32.480 ;
        RECT 22.520 31.800 58.400 32.280 ;
        RECT 23.970 31.400 24.290 31.660 ;
        RECT 40.990 31.600 41.310 31.660 ;
        RECT 42.385 31.600 42.675 31.645 ;
        RECT 40.990 31.460 42.675 31.600 ;
        RECT 40.990 31.400 41.310 31.460 ;
        RECT 42.385 31.415 42.675 31.460 ;
        RECT 50.205 31.600 50.495 31.645 ;
        RECT 52.490 31.600 52.810 31.660 ;
        RECT 50.205 31.460 52.810 31.600 ;
        RECT 50.205 31.415 50.495 31.460 ;
        RECT 52.490 31.400 52.810 31.460 ;
        RECT 53.425 31.600 53.715 31.645 ;
        RECT 53.870 31.600 54.190 31.660 ;
        RECT 53.425 31.460 54.190 31.600 ;
        RECT 75.000 31.535 75.875 33.265 ;
        RECT 76.240 32.990 77.385 33.265 ;
        RECT 79.570 33.105 79.975 33.735 ;
        RECT 88.575 33.235 90.580 33.770 ;
        RECT 76.240 32.925 78.490 32.990 ;
        RECT 76.680 32.760 78.490 32.925 ;
        RECT 76.165 32.570 76.415 32.595 ;
        RECT 76.165 32.280 76.435 32.570 ;
        RECT 76.595 32.530 78.595 32.760 ;
        RECT 79.555 32.740 79.980 33.105 ;
        RECT 81.220 33.090 90.580 33.235 ;
        RECT 81.220 32.845 89.075 33.090 ;
        RECT 76.165 32.260 76.415 32.280 ;
        RECT 76.595 32.090 78.595 32.320 ;
        RECT 78.745 32.230 80.935 32.740 ;
        RECT 81.125 32.615 89.125 32.845 ;
        RECT 89.355 32.655 89.605 32.670 ;
        RECT 78.745 32.225 79.445 32.230 ;
        RECT 80.445 32.225 80.935 32.230 ;
        RECT 81.125 32.175 89.125 32.405 ;
        RECT 89.330 32.365 89.605 32.655 ;
        RECT 89.355 32.335 89.605 32.365 ;
        RECT 76.665 31.925 78.530 32.090 ;
        RECT 79.415 31.925 80.415 32.000 ;
        RECT 81.200 31.925 89.050 32.175 ;
        RECT 76.665 31.630 89.050 31.925 ;
        RECT 89.880 31.690 90.580 33.090 ;
        RECT 92.000 58.025 92.875 58.140 ;
        RECT 92.000 57.665 98.445 58.025 ;
        RECT 92.000 57.530 105.975 57.665 ;
        RECT 92.000 57.085 92.875 57.530 ;
        RECT 98.015 57.435 105.975 57.530 ;
        RECT 92.000 56.860 92.885 57.085 ;
        RECT 93.595 57.000 94.815 57.085 ;
        RECT 93.595 56.945 94.830 57.000 ;
        RECT 92.000 52.185 92.875 56.860 ;
        RECT 93.585 56.715 95.585 56.945 ;
        RECT 93.195 55.465 93.425 56.665 ;
        RECT 93.970 55.465 95.135 56.715 ;
        RECT 95.745 55.465 95.975 56.665 ;
        RECT 93.195 54.675 95.975 55.465 ;
        RECT 97.735 56.510 97.965 57.230 ;
        RECT 97.735 56.485 98.100 56.510 ;
        RECT 98.260 56.485 98.580 56.540 ;
        RECT 97.735 56.335 98.580 56.485 ;
        RECT 97.735 56.305 98.100 56.335 ;
        RECT 97.735 55.230 97.965 56.305 ;
        RECT 98.260 56.280 98.580 56.335 ;
        RECT 100.865 55.055 102.680 57.435 ;
        RECT 106.025 57.195 106.255 57.230 ;
        RECT 106.880 57.195 107.580 58.165 ;
        RECT 106.025 55.285 107.580 57.195 ;
        RECT 106.025 55.230 106.255 55.285 ;
        RECT 98.265 55.025 105.895 55.055 ;
        RECT 98.015 54.795 105.975 55.025 ;
        RECT 93.195 52.705 93.425 54.675 ;
        RECT 95.745 54.005 95.975 54.675 ;
        RECT 95.745 53.725 98.610 54.005 ;
        RECT 95.745 53.635 106.030 53.725 ;
        RECT 95.745 52.705 95.975 53.635 ;
        RECT 98.170 53.485 106.030 53.635 ;
        RECT 98.110 53.255 106.110 53.485 ;
        RECT 97.675 52.765 97.905 53.205 ;
        RECT 106.315 53.195 106.545 53.205 ;
        RECT 98.395 52.765 99.395 52.835 ;
        RECT 106.315 52.765 106.550 53.195 ;
        RECT 93.585 52.425 95.585 52.655 ;
        RECT 93.675 52.185 95.500 52.425 ;
        RECT 92.000 51.695 95.500 52.185 ;
        RECT 92.000 46.860 92.875 51.695 ;
        RECT 93.675 51.515 95.500 51.695 ;
        RECT 97.675 51.875 106.550 52.765 ;
        RECT 93.585 51.285 95.585 51.515 ;
        RECT 97.675 51.245 97.905 51.875 ;
        RECT 98.395 51.820 99.395 51.875 ;
        RECT 106.315 51.310 106.550 51.875 ;
        RECT 106.315 51.245 106.545 51.310 ;
        RECT 93.195 49.800 93.425 51.235 ;
        RECT 95.745 49.800 95.975 51.235 ;
        RECT 98.110 50.965 106.110 51.195 ;
        RECT 98.180 50.840 106.010 50.965 ;
        RECT 98.200 50.055 106.000 50.840 ;
        RECT 98.110 49.825 106.110 50.055 ;
        RECT 93.195 48.460 95.975 49.800 ;
        RECT 97.675 49.750 97.905 49.775 ;
        RECT 93.195 47.275 93.425 48.460 ;
        RECT 93.770 47.225 95.365 48.460 ;
        RECT 95.745 47.570 95.975 48.460 ;
        RECT 97.670 49.305 97.905 49.750 ;
        RECT 106.315 49.750 106.545 49.775 ;
        RECT 97.670 49.295 98.085 49.305 ;
        RECT 98.225 49.295 99.225 49.365 ;
        RECT 97.670 49.290 99.225 49.295 ;
        RECT 99.635 49.290 101.255 49.295 ;
        RECT 106.315 49.290 106.550 49.750 ;
        RECT 97.670 48.400 106.550 49.290 ;
        RECT 97.670 48.385 99.225 48.400 ;
        RECT 99.635 48.395 101.255 48.400 ;
        RECT 97.670 48.295 98.085 48.385 ;
        RECT 98.225 48.335 99.225 48.385 ;
        RECT 97.670 47.865 97.905 48.295 ;
        RECT 97.675 47.815 97.905 47.865 ;
        RECT 106.315 47.865 106.550 48.400 ;
        RECT 106.315 47.815 106.545 47.865 ;
        RECT 98.110 47.570 106.110 47.765 ;
        RECT 95.745 47.535 106.110 47.570 ;
        RECT 95.745 47.390 106.030 47.535 ;
        RECT 95.745 47.375 98.245 47.390 ;
        RECT 95.745 47.275 95.975 47.375 ;
        RECT 93.585 46.995 95.585 47.225 ;
        RECT 106.880 47.115 107.580 55.285 ;
        RECT 101.955 46.985 102.230 47.055 ;
        RECT 96.260 46.860 102.230 46.985 ;
        RECT 92.000 46.845 93.405 46.860 ;
        RECT 95.750 46.845 102.230 46.860 ;
        RECT 92.000 46.795 102.230 46.845 ;
        RECT 92.000 46.670 96.450 46.795 ;
        RECT 101.955 46.720 102.230 46.795 ;
        RECT 92.000 41.390 92.875 46.670 ;
        RECT 94.825 46.365 98.610 46.370 ;
        RECT 94.825 46.300 102.060 46.365 ;
        RECT 93.645 46.175 102.060 46.300 ;
        RECT 93.645 46.085 102.105 46.175 ;
        RECT 93.585 46.075 102.105 46.085 ;
        RECT 93.585 45.855 95.585 46.075 ;
        RECT 98.105 45.945 102.105 46.075 ;
        RECT 93.195 44.425 93.425 45.805 ;
        RECT 95.745 44.425 95.975 45.805 ;
        RECT 93.195 43.470 95.975 44.425 ;
        RECT 93.195 41.845 93.425 43.470 ;
        RECT 95.745 41.845 95.975 43.470 ;
        RECT 97.670 44.640 97.900 45.895 ;
        RECT 99.340 44.640 100.725 45.945 ;
        RECT 102.310 44.640 102.540 45.895 ;
        RECT 102.905 45.435 107.580 47.115 ;
        RECT 104.265 45.095 104.540 45.125 ;
        RECT 104.250 44.840 104.580 45.095 ;
        RECT 104.265 44.820 104.555 44.840 ;
        RECT 104.265 44.790 104.540 44.820 ;
        RECT 97.670 44.570 102.540 44.640 ;
        RECT 104.075 44.570 104.305 44.615 ;
        RECT 97.670 43.295 102.545 44.570 ;
        RECT 97.670 41.935 97.900 43.295 ;
        RECT 102.310 41.935 102.545 43.295 ;
        RECT 93.585 41.565 95.585 41.795 ;
        RECT 93.650 41.390 95.520 41.565 ;
        RECT 92.000 40.835 95.520 41.390 ;
        RECT 92.000 35.730 92.875 40.835 ;
        RECT 93.650 40.655 95.520 40.835 ;
        RECT 93.585 40.425 95.585 40.655 ;
        RECT 97.710 40.465 97.870 41.935 ;
        RECT 102.340 41.925 102.545 41.935 ;
        RECT 98.105 41.655 102.105 41.885 ;
        RECT 98.185 41.410 102.010 41.655 ;
        RECT 104.065 41.410 104.305 44.570 ;
        RECT 98.185 40.920 104.305 41.410 ;
        RECT 98.185 40.745 102.010 40.920 ;
        RECT 98.105 40.515 102.105 40.745 ;
        RECT 93.195 38.980 93.425 40.375 ;
        RECT 95.745 38.980 95.975 40.375 ;
        RECT 93.195 38.025 95.975 38.980 ;
        RECT 93.195 36.415 93.425 38.025 ;
        RECT 95.745 36.415 95.975 38.025 ;
        RECT 97.670 39.090 97.900 40.465 ;
        RECT 102.310 40.350 102.540 40.465 ;
        RECT 102.310 39.715 102.545 40.350 ;
        RECT 104.065 39.715 104.305 40.920 ;
        RECT 102.310 39.090 102.540 39.715 ;
        RECT 104.075 39.615 104.305 39.715 ;
        RECT 104.515 44.600 104.745 44.615 ;
        RECT 105.165 44.600 105.645 45.435 ;
        RECT 104.515 39.675 105.655 44.600 ;
        RECT 104.515 39.615 104.745 39.675 ;
        RECT 104.265 39.405 104.555 39.410 ;
        RECT 104.250 39.150 104.580 39.405 ;
        RECT 97.670 37.745 102.540 39.090 ;
        RECT 97.670 36.505 97.900 37.745 ;
        RECT 102.310 36.505 102.540 37.745 ;
        RECT 93.585 36.340 95.585 36.365 ;
        RECT 98.105 36.340 102.105 36.455 ;
        RECT 93.585 36.265 95.590 36.340 ;
        RECT 96.125 36.265 102.105 36.340 ;
        RECT 93.585 36.225 102.105 36.265 ;
        RECT 93.585 36.135 102.040 36.225 ;
        RECT 93.640 36.000 102.040 36.135 ;
        RECT 92.000 35.290 93.860 35.730 ;
        RECT 92.000 35.280 94.850 35.290 ;
        RECT 92.000 34.935 95.520 35.280 ;
        RECT 92.000 33.310 93.860 34.935 ;
        RECT 94.660 34.785 95.520 34.935 ;
        RECT 94.155 34.595 94.405 34.610 ;
        RECT 94.155 34.305 94.430 34.595 ;
        RECT 94.590 34.555 95.590 34.785 ;
        RECT 96.010 34.690 96.280 36.000 ;
        RECT 106.880 35.570 107.580 45.435 ;
        RECT 101.300 35.235 107.580 35.570 ;
        RECT 98.185 35.095 107.580 35.235 ;
        RECT 98.185 34.870 102.045 35.095 ;
        RECT 94.155 34.275 94.405 34.305 ;
        RECT 94.590 34.115 95.590 34.345 ;
        RECT 95.735 34.270 97.925 34.690 ;
        RECT 98.120 34.640 102.120 34.870 ;
        RECT 102.355 34.680 102.605 34.700 ;
        RECT 98.120 34.200 102.120 34.430 ;
        RECT 102.325 34.390 102.605 34.680 ;
        RECT 102.355 34.365 102.605 34.390 ;
        RECT 94.660 33.975 95.545 34.115 ;
        RECT 98.170 34.035 102.095 34.200 ;
        RECT 95.730 33.975 102.095 34.035 ;
        RECT 94.660 33.920 102.095 33.975 ;
        RECT 94.660 33.850 98.540 33.920 ;
        RECT 95.215 33.735 98.540 33.850 ;
        RECT 106.880 33.770 107.580 35.095 ;
        RECT 92.000 33.265 94.385 33.310 ;
        RECT 89.920 31.675 90.395 31.690 ;
        RECT 76.665 31.560 81.730 31.630 ;
        RECT 78.205 31.555 81.730 31.560 ;
        RECT 53.425 31.415 53.715 31.460 ;
        RECT 53.870 31.400 54.190 31.460 ;
        RECT 63.290 31.340 63.610 31.380 ;
        RECT 79.415 31.340 80.415 31.555 ;
        RECT 92.000 31.535 92.875 33.265 ;
        RECT 93.240 32.990 94.385 33.265 ;
        RECT 96.570 33.105 96.975 33.735 ;
        RECT 105.575 33.235 107.580 33.770 ;
        RECT 93.240 32.925 95.490 32.990 ;
        RECT 93.680 32.760 95.490 32.925 ;
        RECT 93.165 32.570 93.415 32.595 ;
        RECT 93.165 32.280 93.435 32.570 ;
        RECT 93.595 32.530 95.595 32.760 ;
        RECT 96.555 32.740 96.980 33.105 ;
        RECT 98.220 33.090 107.580 33.235 ;
        RECT 98.220 32.845 106.075 33.090 ;
        RECT 93.165 32.260 93.415 32.280 ;
        RECT 93.595 32.090 95.595 32.320 ;
        RECT 95.745 32.230 97.935 32.740 ;
        RECT 98.125 32.615 106.125 32.845 ;
        RECT 106.355 32.655 106.605 32.670 ;
        RECT 95.745 32.225 96.445 32.230 ;
        RECT 97.445 32.225 97.935 32.230 ;
        RECT 98.125 32.175 106.125 32.405 ;
        RECT 106.330 32.365 106.605 32.655 ;
        RECT 106.355 32.335 106.605 32.365 ;
        RECT 93.665 31.925 95.530 32.090 ;
        RECT 96.415 31.925 97.415 32.000 ;
        RECT 98.200 31.925 106.050 32.175 ;
        RECT 93.665 31.630 106.050 31.925 ;
        RECT 106.880 31.690 107.580 33.090 ;
        RECT 93.665 31.560 98.730 31.630 ;
        RECT 106.960 31.580 107.580 31.690 ;
        RECT 109.000 58.025 109.875 58.140 ;
        RECT 109.000 57.665 115.445 58.025 ;
        RECT 109.000 57.530 122.975 57.665 ;
        RECT 109.000 57.085 109.875 57.530 ;
        RECT 115.015 57.435 122.975 57.530 ;
        RECT 109.000 56.860 109.885 57.085 ;
        RECT 110.595 57.000 111.815 57.085 ;
        RECT 110.595 56.945 111.830 57.000 ;
        RECT 109.000 52.185 109.875 56.860 ;
        RECT 110.585 56.715 112.585 56.945 ;
        RECT 110.195 55.465 110.425 56.665 ;
        RECT 110.970 55.465 112.135 56.715 ;
        RECT 112.745 55.465 112.975 56.665 ;
        RECT 110.195 54.675 112.975 55.465 ;
        RECT 114.735 56.510 114.965 57.230 ;
        RECT 114.735 56.485 115.100 56.510 ;
        RECT 115.260 56.485 115.580 56.540 ;
        RECT 114.735 56.335 115.580 56.485 ;
        RECT 114.735 56.305 115.100 56.335 ;
        RECT 114.735 55.230 114.965 56.305 ;
        RECT 115.260 56.280 115.580 56.335 ;
        RECT 117.865 55.055 119.680 57.435 ;
        RECT 123.025 57.195 123.255 57.230 ;
        RECT 123.880 57.195 124.580 58.165 ;
        RECT 123.025 55.285 124.580 57.195 ;
        RECT 123.025 55.230 123.255 55.285 ;
        RECT 115.265 55.025 122.895 55.055 ;
        RECT 115.015 54.795 122.975 55.025 ;
        RECT 110.195 52.705 110.425 54.675 ;
        RECT 112.745 54.005 112.975 54.675 ;
        RECT 112.745 53.725 115.610 54.005 ;
        RECT 112.745 53.635 123.030 53.725 ;
        RECT 112.745 52.705 112.975 53.635 ;
        RECT 115.170 53.485 123.030 53.635 ;
        RECT 115.110 53.255 123.110 53.485 ;
        RECT 114.675 52.765 114.905 53.205 ;
        RECT 123.315 53.195 123.545 53.205 ;
        RECT 115.395 52.765 116.395 52.835 ;
        RECT 123.315 52.765 123.550 53.195 ;
        RECT 110.585 52.425 112.585 52.655 ;
        RECT 110.675 52.185 112.500 52.425 ;
        RECT 109.000 51.695 112.500 52.185 ;
        RECT 109.000 46.860 109.875 51.695 ;
        RECT 110.675 51.515 112.500 51.695 ;
        RECT 114.675 51.875 123.550 52.765 ;
        RECT 110.585 51.285 112.585 51.515 ;
        RECT 114.675 51.245 114.905 51.875 ;
        RECT 115.395 51.820 116.395 51.875 ;
        RECT 123.315 51.310 123.550 51.875 ;
        RECT 123.315 51.245 123.545 51.310 ;
        RECT 110.195 49.800 110.425 51.235 ;
        RECT 112.745 49.800 112.975 51.235 ;
        RECT 115.110 50.965 123.110 51.195 ;
        RECT 115.180 50.840 123.010 50.965 ;
        RECT 115.200 50.055 123.000 50.840 ;
        RECT 115.110 49.825 123.110 50.055 ;
        RECT 110.195 48.460 112.975 49.800 ;
        RECT 114.675 49.750 114.905 49.775 ;
        RECT 110.195 47.275 110.425 48.460 ;
        RECT 110.770 47.225 112.365 48.460 ;
        RECT 112.745 47.570 112.975 48.460 ;
        RECT 114.670 49.305 114.905 49.750 ;
        RECT 123.315 49.750 123.545 49.775 ;
        RECT 114.670 49.295 115.085 49.305 ;
        RECT 115.225 49.295 116.225 49.365 ;
        RECT 114.670 49.290 116.225 49.295 ;
        RECT 116.635 49.290 118.255 49.295 ;
        RECT 123.315 49.290 123.550 49.750 ;
        RECT 114.670 48.400 123.550 49.290 ;
        RECT 114.670 48.385 116.225 48.400 ;
        RECT 116.635 48.395 118.255 48.400 ;
        RECT 114.670 48.295 115.085 48.385 ;
        RECT 115.225 48.335 116.225 48.385 ;
        RECT 114.670 47.865 114.905 48.295 ;
        RECT 114.675 47.815 114.905 47.865 ;
        RECT 123.315 47.865 123.550 48.400 ;
        RECT 123.315 47.815 123.545 47.865 ;
        RECT 115.110 47.570 123.110 47.765 ;
        RECT 112.745 47.535 123.110 47.570 ;
        RECT 112.745 47.390 123.030 47.535 ;
        RECT 112.745 47.375 115.245 47.390 ;
        RECT 112.745 47.275 112.975 47.375 ;
        RECT 110.585 46.995 112.585 47.225 ;
        RECT 123.880 47.115 124.580 55.285 ;
        RECT 118.955 46.985 119.230 47.055 ;
        RECT 113.260 46.860 119.230 46.985 ;
        RECT 109.000 46.845 110.405 46.860 ;
        RECT 112.750 46.845 119.230 46.860 ;
        RECT 109.000 46.795 119.230 46.845 ;
        RECT 109.000 46.670 113.450 46.795 ;
        RECT 118.955 46.720 119.230 46.795 ;
        RECT 109.000 41.390 109.875 46.670 ;
        RECT 111.825 46.365 115.610 46.370 ;
        RECT 111.825 46.300 119.060 46.365 ;
        RECT 110.645 46.175 119.060 46.300 ;
        RECT 110.645 46.085 119.105 46.175 ;
        RECT 110.585 46.075 119.105 46.085 ;
        RECT 110.585 45.855 112.585 46.075 ;
        RECT 115.105 45.945 119.105 46.075 ;
        RECT 110.195 44.425 110.425 45.805 ;
        RECT 112.745 44.425 112.975 45.805 ;
        RECT 110.195 43.470 112.975 44.425 ;
        RECT 110.195 41.845 110.425 43.470 ;
        RECT 112.745 41.845 112.975 43.470 ;
        RECT 114.670 44.640 114.900 45.895 ;
        RECT 116.340 44.640 117.725 45.945 ;
        RECT 119.310 44.640 119.540 45.895 ;
        RECT 119.905 45.435 124.580 47.115 ;
        RECT 121.265 45.095 121.540 45.125 ;
        RECT 121.250 44.840 121.580 45.095 ;
        RECT 121.265 44.820 121.555 44.840 ;
        RECT 121.265 44.790 121.540 44.820 ;
        RECT 114.670 44.570 119.540 44.640 ;
        RECT 121.075 44.570 121.305 44.615 ;
        RECT 114.670 43.295 119.545 44.570 ;
        RECT 114.670 41.935 114.900 43.295 ;
        RECT 119.310 41.935 119.545 43.295 ;
        RECT 110.585 41.565 112.585 41.795 ;
        RECT 110.650 41.390 112.520 41.565 ;
        RECT 109.000 40.835 112.520 41.390 ;
        RECT 109.000 35.730 109.875 40.835 ;
        RECT 110.650 40.655 112.520 40.835 ;
        RECT 110.585 40.425 112.585 40.655 ;
        RECT 114.710 40.465 114.870 41.935 ;
        RECT 119.340 41.925 119.545 41.935 ;
        RECT 115.105 41.655 119.105 41.885 ;
        RECT 115.185 41.410 119.010 41.655 ;
        RECT 121.065 41.410 121.305 44.570 ;
        RECT 115.185 40.920 121.305 41.410 ;
        RECT 115.185 40.745 119.010 40.920 ;
        RECT 115.105 40.515 119.105 40.745 ;
        RECT 110.195 38.980 110.425 40.375 ;
        RECT 112.745 38.980 112.975 40.375 ;
        RECT 110.195 38.025 112.975 38.980 ;
        RECT 110.195 36.415 110.425 38.025 ;
        RECT 112.745 36.415 112.975 38.025 ;
        RECT 114.670 39.090 114.900 40.465 ;
        RECT 119.310 40.350 119.540 40.465 ;
        RECT 119.310 39.715 119.545 40.350 ;
        RECT 121.065 39.715 121.305 40.920 ;
        RECT 119.310 39.090 119.540 39.715 ;
        RECT 121.075 39.615 121.305 39.715 ;
        RECT 121.515 44.600 121.745 44.615 ;
        RECT 122.165 44.600 122.645 45.435 ;
        RECT 121.515 39.675 122.655 44.600 ;
        RECT 121.515 39.615 121.745 39.675 ;
        RECT 121.265 39.405 121.555 39.410 ;
        RECT 121.250 39.150 121.580 39.405 ;
        RECT 114.670 37.745 119.540 39.090 ;
        RECT 114.670 36.505 114.900 37.745 ;
        RECT 119.310 36.505 119.540 37.745 ;
        RECT 110.585 36.340 112.585 36.365 ;
        RECT 115.105 36.340 119.105 36.455 ;
        RECT 110.585 36.265 112.590 36.340 ;
        RECT 113.125 36.265 119.105 36.340 ;
        RECT 110.585 36.225 119.105 36.265 ;
        RECT 110.585 36.135 119.040 36.225 ;
        RECT 110.640 36.000 119.040 36.135 ;
        RECT 109.000 35.290 110.860 35.730 ;
        RECT 109.000 35.280 111.850 35.290 ;
        RECT 109.000 34.935 112.520 35.280 ;
        RECT 109.000 33.310 110.860 34.935 ;
        RECT 111.660 34.785 112.520 34.935 ;
        RECT 111.155 34.595 111.405 34.610 ;
        RECT 111.155 34.305 111.430 34.595 ;
        RECT 111.590 34.555 112.590 34.785 ;
        RECT 113.010 34.690 113.280 36.000 ;
        RECT 123.880 35.570 124.580 45.435 ;
        RECT 118.300 35.235 124.580 35.570 ;
        RECT 115.185 35.095 124.580 35.235 ;
        RECT 115.185 34.870 119.045 35.095 ;
        RECT 111.155 34.275 111.405 34.305 ;
        RECT 111.590 34.115 112.590 34.345 ;
        RECT 112.735 34.270 114.925 34.690 ;
        RECT 115.120 34.640 119.120 34.870 ;
        RECT 119.355 34.680 119.605 34.700 ;
        RECT 115.120 34.200 119.120 34.430 ;
        RECT 119.325 34.390 119.605 34.680 ;
        RECT 119.355 34.365 119.605 34.390 ;
        RECT 111.660 33.975 112.545 34.115 ;
        RECT 115.170 34.035 119.095 34.200 ;
        RECT 112.730 33.975 119.095 34.035 ;
        RECT 111.660 33.920 119.095 33.975 ;
        RECT 111.660 33.850 115.540 33.920 ;
        RECT 112.215 33.735 115.540 33.850 ;
        RECT 123.880 33.770 124.580 35.095 ;
        RECT 109.000 33.265 111.385 33.310 ;
        RECT 95.205 31.555 98.730 31.560 ;
        RECT 26.730 31.260 27.020 31.305 ;
        RECT 28.300 31.260 28.590 31.305 ;
        RECT 30.400 31.260 30.690 31.305 ;
        RECT 26.730 31.120 30.690 31.260 ;
        RECT 26.730 31.075 27.020 31.120 ;
        RECT 28.300 31.075 28.590 31.120 ;
        RECT 30.400 31.075 30.690 31.120 ;
        RECT 47.445 31.260 47.735 31.305 ;
        RECT 52.950 31.260 53.270 31.320 ;
        RECT 47.445 31.120 53.270 31.260 ;
        RECT 47.445 31.075 47.735 31.120 ;
        RECT 52.950 31.060 53.270 31.120 ;
        RECT 62.605 31.040 62.865 31.220 ;
        RECT 63.290 31.160 80.415 31.340 ;
        RECT 63.290 31.120 63.610 31.160 ;
        RECT 26.295 30.920 26.585 30.965 ;
        RECT 28.815 30.920 29.105 30.965 ;
        RECT 30.005 30.920 30.295 30.965 ;
        RECT 26.295 30.780 30.295 30.920 ;
        RECT 26.295 30.735 26.585 30.780 ;
        RECT 28.815 30.735 29.105 30.780 ;
        RECT 30.005 30.735 30.295 30.780 ;
        RECT 30.870 30.720 31.190 30.980 ;
        RECT 56.170 30.920 56.490 30.980 ;
        RECT 46.600 30.780 56.490 30.920 ;
        RECT 62.605 30.900 62.880 31.040 ;
        RECT 79.415 31.000 80.415 31.160 ;
        RECT 96.415 31.000 97.415 31.555 ;
        RECT 109.000 31.535 109.875 33.265 ;
        RECT 110.240 32.990 111.385 33.265 ;
        RECT 113.570 33.105 113.975 33.735 ;
        RECT 122.575 33.235 124.580 33.770 ;
        RECT 110.240 32.925 112.490 32.990 ;
        RECT 110.680 32.760 112.490 32.925 ;
        RECT 110.165 32.570 110.415 32.595 ;
        RECT 110.165 32.280 110.435 32.570 ;
        RECT 110.595 32.530 112.595 32.760 ;
        RECT 113.555 32.740 113.980 33.105 ;
        RECT 115.220 33.090 124.580 33.235 ;
        RECT 115.220 32.845 123.075 33.090 ;
        RECT 110.165 32.260 110.415 32.280 ;
        RECT 110.595 32.090 112.595 32.320 ;
        RECT 112.745 32.230 114.935 32.740 ;
        RECT 115.125 32.615 123.125 32.845 ;
        RECT 123.355 32.655 123.605 32.670 ;
        RECT 112.745 32.225 113.445 32.230 ;
        RECT 114.445 32.225 114.935 32.230 ;
        RECT 115.125 32.175 123.125 32.405 ;
        RECT 123.330 32.365 123.605 32.655 ;
        RECT 123.355 32.335 123.605 32.365 ;
        RECT 110.665 31.925 112.530 32.090 ;
        RECT 113.415 31.925 114.415 32.000 ;
        RECT 115.200 31.925 123.050 32.175 ;
        RECT 110.665 31.630 123.050 31.925 ;
        RECT 123.880 31.690 124.580 33.090 ;
        RECT 126.000 58.025 126.875 58.140 ;
        RECT 126.000 57.665 132.445 58.025 ;
        RECT 126.000 57.530 139.975 57.665 ;
        RECT 126.000 57.085 126.875 57.530 ;
        RECT 132.015 57.435 139.975 57.530 ;
        RECT 126.000 56.860 126.885 57.085 ;
        RECT 127.595 57.000 128.815 57.085 ;
        RECT 127.595 56.945 128.830 57.000 ;
        RECT 126.000 52.185 126.875 56.860 ;
        RECT 127.585 56.715 129.585 56.945 ;
        RECT 127.195 55.465 127.425 56.665 ;
        RECT 127.970 55.465 129.135 56.715 ;
        RECT 129.745 55.465 129.975 56.665 ;
        RECT 127.195 54.675 129.975 55.465 ;
        RECT 131.735 56.510 131.965 57.230 ;
        RECT 131.735 56.485 132.100 56.510 ;
        RECT 132.260 56.485 132.580 56.540 ;
        RECT 131.735 56.335 132.580 56.485 ;
        RECT 131.735 56.305 132.100 56.335 ;
        RECT 131.735 55.230 131.965 56.305 ;
        RECT 132.260 56.280 132.580 56.335 ;
        RECT 134.865 55.055 136.680 57.435 ;
        RECT 140.025 57.195 140.255 57.230 ;
        RECT 140.880 57.195 141.580 58.165 ;
        RECT 140.025 55.285 141.580 57.195 ;
        RECT 140.025 55.230 140.255 55.285 ;
        RECT 132.265 55.025 139.895 55.055 ;
        RECT 132.015 54.795 139.975 55.025 ;
        RECT 127.195 52.705 127.425 54.675 ;
        RECT 129.745 54.005 129.975 54.675 ;
        RECT 129.745 53.725 132.610 54.005 ;
        RECT 129.745 53.635 140.030 53.725 ;
        RECT 129.745 52.705 129.975 53.635 ;
        RECT 132.170 53.485 140.030 53.635 ;
        RECT 132.110 53.255 140.110 53.485 ;
        RECT 131.675 52.765 131.905 53.205 ;
        RECT 140.315 53.195 140.545 53.205 ;
        RECT 132.395 52.765 133.395 52.835 ;
        RECT 140.315 52.765 140.550 53.195 ;
        RECT 127.585 52.425 129.585 52.655 ;
        RECT 127.675 52.185 129.500 52.425 ;
        RECT 126.000 51.695 129.500 52.185 ;
        RECT 126.000 46.860 126.875 51.695 ;
        RECT 127.675 51.515 129.500 51.695 ;
        RECT 131.675 51.875 140.550 52.765 ;
        RECT 127.585 51.285 129.585 51.515 ;
        RECT 131.675 51.245 131.905 51.875 ;
        RECT 132.395 51.820 133.395 51.875 ;
        RECT 140.315 51.310 140.550 51.875 ;
        RECT 140.315 51.245 140.545 51.310 ;
        RECT 127.195 49.800 127.425 51.235 ;
        RECT 129.745 49.800 129.975 51.235 ;
        RECT 132.110 50.965 140.110 51.195 ;
        RECT 132.180 50.840 140.010 50.965 ;
        RECT 132.200 50.055 140.000 50.840 ;
        RECT 132.110 49.825 140.110 50.055 ;
        RECT 127.195 48.460 129.975 49.800 ;
        RECT 131.675 49.750 131.905 49.775 ;
        RECT 127.195 47.275 127.425 48.460 ;
        RECT 127.770 47.225 129.365 48.460 ;
        RECT 129.745 47.570 129.975 48.460 ;
        RECT 131.670 49.305 131.905 49.750 ;
        RECT 140.315 49.750 140.545 49.775 ;
        RECT 131.670 49.295 132.085 49.305 ;
        RECT 132.225 49.295 133.225 49.365 ;
        RECT 131.670 49.290 133.225 49.295 ;
        RECT 133.635 49.290 135.255 49.295 ;
        RECT 140.315 49.290 140.550 49.750 ;
        RECT 131.670 48.400 140.550 49.290 ;
        RECT 131.670 48.385 133.225 48.400 ;
        RECT 133.635 48.395 135.255 48.400 ;
        RECT 131.670 48.295 132.085 48.385 ;
        RECT 132.225 48.335 133.225 48.385 ;
        RECT 131.670 47.865 131.905 48.295 ;
        RECT 131.675 47.815 131.905 47.865 ;
        RECT 140.315 47.865 140.550 48.400 ;
        RECT 140.315 47.815 140.545 47.865 ;
        RECT 132.110 47.570 140.110 47.765 ;
        RECT 129.745 47.535 140.110 47.570 ;
        RECT 129.745 47.390 140.030 47.535 ;
        RECT 129.745 47.375 132.245 47.390 ;
        RECT 129.745 47.275 129.975 47.375 ;
        RECT 127.585 46.995 129.585 47.225 ;
        RECT 140.880 47.115 141.580 55.285 ;
        RECT 135.955 46.985 136.230 47.055 ;
        RECT 130.260 46.860 136.230 46.985 ;
        RECT 126.000 46.845 127.405 46.860 ;
        RECT 129.750 46.845 136.230 46.860 ;
        RECT 126.000 46.795 136.230 46.845 ;
        RECT 126.000 46.670 130.450 46.795 ;
        RECT 135.955 46.720 136.230 46.795 ;
        RECT 126.000 41.390 126.875 46.670 ;
        RECT 128.825 46.365 132.610 46.370 ;
        RECT 128.825 46.300 136.060 46.365 ;
        RECT 127.645 46.175 136.060 46.300 ;
        RECT 127.645 46.085 136.105 46.175 ;
        RECT 127.585 46.075 136.105 46.085 ;
        RECT 127.585 45.855 129.585 46.075 ;
        RECT 132.105 45.945 136.105 46.075 ;
        RECT 127.195 44.425 127.425 45.805 ;
        RECT 129.745 44.425 129.975 45.805 ;
        RECT 127.195 43.470 129.975 44.425 ;
        RECT 127.195 41.845 127.425 43.470 ;
        RECT 129.745 41.845 129.975 43.470 ;
        RECT 131.670 44.640 131.900 45.895 ;
        RECT 133.340 44.640 134.725 45.945 ;
        RECT 136.310 44.640 136.540 45.895 ;
        RECT 136.905 45.435 141.580 47.115 ;
        RECT 138.265 45.095 138.540 45.125 ;
        RECT 138.250 44.840 138.580 45.095 ;
        RECT 138.265 44.820 138.555 44.840 ;
        RECT 138.265 44.790 138.540 44.820 ;
        RECT 131.670 44.570 136.540 44.640 ;
        RECT 138.075 44.570 138.305 44.615 ;
        RECT 131.670 43.295 136.545 44.570 ;
        RECT 131.670 41.935 131.900 43.295 ;
        RECT 136.310 41.935 136.545 43.295 ;
        RECT 127.585 41.565 129.585 41.795 ;
        RECT 127.650 41.390 129.520 41.565 ;
        RECT 126.000 40.835 129.520 41.390 ;
        RECT 126.000 35.730 126.875 40.835 ;
        RECT 127.650 40.655 129.520 40.835 ;
        RECT 127.585 40.425 129.585 40.655 ;
        RECT 131.710 40.465 131.870 41.935 ;
        RECT 136.340 41.925 136.545 41.935 ;
        RECT 132.105 41.655 136.105 41.885 ;
        RECT 132.185 41.410 136.010 41.655 ;
        RECT 138.065 41.410 138.305 44.570 ;
        RECT 132.185 40.920 138.305 41.410 ;
        RECT 132.185 40.745 136.010 40.920 ;
        RECT 132.105 40.515 136.105 40.745 ;
        RECT 127.195 38.980 127.425 40.375 ;
        RECT 129.745 38.980 129.975 40.375 ;
        RECT 127.195 38.025 129.975 38.980 ;
        RECT 127.195 36.415 127.425 38.025 ;
        RECT 129.745 36.415 129.975 38.025 ;
        RECT 131.670 39.090 131.900 40.465 ;
        RECT 136.310 40.350 136.540 40.465 ;
        RECT 136.310 39.715 136.545 40.350 ;
        RECT 138.065 39.715 138.305 40.920 ;
        RECT 136.310 39.090 136.540 39.715 ;
        RECT 138.075 39.615 138.305 39.715 ;
        RECT 138.515 44.600 138.745 44.615 ;
        RECT 139.165 44.600 139.645 45.435 ;
        RECT 138.515 39.675 139.655 44.600 ;
        RECT 138.515 39.615 138.745 39.675 ;
        RECT 138.265 39.405 138.555 39.410 ;
        RECT 138.250 39.150 138.580 39.405 ;
        RECT 131.670 37.745 136.540 39.090 ;
        RECT 131.670 36.505 131.900 37.745 ;
        RECT 136.310 36.505 136.540 37.745 ;
        RECT 127.585 36.340 129.585 36.365 ;
        RECT 132.105 36.340 136.105 36.455 ;
        RECT 127.585 36.265 129.590 36.340 ;
        RECT 130.125 36.265 136.105 36.340 ;
        RECT 127.585 36.225 136.105 36.265 ;
        RECT 127.585 36.135 136.040 36.225 ;
        RECT 127.640 36.000 136.040 36.135 ;
        RECT 126.000 35.290 127.860 35.730 ;
        RECT 126.000 35.280 128.850 35.290 ;
        RECT 126.000 34.935 129.520 35.280 ;
        RECT 126.000 33.310 127.860 34.935 ;
        RECT 128.660 34.785 129.520 34.935 ;
        RECT 128.155 34.595 128.405 34.610 ;
        RECT 128.155 34.305 128.430 34.595 ;
        RECT 128.590 34.555 129.590 34.785 ;
        RECT 130.010 34.690 130.280 36.000 ;
        RECT 140.880 35.570 141.580 45.435 ;
        RECT 135.300 35.235 141.580 35.570 ;
        RECT 132.185 35.095 141.580 35.235 ;
        RECT 132.185 34.870 136.045 35.095 ;
        RECT 128.155 34.275 128.405 34.305 ;
        RECT 128.590 34.115 129.590 34.345 ;
        RECT 129.735 34.270 131.925 34.690 ;
        RECT 132.120 34.640 136.120 34.870 ;
        RECT 136.355 34.680 136.605 34.700 ;
        RECT 132.120 34.200 136.120 34.430 ;
        RECT 136.325 34.390 136.605 34.680 ;
        RECT 136.355 34.365 136.605 34.390 ;
        RECT 128.660 33.975 129.545 34.115 ;
        RECT 132.170 34.035 136.095 34.200 ;
        RECT 129.730 33.975 136.095 34.035 ;
        RECT 128.660 33.920 136.095 33.975 ;
        RECT 128.660 33.850 132.540 33.920 ;
        RECT 129.215 33.735 132.540 33.850 ;
        RECT 140.880 33.770 141.580 35.095 ;
        RECT 126.000 33.265 128.385 33.310 ;
        RECT 110.665 31.560 115.730 31.630 ;
        RECT 112.205 31.555 115.730 31.560 ;
        RECT 113.415 31.000 114.415 31.555 ;
        RECT 126.000 31.535 126.875 33.265 ;
        RECT 127.240 32.990 128.385 33.265 ;
        RECT 130.570 33.105 130.975 33.735 ;
        RECT 139.575 33.235 141.580 33.770 ;
        RECT 127.240 32.925 129.490 32.990 ;
        RECT 127.680 32.760 129.490 32.925 ;
        RECT 127.165 32.570 127.415 32.595 ;
        RECT 127.165 32.280 127.435 32.570 ;
        RECT 127.595 32.530 129.595 32.760 ;
        RECT 130.555 32.740 130.980 33.105 ;
        RECT 132.220 33.090 141.580 33.235 ;
        RECT 132.220 32.845 140.075 33.090 ;
        RECT 127.165 32.260 127.415 32.280 ;
        RECT 127.595 32.090 129.595 32.320 ;
        RECT 129.745 32.230 131.935 32.740 ;
        RECT 132.125 32.615 140.125 32.845 ;
        RECT 140.355 32.655 140.605 32.670 ;
        RECT 129.745 32.225 130.445 32.230 ;
        RECT 131.445 32.225 131.935 32.230 ;
        RECT 132.125 32.175 140.125 32.405 ;
        RECT 140.330 32.365 140.605 32.655 ;
        RECT 140.355 32.335 140.605 32.365 ;
        RECT 127.665 31.925 129.530 32.090 ;
        RECT 130.415 31.925 131.415 32.000 ;
        RECT 132.200 31.925 140.050 32.175 ;
        RECT 127.665 31.630 140.050 31.925 ;
        RECT 140.880 31.690 141.580 33.090 ;
        RECT 143.000 58.025 143.875 58.140 ;
        RECT 143.000 57.665 149.445 58.025 ;
        RECT 143.000 57.530 156.975 57.665 ;
        RECT 143.000 57.085 143.875 57.530 ;
        RECT 149.015 57.435 156.975 57.530 ;
        RECT 143.000 56.860 143.885 57.085 ;
        RECT 144.595 57.000 145.815 57.085 ;
        RECT 144.595 56.945 145.830 57.000 ;
        RECT 143.000 52.185 143.875 56.860 ;
        RECT 144.585 56.715 146.585 56.945 ;
        RECT 144.195 55.465 144.425 56.665 ;
        RECT 144.970 55.465 146.135 56.715 ;
        RECT 146.745 55.465 146.975 56.665 ;
        RECT 144.195 54.675 146.975 55.465 ;
        RECT 148.735 56.510 148.965 57.230 ;
        RECT 148.735 56.485 149.100 56.510 ;
        RECT 149.260 56.485 149.580 56.540 ;
        RECT 148.735 56.335 149.580 56.485 ;
        RECT 148.735 56.305 149.100 56.335 ;
        RECT 148.735 55.230 148.965 56.305 ;
        RECT 149.260 56.280 149.580 56.335 ;
        RECT 151.865 55.055 153.680 57.435 ;
        RECT 157.025 57.195 157.255 57.230 ;
        RECT 157.880 57.195 158.580 58.165 ;
        RECT 157.025 55.285 158.580 57.195 ;
        RECT 157.025 55.230 157.255 55.285 ;
        RECT 149.265 55.025 156.895 55.055 ;
        RECT 149.015 54.795 156.975 55.025 ;
        RECT 144.195 52.705 144.425 54.675 ;
        RECT 146.745 54.005 146.975 54.675 ;
        RECT 146.745 53.725 149.610 54.005 ;
        RECT 146.745 53.635 157.030 53.725 ;
        RECT 146.745 52.705 146.975 53.635 ;
        RECT 149.170 53.485 157.030 53.635 ;
        RECT 149.110 53.255 157.110 53.485 ;
        RECT 148.675 52.765 148.905 53.205 ;
        RECT 157.315 53.195 157.545 53.205 ;
        RECT 149.395 52.765 150.395 52.835 ;
        RECT 157.315 52.765 157.550 53.195 ;
        RECT 144.585 52.425 146.585 52.655 ;
        RECT 144.675 52.185 146.500 52.425 ;
        RECT 143.000 51.695 146.500 52.185 ;
        RECT 143.000 46.860 143.875 51.695 ;
        RECT 144.675 51.515 146.500 51.695 ;
        RECT 148.675 51.875 157.550 52.765 ;
        RECT 144.585 51.285 146.585 51.515 ;
        RECT 148.675 51.245 148.905 51.875 ;
        RECT 149.395 51.820 150.395 51.875 ;
        RECT 157.315 51.310 157.550 51.875 ;
        RECT 157.315 51.245 157.545 51.310 ;
        RECT 144.195 49.800 144.425 51.235 ;
        RECT 146.745 49.800 146.975 51.235 ;
        RECT 149.110 50.965 157.110 51.195 ;
        RECT 149.180 50.840 157.010 50.965 ;
        RECT 149.200 50.055 157.000 50.840 ;
        RECT 149.110 49.825 157.110 50.055 ;
        RECT 144.195 48.460 146.975 49.800 ;
        RECT 148.675 49.750 148.905 49.775 ;
        RECT 144.195 47.275 144.425 48.460 ;
        RECT 144.770 47.225 146.365 48.460 ;
        RECT 146.745 47.570 146.975 48.460 ;
        RECT 148.670 49.305 148.905 49.750 ;
        RECT 157.315 49.750 157.545 49.775 ;
        RECT 148.670 49.295 149.085 49.305 ;
        RECT 149.225 49.295 150.225 49.365 ;
        RECT 148.670 49.290 150.225 49.295 ;
        RECT 150.635 49.290 152.255 49.295 ;
        RECT 157.315 49.290 157.550 49.750 ;
        RECT 148.670 48.400 157.550 49.290 ;
        RECT 148.670 48.385 150.225 48.400 ;
        RECT 150.635 48.395 152.255 48.400 ;
        RECT 148.670 48.295 149.085 48.385 ;
        RECT 149.225 48.335 150.225 48.385 ;
        RECT 148.670 47.865 148.905 48.295 ;
        RECT 148.675 47.815 148.905 47.865 ;
        RECT 157.315 47.865 157.550 48.400 ;
        RECT 157.315 47.815 157.545 47.865 ;
        RECT 149.110 47.570 157.110 47.765 ;
        RECT 146.745 47.535 157.110 47.570 ;
        RECT 146.745 47.390 157.030 47.535 ;
        RECT 146.745 47.375 149.245 47.390 ;
        RECT 146.745 47.275 146.975 47.375 ;
        RECT 144.585 46.995 146.585 47.225 ;
        RECT 157.880 47.115 158.580 55.285 ;
        RECT 152.955 46.985 153.230 47.055 ;
        RECT 147.260 46.860 153.230 46.985 ;
        RECT 143.000 46.845 144.405 46.860 ;
        RECT 146.750 46.845 153.230 46.860 ;
        RECT 143.000 46.795 153.230 46.845 ;
        RECT 143.000 46.670 147.450 46.795 ;
        RECT 152.955 46.720 153.230 46.795 ;
        RECT 143.000 41.390 143.875 46.670 ;
        RECT 145.825 46.365 149.610 46.370 ;
        RECT 145.825 46.300 153.060 46.365 ;
        RECT 144.645 46.175 153.060 46.300 ;
        RECT 144.645 46.085 153.105 46.175 ;
        RECT 144.585 46.075 153.105 46.085 ;
        RECT 144.585 45.855 146.585 46.075 ;
        RECT 149.105 45.945 153.105 46.075 ;
        RECT 144.195 44.425 144.425 45.805 ;
        RECT 146.745 44.425 146.975 45.805 ;
        RECT 144.195 43.470 146.975 44.425 ;
        RECT 144.195 41.845 144.425 43.470 ;
        RECT 146.745 41.845 146.975 43.470 ;
        RECT 148.670 44.640 148.900 45.895 ;
        RECT 150.340 44.640 151.725 45.945 ;
        RECT 153.310 44.640 153.540 45.895 ;
        RECT 153.905 45.435 158.580 47.115 ;
        RECT 155.265 45.095 155.540 45.125 ;
        RECT 155.250 44.840 155.580 45.095 ;
        RECT 155.265 44.820 155.555 44.840 ;
        RECT 155.265 44.790 155.540 44.820 ;
        RECT 148.670 44.570 153.540 44.640 ;
        RECT 155.075 44.570 155.305 44.615 ;
        RECT 148.670 43.295 153.545 44.570 ;
        RECT 148.670 41.935 148.900 43.295 ;
        RECT 153.310 41.935 153.545 43.295 ;
        RECT 144.585 41.565 146.585 41.795 ;
        RECT 144.650 41.390 146.520 41.565 ;
        RECT 143.000 40.835 146.520 41.390 ;
        RECT 143.000 35.730 143.875 40.835 ;
        RECT 144.650 40.655 146.520 40.835 ;
        RECT 144.585 40.425 146.585 40.655 ;
        RECT 148.710 40.465 148.870 41.935 ;
        RECT 153.340 41.925 153.545 41.935 ;
        RECT 149.105 41.655 153.105 41.885 ;
        RECT 149.185 41.410 153.010 41.655 ;
        RECT 155.065 41.410 155.305 44.570 ;
        RECT 149.185 40.920 155.305 41.410 ;
        RECT 149.185 40.745 153.010 40.920 ;
        RECT 149.105 40.515 153.105 40.745 ;
        RECT 144.195 38.980 144.425 40.375 ;
        RECT 146.745 38.980 146.975 40.375 ;
        RECT 144.195 38.025 146.975 38.980 ;
        RECT 144.195 36.415 144.425 38.025 ;
        RECT 146.745 36.415 146.975 38.025 ;
        RECT 148.670 39.090 148.900 40.465 ;
        RECT 153.310 40.350 153.540 40.465 ;
        RECT 153.310 39.715 153.545 40.350 ;
        RECT 155.065 39.715 155.305 40.920 ;
        RECT 153.310 39.090 153.540 39.715 ;
        RECT 155.075 39.615 155.305 39.715 ;
        RECT 155.515 44.600 155.745 44.615 ;
        RECT 156.165 44.600 156.645 45.435 ;
        RECT 155.515 39.675 156.655 44.600 ;
        RECT 155.515 39.615 155.745 39.675 ;
        RECT 155.265 39.405 155.555 39.410 ;
        RECT 155.250 39.150 155.580 39.405 ;
        RECT 148.670 37.745 153.540 39.090 ;
        RECT 148.670 36.505 148.900 37.745 ;
        RECT 153.310 36.505 153.540 37.745 ;
        RECT 144.585 36.340 146.585 36.365 ;
        RECT 149.105 36.340 153.105 36.455 ;
        RECT 144.585 36.265 146.590 36.340 ;
        RECT 147.125 36.265 153.105 36.340 ;
        RECT 144.585 36.225 153.105 36.265 ;
        RECT 144.585 36.135 153.040 36.225 ;
        RECT 144.640 36.000 153.040 36.135 ;
        RECT 143.000 35.290 144.860 35.730 ;
        RECT 143.000 35.280 145.850 35.290 ;
        RECT 143.000 34.935 146.520 35.280 ;
        RECT 143.000 33.310 144.860 34.935 ;
        RECT 145.660 34.785 146.520 34.935 ;
        RECT 145.155 34.595 145.405 34.610 ;
        RECT 145.155 34.305 145.430 34.595 ;
        RECT 145.590 34.555 146.590 34.785 ;
        RECT 147.010 34.690 147.280 36.000 ;
        RECT 157.880 35.570 158.580 45.435 ;
        RECT 152.300 35.235 158.580 35.570 ;
        RECT 149.185 35.095 158.580 35.235 ;
        RECT 149.185 34.870 153.045 35.095 ;
        RECT 145.155 34.275 145.405 34.305 ;
        RECT 145.590 34.115 146.590 34.345 ;
        RECT 146.735 34.270 148.925 34.690 ;
        RECT 149.120 34.640 153.120 34.870 ;
        RECT 153.355 34.680 153.605 34.700 ;
        RECT 149.120 34.200 153.120 34.430 ;
        RECT 153.325 34.390 153.605 34.680 ;
        RECT 153.355 34.365 153.605 34.390 ;
        RECT 145.660 33.975 146.545 34.115 ;
        RECT 149.170 34.035 153.095 34.200 ;
        RECT 146.730 33.975 153.095 34.035 ;
        RECT 145.660 33.920 153.095 33.975 ;
        RECT 145.660 33.850 149.540 33.920 ;
        RECT 146.215 33.735 149.540 33.850 ;
        RECT 157.880 33.770 158.580 35.095 ;
        RECT 143.000 33.265 145.385 33.310 ;
        RECT 127.665 31.560 132.730 31.630 ;
        RECT 129.205 31.555 132.730 31.560 ;
        RECT 130.415 31.000 131.415 31.555 ;
        RECT 143.000 31.535 143.875 33.265 ;
        RECT 144.240 32.990 145.385 33.265 ;
        RECT 147.570 33.105 147.975 33.735 ;
        RECT 156.575 33.235 158.580 33.770 ;
        RECT 144.240 32.925 146.490 32.990 ;
        RECT 144.680 32.760 146.490 32.925 ;
        RECT 144.165 32.570 144.415 32.595 ;
        RECT 144.165 32.280 144.435 32.570 ;
        RECT 144.595 32.530 146.595 32.760 ;
        RECT 147.555 32.740 147.980 33.105 ;
        RECT 149.220 33.090 158.580 33.235 ;
        RECT 149.220 32.845 157.075 33.090 ;
        RECT 144.165 32.260 144.415 32.280 ;
        RECT 144.595 32.090 146.595 32.320 ;
        RECT 146.745 32.230 148.935 32.740 ;
        RECT 149.125 32.615 157.125 32.845 ;
        RECT 157.355 32.655 157.605 32.670 ;
        RECT 146.745 32.225 147.445 32.230 ;
        RECT 148.445 32.225 148.935 32.230 ;
        RECT 149.125 32.175 157.125 32.405 ;
        RECT 157.330 32.365 157.605 32.655 ;
        RECT 157.355 32.335 157.605 32.365 ;
        RECT 144.665 31.925 146.530 32.090 ;
        RECT 147.415 31.925 148.415 32.000 ;
        RECT 149.200 31.925 157.050 32.175 ;
        RECT 144.665 31.630 157.050 31.925 ;
        RECT 157.880 31.690 158.580 33.090 ;
        RECT 144.665 31.560 149.730 31.630 ;
        RECT 146.205 31.555 149.730 31.560 ;
        RECT 143.085 31.395 143.705 31.535 ;
        RECT 147.415 31.000 148.415 31.555 ;
        RECT 35.945 30.580 36.235 30.625 ;
        RECT 40.530 30.580 40.850 30.640 ;
        RECT 46.600 30.625 46.740 30.780 ;
        RECT 56.170 30.720 56.490 30.780 ;
        RECT 62.650 30.855 62.880 30.900 ;
        RECT 96.835 30.855 97.000 31.000 ;
        RECT 62.650 30.690 97.000 30.855 ;
        RECT 35.945 30.440 40.850 30.580 ;
        RECT 35.945 30.395 36.235 30.440 ;
        RECT 40.530 30.380 40.850 30.440 ;
        RECT 46.525 30.395 46.815 30.625 ;
        RECT 47.890 30.380 48.210 30.640 ;
        RECT 49.270 30.380 49.590 30.640 ;
        RECT 50.650 30.380 50.970 30.640 ;
        RECT 52.045 30.395 52.335 30.625 ;
        RECT 52.965 30.580 53.255 30.625 ;
        RECT 53.410 30.580 53.730 30.640 ;
        RECT 52.965 30.440 53.730 30.580 ;
        RECT 52.965 30.395 53.255 30.440 ;
        RECT 26.730 30.240 27.050 30.300 ;
        RECT 29.550 30.240 29.840 30.285 ;
        RECT 52.120 30.240 52.260 30.395 ;
        RECT 53.410 30.380 53.730 30.440 ;
        RECT 54.330 30.380 54.650 30.640 ;
        RECT 55.710 30.380 56.030 30.640 ;
        RECT 56.630 30.380 56.950 30.640 ;
        RECT 61.950 30.565 62.270 30.580 ;
        RECT 113.800 30.565 114.030 31.000 ;
        RECT 61.950 30.550 62.490 30.565 ;
        RECT 98.090 30.550 114.030 30.565 ;
        RECT 54.420 30.240 54.560 30.380 ;
        RECT 61.950 30.335 114.030 30.550 ;
        RECT 61.950 30.320 62.270 30.335 ;
        RECT 26.730 30.100 29.840 30.240 ;
        RECT 26.730 30.040 27.050 30.100 ;
        RECT 29.550 30.055 29.840 30.100 ;
        RECT 48.900 30.100 54.560 30.240 ;
        RECT 48.900 29.945 49.040 30.100 ;
        RECT 61.055 30.085 61.375 30.095 ;
        RECT 130.795 30.085 131.040 31.000 ;
        RECT 48.825 29.715 49.115 29.945 ;
        RECT 51.585 29.900 51.875 29.945 ;
        RECT 52.030 29.900 52.350 29.960 ;
        RECT 51.585 29.760 52.350 29.900 ;
        RECT 51.585 29.715 51.875 29.760 ;
        RECT 52.030 29.700 52.350 29.760 ;
        RECT 52.490 29.700 52.810 29.960 ;
        RECT 61.055 29.840 131.040 30.085 ;
        RECT 61.055 29.835 61.375 29.840 ;
        RECT 60.270 29.635 60.590 29.650 ;
        RECT 147.800 29.635 148.030 31.000 ;
        RECT 22.520 29.080 58.400 29.560 ;
        RECT 60.270 29.405 148.030 29.635 ;
        RECT 60.270 29.390 60.590 29.405 ;
        RECT 75.000 29.025 75.875 29.140 ;
        RECT 26.730 28.680 27.050 28.940 ;
        RECT 28.570 28.680 28.890 28.940 ;
        RECT 29.030 28.680 29.350 28.940 ;
        RECT 31.330 28.880 31.650 28.940 ;
        RECT 33.630 28.880 33.950 28.940 ;
        RECT 35.945 28.880 36.235 28.925 ;
        RECT 31.330 28.740 36.235 28.880 ;
        RECT 31.330 28.680 31.650 28.740 ;
        RECT 33.630 28.680 33.950 28.740 ;
        RECT 35.945 28.695 36.235 28.740 ;
        RECT 40.070 28.680 40.390 28.940 ;
        RECT 45.590 28.680 45.910 28.940 ;
        RECT 55.250 28.880 55.570 28.940 ;
        RECT 55.725 28.880 56.015 28.925 ;
        RECT 55.250 28.740 56.015 28.880 ;
        RECT 55.250 28.680 55.570 28.740 ;
        RECT 55.725 28.695 56.015 28.740 ;
        RECT 23.970 28.200 24.290 28.260 ;
        RECT 25.365 28.200 25.655 28.245 ;
        RECT 23.970 28.060 25.655 28.200 ;
        RECT 40.160 28.200 40.300 28.680 ;
        RECT 75.000 28.665 81.445 29.025 ;
        RECT 40.990 28.540 41.310 28.600 ;
        RECT 40.990 28.400 43.060 28.540 ;
        RECT 40.990 28.340 41.310 28.400 ;
        RECT 42.920 28.245 43.060 28.400 ;
        RECT 75.000 28.530 88.975 28.665 ;
        RECT 41.510 28.200 41.800 28.245 ;
        RECT 40.160 28.060 41.800 28.200 ;
        RECT 23.970 28.000 24.290 28.060 ;
        RECT 25.365 28.015 25.655 28.060 ;
        RECT 41.510 28.015 41.800 28.060 ;
        RECT 42.845 28.015 43.135 28.245 ;
        RECT 45.145 28.200 45.435 28.245 ;
        RECT 48.825 28.200 49.115 28.245 ;
        RECT 45.145 28.060 49.115 28.200 ;
        RECT 45.145 28.015 45.435 28.060 ;
        RECT 48.825 28.015 49.115 28.060 ;
        RECT 52.490 28.200 52.810 28.260 ;
        RECT 54.805 28.200 55.095 28.245 ;
        RECT 52.490 28.060 55.095 28.200 ;
        RECT 52.490 28.000 52.810 28.060 ;
        RECT 54.805 28.015 55.095 28.060 ;
        RECT 75.000 28.085 75.875 28.530 ;
        RECT 81.015 28.435 88.975 28.530 ;
        RECT 29.965 27.860 30.255 27.905 ;
        RECT 35.470 27.860 35.790 27.920 ;
        RECT 29.965 27.720 35.790 27.860 ;
        RECT 29.965 27.675 30.255 27.720 ;
        RECT 35.470 27.660 35.790 27.720 ;
        RECT 38.255 27.860 38.545 27.905 ;
        RECT 40.775 27.860 41.065 27.905 ;
        RECT 41.965 27.860 42.255 27.905 ;
        RECT 38.255 27.720 42.255 27.860 ;
        RECT 38.255 27.675 38.545 27.720 ;
        RECT 40.775 27.675 41.065 27.720 ;
        RECT 41.965 27.675 42.255 27.720 ;
        RECT 46.510 27.660 46.830 27.920 ;
        RECT 46.970 27.860 47.290 27.920 ;
        RECT 51.585 27.860 51.875 27.905 ;
        RECT 46.970 27.720 51.875 27.860 ;
        RECT 46.970 27.660 47.290 27.720 ;
        RECT 51.585 27.675 51.875 27.720 ;
        RECT 52.030 27.860 52.350 27.920 ;
        RECT 53.425 27.860 53.715 27.905 ;
        RECT 52.030 27.720 53.715 27.860 ;
        RECT 52.030 27.660 52.350 27.720 ;
        RECT 53.425 27.675 53.715 27.720 ;
        RECT 53.885 27.860 54.175 27.905 ;
        RECT 56.630 27.860 56.950 27.920 ;
        RECT 53.885 27.720 56.950 27.860 ;
        RECT 53.885 27.675 54.175 27.720 ;
        RECT 56.630 27.660 56.950 27.720 ;
        RECT 75.000 27.860 75.885 28.085 ;
        RECT 76.595 28.000 77.815 28.085 ;
        RECT 76.595 27.945 77.830 28.000 ;
        RECT 21.210 27.520 21.530 27.580 ;
        RECT 24.445 27.520 24.735 27.565 ;
        RECT 21.210 27.380 24.735 27.520 ;
        RECT 21.210 27.320 21.530 27.380 ;
        RECT 24.445 27.335 24.735 27.380 ;
        RECT 38.690 27.520 38.980 27.565 ;
        RECT 40.260 27.520 40.550 27.565 ;
        RECT 42.360 27.520 42.650 27.565 ;
        RECT 38.690 27.380 42.650 27.520 ;
        RECT 38.690 27.335 38.980 27.380 ;
        RECT 40.260 27.335 40.550 27.380 ;
        RECT 42.360 27.335 42.650 27.380 ;
        RECT 40.990 27.180 41.310 27.240 ;
        RECT 43.305 27.180 43.595 27.225 ;
        RECT 40.990 27.040 43.595 27.180 ;
        RECT 40.990 26.980 41.310 27.040 ;
        RECT 43.305 26.995 43.595 27.040 ;
        RECT 22.520 26.360 58.400 26.840 ;
        RECT 43.750 26.160 44.070 26.220 ;
        RECT 37.860 26.020 44.070 26.160 ;
        RECT 33.630 24.940 33.950 25.200 ;
        RECT 37.860 25.185 38.000 26.020 ;
        RECT 43.750 25.960 44.070 26.020 ;
        RECT 51.585 26.160 51.875 26.205 ;
        RECT 53.410 26.160 53.730 26.220 ;
        RECT 51.585 26.020 53.730 26.160 ;
        RECT 51.585 25.975 51.875 26.020 ;
        RECT 53.410 25.960 53.730 26.020 ;
        RECT 55.710 26.160 56.030 26.220 ;
        RECT 56.185 26.160 56.475 26.205 ;
        RECT 55.710 26.020 56.475 26.160 ;
        RECT 55.710 25.960 56.030 26.020 ;
        RECT 56.185 25.975 56.475 26.020 ;
        RECT 38.730 25.820 39.020 25.865 ;
        RECT 40.830 25.820 41.120 25.865 ;
        RECT 42.400 25.820 42.690 25.865 ;
        RECT 38.730 25.680 42.690 25.820 ;
        RECT 38.730 25.635 39.020 25.680 ;
        RECT 40.830 25.635 41.120 25.680 ;
        RECT 42.400 25.635 42.690 25.680 ;
        RECT 45.145 25.820 45.435 25.865 ;
        RECT 46.970 25.820 47.290 25.880 ;
        RECT 45.145 25.680 47.290 25.820 ;
        RECT 45.145 25.635 45.435 25.680 ;
        RECT 46.970 25.620 47.290 25.680 ;
        RECT 52.950 25.820 53.270 25.880 ;
        RECT 55.265 25.820 55.555 25.865 ;
        RECT 52.950 25.680 55.555 25.820 ;
        RECT 52.950 25.620 53.270 25.680 ;
        RECT 55.265 25.635 55.555 25.680 ;
        RECT 39.125 25.480 39.415 25.525 ;
        RECT 40.315 25.480 40.605 25.525 ;
        RECT 42.835 25.480 43.125 25.525 ;
        RECT 39.125 25.340 43.125 25.480 ;
        RECT 39.125 25.295 39.415 25.340 ;
        RECT 40.315 25.295 40.605 25.340 ;
        RECT 42.835 25.295 43.125 25.340 ;
        RECT 52.030 25.480 52.350 25.540 ;
        RECT 53.885 25.480 54.175 25.525 ;
        RECT 52.030 25.340 54.175 25.480 ;
        RECT 52.030 25.280 52.350 25.340 ;
        RECT 53.885 25.295 54.175 25.340 ;
        RECT 37.785 24.955 38.075 25.185 ;
        RECT 38.245 25.140 38.535 25.185 ;
        RECT 38.690 25.140 39.010 25.200 ;
        RECT 38.245 25.000 39.010 25.140 ;
        RECT 38.245 24.955 38.535 25.000 ;
        RECT 38.690 24.940 39.010 25.000 ;
        RECT 46.970 24.940 47.290 25.200 ;
        RECT 49.730 24.940 50.050 25.200 ;
        RECT 52.490 24.940 52.810 25.200 ;
        RECT 39.580 24.800 39.870 24.845 ;
        RECT 40.990 24.800 41.310 24.860 ;
        RECT 39.580 24.660 41.310 24.800 ;
        RECT 39.580 24.615 39.870 24.660 ;
        RECT 40.990 24.600 41.310 24.660 ;
        RECT 43.380 24.660 46.280 24.800 ;
        RECT 43.380 24.520 43.520 24.660 ;
        RECT 34.565 24.460 34.855 24.505 ;
        RECT 36.390 24.460 36.710 24.520 ;
        RECT 34.565 24.320 36.710 24.460 ;
        RECT 34.565 24.275 34.855 24.320 ;
        RECT 36.390 24.260 36.710 24.320 ;
        RECT 36.865 24.460 37.155 24.505 ;
        RECT 39.150 24.460 39.470 24.520 ;
        RECT 36.865 24.320 39.470 24.460 ;
        RECT 36.865 24.275 37.155 24.320 ;
        RECT 39.150 24.260 39.470 24.320 ;
        RECT 43.290 24.260 43.610 24.520 ;
        RECT 46.140 24.505 46.280 24.660 ;
        RECT 46.065 24.275 46.355 24.505 ;
        RECT 49.270 24.460 49.590 24.520 ;
        RECT 50.665 24.460 50.955 24.505 ;
        RECT 49.270 24.320 50.955 24.460 ;
        RECT 49.270 24.260 49.590 24.320 ;
        RECT 50.665 24.275 50.955 24.320 ;
        RECT 22.520 23.640 58.400 24.120 ;
        RECT 37.235 23.105 37.495 23.195 ;
        RECT 35.695 23.060 37.495 23.105 ;
        RECT 35.635 22.965 37.495 23.060 ;
        RECT 35.635 22.740 35.895 22.965 ;
        RECT 37.235 22.875 37.495 22.965 ;
        RECT 75.000 23.185 75.875 27.860 ;
        RECT 76.585 27.715 78.585 27.945 ;
        RECT 76.195 26.465 76.425 27.665 ;
        RECT 76.970 26.465 78.135 27.715 ;
        RECT 78.745 26.465 78.975 27.665 ;
        RECT 76.195 25.675 78.975 26.465 ;
        RECT 80.735 27.510 80.965 28.230 ;
        RECT 80.735 27.485 81.100 27.510 ;
        RECT 81.260 27.485 81.580 27.540 ;
        RECT 80.735 27.335 81.580 27.485 ;
        RECT 80.735 27.305 81.100 27.335 ;
        RECT 80.735 26.230 80.965 27.305 ;
        RECT 81.260 27.280 81.580 27.335 ;
        RECT 83.865 26.055 85.680 28.435 ;
        RECT 89.025 28.195 89.255 28.230 ;
        RECT 89.880 28.195 90.580 29.165 ;
        RECT 89.025 26.285 90.580 28.195 ;
        RECT 89.025 26.230 89.255 26.285 ;
        RECT 81.265 26.025 88.895 26.055 ;
        RECT 81.015 25.795 88.975 26.025 ;
        RECT 76.195 23.705 76.425 25.675 ;
        RECT 78.745 25.005 78.975 25.675 ;
        RECT 78.745 24.725 81.610 25.005 ;
        RECT 78.745 24.635 89.030 24.725 ;
        RECT 78.745 23.705 78.975 24.635 ;
        RECT 81.170 24.485 89.030 24.635 ;
        RECT 81.110 24.255 89.110 24.485 ;
        RECT 80.675 23.765 80.905 24.205 ;
        RECT 89.315 24.195 89.545 24.205 ;
        RECT 81.395 23.765 82.395 23.835 ;
        RECT 89.315 23.765 89.550 24.195 ;
        RECT 76.585 23.425 78.585 23.655 ;
        RECT 76.675 23.185 78.500 23.425 ;
        RECT 75.000 22.695 78.500 23.185 ;
        RECT 34.690 22.510 35.010 22.570 ;
        RECT 40.960 22.510 41.220 22.600 ;
        RECT 34.690 22.370 41.220 22.510 ;
        RECT 34.690 22.310 35.010 22.370 ;
        RECT 40.960 22.280 41.220 22.370 ;
        RECT 31.885 22.115 32.205 22.175 ;
        RECT 44.170 22.115 44.430 22.205 ;
        RECT 31.885 21.975 44.430 22.115 ;
        RECT 31.885 21.915 32.205 21.975 ;
        RECT 44.170 21.885 44.430 21.975 ;
        RECT 75.000 17.860 75.875 22.695 ;
        RECT 76.675 22.515 78.500 22.695 ;
        RECT 80.675 22.875 89.550 23.765 ;
        RECT 76.585 22.285 78.585 22.515 ;
        RECT 80.675 22.245 80.905 22.875 ;
        RECT 81.395 22.820 82.395 22.875 ;
        RECT 89.315 22.310 89.550 22.875 ;
        RECT 89.315 22.245 89.545 22.310 ;
        RECT 76.195 20.800 76.425 22.235 ;
        RECT 78.745 20.800 78.975 22.235 ;
        RECT 81.110 21.965 89.110 22.195 ;
        RECT 81.180 21.840 89.010 21.965 ;
        RECT 81.200 21.055 89.000 21.840 ;
        RECT 81.110 20.825 89.110 21.055 ;
        RECT 76.195 19.460 78.975 20.800 ;
        RECT 80.675 20.750 80.905 20.775 ;
        RECT 76.195 18.275 76.425 19.460 ;
        RECT 76.770 18.225 78.365 19.460 ;
        RECT 78.745 18.570 78.975 19.460 ;
        RECT 80.670 20.305 80.905 20.750 ;
        RECT 89.315 20.750 89.545 20.775 ;
        RECT 80.670 20.295 81.085 20.305 ;
        RECT 81.225 20.295 82.225 20.365 ;
        RECT 80.670 20.290 82.225 20.295 ;
        RECT 82.635 20.290 84.255 20.295 ;
        RECT 89.315 20.290 89.550 20.750 ;
        RECT 80.670 19.400 89.550 20.290 ;
        RECT 80.670 19.385 82.225 19.400 ;
        RECT 82.635 19.395 84.255 19.400 ;
        RECT 80.670 19.295 81.085 19.385 ;
        RECT 81.225 19.335 82.225 19.385 ;
        RECT 80.670 18.865 80.905 19.295 ;
        RECT 80.675 18.815 80.905 18.865 ;
        RECT 89.315 18.865 89.550 19.400 ;
        RECT 89.315 18.815 89.545 18.865 ;
        RECT 81.110 18.570 89.110 18.765 ;
        RECT 78.745 18.535 89.110 18.570 ;
        RECT 78.745 18.390 89.030 18.535 ;
        RECT 78.745 18.375 81.245 18.390 ;
        RECT 78.745 18.275 78.975 18.375 ;
        RECT 76.585 17.995 78.585 18.225 ;
        RECT 89.880 18.115 90.580 26.285 ;
        RECT 84.955 17.985 85.230 18.055 ;
        RECT 79.260 17.860 85.230 17.985 ;
        RECT 75.000 17.845 76.405 17.860 ;
        RECT 78.750 17.845 85.230 17.860 ;
        RECT 75.000 17.795 85.230 17.845 ;
        RECT 75.000 17.670 79.450 17.795 ;
        RECT 84.955 17.720 85.230 17.795 ;
        RECT 75.000 12.390 75.875 17.670 ;
        RECT 77.825 17.365 81.610 17.370 ;
        RECT 77.825 17.300 85.060 17.365 ;
        RECT 76.645 17.175 85.060 17.300 ;
        RECT 76.645 17.085 85.105 17.175 ;
        RECT 76.585 17.075 85.105 17.085 ;
        RECT 76.585 16.855 78.585 17.075 ;
        RECT 81.105 16.945 85.105 17.075 ;
        RECT 76.195 15.425 76.425 16.805 ;
        RECT 78.745 15.425 78.975 16.805 ;
        RECT 76.195 14.470 78.975 15.425 ;
        RECT 76.195 12.845 76.425 14.470 ;
        RECT 78.745 12.845 78.975 14.470 ;
        RECT 80.670 15.640 80.900 16.895 ;
        RECT 82.340 15.640 83.725 16.945 ;
        RECT 85.310 15.640 85.540 16.895 ;
        RECT 85.905 16.435 90.580 18.115 ;
        RECT 87.265 16.095 87.540 16.125 ;
        RECT 87.250 15.840 87.580 16.095 ;
        RECT 87.265 15.820 87.555 15.840 ;
        RECT 87.265 15.790 87.540 15.820 ;
        RECT 80.670 15.570 85.540 15.640 ;
        RECT 87.075 15.570 87.305 15.615 ;
        RECT 80.670 14.295 85.545 15.570 ;
        RECT 80.670 12.935 80.900 14.295 ;
        RECT 85.310 12.935 85.545 14.295 ;
        RECT 76.585 12.565 78.585 12.795 ;
        RECT 76.650 12.390 78.520 12.565 ;
        RECT 75.000 11.835 78.520 12.390 ;
        RECT 75.000 6.730 75.875 11.835 ;
        RECT 76.650 11.655 78.520 11.835 ;
        RECT 76.585 11.425 78.585 11.655 ;
        RECT 80.710 11.465 80.870 12.935 ;
        RECT 85.340 12.925 85.545 12.935 ;
        RECT 81.105 12.655 85.105 12.885 ;
        RECT 81.185 12.410 85.010 12.655 ;
        RECT 87.065 12.410 87.305 15.570 ;
        RECT 81.185 11.920 87.305 12.410 ;
        RECT 81.185 11.745 85.010 11.920 ;
        RECT 81.105 11.515 85.105 11.745 ;
        RECT 76.195 9.980 76.425 11.375 ;
        RECT 78.745 9.980 78.975 11.375 ;
        RECT 76.195 9.025 78.975 9.980 ;
        RECT 76.195 7.415 76.425 9.025 ;
        RECT 78.745 7.415 78.975 9.025 ;
        RECT 80.670 10.090 80.900 11.465 ;
        RECT 85.310 11.350 85.540 11.465 ;
        RECT 85.310 10.715 85.545 11.350 ;
        RECT 87.065 10.715 87.305 11.920 ;
        RECT 85.310 10.090 85.540 10.715 ;
        RECT 87.075 10.615 87.305 10.715 ;
        RECT 87.515 15.600 87.745 15.615 ;
        RECT 88.165 15.600 88.645 16.435 ;
        RECT 87.515 10.675 88.655 15.600 ;
        RECT 89.880 12.535 90.580 16.435 ;
        RECT 92.000 29.025 92.875 29.140 ;
        RECT 92.000 28.665 98.445 29.025 ;
        RECT 92.000 28.530 105.975 28.665 ;
        RECT 92.000 28.085 92.875 28.530 ;
        RECT 98.015 28.435 105.975 28.530 ;
        RECT 92.000 27.860 92.885 28.085 ;
        RECT 93.595 28.000 94.815 28.085 ;
        RECT 93.595 27.945 94.830 28.000 ;
        RECT 92.000 23.185 92.875 27.860 ;
        RECT 93.585 27.715 95.585 27.945 ;
        RECT 93.195 26.465 93.425 27.665 ;
        RECT 93.970 26.465 95.135 27.715 ;
        RECT 95.745 26.465 95.975 27.665 ;
        RECT 93.195 25.675 95.975 26.465 ;
        RECT 97.735 27.510 97.965 28.230 ;
        RECT 97.735 27.485 98.100 27.510 ;
        RECT 98.260 27.485 98.580 27.540 ;
        RECT 97.735 27.335 98.580 27.485 ;
        RECT 97.735 27.305 98.100 27.335 ;
        RECT 97.735 26.230 97.965 27.305 ;
        RECT 98.260 27.280 98.580 27.335 ;
        RECT 100.865 26.055 102.680 28.435 ;
        RECT 106.025 28.195 106.255 28.230 ;
        RECT 106.880 28.195 107.580 29.165 ;
        RECT 106.025 26.285 107.580 28.195 ;
        RECT 106.025 26.230 106.255 26.285 ;
        RECT 98.265 26.025 105.895 26.055 ;
        RECT 98.015 25.795 105.975 26.025 ;
        RECT 93.195 23.705 93.425 25.675 ;
        RECT 95.745 25.005 95.975 25.675 ;
        RECT 95.745 24.725 98.610 25.005 ;
        RECT 95.745 24.635 106.030 24.725 ;
        RECT 95.745 23.705 95.975 24.635 ;
        RECT 98.170 24.485 106.030 24.635 ;
        RECT 98.110 24.255 106.110 24.485 ;
        RECT 97.675 23.765 97.905 24.205 ;
        RECT 106.315 24.195 106.545 24.205 ;
        RECT 98.395 23.765 99.395 23.835 ;
        RECT 106.315 23.765 106.550 24.195 ;
        RECT 93.585 23.425 95.585 23.655 ;
        RECT 93.675 23.185 95.500 23.425 ;
        RECT 92.000 22.695 95.500 23.185 ;
        RECT 92.000 17.860 92.875 22.695 ;
        RECT 93.675 22.515 95.500 22.695 ;
        RECT 97.675 22.875 106.550 23.765 ;
        RECT 93.585 22.285 95.585 22.515 ;
        RECT 97.675 22.245 97.905 22.875 ;
        RECT 98.395 22.820 99.395 22.875 ;
        RECT 106.315 22.310 106.550 22.875 ;
        RECT 106.315 22.245 106.545 22.310 ;
        RECT 93.195 20.800 93.425 22.235 ;
        RECT 95.745 20.800 95.975 22.235 ;
        RECT 98.110 21.965 106.110 22.195 ;
        RECT 98.180 21.840 106.010 21.965 ;
        RECT 98.200 21.055 106.000 21.840 ;
        RECT 98.110 20.825 106.110 21.055 ;
        RECT 93.195 19.460 95.975 20.800 ;
        RECT 97.675 20.750 97.905 20.775 ;
        RECT 93.195 18.275 93.425 19.460 ;
        RECT 93.770 18.225 95.365 19.460 ;
        RECT 95.745 18.570 95.975 19.460 ;
        RECT 97.670 20.305 97.905 20.750 ;
        RECT 106.315 20.750 106.545 20.775 ;
        RECT 97.670 20.295 98.085 20.305 ;
        RECT 98.225 20.295 99.225 20.365 ;
        RECT 97.670 20.290 99.225 20.295 ;
        RECT 99.635 20.290 101.255 20.295 ;
        RECT 106.315 20.290 106.550 20.750 ;
        RECT 97.670 19.400 106.550 20.290 ;
        RECT 97.670 19.385 99.225 19.400 ;
        RECT 99.635 19.395 101.255 19.400 ;
        RECT 97.670 19.295 98.085 19.385 ;
        RECT 98.225 19.335 99.225 19.385 ;
        RECT 97.670 18.865 97.905 19.295 ;
        RECT 97.675 18.815 97.905 18.865 ;
        RECT 106.315 18.865 106.550 19.400 ;
        RECT 106.315 18.815 106.545 18.865 ;
        RECT 98.110 18.570 106.110 18.765 ;
        RECT 95.745 18.535 106.110 18.570 ;
        RECT 95.745 18.390 106.030 18.535 ;
        RECT 95.745 18.375 98.245 18.390 ;
        RECT 95.745 18.275 95.975 18.375 ;
        RECT 93.585 17.995 95.585 18.225 ;
        RECT 106.880 18.115 107.580 26.285 ;
        RECT 101.955 17.985 102.230 18.055 ;
        RECT 96.260 17.860 102.230 17.985 ;
        RECT 92.000 17.845 93.405 17.860 ;
        RECT 95.750 17.845 102.230 17.860 ;
        RECT 92.000 17.795 102.230 17.845 ;
        RECT 92.000 17.670 96.450 17.795 ;
        RECT 101.955 17.720 102.230 17.795 ;
        RECT 89.795 11.700 90.660 12.535 ;
        RECT 92.000 12.390 92.875 17.670 ;
        RECT 94.825 17.365 98.610 17.370 ;
        RECT 94.825 17.300 102.060 17.365 ;
        RECT 93.645 17.175 102.060 17.300 ;
        RECT 93.645 17.085 102.105 17.175 ;
        RECT 93.585 17.075 102.105 17.085 ;
        RECT 93.585 16.855 95.585 17.075 ;
        RECT 98.105 16.945 102.105 17.075 ;
        RECT 93.195 15.425 93.425 16.805 ;
        RECT 95.745 15.425 95.975 16.805 ;
        RECT 93.195 14.470 95.975 15.425 ;
        RECT 93.195 12.845 93.425 14.470 ;
        RECT 95.745 12.845 95.975 14.470 ;
        RECT 97.670 15.640 97.900 16.895 ;
        RECT 99.340 15.640 100.725 16.945 ;
        RECT 102.310 15.640 102.540 16.895 ;
        RECT 102.905 16.435 107.580 18.115 ;
        RECT 104.265 16.095 104.540 16.125 ;
        RECT 104.250 15.840 104.580 16.095 ;
        RECT 104.265 15.820 104.555 15.840 ;
        RECT 104.265 15.790 104.540 15.820 ;
        RECT 97.670 15.570 102.540 15.640 ;
        RECT 104.075 15.570 104.305 15.615 ;
        RECT 97.670 14.295 102.545 15.570 ;
        RECT 97.670 12.935 97.900 14.295 ;
        RECT 102.310 12.935 102.545 14.295 ;
        RECT 93.585 12.565 95.585 12.795 ;
        RECT 93.650 12.390 95.520 12.565 ;
        RECT 92.000 11.835 95.520 12.390 ;
        RECT 87.515 10.615 87.745 10.675 ;
        RECT 87.265 10.405 87.555 10.410 ;
        RECT 87.250 10.150 87.580 10.405 ;
        RECT 80.670 8.745 85.540 10.090 ;
        RECT 80.670 7.505 80.900 8.745 ;
        RECT 85.310 7.505 85.540 8.745 ;
        RECT 76.585 7.340 78.585 7.365 ;
        RECT 81.105 7.340 85.105 7.455 ;
        RECT 76.585 7.265 78.590 7.340 ;
        RECT 79.125 7.265 85.105 7.340 ;
        RECT 76.585 7.225 85.105 7.265 ;
        RECT 76.585 7.135 85.040 7.225 ;
        RECT 76.640 7.000 85.040 7.135 ;
        RECT 75.000 6.290 76.860 6.730 ;
        RECT 75.000 6.280 77.850 6.290 ;
        RECT 75.000 5.935 78.520 6.280 ;
        RECT 75.000 4.310 76.860 5.935 ;
        RECT 77.660 5.785 78.520 5.935 ;
        RECT 77.155 5.595 77.405 5.610 ;
        RECT 77.155 5.305 77.430 5.595 ;
        RECT 77.590 5.555 78.590 5.785 ;
        RECT 79.010 5.690 79.280 7.000 ;
        RECT 89.880 6.570 90.580 11.700 ;
        RECT 84.300 6.235 90.580 6.570 ;
        RECT 81.185 6.095 90.580 6.235 ;
        RECT 81.185 5.870 85.045 6.095 ;
        RECT 77.155 5.275 77.405 5.305 ;
        RECT 77.590 5.115 78.590 5.345 ;
        RECT 78.735 5.270 80.925 5.690 ;
        RECT 81.120 5.640 85.120 5.870 ;
        RECT 85.355 5.680 85.605 5.700 ;
        RECT 81.120 5.200 85.120 5.430 ;
        RECT 85.325 5.390 85.605 5.680 ;
        RECT 85.355 5.365 85.605 5.390 ;
        RECT 77.660 4.975 78.545 5.115 ;
        RECT 81.170 5.035 85.095 5.200 ;
        RECT 78.730 4.975 85.095 5.035 ;
        RECT 77.660 4.920 85.095 4.975 ;
        RECT 77.660 4.850 81.540 4.920 ;
        RECT 78.215 4.735 81.540 4.850 ;
        RECT 89.880 4.770 90.580 6.095 ;
        RECT 75.000 4.265 77.385 4.310 ;
        RECT 75.000 2.535 75.875 4.265 ;
        RECT 76.240 3.990 77.385 4.265 ;
        RECT 79.570 4.105 79.975 4.735 ;
        RECT 88.575 4.235 90.580 4.770 ;
        RECT 76.240 3.925 78.490 3.990 ;
        RECT 76.680 3.760 78.490 3.925 ;
        RECT 76.165 3.570 76.415 3.595 ;
        RECT 76.165 3.280 76.435 3.570 ;
        RECT 76.595 3.530 78.595 3.760 ;
        RECT 79.555 3.740 79.980 4.105 ;
        RECT 81.220 4.090 90.580 4.235 ;
        RECT 81.220 3.845 89.075 4.090 ;
        RECT 76.165 3.260 76.415 3.280 ;
        RECT 76.595 3.090 78.595 3.320 ;
        RECT 78.745 3.230 80.935 3.740 ;
        RECT 81.125 3.615 89.125 3.845 ;
        RECT 89.355 3.655 89.605 3.670 ;
        RECT 78.745 3.225 79.445 3.230 ;
        RECT 80.445 3.225 80.935 3.230 ;
        RECT 81.125 3.175 89.125 3.405 ;
        RECT 89.330 3.365 89.605 3.655 ;
        RECT 89.355 3.335 89.605 3.365 ;
        RECT 76.665 2.925 78.530 3.090 ;
        RECT 79.415 2.925 80.415 3.000 ;
        RECT 81.200 2.925 89.050 3.175 ;
        RECT 76.665 2.630 89.050 2.925 ;
        RECT 89.880 2.690 90.580 4.090 ;
        RECT 92.000 6.730 92.875 11.835 ;
        RECT 93.650 11.655 95.520 11.835 ;
        RECT 93.585 11.425 95.585 11.655 ;
        RECT 97.710 11.465 97.870 12.935 ;
        RECT 102.340 12.925 102.545 12.935 ;
        RECT 98.105 12.655 102.105 12.885 ;
        RECT 98.185 12.410 102.010 12.655 ;
        RECT 104.065 12.410 104.305 15.570 ;
        RECT 98.185 11.920 104.305 12.410 ;
        RECT 98.185 11.745 102.010 11.920 ;
        RECT 98.105 11.515 102.105 11.745 ;
        RECT 93.195 9.980 93.425 11.375 ;
        RECT 95.745 9.980 95.975 11.375 ;
        RECT 93.195 9.025 95.975 9.980 ;
        RECT 93.195 7.415 93.425 9.025 ;
        RECT 95.745 7.415 95.975 9.025 ;
        RECT 97.670 10.090 97.900 11.465 ;
        RECT 102.310 11.350 102.540 11.465 ;
        RECT 102.310 10.715 102.545 11.350 ;
        RECT 104.065 10.715 104.305 11.920 ;
        RECT 102.310 10.090 102.540 10.715 ;
        RECT 104.075 10.615 104.305 10.715 ;
        RECT 104.515 15.600 104.745 15.615 ;
        RECT 105.165 15.600 105.645 16.435 ;
        RECT 104.515 10.675 105.655 15.600 ;
        RECT 106.880 12.500 107.580 16.435 ;
        RECT 109.000 29.025 109.875 29.140 ;
        RECT 109.000 28.665 115.445 29.025 ;
        RECT 109.000 28.530 122.975 28.665 ;
        RECT 109.000 28.085 109.875 28.530 ;
        RECT 115.015 28.435 122.975 28.530 ;
        RECT 109.000 27.860 109.885 28.085 ;
        RECT 110.595 28.000 111.815 28.085 ;
        RECT 110.595 27.945 111.830 28.000 ;
        RECT 109.000 23.185 109.875 27.860 ;
        RECT 110.585 27.715 112.585 27.945 ;
        RECT 110.195 26.465 110.425 27.665 ;
        RECT 110.970 26.465 112.135 27.715 ;
        RECT 112.745 26.465 112.975 27.665 ;
        RECT 110.195 25.675 112.975 26.465 ;
        RECT 114.735 27.510 114.965 28.230 ;
        RECT 114.735 27.485 115.100 27.510 ;
        RECT 115.260 27.485 115.580 27.540 ;
        RECT 114.735 27.335 115.580 27.485 ;
        RECT 114.735 27.305 115.100 27.335 ;
        RECT 114.735 26.230 114.965 27.305 ;
        RECT 115.260 27.280 115.580 27.335 ;
        RECT 117.865 26.055 119.680 28.435 ;
        RECT 123.025 28.195 123.255 28.230 ;
        RECT 123.880 28.195 124.580 29.165 ;
        RECT 123.025 26.285 124.580 28.195 ;
        RECT 123.025 26.230 123.255 26.285 ;
        RECT 115.265 26.025 122.895 26.055 ;
        RECT 115.015 25.795 122.975 26.025 ;
        RECT 110.195 23.705 110.425 25.675 ;
        RECT 112.745 25.005 112.975 25.675 ;
        RECT 112.745 24.725 115.610 25.005 ;
        RECT 112.745 24.635 123.030 24.725 ;
        RECT 112.745 23.705 112.975 24.635 ;
        RECT 115.170 24.485 123.030 24.635 ;
        RECT 115.110 24.255 123.110 24.485 ;
        RECT 114.675 23.765 114.905 24.205 ;
        RECT 123.315 24.195 123.545 24.205 ;
        RECT 115.395 23.765 116.395 23.835 ;
        RECT 123.315 23.765 123.550 24.195 ;
        RECT 110.585 23.425 112.585 23.655 ;
        RECT 110.675 23.185 112.500 23.425 ;
        RECT 109.000 22.695 112.500 23.185 ;
        RECT 109.000 17.860 109.875 22.695 ;
        RECT 110.675 22.515 112.500 22.695 ;
        RECT 114.675 22.875 123.550 23.765 ;
        RECT 110.585 22.285 112.585 22.515 ;
        RECT 114.675 22.245 114.905 22.875 ;
        RECT 115.395 22.820 116.395 22.875 ;
        RECT 123.315 22.310 123.550 22.875 ;
        RECT 123.315 22.245 123.545 22.310 ;
        RECT 110.195 20.800 110.425 22.235 ;
        RECT 112.745 20.800 112.975 22.235 ;
        RECT 115.110 21.965 123.110 22.195 ;
        RECT 115.180 21.840 123.010 21.965 ;
        RECT 115.200 21.055 123.000 21.840 ;
        RECT 115.110 20.825 123.110 21.055 ;
        RECT 110.195 19.460 112.975 20.800 ;
        RECT 114.675 20.750 114.905 20.775 ;
        RECT 110.195 18.275 110.425 19.460 ;
        RECT 110.770 18.225 112.365 19.460 ;
        RECT 112.745 18.570 112.975 19.460 ;
        RECT 114.670 20.305 114.905 20.750 ;
        RECT 123.315 20.750 123.545 20.775 ;
        RECT 114.670 20.295 115.085 20.305 ;
        RECT 115.225 20.295 116.225 20.365 ;
        RECT 114.670 20.290 116.225 20.295 ;
        RECT 116.635 20.290 118.255 20.295 ;
        RECT 123.315 20.290 123.550 20.750 ;
        RECT 114.670 19.400 123.550 20.290 ;
        RECT 114.670 19.385 116.225 19.400 ;
        RECT 116.635 19.395 118.255 19.400 ;
        RECT 114.670 19.295 115.085 19.385 ;
        RECT 115.225 19.335 116.225 19.385 ;
        RECT 114.670 18.865 114.905 19.295 ;
        RECT 114.675 18.815 114.905 18.865 ;
        RECT 123.315 18.865 123.550 19.400 ;
        RECT 123.315 18.815 123.545 18.865 ;
        RECT 115.110 18.570 123.110 18.765 ;
        RECT 112.745 18.535 123.110 18.570 ;
        RECT 112.745 18.390 123.030 18.535 ;
        RECT 112.745 18.375 115.245 18.390 ;
        RECT 112.745 18.275 112.975 18.375 ;
        RECT 110.585 17.995 112.585 18.225 ;
        RECT 123.880 18.115 124.580 26.285 ;
        RECT 118.955 17.985 119.230 18.055 ;
        RECT 113.260 17.860 119.230 17.985 ;
        RECT 109.000 17.845 110.405 17.860 ;
        RECT 112.750 17.845 119.230 17.860 ;
        RECT 109.000 17.795 119.230 17.845 ;
        RECT 109.000 17.670 113.450 17.795 ;
        RECT 118.955 17.720 119.230 17.795 ;
        RECT 106.820 11.725 107.595 12.500 ;
        RECT 109.000 12.390 109.875 17.670 ;
        RECT 111.825 17.365 115.610 17.370 ;
        RECT 111.825 17.300 119.060 17.365 ;
        RECT 110.645 17.175 119.060 17.300 ;
        RECT 110.645 17.085 119.105 17.175 ;
        RECT 110.585 17.075 119.105 17.085 ;
        RECT 110.585 16.855 112.585 17.075 ;
        RECT 115.105 16.945 119.105 17.075 ;
        RECT 110.195 15.425 110.425 16.805 ;
        RECT 112.745 15.425 112.975 16.805 ;
        RECT 110.195 14.470 112.975 15.425 ;
        RECT 110.195 12.845 110.425 14.470 ;
        RECT 112.745 12.845 112.975 14.470 ;
        RECT 114.670 15.640 114.900 16.895 ;
        RECT 116.340 15.640 117.725 16.945 ;
        RECT 119.310 15.640 119.540 16.895 ;
        RECT 119.905 16.435 124.580 18.115 ;
        RECT 121.265 16.095 121.540 16.125 ;
        RECT 121.250 15.840 121.580 16.095 ;
        RECT 121.265 15.820 121.555 15.840 ;
        RECT 121.265 15.790 121.540 15.820 ;
        RECT 114.670 15.570 119.540 15.640 ;
        RECT 121.075 15.570 121.305 15.615 ;
        RECT 114.670 14.295 119.545 15.570 ;
        RECT 114.670 12.935 114.900 14.295 ;
        RECT 119.310 12.935 119.545 14.295 ;
        RECT 110.585 12.565 112.585 12.795 ;
        RECT 110.650 12.390 112.520 12.565 ;
        RECT 109.000 11.835 112.520 12.390 ;
        RECT 104.515 10.615 104.745 10.675 ;
        RECT 104.265 10.405 104.555 10.410 ;
        RECT 104.250 10.150 104.580 10.405 ;
        RECT 97.670 8.745 102.540 10.090 ;
        RECT 97.670 7.505 97.900 8.745 ;
        RECT 102.310 7.505 102.540 8.745 ;
        RECT 93.585 7.340 95.585 7.365 ;
        RECT 98.105 7.340 102.105 7.455 ;
        RECT 93.585 7.265 95.590 7.340 ;
        RECT 96.125 7.265 102.105 7.340 ;
        RECT 93.585 7.225 102.105 7.265 ;
        RECT 93.585 7.135 102.040 7.225 ;
        RECT 93.640 7.000 102.040 7.135 ;
        RECT 92.000 6.290 93.860 6.730 ;
        RECT 92.000 6.280 94.850 6.290 ;
        RECT 92.000 5.935 95.520 6.280 ;
        RECT 92.000 4.310 93.860 5.935 ;
        RECT 94.660 5.785 95.520 5.935 ;
        RECT 94.155 5.595 94.405 5.610 ;
        RECT 94.155 5.305 94.430 5.595 ;
        RECT 94.590 5.555 95.590 5.785 ;
        RECT 96.010 5.690 96.280 7.000 ;
        RECT 106.880 6.570 107.580 11.725 ;
        RECT 101.300 6.235 107.580 6.570 ;
        RECT 98.185 6.095 107.580 6.235 ;
        RECT 98.185 5.870 102.045 6.095 ;
        RECT 94.155 5.275 94.405 5.305 ;
        RECT 94.590 5.115 95.590 5.345 ;
        RECT 95.735 5.270 97.925 5.690 ;
        RECT 98.120 5.640 102.120 5.870 ;
        RECT 102.355 5.680 102.605 5.700 ;
        RECT 98.120 5.200 102.120 5.430 ;
        RECT 102.325 5.390 102.605 5.680 ;
        RECT 102.355 5.365 102.605 5.390 ;
        RECT 94.660 4.975 95.545 5.115 ;
        RECT 98.170 5.035 102.095 5.200 ;
        RECT 95.730 4.975 102.095 5.035 ;
        RECT 94.660 4.920 102.095 4.975 ;
        RECT 94.660 4.850 98.540 4.920 ;
        RECT 95.215 4.735 98.540 4.850 ;
        RECT 106.880 4.770 107.580 6.095 ;
        RECT 92.000 4.265 94.385 4.310 ;
        RECT 76.665 2.560 81.730 2.630 ;
        RECT 78.205 2.555 81.730 2.560 ;
        RECT 60.850 2.190 61.170 2.210 ;
        RECT 79.415 2.190 80.415 2.555 ;
        RECT 92.000 2.535 92.875 4.265 ;
        RECT 93.240 3.990 94.385 4.265 ;
        RECT 96.570 4.105 96.975 4.735 ;
        RECT 105.575 4.235 107.580 4.770 ;
        RECT 93.240 3.925 95.490 3.990 ;
        RECT 93.680 3.760 95.490 3.925 ;
        RECT 93.165 3.570 93.415 3.595 ;
        RECT 93.165 3.280 93.435 3.570 ;
        RECT 93.595 3.530 95.595 3.760 ;
        RECT 96.555 3.740 96.980 4.105 ;
        RECT 98.220 4.090 107.580 4.235 ;
        RECT 98.220 3.845 106.075 4.090 ;
        RECT 93.165 3.260 93.415 3.280 ;
        RECT 93.595 3.090 95.595 3.320 ;
        RECT 95.745 3.230 97.935 3.740 ;
        RECT 98.125 3.615 106.125 3.845 ;
        RECT 106.355 3.655 106.605 3.670 ;
        RECT 95.745 3.225 96.445 3.230 ;
        RECT 97.445 3.225 97.935 3.230 ;
        RECT 98.125 3.175 106.125 3.405 ;
        RECT 106.330 3.365 106.605 3.655 ;
        RECT 106.355 3.335 106.605 3.365 ;
        RECT 93.665 2.925 95.530 3.090 ;
        RECT 96.415 2.925 97.415 3.000 ;
        RECT 98.200 2.925 106.050 3.175 ;
        RECT 93.665 2.630 106.050 2.925 ;
        RECT 106.880 2.690 107.580 4.090 ;
        RECT 109.000 6.730 109.875 11.835 ;
        RECT 110.650 11.655 112.520 11.835 ;
        RECT 110.585 11.425 112.585 11.655 ;
        RECT 114.710 11.465 114.870 12.935 ;
        RECT 119.340 12.925 119.545 12.935 ;
        RECT 115.105 12.655 119.105 12.885 ;
        RECT 115.185 12.410 119.010 12.655 ;
        RECT 121.065 12.410 121.305 15.570 ;
        RECT 115.185 11.920 121.305 12.410 ;
        RECT 115.185 11.745 119.010 11.920 ;
        RECT 115.105 11.515 119.105 11.745 ;
        RECT 110.195 9.980 110.425 11.375 ;
        RECT 112.745 9.980 112.975 11.375 ;
        RECT 110.195 9.025 112.975 9.980 ;
        RECT 110.195 7.415 110.425 9.025 ;
        RECT 112.745 7.415 112.975 9.025 ;
        RECT 114.670 10.090 114.900 11.465 ;
        RECT 119.310 11.350 119.540 11.465 ;
        RECT 119.310 10.715 119.545 11.350 ;
        RECT 121.065 10.715 121.305 11.920 ;
        RECT 119.310 10.090 119.540 10.715 ;
        RECT 121.075 10.615 121.305 10.715 ;
        RECT 121.515 15.600 121.745 15.615 ;
        RECT 122.165 15.600 122.645 16.435 ;
        RECT 121.515 10.675 122.655 15.600 ;
        RECT 123.880 12.530 124.580 16.435 ;
        RECT 123.715 11.710 124.580 12.530 ;
        RECT 121.515 10.615 121.745 10.675 ;
        RECT 121.265 10.405 121.555 10.410 ;
        RECT 121.250 10.150 121.580 10.405 ;
        RECT 114.670 8.745 119.540 10.090 ;
        RECT 114.670 7.505 114.900 8.745 ;
        RECT 119.310 7.505 119.540 8.745 ;
        RECT 110.585 7.340 112.585 7.365 ;
        RECT 115.105 7.340 119.105 7.455 ;
        RECT 110.585 7.265 112.590 7.340 ;
        RECT 113.125 7.265 119.105 7.340 ;
        RECT 110.585 7.225 119.105 7.265 ;
        RECT 110.585 7.135 119.040 7.225 ;
        RECT 110.640 7.000 119.040 7.135 ;
        RECT 109.000 6.290 110.860 6.730 ;
        RECT 109.000 6.280 111.850 6.290 ;
        RECT 109.000 5.935 112.520 6.280 ;
        RECT 109.000 4.310 110.860 5.935 ;
        RECT 111.660 5.785 112.520 5.935 ;
        RECT 111.155 5.595 111.405 5.610 ;
        RECT 111.155 5.305 111.430 5.595 ;
        RECT 111.590 5.555 112.590 5.785 ;
        RECT 113.010 5.690 113.280 7.000 ;
        RECT 123.880 6.570 124.580 11.710 ;
        RECT 118.300 6.235 124.580 6.570 ;
        RECT 115.185 6.095 124.580 6.235 ;
        RECT 115.185 5.870 119.045 6.095 ;
        RECT 111.155 5.275 111.405 5.305 ;
        RECT 111.590 5.115 112.590 5.345 ;
        RECT 112.735 5.270 114.925 5.690 ;
        RECT 115.120 5.640 119.120 5.870 ;
        RECT 119.355 5.680 119.605 5.700 ;
        RECT 115.120 5.200 119.120 5.430 ;
        RECT 119.325 5.390 119.605 5.680 ;
        RECT 119.355 5.365 119.605 5.390 ;
        RECT 111.660 4.975 112.545 5.115 ;
        RECT 115.170 5.035 119.095 5.200 ;
        RECT 112.730 4.975 119.095 5.035 ;
        RECT 111.660 4.920 119.095 4.975 ;
        RECT 111.660 4.850 115.540 4.920 ;
        RECT 112.215 4.735 115.540 4.850 ;
        RECT 123.880 4.770 124.580 6.095 ;
        RECT 109.000 4.265 111.385 4.310 ;
        RECT 93.665 2.560 98.730 2.630 ;
        RECT 95.205 2.555 98.730 2.560 ;
        RECT 60.850 2.000 80.415 2.190 ;
        RECT 96.415 2.000 97.415 2.555 ;
        RECT 109.000 2.535 109.875 4.265 ;
        RECT 110.240 3.990 111.385 4.265 ;
        RECT 113.570 4.105 113.975 4.735 ;
        RECT 122.575 4.235 124.580 4.770 ;
        RECT 110.240 3.925 112.490 3.990 ;
        RECT 110.680 3.760 112.490 3.925 ;
        RECT 110.165 3.570 110.415 3.595 ;
        RECT 110.165 3.280 110.435 3.570 ;
        RECT 110.595 3.530 112.595 3.760 ;
        RECT 113.555 3.740 113.980 4.105 ;
        RECT 115.220 4.090 124.580 4.235 ;
        RECT 115.220 3.845 123.075 4.090 ;
        RECT 110.165 3.260 110.415 3.280 ;
        RECT 110.595 3.090 112.595 3.320 ;
        RECT 112.745 3.230 114.935 3.740 ;
        RECT 115.125 3.615 123.125 3.845 ;
        RECT 123.355 3.655 123.605 3.670 ;
        RECT 112.745 3.225 113.445 3.230 ;
        RECT 114.445 3.225 114.935 3.230 ;
        RECT 115.125 3.175 123.125 3.405 ;
        RECT 123.330 3.365 123.605 3.655 ;
        RECT 123.355 3.335 123.605 3.365 ;
        RECT 110.665 2.925 112.530 3.090 ;
        RECT 113.415 2.925 114.415 3.000 ;
        RECT 115.200 2.925 123.050 3.175 ;
        RECT 110.665 2.630 123.050 2.925 ;
        RECT 123.880 2.690 124.580 4.090 ;
        RECT 126.000 29.025 126.875 29.140 ;
        RECT 126.000 28.665 132.445 29.025 ;
        RECT 126.000 28.530 139.975 28.665 ;
        RECT 126.000 28.085 126.875 28.530 ;
        RECT 132.015 28.435 139.975 28.530 ;
        RECT 126.000 27.860 126.885 28.085 ;
        RECT 127.595 28.000 128.815 28.085 ;
        RECT 127.595 27.945 128.830 28.000 ;
        RECT 126.000 23.185 126.875 27.860 ;
        RECT 127.585 27.715 129.585 27.945 ;
        RECT 127.195 26.465 127.425 27.665 ;
        RECT 127.970 26.465 129.135 27.715 ;
        RECT 129.745 26.465 129.975 27.665 ;
        RECT 127.195 25.675 129.975 26.465 ;
        RECT 131.735 27.510 131.965 28.230 ;
        RECT 131.735 27.485 132.100 27.510 ;
        RECT 132.260 27.485 132.580 27.540 ;
        RECT 131.735 27.335 132.580 27.485 ;
        RECT 131.735 27.305 132.100 27.335 ;
        RECT 131.735 26.230 131.965 27.305 ;
        RECT 132.260 27.280 132.580 27.335 ;
        RECT 134.865 26.055 136.680 28.435 ;
        RECT 140.025 28.195 140.255 28.230 ;
        RECT 140.880 28.195 141.580 29.165 ;
        RECT 140.025 26.285 141.580 28.195 ;
        RECT 140.025 26.230 140.255 26.285 ;
        RECT 140.815 26.175 141.580 26.285 ;
        RECT 132.265 26.025 139.895 26.055 ;
        RECT 132.015 25.795 139.975 26.025 ;
        RECT 127.195 23.705 127.425 25.675 ;
        RECT 129.745 25.005 129.975 25.675 ;
        RECT 129.745 24.725 132.610 25.005 ;
        RECT 129.745 24.635 140.030 24.725 ;
        RECT 129.745 23.705 129.975 24.635 ;
        RECT 132.170 24.485 140.030 24.635 ;
        RECT 132.110 24.255 140.110 24.485 ;
        RECT 131.675 23.765 131.905 24.205 ;
        RECT 140.315 24.195 140.545 24.205 ;
        RECT 132.395 23.765 133.395 23.835 ;
        RECT 140.315 23.765 140.550 24.195 ;
        RECT 127.585 23.425 129.585 23.655 ;
        RECT 127.675 23.185 129.500 23.425 ;
        RECT 126.000 22.695 129.500 23.185 ;
        RECT 126.000 17.860 126.875 22.695 ;
        RECT 127.675 22.515 129.500 22.695 ;
        RECT 131.675 22.875 140.550 23.765 ;
        RECT 127.585 22.285 129.585 22.515 ;
        RECT 131.675 22.245 131.905 22.875 ;
        RECT 132.395 22.820 133.395 22.875 ;
        RECT 140.315 22.310 140.550 22.875 ;
        RECT 140.315 22.245 140.545 22.310 ;
        RECT 127.195 20.800 127.425 22.235 ;
        RECT 129.745 20.800 129.975 22.235 ;
        RECT 132.110 21.965 140.110 22.195 ;
        RECT 132.180 21.840 140.010 21.965 ;
        RECT 132.200 21.055 140.000 21.840 ;
        RECT 132.110 20.825 140.110 21.055 ;
        RECT 127.195 19.460 129.975 20.800 ;
        RECT 131.675 20.750 131.905 20.775 ;
        RECT 127.195 18.275 127.425 19.460 ;
        RECT 127.770 18.225 129.365 19.460 ;
        RECT 129.745 18.570 129.975 19.460 ;
        RECT 131.670 20.305 131.905 20.750 ;
        RECT 140.315 20.750 140.545 20.775 ;
        RECT 131.670 20.295 132.085 20.305 ;
        RECT 132.225 20.295 133.225 20.365 ;
        RECT 131.670 20.290 133.225 20.295 ;
        RECT 133.635 20.290 135.255 20.295 ;
        RECT 140.315 20.290 140.550 20.750 ;
        RECT 131.670 19.400 140.550 20.290 ;
        RECT 131.670 19.385 133.225 19.400 ;
        RECT 133.635 19.395 135.255 19.400 ;
        RECT 131.670 19.295 132.085 19.385 ;
        RECT 132.225 19.335 133.225 19.385 ;
        RECT 131.670 18.865 131.905 19.295 ;
        RECT 131.675 18.815 131.905 18.865 ;
        RECT 140.315 18.865 140.550 19.400 ;
        RECT 140.315 18.815 140.545 18.865 ;
        RECT 132.110 18.570 140.110 18.765 ;
        RECT 129.745 18.535 140.110 18.570 ;
        RECT 129.745 18.390 140.030 18.535 ;
        RECT 129.745 18.375 132.245 18.390 ;
        RECT 129.745 18.275 129.975 18.375 ;
        RECT 127.585 17.995 129.585 18.225 ;
        RECT 140.880 18.115 141.580 26.175 ;
        RECT 135.955 17.985 136.230 18.055 ;
        RECT 130.260 17.860 136.230 17.985 ;
        RECT 126.000 17.845 127.405 17.860 ;
        RECT 129.750 17.845 136.230 17.860 ;
        RECT 126.000 17.795 136.230 17.845 ;
        RECT 126.000 17.670 130.450 17.795 ;
        RECT 135.955 17.720 136.230 17.795 ;
        RECT 126.000 12.390 126.875 17.670 ;
        RECT 128.825 17.365 132.610 17.370 ;
        RECT 128.825 17.300 136.060 17.365 ;
        RECT 127.645 17.175 136.060 17.300 ;
        RECT 127.645 17.085 136.105 17.175 ;
        RECT 127.585 17.075 136.105 17.085 ;
        RECT 127.585 16.855 129.585 17.075 ;
        RECT 132.105 16.945 136.105 17.075 ;
        RECT 127.195 15.425 127.425 16.805 ;
        RECT 129.745 15.425 129.975 16.805 ;
        RECT 127.195 14.470 129.975 15.425 ;
        RECT 127.195 12.845 127.425 14.470 ;
        RECT 129.745 12.845 129.975 14.470 ;
        RECT 131.670 15.640 131.900 16.895 ;
        RECT 133.340 15.640 134.725 16.945 ;
        RECT 136.310 15.640 136.540 16.895 ;
        RECT 136.905 16.435 141.580 18.115 ;
        RECT 138.265 16.095 138.540 16.125 ;
        RECT 138.250 15.840 138.580 16.095 ;
        RECT 138.265 15.820 138.555 15.840 ;
        RECT 138.265 15.790 138.540 15.820 ;
        RECT 131.670 15.570 136.540 15.640 ;
        RECT 138.075 15.570 138.305 15.615 ;
        RECT 131.670 14.295 136.545 15.570 ;
        RECT 131.670 12.935 131.900 14.295 ;
        RECT 136.310 12.935 136.545 14.295 ;
        RECT 127.585 12.565 129.585 12.795 ;
        RECT 127.650 12.390 129.520 12.565 ;
        RECT 126.000 11.835 129.520 12.390 ;
        RECT 126.000 6.730 126.875 11.835 ;
        RECT 127.650 11.655 129.520 11.835 ;
        RECT 127.585 11.425 129.585 11.655 ;
        RECT 131.710 11.465 131.870 12.935 ;
        RECT 136.340 12.925 136.545 12.935 ;
        RECT 132.105 12.655 136.105 12.885 ;
        RECT 132.185 12.410 136.010 12.655 ;
        RECT 138.065 12.410 138.305 15.570 ;
        RECT 132.185 11.920 138.305 12.410 ;
        RECT 132.185 11.745 136.010 11.920 ;
        RECT 132.105 11.515 136.105 11.745 ;
        RECT 127.195 9.980 127.425 11.375 ;
        RECT 129.745 9.980 129.975 11.375 ;
        RECT 127.195 9.025 129.975 9.980 ;
        RECT 127.195 7.415 127.425 9.025 ;
        RECT 129.745 7.415 129.975 9.025 ;
        RECT 131.670 10.090 131.900 11.465 ;
        RECT 136.310 11.350 136.540 11.465 ;
        RECT 136.310 10.715 136.545 11.350 ;
        RECT 138.065 10.715 138.305 11.920 ;
        RECT 136.310 10.090 136.540 10.715 ;
        RECT 138.075 10.615 138.305 10.715 ;
        RECT 138.515 15.600 138.745 15.615 ;
        RECT 139.165 15.600 139.645 16.435 ;
        RECT 138.515 10.675 139.655 15.600 ;
        RECT 140.880 12.535 141.580 16.435 ;
        RECT 140.680 11.715 141.580 12.535 ;
        RECT 138.515 10.615 138.745 10.675 ;
        RECT 138.265 10.405 138.555 10.410 ;
        RECT 138.250 10.150 138.580 10.405 ;
        RECT 131.670 8.745 136.540 10.090 ;
        RECT 131.670 7.505 131.900 8.745 ;
        RECT 136.310 7.505 136.540 8.745 ;
        RECT 127.585 7.340 129.585 7.365 ;
        RECT 132.105 7.340 136.105 7.455 ;
        RECT 127.585 7.265 129.590 7.340 ;
        RECT 130.125 7.265 136.105 7.340 ;
        RECT 127.585 7.225 136.105 7.265 ;
        RECT 127.585 7.135 136.040 7.225 ;
        RECT 127.640 7.000 136.040 7.135 ;
        RECT 126.000 6.290 127.860 6.730 ;
        RECT 126.000 6.280 128.850 6.290 ;
        RECT 126.000 5.935 129.520 6.280 ;
        RECT 126.000 4.310 127.860 5.935 ;
        RECT 128.660 5.785 129.520 5.935 ;
        RECT 128.155 5.595 128.405 5.610 ;
        RECT 128.155 5.305 128.430 5.595 ;
        RECT 128.590 5.555 129.590 5.785 ;
        RECT 130.010 5.690 130.280 7.000 ;
        RECT 140.880 6.570 141.580 11.715 ;
        RECT 135.300 6.235 141.580 6.570 ;
        RECT 132.185 6.095 141.580 6.235 ;
        RECT 132.185 5.870 136.045 6.095 ;
        RECT 128.155 5.275 128.405 5.305 ;
        RECT 128.590 5.115 129.590 5.345 ;
        RECT 129.735 5.270 131.925 5.690 ;
        RECT 132.120 5.640 136.120 5.870 ;
        RECT 136.355 5.680 136.605 5.700 ;
        RECT 132.120 5.200 136.120 5.430 ;
        RECT 136.325 5.390 136.605 5.680 ;
        RECT 136.355 5.365 136.605 5.390 ;
        RECT 128.660 4.975 129.545 5.115 ;
        RECT 132.170 5.035 136.095 5.200 ;
        RECT 129.730 4.975 136.095 5.035 ;
        RECT 128.660 4.920 136.095 4.975 ;
        RECT 128.660 4.850 132.540 4.920 ;
        RECT 129.215 4.735 132.540 4.850 ;
        RECT 140.880 4.770 141.580 6.095 ;
        RECT 126.000 4.265 128.385 4.310 ;
        RECT 110.665 2.560 115.730 2.630 ;
        RECT 112.205 2.555 115.730 2.560 ;
        RECT 113.415 2.000 114.415 2.555 ;
        RECT 126.000 2.535 126.875 4.265 ;
        RECT 127.240 3.990 128.385 4.265 ;
        RECT 130.570 4.105 130.975 4.735 ;
        RECT 139.575 4.235 141.580 4.770 ;
        RECT 127.240 3.925 129.490 3.990 ;
        RECT 127.680 3.760 129.490 3.925 ;
        RECT 127.165 3.570 127.415 3.595 ;
        RECT 127.165 3.280 127.435 3.570 ;
        RECT 127.595 3.530 129.595 3.760 ;
        RECT 130.555 3.740 130.980 4.105 ;
        RECT 132.220 4.090 141.580 4.235 ;
        RECT 132.220 3.845 140.075 4.090 ;
        RECT 127.165 3.260 127.415 3.280 ;
        RECT 127.595 3.090 129.595 3.320 ;
        RECT 129.745 3.230 131.935 3.740 ;
        RECT 132.125 3.615 140.125 3.845 ;
        RECT 140.355 3.655 140.605 3.670 ;
        RECT 129.745 3.225 130.445 3.230 ;
        RECT 131.445 3.225 131.935 3.230 ;
        RECT 132.125 3.175 140.125 3.405 ;
        RECT 140.330 3.365 140.605 3.655 ;
        RECT 140.355 3.335 140.605 3.365 ;
        RECT 127.665 2.925 129.530 3.090 ;
        RECT 130.415 2.925 131.415 3.000 ;
        RECT 132.200 2.925 140.050 3.175 ;
        RECT 127.665 2.630 140.050 2.925 ;
        RECT 140.880 2.690 141.580 4.090 ;
        RECT 143.000 29.025 143.875 29.140 ;
        RECT 143.000 28.665 149.445 29.025 ;
        RECT 143.000 28.530 156.975 28.665 ;
        RECT 143.000 28.085 143.875 28.530 ;
        RECT 149.015 28.435 156.975 28.530 ;
        RECT 143.000 27.860 143.885 28.085 ;
        RECT 144.595 28.000 145.815 28.085 ;
        RECT 144.595 27.945 145.830 28.000 ;
        RECT 143.000 23.185 143.875 27.860 ;
        RECT 144.585 27.715 146.585 27.945 ;
        RECT 144.195 26.465 144.425 27.665 ;
        RECT 144.970 26.465 146.135 27.715 ;
        RECT 146.745 26.465 146.975 27.665 ;
        RECT 144.195 25.675 146.975 26.465 ;
        RECT 148.735 27.510 148.965 28.230 ;
        RECT 148.735 27.485 149.100 27.510 ;
        RECT 149.260 27.485 149.580 27.540 ;
        RECT 148.735 27.335 149.580 27.485 ;
        RECT 148.735 27.305 149.100 27.335 ;
        RECT 148.735 26.230 148.965 27.305 ;
        RECT 149.260 27.280 149.580 27.335 ;
        RECT 151.865 26.055 153.680 28.435 ;
        RECT 157.025 28.195 157.255 28.230 ;
        RECT 157.880 28.195 158.580 29.165 ;
        RECT 157.025 26.285 158.580 28.195 ;
        RECT 157.025 26.230 157.255 26.285 ;
        RECT 149.265 26.025 156.895 26.055 ;
        RECT 149.015 25.795 156.975 26.025 ;
        RECT 144.195 23.705 144.425 25.675 ;
        RECT 146.745 25.005 146.975 25.675 ;
        RECT 146.745 24.725 149.610 25.005 ;
        RECT 146.745 24.635 157.030 24.725 ;
        RECT 146.745 23.705 146.975 24.635 ;
        RECT 149.170 24.485 157.030 24.635 ;
        RECT 149.110 24.255 157.110 24.485 ;
        RECT 148.675 23.765 148.905 24.205 ;
        RECT 157.315 24.195 157.545 24.205 ;
        RECT 149.395 23.765 150.395 23.835 ;
        RECT 157.315 23.765 157.550 24.195 ;
        RECT 144.585 23.425 146.585 23.655 ;
        RECT 144.675 23.185 146.500 23.425 ;
        RECT 143.000 22.695 146.500 23.185 ;
        RECT 143.000 17.860 143.875 22.695 ;
        RECT 144.675 22.515 146.500 22.695 ;
        RECT 148.675 22.875 157.550 23.765 ;
        RECT 144.585 22.285 146.585 22.515 ;
        RECT 148.675 22.245 148.905 22.875 ;
        RECT 149.395 22.820 150.395 22.875 ;
        RECT 157.315 22.310 157.550 22.875 ;
        RECT 157.315 22.245 157.545 22.310 ;
        RECT 144.195 20.800 144.425 22.235 ;
        RECT 146.745 20.800 146.975 22.235 ;
        RECT 149.110 21.965 157.110 22.195 ;
        RECT 149.180 21.840 157.010 21.965 ;
        RECT 149.200 21.055 157.000 21.840 ;
        RECT 149.110 20.825 157.110 21.055 ;
        RECT 144.195 19.460 146.975 20.800 ;
        RECT 148.675 20.750 148.905 20.775 ;
        RECT 144.195 18.275 144.425 19.460 ;
        RECT 144.770 18.225 146.365 19.460 ;
        RECT 146.745 18.570 146.975 19.460 ;
        RECT 148.670 20.305 148.905 20.750 ;
        RECT 157.315 20.750 157.545 20.775 ;
        RECT 148.670 20.295 149.085 20.305 ;
        RECT 149.225 20.295 150.225 20.365 ;
        RECT 148.670 20.290 150.225 20.295 ;
        RECT 150.635 20.290 152.255 20.295 ;
        RECT 157.315 20.290 157.550 20.750 ;
        RECT 148.670 19.400 157.550 20.290 ;
        RECT 148.670 19.385 150.225 19.400 ;
        RECT 150.635 19.395 152.255 19.400 ;
        RECT 148.670 19.295 149.085 19.385 ;
        RECT 149.225 19.335 150.225 19.385 ;
        RECT 148.670 18.865 148.905 19.295 ;
        RECT 148.675 18.815 148.905 18.865 ;
        RECT 157.315 18.865 157.550 19.400 ;
        RECT 157.315 18.815 157.545 18.865 ;
        RECT 149.110 18.570 157.110 18.765 ;
        RECT 146.745 18.535 157.110 18.570 ;
        RECT 146.745 18.390 157.030 18.535 ;
        RECT 146.745 18.375 149.245 18.390 ;
        RECT 146.745 18.275 146.975 18.375 ;
        RECT 144.585 17.995 146.585 18.225 ;
        RECT 157.880 18.115 158.580 26.285 ;
        RECT 152.955 17.985 153.230 18.055 ;
        RECT 147.260 17.860 153.230 17.985 ;
        RECT 143.000 17.845 144.405 17.860 ;
        RECT 146.750 17.845 153.230 17.860 ;
        RECT 143.000 17.795 153.230 17.845 ;
        RECT 143.000 17.670 147.450 17.795 ;
        RECT 152.955 17.720 153.230 17.795 ;
        RECT 143.000 12.390 143.875 17.670 ;
        RECT 145.825 17.365 149.610 17.370 ;
        RECT 145.825 17.300 153.060 17.365 ;
        RECT 144.645 17.175 153.060 17.300 ;
        RECT 144.645 17.085 153.105 17.175 ;
        RECT 144.585 17.075 153.105 17.085 ;
        RECT 144.585 16.855 146.585 17.075 ;
        RECT 149.105 16.945 153.105 17.075 ;
        RECT 144.195 15.425 144.425 16.805 ;
        RECT 146.745 15.425 146.975 16.805 ;
        RECT 144.195 14.470 146.975 15.425 ;
        RECT 144.195 12.845 144.425 14.470 ;
        RECT 146.745 12.845 146.975 14.470 ;
        RECT 148.670 15.640 148.900 16.895 ;
        RECT 150.340 15.640 151.725 16.945 ;
        RECT 153.310 15.640 153.540 16.895 ;
        RECT 153.905 16.435 158.580 18.115 ;
        RECT 155.265 16.095 155.540 16.125 ;
        RECT 155.250 15.840 155.580 16.095 ;
        RECT 155.265 15.820 155.555 15.840 ;
        RECT 155.265 15.790 155.540 15.820 ;
        RECT 148.670 15.570 153.540 15.640 ;
        RECT 155.075 15.570 155.305 15.615 ;
        RECT 148.670 14.295 153.545 15.570 ;
        RECT 148.670 12.935 148.900 14.295 ;
        RECT 153.310 12.935 153.545 14.295 ;
        RECT 144.585 12.565 146.585 12.795 ;
        RECT 144.650 12.390 146.520 12.565 ;
        RECT 143.000 11.835 146.520 12.390 ;
        RECT 143.000 6.730 143.875 11.835 ;
        RECT 144.650 11.655 146.520 11.835 ;
        RECT 144.585 11.425 146.585 11.655 ;
        RECT 148.710 11.465 148.870 12.935 ;
        RECT 153.340 12.925 153.545 12.935 ;
        RECT 149.105 12.655 153.105 12.885 ;
        RECT 149.185 12.410 153.010 12.655 ;
        RECT 155.065 12.410 155.305 15.570 ;
        RECT 149.185 11.920 155.305 12.410 ;
        RECT 149.185 11.745 153.010 11.920 ;
        RECT 149.105 11.515 153.105 11.745 ;
        RECT 144.195 9.980 144.425 11.375 ;
        RECT 146.745 9.980 146.975 11.375 ;
        RECT 144.195 9.025 146.975 9.980 ;
        RECT 144.195 7.415 144.425 9.025 ;
        RECT 146.745 7.415 146.975 9.025 ;
        RECT 148.670 10.090 148.900 11.465 ;
        RECT 153.310 11.350 153.540 11.465 ;
        RECT 153.310 10.715 153.545 11.350 ;
        RECT 155.065 10.715 155.305 11.920 ;
        RECT 153.310 10.090 153.540 10.715 ;
        RECT 155.075 10.615 155.305 10.715 ;
        RECT 155.515 15.600 155.745 15.615 ;
        RECT 156.165 15.600 156.645 16.435 ;
        RECT 155.515 10.675 156.655 15.600 ;
        RECT 157.880 12.510 158.580 16.435 ;
        RECT 157.420 12.460 158.580 12.510 ;
        RECT 157.420 11.775 158.620 12.460 ;
        RECT 157.420 11.690 158.580 11.775 ;
        RECT 155.515 10.615 155.745 10.675 ;
        RECT 155.265 10.405 155.555 10.410 ;
        RECT 155.250 10.150 155.580 10.405 ;
        RECT 148.670 8.745 153.540 10.090 ;
        RECT 148.670 7.505 148.900 8.745 ;
        RECT 153.310 7.505 153.540 8.745 ;
        RECT 144.585 7.340 146.585 7.365 ;
        RECT 149.105 7.340 153.105 7.455 ;
        RECT 144.585 7.265 146.590 7.340 ;
        RECT 147.125 7.265 153.105 7.340 ;
        RECT 144.585 7.225 153.105 7.265 ;
        RECT 144.585 7.135 153.040 7.225 ;
        RECT 144.640 7.000 153.040 7.135 ;
        RECT 143.000 6.290 144.860 6.730 ;
        RECT 143.000 6.280 145.850 6.290 ;
        RECT 143.000 5.935 146.520 6.280 ;
        RECT 143.000 4.310 144.860 5.935 ;
        RECT 145.660 5.785 146.520 5.935 ;
        RECT 145.155 5.595 145.405 5.610 ;
        RECT 145.155 5.305 145.430 5.595 ;
        RECT 145.590 5.555 146.590 5.785 ;
        RECT 147.010 5.690 147.280 7.000 ;
        RECT 157.880 6.570 158.580 11.690 ;
        RECT 152.300 6.235 158.580 6.570 ;
        RECT 149.185 6.095 158.580 6.235 ;
        RECT 149.185 5.870 153.045 6.095 ;
        RECT 145.155 5.275 145.405 5.305 ;
        RECT 145.590 5.115 146.590 5.345 ;
        RECT 146.735 5.270 148.925 5.690 ;
        RECT 149.120 5.640 153.120 5.870 ;
        RECT 153.355 5.680 153.605 5.700 ;
        RECT 149.120 5.200 153.120 5.430 ;
        RECT 153.325 5.390 153.605 5.680 ;
        RECT 153.355 5.365 153.605 5.390 ;
        RECT 145.660 4.975 146.545 5.115 ;
        RECT 149.170 5.035 153.095 5.200 ;
        RECT 146.730 4.975 153.095 5.035 ;
        RECT 145.660 4.920 153.095 4.975 ;
        RECT 145.660 4.850 149.540 4.920 ;
        RECT 146.215 4.735 149.540 4.850 ;
        RECT 157.880 4.770 158.580 6.095 ;
        RECT 143.000 4.265 145.385 4.310 ;
        RECT 127.665 2.560 132.730 2.630 ;
        RECT 129.205 2.555 132.730 2.560 ;
        RECT 130.415 2.000 131.415 2.555 ;
        RECT 143.000 2.535 143.875 4.265 ;
        RECT 144.240 3.990 145.385 4.265 ;
        RECT 147.570 4.105 147.975 4.735 ;
        RECT 156.575 4.235 158.580 4.770 ;
        RECT 144.240 3.925 146.490 3.990 ;
        RECT 144.680 3.760 146.490 3.925 ;
        RECT 144.165 3.570 144.415 3.595 ;
        RECT 144.165 3.280 144.435 3.570 ;
        RECT 144.595 3.530 146.595 3.760 ;
        RECT 147.555 3.740 147.980 4.105 ;
        RECT 149.220 4.090 158.580 4.235 ;
        RECT 149.220 3.845 157.075 4.090 ;
        RECT 144.165 3.260 144.415 3.280 ;
        RECT 144.595 3.090 146.595 3.320 ;
        RECT 146.745 3.230 148.935 3.740 ;
        RECT 149.125 3.615 157.125 3.845 ;
        RECT 157.355 3.655 157.605 3.670 ;
        RECT 146.745 3.225 147.445 3.230 ;
        RECT 148.445 3.225 148.935 3.230 ;
        RECT 149.125 3.175 157.125 3.405 ;
        RECT 157.330 3.365 157.605 3.655 ;
        RECT 157.355 3.335 157.605 3.365 ;
        RECT 144.665 2.925 146.530 3.090 ;
        RECT 147.415 2.925 148.415 3.000 ;
        RECT 149.200 2.925 157.050 3.175 ;
        RECT 144.665 2.630 157.050 2.925 ;
        RECT 157.880 2.690 158.580 4.090 ;
        RECT 144.665 2.560 149.730 2.630 ;
        RECT 146.205 2.555 149.730 2.560 ;
        RECT 147.415 2.000 148.415 2.555 ;
        RECT 60.850 1.970 80.025 2.000 ;
        RECT 60.850 1.950 61.170 1.970 ;
        RECT 56.085 1.510 56.345 1.830 ;
        RECT 58.955 1.605 59.215 1.925 ;
        RECT 60.245 1.770 60.625 1.935 ;
        RECT 60.225 1.635 60.625 1.770 ;
        RECT 96.815 1.635 97.020 2.000 ;
        RECT 56.120 0.510 56.310 1.510 ;
        RECT 59.000 0.875 59.170 1.605 ;
        RECT 59.575 1.215 59.835 1.475 ;
        RECT 60.225 1.450 97.020 1.635 ;
        RECT 60.245 1.430 97.020 1.450 ;
        RECT 113.825 1.215 114.010 2.000 ;
        RECT 59.575 1.155 114.010 1.215 ;
        RECT 59.610 1.030 114.010 1.155 ;
        RECT 130.830 0.875 131.000 2.000 ;
        RECT 59.000 0.705 131.000 0.875 ;
        RECT 147.820 0.510 148.010 2.000 ;
        RECT 56.120 0.320 148.010 0.510 ;
      LAYER met2 ;
        RECT 21.600 224.290 144.190 224.300 ;
        RECT 21.565 224.010 144.190 224.290 ;
        RECT 21.600 224.000 144.190 224.010 ;
        RECT 22.255 223.420 94.425 223.430 ;
        RECT 22.220 223.140 94.425 223.420 ;
        RECT 138.760 223.270 157.465 223.460 ;
        RECT 22.255 223.130 94.425 223.140 ;
        RECT 135.500 223.050 135.890 223.095 ;
        RECT 135.500 222.835 157.020 223.050 ;
        RECT 135.500 222.795 135.890 222.835 ;
        RECT 23.125 222.625 91.695 222.635 ;
        RECT 23.090 222.345 91.695 222.625 ;
        RECT 132.730 222.595 133.120 222.645 ;
        RECT 132.730 222.395 156.565 222.595 ;
        RECT 132.730 222.345 133.120 222.395 ;
        RECT 23.125 222.335 91.695 222.345 ;
        RECT 129.915 222.165 130.305 222.195 ;
        RECT 20.755 221.950 88.945 221.960 ;
        RECT 20.720 221.670 88.945 221.950 ;
        RECT 129.915 221.925 156.095 222.165 ;
        RECT 129.915 221.895 130.305 221.925 ;
        RECT 20.755 221.660 88.945 221.670 ;
        RECT 127.235 221.645 127.625 221.690 ;
        RECT 127.235 221.435 155.630 221.645 ;
        RECT 127.235 221.390 127.625 221.435 ;
        RECT 19.995 221.195 86.155 221.205 ;
        RECT 19.960 220.915 86.155 221.195 ;
        RECT 124.485 221.180 124.875 221.230 ;
        RECT 124.485 220.980 155.205 221.180 ;
        RECT 124.485 220.930 124.875 220.980 ;
        RECT 19.995 220.905 86.155 220.915 ;
        RECT 121.720 220.760 122.020 220.840 ;
        RECT 23.995 220.640 83.400 220.650 ;
        RECT 23.960 220.360 83.400 220.640 ;
        RECT 121.720 220.525 154.810 220.760 ;
        RECT 121.720 220.450 122.020 220.525 ;
        RECT 23.995 220.350 83.400 220.360 ;
        RECT 118.960 220.290 119.350 220.320 ;
        RECT 118.960 220.050 154.340 220.290 ;
        RECT 19.215 220.015 20.605 220.040 ;
        RECT 19.190 219.990 20.605 220.015 ;
        RECT 80.235 219.990 80.625 220.025 ;
        RECT 118.960 220.020 119.350 220.050 ;
        RECT 19.190 219.760 80.625 219.990 ;
        RECT 19.190 219.735 20.605 219.760 ;
        RECT 19.215 219.715 20.605 219.735 ;
        RECT 80.235 219.725 80.625 219.760 ;
        RECT 105.095 219.700 105.485 219.765 ;
        RECT 105.095 219.530 153.815 219.700 ;
        RECT 105.095 219.465 105.485 219.530 ;
        RECT 18.570 219.395 19.920 219.405 ;
        RECT 18.535 219.370 19.920 219.395 ;
        RECT 77.495 219.370 77.885 219.405 ;
        RECT 18.535 219.140 77.885 219.370 ;
        RECT 18.535 219.115 19.920 219.140 ;
        RECT 18.570 219.105 19.920 219.115 ;
        RECT 77.495 219.105 77.885 219.140 ;
        RECT 102.365 219.240 102.755 219.305 ;
        RECT 102.365 219.070 153.345 219.240 ;
        RECT 102.365 219.005 102.755 219.070 ;
        RECT 17.785 218.910 18.425 218.925 ;
        RECT 17.755 218.895 18.425 218.910 ;
        RECT 74.765 218.895 75.155 218.925 ;
        RECT 17.755 218.650 75.155 218.895 ;
        RECT 17.755 218.630 18.425 218.650 ;
        RECT 17.785 218.615 18.425 218.630 ;
        RECT 74.765 218.625 75.155 218.650 ;
        RECT 24.730 218.325 25.680 218.335 ;
        RECT 24.695 218.300 25.680 218.325 ;
        RECT 72.030 218.300 72.420 218.340 ;
        RECT 24.695 218.075 72.420 218.300 ;
        RECT 24.695 218.045 25.680 218.075 ;
        RECT 24.730 218.035 25.680 218.045 ;
        RECT 72.030 218.040 72.420 218.075 ;
        RECT 25.385 217.725 69.640 217.735 ;
        RECT 25.350 217.445 69.640 217.725 ;
        RECT 25.385 217.435 69.640 217.445 ;
        RECT 17.115 217.320 17.395 217.355 ;
        RECT 17.105 217.285 18.555 217.320 ;
        RECT 17.105 217.055 66.810 217.285 ;
        RECT 17.105 217.020 18.555 217.055 ;
        RECT 17.115 216.985 17.395 217.020 ;
        RECT 66.350 216.995 66.810 217.055 ;
        RECT 66.350 216.875 66.845 216.995 ;
        RECT 16.425 216.715 64.155 216.725 ;
        RECT 16.390 216.435 64.155 216.715 ;
        RECT 66.545 216.605 66.845 216.875 ;
        RECT 16.425 216.425 64.155 216.435 ;
        RECT 153.175 131.150 153.345 219.070 ;
        RECT 130.180 130.980 153.345 131.150 ;
        RECT 74.790 119.960 75.110 120.830 ;
        RECT 74.780 118.930 75.110 119.960 ;
        RECT 76.460 119.940 76.780 120.820 ;
        RECT 74.780 117.170 75.090 118.930 ;
        RECT 76.440 118.920 76.780 119.940 ;
        RECT 78.020 118.920 78.340 120.820 ;
        RECT 79.560 119.930 79.880 120.830 ;
        RECT 79.540 118.930 79.880 119.930 ;
        RECT 81.150 119.740 81.470 120.850 ;
        RECT 76.440 117.280 76.750 118.920 ;
        RECT 74.780 117.010 75.000 117.170 ;
        RECT 75.250 117.010 75.790 117.150 ;
        RECT 74.780 114.920 75.790 117.010 ;
        RECT 74.820 114.900 75.790 114.920 ;
        RECT 76.440 116.960 77.250 117.280 ;
        RECT 78.020 117.150 78.330 118.920 ;
        RECT 76.440 114.900 77.170 116.960 ;
        RECT 75.180 114.810 75.790 114.900 ;
        RECT 76.720 114.870 77.170 114.900 ;
        RECT 76.750 114.840 77.120 114.870 ;
        RECT 78.020 114.860 78.690 117.150 ;
        RECT 79.540 117.130 79.850 118.930 ;
        RECT 81.110 117.160 81.480 119.740 ;
        RECT 82.710 119.730 83.030 120.820 ;
        RECT 84.300 119.770 84.620 120.840 ;
        RECT 85.900 120.080 86.180 120.830 ;
        RECT 82.690 117.190 83.060 119.730 ;
        RECT 79.540 114.890 80.200 117.130 ;
        RECT 78.140 114.800 78.690 114.860 ;
        RECT 79.650 114.780 80.200 114.890 ;
        RECT 81.110 114.810 81.660 117.160 ;
        RECT 82.590 114.840 83.140 117.190 ;
        RECT 84.300 117.180 84.650 119.770 ;
        RECT 85.880 117.190 86.180 120.080 ;
        RECT 130.180 118.075 130.350 130.980 ;
        RECT 153.645 130.705 153.815 219.530 ;
        RECT 136.655 130.535 153.815 130.705 ;
        RECT 136.655 118.105 136.825 130.535 ;
        RECT 154.100 130.340 154.340 220.050 ;
        RECT 146.230 130.100 154.340 130.340 ;
        RECT 146.230 119.120 146.470 130.100 ;
        RECT 154.575 129.790 154.810 220.525 ;
        RECT 147.735 129.555 154.810 129.790 ;
        RECT 147.735 119.170 147.970 129.555 ;
        RECT 155.005 129.315 155.205 220.980 ;
        RECT 149.260 129.115 155.205 129.315 ;
        RECT 149.260 119.170 149.460 129.115 ;
        RECT 155.420 128.895 155.630 221.435 ;
        RECT 150.865 128.685 155.630 128.895 ;
        RECT 150.865 119.200 151.075 128.685 ;
        RECT 155.855 128.490 156.095 221.925 ;
        RECT 152.400 128.250 156.095 128.490 ;
        RECT 145.820 118.860 146.880 119.120 ;
        RECT 147.320 118.910 148.380 119.170 ;
        RECT 148.830 118.910 149.890 119.170 ;
        RECT 150.440 118.940 151.500 119.200 ;
        RECT 152.400 119.170 152.640 128.250 ;
        RECT 156.365 128.100 156.565 222.395 ;
        RECT 154.040 127.900 156.565 128.100 ;
        RECT 154.040 119.200 154.240 127.900 ;
        RECT 156.805 127.720 157.020 222.835 ;
        RECT 155.605 127.505 157.020 127.720 ;
        RECT 151.990 118.910 153.050 119.170 ;
        RECT 153.610 118.940 154.670 119.200 ;
        RECT 155.605 119.170 155.820 127.505 ;
        RECT 157.275 119.190 157.465 223.270 ;
        RECT 155.180 118.910 156.240 119.170 ;
        RECT 156.840 118.930 157.900 119.190 ;
        RECT 84.040 114.930 84.650 117.180 ;
        RECT 84.040 114.830 84.590 114.930 ;
        RECT 85.540 114.900 86.180 117.190 ;
        RECT 120.375 117.905 130.350 118.075 ;
        RECT 85.540 114.840 86.090 114.900 ;
        RECT 120.375 104.425 120.545 117.905 ;
        RECT 130.180 117.840 130.350 117.905 ;
        RECT 132.745 117.935 136.825 118.105 ;
        RECT 123.570 115.565 124.045 115.595 ;
        RECT 126.360 115.565 126.680 115.595 ;
        RECT 129.120 115.565 129.440 115.595 ;
        RECT 123.570 115.365 129.440 115.565 ;
        RECT 123.570 115.335 124.045 115.365 ;
        RECT 126.360 115.335 126.680 115.365 ;
        RECT 129.120 115.335 129.440 115.365 ;
        RECT 123.685 105.850 123.945 106.170 ;
        RECT 124.775 105.895 125.035 106.215 ;
        RECT 121.880 104.425 122.200 104.470 ;
        RECT 120.375 104.255 122.200 104.425 ;
        RECT 121.880 104.210 122.200 104.255 ;
        RECT 123.710 103.075 123.920 105.850 ;
        RECT 124.780 103.115 125.030 105.895 ;
        RECT 126.350 105.885 126.610 106.205 ;
        RECT 127.915 105.930 128.175 106.250 ;
        RECT 126.350 103.140 126.605 105.885 ;
        RECT 127.930 104.590 128.155 105.930 ;
        RECT 129.090 105.780 129.350 106.100 ;
        RECT 127.865 104.230 128.245 104.590 ;
        RECT 123.590 102.815 124.045 103.075 ;
        RECT 124.255 102.855 125.560 103.115 ;
        RECT 125.825 102.880 127.130 103.140 ;
        RECT 127.930 103.095 128.155 104.230 ;
        RECT 129.105 103.145 129.330 105.780 ;
        RECT 130.330 105.265 130.650 105.280 ;
        RECT 130.330 105.035 132.195 105.265 ;
        RECT 130.330 105.020 130.650 105.035 ;
        RECT 127.390 102.835 128.695 103.095 ;
        RECT 129.005 102.885 129.430 103.145 ;
        RECT 123.590 98.590 124.045 98.615 ;
        RECT 126.315 98.590 126.635 98.615 ;
        RECT 129.090 98.590 129.410 98.615 ;
        RECT 123.590 98.380 129.410 98.590 ;
        RECT 123.590 98.355 124.045 98.380 ;
        RECT 126.315 98.355 126.635 98.380 ;
        RECT 129.090 98.355 129.410 98.380 ;
        RECT 130.190 95.920 130.470 103.630 ;
        RECT 131.965 96.670 132.195 105.035 ;
        RECT 132.745 104.455 132.915 117.935 ;
        RECT 136.655 117.840 136.825 117.935 ;
        RECT 134.290 104.455 134.610 104.500 ;
        RECT 132.745 104.285 134.610 104.455 ;
        RECT 134.290 104.240 134.610 104.285 ;
        RECT 142.790 103.270 143.050 103.590 ;
        RECT 142.805 96.670 143.035 103.270 ;
        RECT 143.870 99.550 144.670 114.830 ;
        RECT 143.840 98.750 144.700 99.550 ;
        RECT 150.075 98.560 150.645 98.840 ;
        RECT 150.075 98.280 158.800 98.560 ;
        RECT 150.075 98.060 150.645 98.280 ;
        RECT 131.965 96.440 152.375 96.670 ;
        RECT 130.190 95.640 150.070 95.920 ;
        RECT 117.325 95.350 117.715 95.390 ;
        RECT 117.325 95.130 148.455 95.350 ;
        RECT 117.325 95.090 117.715 95.130 ;
        RECT 118.300 94.555 147.040 94.900 ;
        RECT 119.225 94.215 119.615 94.245 ;
        RECT 119.225 93.970 145.550 94.215 ;
        RECT 119.225 93.945 119.615 93.970 ;
        RECT 120.330 93.765 120.720 93.810 ;
        RECT 120.330 93.555 141.040 93.765 ;
        RECT 120.330 93.510 120.720 93.555 ;
        RECT 121.235 93.270 121.625 93.295 ;
        RECT 121.235 93.020 139.605 93.270 ;
        RECT 121.235 92.995 121.625 93.020 ;
        RECT 122.075 92.825 122.465 92.830 ;
        RECT 122.075 92.535 138.130 92.825 ;
        RECT 122.075 92.530 122.465 92.535 ;
        RECT 127.300 92.075 127.900 92.200 ;
        RECT 127.200 91.700 127.900 92.075 ;
        RECT 130.300 92.005 130.800 92.200 ;
        RECT 130.190 91.700 130.800 92.005 ;
        RECT 133.300 91.985 133.800 92.200 ;
        RECT 133.205 91.700 133.800 91.985 ;
        RECT 136.200 91.905 136.700 92.100 ;
        RECT 127.200 91.685 127.500 91.700 ;
        RECT 69.130 89.040 70.440 90.340 ;
        RECT 130.190 90.270 130.515 91.700 ;
        RECT 133.205 91.695 133.750 91.700 ;
        RECT 133.360 91.690 133.750 91.695 ;
        RECT 136.135 91.670 136.700 91.905 ;
        RECT 136.200 91.600 136.700 91.670 ;
        RECT 136.360 90.600 136.595 91.600 ;
        RECT 125.120 89.945 130.515 90.270 ;
        RECT 134.020 90.365 136.595 90.600 ;
        RECT 128.800 89.370 129.300 89.500 ;
        RECT 126.215 89.070 129.300 89.370 ;
        RECT 131.800 89.075 132.300 89.300 ;
        RECT 128.800 89.000 129.300 89.070 ;
        RECT 131.710 88.800 132.300 89.075 ;
        RECT 124.025 88.505 124.415 88.515 ;
        RECT 131.710 88.505 131.990 88.800 ;
        RECT 124.025 88.225 131.990 88.505 ;
        RECT 124.025 88.215 124.415 88.225 ;
        RECT 134.020 87.300 134.255 90.365 ;
        RECT 134.800 89.000 135.300 89.500 ;
        RECT 137.840 89.400 138.130 92.535 ;
        RECT 139.355 92.100 139.605 93.020 ;
        RECT 139.200 91.600 139.700 92.100 ;
        RECT 134.900 88.115 135.150 89.000 ;
        RECT 137.700 88.900 138.200 89.400 ;
        RECT 140.830 89.300 141.040 93.555 ;
        RECT 145.305 92.100 145.550 93.970 ;
        RECT 142.200 91.600 142.700 92.100 ;
        RECT 145.200 91.600 145.700 92.100 ;
        RECT 137.840 88.895 138.130 88.900 ;
        RECT 140.700 88.800 141.200 89.300 ;
        RECT 134.875 87.725 135.175 88.115 ;
        RECT 133.990 86.910 134.290 87.300 ;
        RECT 81.290 85.250 81.550 85.570 ;
        RECT 98.290 85.250 98.550 85.570 ;
        RECT 115.290 85.250 115.550 85.570 ;
        RECT 132.290 85.250 132.550 85.570 ;
        RECT 77.650 84.455 77.910 84.775 ;
        RECT 76.880 72.815 77.175 77.320 ;
        RECT 36.410 66.765 36.690 70.765 ;
        RECT 39.630 66.765 39.910 70.765 ;
        RECT 42.850 66.765 43.130 70.765 ;
        RECT 46.070 66.765 46.350 70.765 ;
        RECT 49.290 66.765 49.570 70.765 ;
        RECT 77.675 67.655 77.885 84.455 ;
        RECT 81.345 79.690 81.495 85.250 ;
        RECT 94.650 84.455 94.910 84.775 ;
        RECT 83.570 81.180 83.830 81.500 ;
        RECT 81.290 79.370 81.550 79.690 ;
        RECT 77.650 67.335 77.910 67.655 ;
        RECT 35.700 62.270 36.000 62.515 ;
        RECT 36.480 62.270 36.620 66.765 ;
        RECT 35.700 62.130 36.620 62.270 ;
        RECT 35.700 62.125 36.000 62.130 ;
        RECT 23.125 61.025 23.425 61.375 ;
        RECT 21.745 60.725 23.425 61.025 ;
        RECT 20.710 58.900 21.100 58.980 ;
        RECT 20.710 58.760 21.510 58.900 ;
        RECT 20.710 58.680 21.100 58.760 ;
        RECT 19.950 58.025 21.115 58.325 ;
        RECT 17.745 57.695 18.135 57.760 ;
        RECT 17.745 57.520 18.555 57.695 ;
        RECT 17.745 57.460 18.135 57.520 ;
        RECT 17.060 56.130 17.450 56.210 ;
        RECT 17.060 55.990 17.985 56.130 ;
        RECT 17.060 55.910 17.450 55.990 ;
        RECT 16.380 55.385 16.770 55.465 ;
        RECT 16.380 55.245 17.615 55.385 ;
        RECT 16.380 55.165 16.770 55.245 ;
        RECT 17.475 32.075 17.615 55.245 ;
        RECT 17.845 32.735 17.985 55.990 ;
        RECT 18.380 38.085 18.555 57.520 ;
        RECT 19.220 57.460 19.520 57.505 ;
        RECT 19.220 57.160 20.340 57.460 ;
        RECT 19.220 57.115 19.520 57.160 ;
        RECT 18.715 56.120 19.015 56.510 ;
        RECT 18.795 50.050 18.935 56.120 ;
        RECT 20.040 50.590 20.340 57.160 ;
        RECT 20.050 50.555 20.330 50.590 ;
        RECT 18.795 49.910 20.450 50.050 ;
        RECT 18.315 36.990 18.615 38.085 ;
        RECT 18.325 36.955 18.605 36.990 ;
        RECT 17.845 32.595 20.020 32.735 ;
        RECT 17.475 31.935 19.175 32.075 ;
        RECT 19.035 22.115 19.175 31.935 ;
        RECT 19.880 22.510 20.020 32.595 ;
        RECT 20.310 26.560 20.450 49.910 ;
        RECT 20.815 27.865 21.115 58.025 ;
        RECT 21.370 43.470 21.510 58.760 ;
        RECT 21.745 44.080 22.045 60.725 ;
        RECT 36.480 58.890 36.620 62.130 ;
        RECT 39.700 60.380 39.840 66.765 ;
        RECT 42.035 61.575 42.335 61.855 ;
        RECT 42.025 61.315 42.345 61.575 ;
        RECT 41.060 60.770 41.450 60.850 ;
        RECT 42.920 60.770 43.060 66.765 ;
        RECT 41.060 60.630 43.060 60.770 ;
        RECT 41.060 60.550 41.450 60.630 ;
        RECT 39.620 60.330 39.920 60.380 ;
        RECT 39.620 60.190 40.760 60.330 ;
        RECT 39.620 59.990 39.920 60.190 ;
        RECT 38.070 59.055 39.610 59.425 ;
        RECT 36.420 58.570 36.680 58.890 ;
        RECT 28.140 57.550 28.400 57.870 ;
        RECT 32.740 57.550 33.000 57.870 ;
        RECT 33.200 57.550 33.460 57.870 ;
        RECT 28.200 56.170 28.340 57.550 ;
        RECT 32.800 56.170 32.940 57.550 ;
        RECT 28.140 55.850 28.400 56.170 ;
        RECT 32.740 55.850 33.000 56.170 ;
        RECT 33.260 55.685 33.400 57.550 ;
        RECT 35.040 56.870 35.300 57.190 ;
        RECT 40.100 56.870 40.360 57.190 ;
        RECT 35.100 55.830 35.240 56.870 ;
        RECT 33.190 55.315 33.470 55.685 ;
        RECT 35.040 55.510 35.300 55.830 ;
        RECT 35.960 55.170 36.220 55.490 ;
        RECT 37.330 55.315 37.610 55.685 ;
        RECT 33.660 54.150 33.920 54.470 ;
        RECT 33.720 52.430 33.860 54.150 ;
        RECT 34.570 53.955 34.850 54.325 ;
        RECT 33.660 52.110 33.920 52.430 ;
        RECT 25.840 51.770 26.100 52.090 ;
        RECT 23.530 50.555 23.810 50.925 ;
        RECT 25.900 50.730 26.040 51.770 ;
        RECT 30.900 51.430 31.160 51.750 ;
        RECT 31.360 51.430 31.620 51.750 ;
        RECT 23.540 50.410 23.800 50.555 ;
        RECT 25.840 50.410 26.100 50.730 ;
        RECT 30.960 50.050 31.100 51.430 ;
        RECT 31.420 50.730 31.560 51.430 ;
        RECT 33.720 50.730 33.860 52.110 ;
        RECT 31.360 50.410 31.620 50.730 ;
        RECT 33.660 50.410 33.920 50.730 ;
        RECT 30.900 49.730 31.160 50.050 ;
        RECT 29.520 49.390 29.780 49.710 ;
        RECT 26.300 49.050 26.560 49.370 ;
        RECT 26.360 47.330 26.500 49.050 ;
        RECT 26.300 47.010 26.560 47.330 ;
        RECT 29.580 46.650 29.720 49.390 ;
        RECT 33.720 46.990 33.860 50.410 ;
        RECT 30.900 46.670 31.160 46.990 ;
        RECT 33.660 46.670 33.920 46.990 ;
        RECT 29.520 46.330 29.780 46.650 ;
        RECT 24.000 45.990 24.260 46.310 ;
        RECT 28.600 45.990 28.860 46.310 ;
        RECT 24.060 44.950 24.200 45.990 ;
        RECT 24.000 44.630 24.260 44.950 ;
        RECT 21.710 43.800 22.080 44.080 ;
        RECT 21.745 43.790 22.045 43.800 ;
        RECT 23.530 43.755 23.810 44.125 ;
        RECT 21.370 43.330 22.250 43.470 ;
        RECT 20.815 27.805 21.455 27.865 ;
        RECT 20.815 27.435 21.510 27.805 ;
        RECT 20.815 27.290 21.500 27.435 ;
        RECT 20.815 27.265 21.455 27.290 ;
        RECT 20.310 26.420 21.895 26.560 ;
        RECT 21.755 22.970 21.895 26.420 ;
        RECT 22.110 23.400 22.250 43.330 ;
        RECT 23.600 39.850 23.740 43.755 ;
        RECT 24.000 43.270 24.260 43.590 ;
        RECT 24.060 41.890 24.200 43.270 ;
        RECT 28.660 42.570 28.800 45.990 ;
        RECT 28.600 42.250 28.860 42.570 ;
        RECT 24.000 41.570 24.260 41.890 ;
        RECT 23.540 39.530 23.800 39.850 ;
        RECT 24.060 39.170 24.200 41.570 ;
        RECT 29.060 40.550 29.320 40.870 ;
        RECT 29.120 39.850 29.260 40.550 ;
        RECT 29.060 39.530 29.320 39.850 ;
        RECT 24.000 38.850 24.260 39.170 ;
        RECT 29.580 38.830 29.720 46.330 ;
        RECT 30.960 44.610 31.100 46.670 ;
        RECT 34.640 44.950 34.780 53.955 ;
        RECT 36.020 53.450 36.160 55.170 ;
        RECT 35.960 53.130 36.220 53.450 ;
        RECT 35.960 50.410 36.220 50.730 ;
        RECT 36.880 50.410 37.140 50.730 ;
        RECT 36.020 47.330 36.160 50.410 ;
        RECT 36.940 48.010 37.080 50.410 ;
        RECT 36.880 47.690 37.140 48.010 ;
        RECT 35.960 47.010 36.220 47.330 ;
        RECT 34.580 44.630 34.840 44.950 ;
        RECT 30.900 44.290 31.160 44.610 ;
        RECT 36.940 42.570 37.080 47.690 ;
        RECT 37.400 42.570 37.540 55.315 ;
        RECT 38.070 53.615 39.610 53.985 ;
        RECT 40.160 52.430 40.300 56.870 ;
        RECT 40.620 54.810 40.760 60.190 ;
        RECT 42.920 58.890 43.060 60.630 ;
        RECT 46.140 60.270 46.280 66.765 ;
        RECT 49.360 60.700 49.500 66.765 ;
        RECT 56.650 64.155 56.930 64.525 ;
        RECT 53.890 60.755 54.170 61.125 ;
        RECT 49.090 60.440 49.500 60.700 ;
        RECT 46.110 59.950 46.370 60.270 ;
        RECT 42.860 58.570 43.120 58.890 ;
        RECT 41.020 58.230 41.280 58.550 ;
        RECT 40.560 54.490 40.820 54.810 ;
        RECT 41.080 53.450 41.220 58.230 ;
        RECT 46.140 57.870 46.280 59.950 ;
        RECT 49.360 58.890 49.500 60.440 ;
        RECT 49.300 58.570 49.560 58.890 ;
        RECT 47.920 58.230 48.180 58.550 ;
        RECT 43.320 57.550 43.580 57.870 ;
        RECT 46.080 57.550 46.340 57.870 ;
        RECT 41.370 56.335 42.910 56.705 ;
        RECT 43.380 56.170 43.520 57.550 ;
        RECT 43.780 56.870 44.040 57.190 ;
        RECT 43.320 55.850 43.580 56.170 ;
        RECT 43.840 55.830 43.980 56.870 ;
        RECT 43.780 55.510 44.040 55.830 ;
        RECT 47.980 55.490 48.120 58.230 ;
        RECT 53.960 57.870 54.100 60.755 ;
        RECT 56.720 59.785 56.860 64.155 ;
        RECT 60.730 60.755 61.030 61.145 ;
        RECT 75.085 61.095 75.580 61.645 ;
        RECT 56.720 59.590 58.925 59.785 ;
        RECT 60.775 59.685 60.980 60.755 ;
        RECT 74.260 60.140 75.810 61.095 ;
        RECT 56.720 57.870 56.860 59.590 ;
        RECT 58.730 58.595 58.925 59.590 ;
        RECT 60.065 59.180 60.385 59.440 ;
        RECT 60.745 59.365 61.005 59.685 ;
        RECT 59.360 58.640 59.620 58.960 ;
        RECT 58.695 58.275 58.955 58.595 ;
        RECT 51.140 57.550 51.400 57.870 ;
        RECT 53.900 57.550 54.160 57.870 ;
        RECT 55.280 57.725 55.540 57.870 ;
        RECT 49.760 56.870 50.020 57.190 ;
        RECT 44.700 55.170 44.960 55.490 ;
        RECT 46.080 55.170 46.340 55.490 ;
        RECT 47.920 55.170 48.180 55.490 ;
        RECT 41.480 54.830 41.740 55.150 ;
        RECT 41.020 53.130 41.280 53.450 ;
        RECT 41.540 52.430 41.680 54.830 ;
        RECT 44.240 54.150 44.500 54.470 ;
        RECT 44.300 52.770 44.440 54.150 ;
        RECT 44.240 52.450 44.500 52.770 ;
        RECT 44.760 52.430 44.900 55.170 ;
        RECT 45.620 54.830 45.880 55.150 ;
        RECT 40.100 52.110 40.360 52.430 ;
        RECT 40.560 52.110 40.820 52.430 ;
        RECT 41.480 52.110 41.740 52.430 ;
        RECT 43.320 52.110 43.580 52.430 ;
        RECT 43.780 52.110 44.040 52.430 ;
        RECT 44.700 52.110 44.960 52.430 ;
        RECT 40.100 51.430 40.360 51.750 ;
        RECT 38.070 48.175 39.610 48.545 ;
        RECT 38.070 42.735 39.610 43.105 ;
        RECT 36.880 42.250 37.140 42.570 ;
        RECT 37.340 42.250 37.600 42.570 ;
        RECT 31.820 41.230 32.080 41.550 ;
        RECT 29.060 38.510 29.320 38.830 ;
        RECT 29.520 38.510 29.780 38.830 ;
        RECT 24.000 38.170 24.260 38.490 ;
        RECT 23.530 36.955 23.810 37.325 ;
        RECT 23.600 33.050 23.740 36.955 ;
        RECT 24.060 36.450 24.200 38.170 ;
        RECT 26.300 37.830 26.560 38.150 ;
        RECT 24.000 36.130 24.260 36.450 ;
        RECT 26.360 35.770 26.500 37.830 ;
        RECT 26.300 35.450 26.560 35.770 ;
        RECT 24.000 33.070 24.260 33.390 ;
        RECT 23.540 32.730 23.800 33.050 ;
        RECT 24.060 31.690 24.200 33.070 ;
        RECT 29.120 33.050 29.260 38.510 ;
        RECT 31.880 37.130 32.020 41.230 ;
        RECT 36.940 39.510 37.080 42.250 ;
        RECT 40.160 41.550 40.300 51.430 ;
        RECT 40.620 50.730 40.760 52.110 ;
        RECT 41.370 50.895 42.910 51.265 ;
        RECT 40.560 50.410 40.820 50.730 ;
        RECT 40.560 49.730 40.820 50.050 ;
        RECT 40.620 43.590 40.760 49.730 ;
        RECT 41.020 48.710 41.280 49.030 ;
        RECT 41.080 44.690 41.220 48.710 ;
        RECT 43.380 48.010 43.520 52.110 ;
        RECT 43.320 47.690 43.580 48.010 ;
        RECT 43.840 47.410 43.980 52.110 ;
        RECT 45.680 50.390 45.820 54.830 ;
        RECT 46.140 53.450 46.280 55.170 ;
        RECT 47.000 54.150 47.260 54.470 ;
        RECT 46.080 53.130 46.340 53.450 ;
        RECT 46.140 52.850 46.280 53.130 ;
        RECT 46.140 52.710 46.740 52.850 ;
        RECT 46.080 51.770 46.340 52.090 ;
        RECT 45.620 50.070 45.880 50.390 ;
        RECT 44.240 49.390 44.500 49.710 ;
        RECT 43.380 47.270 43.980 47.410 ;
        RECT 43.380 46.310 43.520 47.270 ;
        RECT 44.300 46.990 44.440 49.390 ;
        RECT 44.700 47.350 44.960 47.670 ;
        RECT 44.240 46.670 44.500 46.990 ;
        RECT 43.780 46.330 44.040 46.650 ;
        RECT 43.320 45.990 43.580 46.310 ;
        RECT 41.370 45.455 42.910 45.825 ;
        RECT 41.080 44.550 41.680 44.690 ;
        RECT 41.020 43.950 41.280 44.270 ;
        RECT 40.560 43.270 40.820 43.590 ;
        RECT 37.340 41.230 37.600 41.550 ;
        RECT 40.100 41.230 40.360 41.550 ;
        RECT 37.400 39.850 37.540 41.230 ;
        RECT 37.340 39.530 37.600 39.850 ;
        RECT 35.500 39.190 35.760 39.510 ;
        RECT 36.880 39.190 37.140 39.510 ;
        RECT 31.820 36.810 32.080 37.130 ;
        RECT 30.900 35.790 31.160 36.110 ;
        RECT 29.060 32.730 29.320 33.050 ;
        RECT 28.600 32.390 28.860 32.710 ;
        RECT 24.000 31.370 24.260 31.690 ;
        RECT 24.060 28.290 24.200 31.370 ;
        RECT 26.760 30.010 27.020 30.330 ;
        RECT 26.820 28.970 26.960 30.010 ;
        RECT 28.660 28.970 28.800 32.390 ;
        RECT 29.120 28.970 29.260 32.730 ;
        RECT 30.960 31.010 31.100 35.790 ;
        RECT 31.880 33.730 32.020 36.810 ;
        RECT 31.820 33.410 32.080 33.730 ;
        RECT 35.560 33.390 35.700 39.190 ;
        RECT 36.880 38.170 37.140 38.490 ;
        RECT 36.940 35.770 37.080 38.170 ;
        RECT 38.070 37.295 39.610 37.665 ;
        RECT 36.880 35.450 37.140 35.770 ;
        RECT 31.360 33.070 31.620 33.390 ;
        RECT 35.500 33.070 35.760 33.390 ;
        RECT 30.900 30.690 31.160 31.010 ;
        RECT 31.420 28.970 31.560 33.070 ;
        RECT 26.760 28.650 27.020 28.970 ;
        RECT 28.600 28.650 28.860 28.970 ;
        RECT 29.060 28.650 29.320 28.970 ;
        RECT 31.360 28.650 31.620 28.970 ;
        RECT 33.660 28.650 33.920 28.970 ;
        RECT 24.000 27.970 24.260 28.290 ;
        RECT 33.720 25.230 33.860 28.650 ;
        RECT 35.560 27.950 35.700 33.070 ;
        RECT 40.100 32.390 40.360 32.710 ;
        RECT 38.070 31.855 39.610 32.225 ;
        RECT 40.160 28.970 40.300 32.390 ;
        RECT 40.620 30.670 40.760 43.270 ;
        RECT 41.080 41.550 41.220 43.950 ;
        RECT 41.540 42.230 41.680 44.550 ;
        RECT 41.480 41.910 41.740 42.230 ;
        RECT 41.020 41.230 41.280 41.550 ;
        RECT 41.370 40.015 42.910 40.385 ;
        RECT 43.380 38.830 43.520 45.990 ;
        RECT 43.840 45.290 43.980 46.330 ;
        RECT 43.780 44.970 44.040 45.290 ;
        RECT 44.760 41.890 44.900 47.350 ;
        RECT 45.160 46.330 45.420 46.650 ;
        RECT 44.700 41.570 44.960 41.890 ;
        RECT 44.240 39.760 44.500 39.850 ;
        RECT 44.760 39.760 44.900 41.570 ;
        RECT 44.240 39.620 44.900 39.760 ;
        RECT 44.240 39.530 44.500 39.620 ;
        RECT 43.320 38.510 43.580 38.830 ;
        RECT 43.780 38.510 44.040 38.830 ;
        RECT 43.840 35.430 43.980 38.510 ;
        RECT 44.760 36.530 44.900 39.620 ;
        RECT 45.220 36.790 45.360 46.330 ;
        RECT 45.680 43.590 45.820 50.070 ;
        RECT 46.140 49.370 46.280 51.770 ;
        RECT 46.080 49.050 46.340 49.370 ;
        RECT 46.140 45.290 46.280 49.050 ;
        RECT 46.080 44.970 46.340 45.290 ;
        RECT 45.620 43.270 45.880 43.590 ;
        RECT 45.680 42.230 45.820 43.270 ;
        RECT 45.620 41.910 45.880 42.230 ;
        RECT 45.620 38.170 45.880 38.490 ;
        RECT 44.300 36.450 44.900 36.530 ;
        RECT 45.160 36.470 45.420 36.790 ;
        RECT 44.240 36.390 44.900 36.450 ;
        RECT 44.240 36.130 44.500 36.390 ;
        RECT 41.020 35.110 41.280 35.430 ;
        RECT 43.780 35.110 44.040 35.430 ;
        RECT 41.080 33.730 41.220 35.110 ;
        RECT 41.370 34.575 42.910 34.945 ;
        RECT 41.020 33.410 41.280 33.730 ;
        RECT 41.080 31.690 41.220 33.410 ;
        RECT 41.020 31.370 41.280 31.690 ;
        RECT 40.560 30.350 40.820 30.670 ;
        RECT 40.100 28.650 40.360 28.970 ;
        RECT 41.080 28.630 41.220 31.370 ;
        RECT 41.370 29.135 42.910 29.505 ;
        RECT 41.020 28.370 41.280 28.630 ;
        RECT 40.160 28.310 41.280 28.370 ;
        RECT 40.160 28.230 41.220 28.310 ;
        RECT 35.500 27.630 35.760 27.950 ;
        RECT 38.070 26.415 39.610 26.785 ;
        RECT 33.660 24.910 33.920 25.230 ;
        RECT 38.720 25.140 38.980 25.230 ;
        RECT 40.160 25.140 40.300 28.230 ;
        RECT 41.020 26.950 41.280 27.270 ;
        RECT 38.720 25.000 40.300 25.140 ;
        RECT 38.720 24.910 38.980 25.000 ;
        RECT 41.080 24.890 41.220 26.950 ;
        RECT 43.840 26.250 43.980 35.110 ;
        RECT 45.680 34.070 45.820 38.170 ;
        RECT 46.600 37.130 46.740 52.710 ;
        RECT 47.060 52.430 47.200 54.150 ;
        RECT 47.000 52.110 47.260 52.430 ;
        RECT 49.820 50.050 49.960 56.870 ;
        RECT 50.670 55.400 50.950 55.685 ;
        RECT 50.280 55.315 50.950 55.400 ;
        RECT 50.280 55.260 50.940 55.315 ;
        RECT 50.280 50.390 50.420 55.260 ;
        RECT 50.680 55.170 50.940 55.260 ;
        RECT 51.200 54.810 51.340 57.550 ;
        RECT 55.270 57.355 55.550 57.725 ;
        RECT 56.660 57.550 56.920 57.870 ;
        RECT 59.390 57.715 59.590 58.640 ;
        RECT 59.340 57.325 59.640 57.715 ;
        RECT 53.440 56.870 53.700 57.190 ;
        RECT 56.200 56.870 56.460 57.190 ;
        RECT 51.140 54.490 51.400 54.810 ;
        RECT 51.200 53.450 51.340 54.490 ;
        RECT 52.980 54.150 53.240 54.470 ;
        RECT 51.140 53.130 51.400 53.450 ;
        RECT 53.040 52.430 53.180 54.150 ;
        RECT 52.980 52.110 53.240 52.430 ;
        RECT 53.500 50.730 53.640 56.870 ;
        RECT 53.900 55.170 54.160 55.490 ;
        RECT 53.960 53.450 54.100 55.170 ;
        RECT 54.360 54.490 54.620 54.810 ;
        RECT 53.900 53.130 54.160 53.450 ;
        RECT 54.420 52.850 54.560 54.490 ;
        RECT 53.960 52.710 54.560 52.850 ;
        RECT 53.440 50.410 53.700 50.730 ;
        RECT 50.220 50.070 50.480 50.390 ;
        RECT 50.680 50.070 50.940 50.390 ;
        RECT 49.760 49.730 50.020 50.050 ;
        RECT 47.920 48.710 48.180 49.030 ;
        RECT 47.980 42.570 48.120 48.710 ;
        RECT 48.840 45.990 49.100 46.310 ;
        RECT 48.900 44.610 49.040 45.990 ;
        RECT 49.820 44.610 49.960 49.730 ;
        RECT 50.740 49.370 50.880 50.070 ;
        RECT 53.500 50.050 53.640 50.410 ;
        RECT 53.440 49.730 53.700 50.050 ;
        RECT 50.680 49.050 50.940 49.370 ;
        RECT 50.740 46.990 50.880 49.050 ;
        RECT 51.600 47.350 51.860 47.670 ;
        RECT 50.680 46.670 50.940 46.990 ;
        RECT 48.840 44.290 49.100 44.610 ;
        RECT 49.760 44.290 50.020 44.610 ;
        RECT 47.920 42.250 48.180 42.570 ;
        RECT 47.460 40.550 47.720 40.870 ;
        RECT 46.540 36.810 46.800 37.130 ;
        RECT 45.620 33.750 45.880 34.070 ;
        RECT 45.680 28.970 45.820 33.750 ;
        RECT 46.600 33.730 46.740 36.810 ;
        RECT 46.540 33.410 46.800 33.730 ;
        RECT 45.620 28.650 45.880 28.970 ;
        RECT 46.600 27.950 46.740 33.410 ;
        RECT 47.520 33.390 47.660 40.550 ;
        RECT 47.980 39.170 48.120 42.250 ;
        RECT 51.660 41.970 51.800 47.350 ;
        RECT 52.520 47.010 52.780 47.330 ;
        RECT 52.060 43.270 52.320 43.590 ;
        RECT 50.740 41.830 51.800 41.970 ;
        RECT 50.740 41.550 50.880 41.830 ;
        RECT 50.680 41.230 50.940 41.550 ;
        RECT 51.600 41.230 51.860 41.550 ;
        RECT 50.220 40.550 50.480 40.870 ;
        RECT 51.660 40.725 51.800 41.230 ;
        RECT 52.120 41.210 52.260 43.270 ;
        RECT 52.060 40.890 52.320 41.210 ;
        RECT 50.280 39.170 50.420 40.550 ;
        RECT 51.590 40.355 51.870 40.725 ;
        RECT 52.120 39.510 52.260 40.890 ;
        RECT 52.060 39.190 52.320 39.510 ;
        RECT 47.920 38.850 48.180 39.170 ;
        RECT 50.220 38.850 50.480 39.170 ;
        RECT 49.290 36.955 49.570 37.325 ;
        RECT 47.460 33.070 47.720 33.390 ;
        RECT 47.520 32.710 47.660 33.070 ;
        RECT 47.460 32.390 47.720 32.710 ;
        RECT 49.360 30.670 49.500 36.955 ;
        RECT 52.120 36.450 52.260 39.190 ;
        RECT 52.580 37.130 52.720 47.010 ;
        RECT 53.500 46.990 53.640 49.730 ;
        RECT 53.960 46.990 54.100 52.710 ;
        RECT 54.360 52.110 54.620 52.430 ;
        RECT 54.420 47.525 54.560 52.110 ;
        RECT 55.280 51.430 55.540 51.750 ;
        RECT 55.740 51.430 56.000 51.750 ;
        RECT 54.820 49.730 55.080 50.050 ;
        RECT 54.880 48.010 55.020 49.730 ;
        RECT 54.820 47.690 55.080 48.010 ;
        RECT 54.350 47.155 54.630 47.525 ;
        RECT 55.340 47.410 55.480 51.430 ;
        RECT 55.800 50.730 55.940 51.430 ;
        RECT 55.740 50.410 56.000 50.730 ;
        RECT 56.260 50.050 56.400 56.870 ;
        RECT 56.660 55.170 56.920 55.490 ;
        RECT 56.720 54.325 56.860 55.170 ;
        RECT 56.650 53.955 56.930 54.325 ;
        RECT 56.660 52.110 56.920 52.430 ;
        RECT 56.720 50.925 56.860 52.110 ;
        RECT 56.650 50.555 56.930 50.925 ;
        RECT 60.155 50.910 60.300 59.180 ;
        RECT 75.085 57.500 75.580 60.140 ;
        RECT 81.290 56.250 81.550 56.570 ;
        RECT 77.650 55.455 77.910 55.775 ;
        RECT 63.300 53.945 63.600 54.335 ;
        RECT 60.080 50.520 60.380 50.910 ;
        RECT 56.200 49.730 56.460 50.050 ;
        RECT 56.260 47.670 56.400 49.730 ;
        RECT 55.340 47.270 55.940 47.410 ;
        RECT 56.200 47.350 56.460 47.670 ;
        RECT 55.800 46.990 55.940 47.270 ;
        RECT 62.590 47.125 62.890 47.515 ;
        RECT 53.440 46.670 53.700 46.990 ;
        RECT 53.900 46.670 54.160 46.990 ;
        RECT 55.280 46.670 55.540 46.990 ;
        RECT 55.740 46.670 56.000 46.990 ;
        RECT 53.960 42.230 54.100 46.670 ;
        RECT 54.360 44.290 54.620 44.610 ;
        RECT 53.900 41.910 54.160 42.230 ;
        RECT 54.420 41.550 54.560 44.290 ;
        RECT 55.340 42.570 55.480 46.670 ;
        RECT 55.800 44.610 55.940 46.670 ;
        RECT 55.740 44.290 56.000 44.610 ;
        RECT 56.660 44.290 56.920 44.610 ;
        RECT 56.720 44.125 56.860 44.290 ;
        RECT 56.650 43.755 56.930 44.125 ;
        RECT 61.960 43.755 62.260 44.145 ;
        RECT 55.280 42.250 55.540 42.570 ;
        RECT 53.900 41.230 54.160 41.550 ;
        RECT 54.360 41.230 54.620 41.550 ;
        RECT 53.960 39.850 54.100 41.230 ;
        RECT 54.820 40.890 55.080 41.210 ;
        RECT 53.900 39.530 54.160 39.850 ;
        RECT 53.440 38.850 53.700 39.170 ;
        RECT 53.900 38.850 54.160 39.170 ;
        RECT 52.520 36.810 52.780 37.130 ;
        RECT 52.060 36.130 52.320 36.450 ;
        RECT 49.760 35.790 50.020 36.110 ;
        RECT 52.520 35.790 52.780 36.110 ;
        RECT 49.820 32.710 49.960 35.790 ;
        RECT 50.680 35.110 50.940 35.430 ;
        RECT 50.740 34.410 50.880 35.110 ;
        RECT 50.680 34.090 50.940 34.410 ;
        RECT 52.580 33.390 52.720 35.790 ;
        RECT 52.970 33.555 53.250 33.925 ;
        RECT 52.980 33.410 53.240 33.555 ;
        RECT 52.520 33.070 52.780 33.390 ;
        RECT 49.760 32.390 50.020 32.710 ;
        RECT 47.920 30.350 48.180 30.670 ;
        RECT 49.300 30.350 49.560 30.670 ;
        RECT 46.540 27.630 46.800 27.950 ;
        RECT 47.000 27.630 47.260 27.950 ;
        RECT 43.780 25.930 44.040 26.250 ;
        RECT 47.060 25.910 47.200 27.630 ;
        RECT 47.980 27.125 48.120 30.350 ;
        RECT 47.910 26.755 48.190 27.125 ;
        RECT 47.000 25.590 47.260 25.910 ;
        RECT 47.060 25.230 47.200 25.590 ;
        RECT 49.820 25.230 49.960 32.390 ;
        RECT 52.580 31.690 52.720 33.070 ;
        RECT 53.500 32.710 53.640 38.850 ;
        RECT 53.440 32.390 53.700 32.710 ;
        RECT 52.520 31.370 52.780 31.690 ;
        RECT 52.980 31.030 53.240 31.350 ;
        RECT 50.680 30.525 50.940 30.670 ;
        RECT 50.670 30.155 50.950 30.525 ;
        RECT 52.060 29.670 52.320 29.990 ;
        RECT 52.520 29.670 52.780 29.990 ;
        RECT 52.120 27.950 52.260 29.670 ;
        RECT 52.580 28.290 52.720 29.670 ;
        RECT 52.520 27.970 52.780 28.290 ;
        RECT 52.060 27.630 52.320 27.950 ;
        RECT 52.120 25.570 52.260 27.630 ;
        RECT 53.040 25.910 53.180 31.030 ;
        RECT 53.500 30.670 53.640 32.390 ;
        RECT 53.960 31.690 54.100 38.850 ;
        RECT 54.360 38.510 54.620 38.830 ;
        RECT 54.420 34.410 54.560 38.510 ;
        RECT 54.880 36.110 55.020 40.890 ;
        RECT 61.070 40.345 61.370 40.735 ;
        RECT 55.740 38.850 56.000 39.170 ;
        RECT 54.820 35.790 55.080 36.110 ;
        RECT 55.280 35.790 55.540 36.110 ;
        RECT 54.360 34.090 54.620 34.410 ;
        RECT 54.880 34.070 55.020 35.790 ;
        RECT 54.820 33.750 55.080 34.070 ;
        RECT 54.360 33.410 54.620 33.730 ;
        RECT 53.900 31.370 54.160 31.690 ;
        RECT 54.420 30.670 54.560 33.410 ;
        RECT 53.440 30.350 53.700 30.670 ;
        RECT 54.360 30.350 54.620 30.670 ;
        RECT 53.500 26.250 53.640 30.350 ;
        RECT 55.340 28.970 55.480 35.790 ;
        RECT 55.800 33.390 55.940 38.850 ;
        RECT 60.280 36.965 60.580 37.355 ;
        RECT 59.560 33.540 59.860 33.930 ;
        RECT 55.740 33.070 56.000 33.390 ;
        RECT 56.660 32.730 56.920 33.050 ;
        RECT 56.200 30.690 56.460 31.010 ;
        RECT 55.740 30.350 56.000 30.670 ;
        RECT 55.280 28.650 55.540 28.970 ;
        RECT 55.800 26.250 55.940 30.350 ;
        RECT 53.440 25.930 53.700 26.250 ;
        RECT 55.740 25.930 56.000 26.250 ;
        RECT 52.980 25.590 53.240 25.910 ;
        RECT 52.060 25.250 52.320 25.570 ;
        RECT 47.000 24.910 47.260 25.230 ;
        RECT 49.760 24.910 50.020 25.230 ;
        RECT 52.520 24.910 52.780 25.230 ;
        RECT 41.020 24.570 41.280 24.890 ;
        RECT 36.420 24.230 36.680 24.550 ;
        RECT 39.180 24.230 39.440 24.550 ;
        RECT 43.320 24.230 43.580 24.550 ;
        RECT 49.300 24.230 49.560 24.550 ;
        RECT 36.480 23.400 36.620 24.230 ;
        RECT 22.110 23.260 36.620 23.400 ;
        RECT 35.605 22.970 35.925 23.030 ;
        RECT 21.755 22.830 35.925 22.970 ;
        RECT 35.605 22.770 35.925 22.830 ;
        RECT 34.720 22.510 34.980 22.600 ;
        RECT 19.880 22.370 34.980 22.510 ;
        RECT 34.720 22.280 34.980 22.370 ;
        RECT 31.915 22.115 32.175 22.205 ;
        RECT 19.035 21.975 32.175 22.115 ;
        RECT 31.915 21.885 32.175 21.975 ;
        RECT 36.480 17.000 36.620 23.260 ;
        RECT 37.205 23.105 37.525 23.165 ;
        RECT 39.240 23.105 39.380 24.230 ;
        RECT 41.370 23.695 42.910 24.065 ;
        RECT 37.205 22.965 39.380 23.105 ;
        RECT 37.205 22.905 37.525 22.965 ;
        RECT 39.240 18.850 39.380 22.965 ;
        RECT 40.930 22.510 41.250 22.570 ;
        RECT 43.380 22.510 43.520 24.230 ;
        RECT 40.930 22.370 43.520 22.510 ;
        RECT 40.930 22.310 41.250 22.370 ;
        RECT 43.380 18.850 43.520 22.370 ;
        RECT 44.140 22.115 44.460 22.175 ;
        RECT 49.360 22.115 49.500 24.230 ;
        RECT 52.580 23.725 52.720 24.910 ;
        RECT 52.510 23.355 52.790 23.725 ;
        RECT 44.140 21.975 49.500 22.115 ;
        RECT 44.140 21.915 44.460 21.975 ;
        RECT 39.240 18.710 39.840 18.850 ;
        RECT 39.700 17.000 39.840 18.710 ;
        RECT 42.920 18.710 43.520 18.850 ;
        RECT 42.920 17.000 43.060 18.710 ;
        RECT 49.360 17.000 49.500 21.975 ;
        RECT 56.260 21.005 56.400 30.690 ;
        RECT 56.720 30.670 56.860 32.730 ;
        RECT 56.660 30.350 56.920 30.670 ;
        RECT 56.720 27.950 56.860 30.350 ;
        RECT 58.935 30.145 59.235 30.535 ;
        RECT 56.660 27.630 56.920 27.950 ;
        RECT 56.120 20.325 56.400 21.005 ;
        RECT 56.120 19.955 56.470 20.325 ;
        RECT 36.410 13.000 36.690 17.000 ;
        RECT 39.630 13.000 39.910 17.000 ;
        RECT 42.850 13.000 43.130 17.000 ;
        RECT 49.290 13.000 49.570 17.000 ;
        RECT 56.120 1.800 56.310 19.955 ;
        RECT 59.000 1.895 59.170 30.145 ;
        RECT 56.055 1.540 56.375 1.800 ;
        RECT 58.925 1.635 59.245 1.895 ;
        RECT 59.615 1.445 59.800 33.540 ;
        RECT 60.315 29.680 60.545 36.965 ;
        RECT 61.095 30.125 61.340 40.345 ;
        RECT 61.995 30.610 62.225 43.755 ;
        RECT 62.655 31.190 62.820 47.125 ;
        RECT 63.360 31.410 63.540 53.945 ;
        RECT 76.880 43.815 77.175 48.320 ;
        RECT 77.675 38.655 77.885 55.455 ;
        RECT 81.345 50.690 81.495 56.250 ;
        RECT 83.585 52.470 83.815 81.180 ;
        RECT 88.070 77.685 88.555 78.150 ;
        RECT 84.925 75.750 87.540 76.025 ;
        RECT 87.265 74.095 87.540 75.750 ;
        RECT 87.235 73.820 87.570 74.095 ;
        RECT 93.880 72.815 94.175 77.320 ;
        RECT 94.675 67.655 94.885 84.455 ;
        RECT 98.345 79.690 98.495 85.250 ;
        RECT 111.650 84.455 111.910 84.775 ;
        RECT 101.160 81.200 101.420 81.520 ;
        RECT 98.290 79.370 98.550 79.690 ;
        RECT 94.650 67.335 94.910 67.655 ;
        RECT 90.030 60.945 90.565 61.420 ;
        RECT 90.060 57.095 90.535 60.945 ;
        RECT 92.225 57.500 92.720 61.710 ;
        RECT 98.290 56.250 98.550 56.570 ;
        RECT 94.650 55.455 94.910 55.775 ;
        RECT 83.570 52.150 83.830 52.470 ;
        RECT 81.290 50.370 81.550 50.690 ;
        RECT 77.650 38.335 77.910 38.655 ;
        RECT 62.575 30.930 62.895 31.190 ;
        RECT 63.320 31.090 63.580 31.410 ;
        RECT 61.980 30.290 62.240 30.610 ;
        RECT 61.085 29.805 61.345 30.125 ;
        RECT 60.300 29.360 60.560 29.680 ;
        RECT 75.280 28.500 75.775 32.635 ;
        RECT 83.585 30.285 83.815 52.150 ;
        RECT 85.400 48.540 85.940 49.050 ;
        RECT 84.925 46.750 87.540 47.025 ;
        RECT 87.265 45.095 87.540 46.750 ;
        RECT 87.235 44.820 87.570 45.095 ;
        RECT 93.880 43.815 94.175 48.320 ;
        RECT 94.675 38.655 94.885 55.455 ;
        RECT 98.345 50.690 98.495 56.250 ;
        RECT 101.175 52.500 101.405 81.200 ;
        RECT 104.935 77.430 105.420 77.895 ;
        RECT 101.925 75.750 104.540 76.025 ;
        RECT 104.265 74.095 104.540 75.750 ;
        RECT 104.235 73.820 104.570 74.095 ;
        RECT 110.880 72.815 111.175 77.320 ;
        RECT 111.675 67.655 111.885 84.455 ;
        RECT 115.345 79.690 115.495 85.250 ;
        RECT 128.650 84.455 128.910 84.775 ;
        RECT 117.690 81.140 117.950 81.460 ;
        RECT 115.290 79.370 115.550 79.690 ;
        RECT 111.650 67.335 111.910 67.655 ;
        RECT 106.980 60.820 107.515 61.295 ;
        RECT 107.010 57.245 107.485 60.820 ;
        RECT 109.110 57.500 109.605 61.355 ;
        RECT 115.290 56.250 115.550 56.570 ;
        RECT 111.650 55.455 111.910 55.775 ;
        RECT 101.160 52.180 101.420 52.500 ;
        RECT 98.290 50.370 98.550 50.690 ;
        RECT 94.650 38.335 94.910 38.655 ;
        RECT 89.850 31.640 90.490 32.260 ;
        RECT 92.145 31.955 92.785 32.575 ;
        RECT 101.175 30.285 101.405 52.180 ;
        RECT 105.225 48.650 105.705 49.100 ;
        RECT 101.925 46.750 104.540 47.025 ;
        RECT 104.265 45.095 104.540 46.750 ;
        RECT 104.235 44.820 104.570 45.095 ;
        RECT 110.880 43.815 111.175 48.320 ;
        RECT 111.675 38.655 111.885 55.455 ;
        RECT 115.345 50.690 115.495 56.250 ;
        RECT 117.705 52.490 117.935 81.140 ;
        RECT 119.185 77.490 119.670 77.955 ;
        RECT 118.925 75.750 121.540 76.025 ;
        RECT 121.265 74.095 121.540 75.750 ;
        RECT 121.235 73.820 121.570 74.095 ;
        RECT 127.880 72.815 128.175 77.320 ;
        RECT 128.675 67.655 128.885 84.455 ;
        RECT 132.345 79.690 132.495 85.250 ;
        RECT 134.710 81.140 134.970 81.460 ;
        RECT 132.290 79.370 132.550 79.690 ;
        RECT 128.650 67.335 128.910 67.655 ;
        RECT 123.905 60.820 124.440 61.295 ;
        RECT 123.935 57.370 124.410 60.820 ;
        RECT 126.230 58.025 126.725 61.415 ;
        RECT 128.595 58.025 129.090 58.055 ;
        RECT 126.230 57.530 129.090 58.025 ;
        RECT 128.595 57.500 129.090 57.530 ;
        RECT 132.290 56.250 132.550 56.570 ;
        RECT 128.650 55.455 128.910 55.775 ;
        RECT 117.690 52.170 117.950 52.490 ;
        RECT 115.290 50.370 115.550 50.690 ;
        RECT 111.650 38.335 111.910 38.655 ;
        RECT 107.010 31.630 107.500 32.110 ;
        RECT 109.015 32.000 109.655 32.620 ;
        RECT 117.705 30.285 117.935 52.170 ;
        RECT 121.835 48.580 122.515 49.050 ;
        RECT 118.925 46.750 121.540 47.025 ;
        RECT 121.265 45.095 121.540 46.750 ;
        RECT 121.235 44.820 121.570 45.095 ;
        RECT 127.880 43.815 128.175 48.320 ;
        RECT 128.675 38.655 128.885 55.455 ;
        RECT 132.345 50.690 132.495 56.250 ;
        RECT 134.725 52.490 134.955 81.140 ;
        RECT 139.750 77.570 140.425 78.040 ;
        RECT 142.300 77.930 142.575 91.600 ;
        RECT 145.305 91.530 145.550 91.600 ;
        RECT 146.695 89.400 147.040 94.555 ;
        RECT 148.235 92.100 148.455 95.130 ;
        RECT 148.100 91.600 148.600 92.100 ;
        RECT 148.235 91.570 148.455 91.600 ;
        RECT 143.700 88.900 144.200 89.400 ;
        RECT 146.600 88.900 147.100 89.400 ;
        RECT 143.795 87.850 144.080 88.900 ;
        RECT 146.695 88.780 147.040 88.900 ;
        RECT 143.745 87.550 144.135 87.850 ;
        RECT 149.290 85.250 149.550 85.570 ;
        RECT 145.650 84.455 145.910 84.775 ;
        RECT 142.290 77.540 142.590 77.930 ;
        RECT 135.925 75.750 138.540 76.025 ;
        RECT 138.265 74.095 138.540 75.750 ;
        RECT 138.235 73.820 138.570 74.095 ;
        RECT 144.880 72.815 145.175 77.320 ;
        RECT 145.675 67.655 145.885 84.455 ;
        RECT 149.345 79.690 149.495 85.250 ;
        RECT 152.145 81.510 152.375 96.440 ;
        RECT 158.520 86.720 158.800 98.280 ;
        RECT 158.085 86.440 158.800 86.720 ;
        RECT 152.130 81.190 152.390 81.510 ;
        RECT 149.290 79.370 149.550 79.690 ;
        RECT 149.630 77.520 150.065 77.955 ;
        RECT 145.650 67.335 145.910 67.655 ;
        RECT 140.955 60.820 141.490 61.295 ;
        RECT 140.985 57.295 141.460 60.820 ;
        RECT 143.170 57.500 143.665 61.420 ;
        RECT 149.290 56.250 149.550 56.570 ;
        RECT 145.650 55.455 145.910 55.775 ;
        RECT 134.710 52.170 134.970 52.490 ;
        RECT 132.290 50.370 132.550 50.690 ;
        RECT 128.650 38.335 128.910 38.655 ;
        RECT 126.055 33.860 128.800 34.355 ;
        RECT 121.605 31.775 124.460 32.250 ;
        RECT 121.605 31.065 122.080 31.775 ;
        RECT 128.305 31.630 128.800 33.860 ;
        RECT 128.305 31.605 129.810 31.630 ;
        RECT 128.305 31.160 129.830 31.605 ;
        RECT 128.305 31.135 129.810 31.160 ;
        RECT 134.725 30.285 134.955 52.170 ;
        RECT 137.950 48.680 138.385 49.115 ;
        RECT 135.925 46.750 138.540 47.025 ;
        RECT 138.265 45.095 138.540 46.750 ;
        RECT 138.235 44.820 138.570 45.095 ;
        RECT 144.880 43.815 145.175 48.320 ;
        RECT 145.675 38.655 145.885 55.455 ;
        RECT 149.345 50.690 149.495 56.250 ;
        RECT 152.145 52.430 152.375 81.190 ;
        RECT 152.925 75.750 155.540 76.025 ;
        RECT 155.265 74.095 155.540 75.750 ;
        RECT 155.235 73.820 155.570 74.095 ;
        RECT 157.950 60.920 158.485 61.395 ;
        RECT 157.980 57.390 158.455 60.920 ;
        RECT 152.130 52.110 152.390 52.430 ;
        RECT 149.290 50.370 149.550 50.690 ;
        RECT 150.785 48.600 151.220 49.035 ;
        RECT 145.650 38.335 145.910 38.655 ;
        RECT 140.930 31.800 142.175 32.275 ;
        RECT 143.060 31.390 143.680 31.985 ;
        RECT 152.145 30.285 152.375 52.110 ;
        RECT 152.925 46.750 155.540 47.025 ;
        RECT 155.265 45.095 155.540 46.750 ;
        RECT 155.235 44.820 155.570 45.095 ;
        RECT 157.940 31.925 158.475 32.400 ;
        RECT 83.585 30.055 152.375 30.285 ;
        RECT 81.290 27.250 81.550 27.570 ;
        RECT 60.210 26.750 60.510 27.140 ;
        RECT 60.255 1.740 60.460 26.750 ;
        RECT 77.650 26.455 77.910 26.775 ;
        RECT 60.860 23.340 61.160 23.730 ;
        RECT 60.900 2.240 61.120 23.340 ;
        RECT 76.880 14.815 77.175 19.320 ;
        RECT 77.675 9.655 77.885 26.455 ;
        RECT 81.345 21.690 81.495 27.250 ;
        RECT 83.585 23.440 83.815 30.055 ;
        RECT 92.200 29.025 92.695 29.055 ;
        RECT 89.835 28.330 90.455 28.900 ;
        RECT 92.155 28.530 92.740 29.025 ;
        RECT 92.200 28.500 92.695 28.530 ;
        RECT 98.290 27.250 98.550 27.570 ;
        RECT 94.650 26.455 94.910 26.775 ;
        RECT 83.570 23.120 83.830 23.440 ;
        RECT 81.290 21.370 81.550 21.690 ;
        RECT 88.070 19.655 88.610 20.165 ;
        RECT 84.925 17.750 87.540 18.025 ;
        RECT 87.265 16.095 87.540 17.750 ;
        RECT 87.235 15.820 87.570 16.095 ;
        RECT 93.880 14.815 94.175 19.320 ;
        RECT 89.795 11.700 90.660 12.535 ;
        RECT 94.675 9.655 94.885 26.455 ;
        RECT 98.345 21.690 98.495 27.250 ;
        RECT 101.175 23.440 101.405 30.055 ;
        RECT 106.985 28.235 107.545 28.795 ;
        RECT 109.025 28.460 109.645 29.095 ;
        RECT 115.290 27.250 115.550 27.570 ;
        RECT 111.650 26.455 111.910 26.775 ;
        RECT 101.160 23.120 101.420 23.440 ;
        RECT 98.290 21.370 98.550 21.690 ;
        RECT 104.865 19.650 105.405 20.160 ;
        RECT 101.925 17.750 104.540 18.025 ;
        RECT 104.265 16.095 104.540 17.750 ;
        RECT 104.235 15.820 104.570 16.095 ;
        RECT 110.880 14.815 111.175 19.320 ;
        RECT 106.820 11.725 107.595 12.500 ;
        RECT 111.675 9.655 111.885 26.455 ;
        RECT 115.345 21.690 115.495 27.250 ;
        RECT 117.705 23.460 117.935 30.055 ;
        RECT 128.590 29.025 129.085 29.055 ;
        RECT 129.315 29.025 129.810 29.430 ;
        RECT 121.605 28.730 124.410 28.755 ;
        RECT 121.585 28.305 124.410 28.730 ;
        RECT 128.590 28.530 129.810 29.025 ;
        RECT 128.590 28.500 129.085 28.530 ;
        RECT 121.605 28.280 124.410 28.305 ;
        RECT 132.290 27.250 132.550 27.570 ;
        RECT 128.650 26.455 128.910 26.775 ;
        RECT 117.690 23.140 117.950 23.460 ;
        RECT 115.290 21.370 115.550 21.690 ;
        RECT 122.360 19.450 122.900 19.960 ;
        RECT 118.925 17.750 121.540 18.025 ;
        RECT 121.265 16.095 121.540 17.750 ;
        RECT 121.235 15.820 121.570 16.095 ;
        RECT 127.880 14.815 128.175 19.320 ;
        RECT 123.715 11.710 124.540 12.530 ;
        RECT 128.675 9.655 128.885 26.455 ;
        RECT 132.345 21.690 132.495 27.250 ;
        RECT 134.715 23.490 134.945 30.055 ;
        RECT 140.870 29.475 141.295 29.495 ;
        RECT 140.845 26.145 141.320 29.475 ;
        RECT 143.135 28.500 143.630 29.480 ;
        RECT 149.290 27.250 149.550 27.570 ;
        RECT 145.650 26.455 145.910 26.775 ;
        RECT 134.700 23.170 134.960 23.490 ;
        RECT 132.290 21.370 132.550 21.690 ;
        RECT 132.575 19.600 133.115 20.110 ;
        RECT 135.925 17.750 138.540 18.025 ;
        RECT 138.265 16.095 138.540 17.750 ;
        RECT 138.235 15.820 138.570 16.095 ;
        RECT 144.880 14.815 145.175 19.320 ;
        RECT 140.680 11.715 141.505 12.535 ;
        RECT 145.675 9.655 145.885 26.455 ;
        RECT 149.345 21.690 149.495 27.250 ;
        RECT 152.145 23.510 152.375 30.055 ;
        RECT 157.970 28.200 158.445 31.925 ;
        RECT 152.130 23.190 152.390 23.510 ;
        RECT 149.290 21.370 149.550 21.690 ;
        RECT 149.445 19.540 149.985 20.050 ;
        RECT 77.650 9.335 77.910 9.655 ;
        RECT 94.650 9.335 94.910 9.655 ;
        RECT 111.650 9.335 111.910 9.655 ;
        RECT 128.650 9.335 128.910 9.655 ;
        RECT 145.650 9.335 145.910 9.655 ;
        RECT 60.880 1.920 61.140 2.240 ;
        RECT 60.195 1.480 60.515 1.740 ;
        RECT 59.545 1.185 59.865 1.445 ;
        RECT 152.145 0.975 152.375 23.190 ;
        RECT 152.925 17.750 155.540 18.025 ;
        RECT 155.265 16.095 155.540 17.750 ;
        RECT 155.235 15.820 155.570 16.095 ;
        RECT 157.420 11.690 158.245 12.510 ;
        RECT 151.795 0.650 152.725 0.975 ;
      LAYER met3 ;
        RECT 63.800 224.860 64.120 225.240 ;
        RECT 66.535 224.915 66.855 225.295 ;
        RECT 69.285 224.920 69.605 225.300 ;
        RECT 72.065 224.925 72.385 225.305 ;
        RECT 21.585 223.985 21.915 224.315 ;
        RECT 20.740 221.645 21.070 221.975 ;
        RECT 19.980 220.890 20.310 221.220 ;
        RECT 19.210 219.710 19.540 220.040 ;
        RECT 18.555 219.090 18.885 219.420 ;
        RECT 17.775 218.605 18.105 218.935 ;
        RECT 17.090 217.005 17.420 217.335 ;
        RECT 16.410 216.410 16.740 216.740 ;
        RECT 16.425 55.490 16.725 216.410 ;
        RECT 17.105 56.235 17.405 217.005 ;
        RECT 17.785 58.380 18.095 218.605 ;
        RECT 17.790 57.785 18.090 58.380 ;
        RECT 17.765 57.435 18.115 57.785 ;
        RECT 18.570 57.275 18.870 219.090 ;
        RECT 19.210 58.245 19.535 219.710 ;
        RECT 19.995 58.350 20.295 220.890 ;
        RECT 20.755 59.005 21.055 221.645 ;
        RECT 20.730 58.655 21.080 59.005 ;
        RECT 19.220 57.485 19.520 58.245 ;
        RECT 19.970 58.000 20.320 58.350 ;
        RECT 18.405 56.975 18.870 57.275 ;
        RECT 19.195 57.135 19.545 57.485 ;
        RECT 18.405 56.490 18.705 56.975 ;
        RECT 17.080 55.885 17.430 56.235 ;
        RECT 18.405 56.165 19.040 56.490 ;
        RECT 18.690 56.140 19.040 56.165 ;
        RECT 16.400 55.140 16.750 55.490 ;
        RECT 17.000 54.290 21.000 54.440 ;
        RECT 21.600 54.290 21.900 223.985 ;
        RECT 22.240 223.115 22.570 223.445 ;
        RECT 22.255 60.335 22.555 223.115 ;
        RECT 23.110 222.320 23.440 222.650 ;
        RECT 23.125 61.355 23.425 222.320 ;
        RECT 23.980 220.335 24.310 220.665 ;
        RECT 23.100 61.005 23.450 61.355 ;
        RECT 23.995 61.070 24.295 220.335 ;
        RECT 24.715 218.020 25.045 218.350 ;
        RECT 24.730 61.810 25.030 218.020 ;
        RECT 25.370 217.420 25.700 217.750 ;
        RECT 25.385 62.470 25.685 217.420 ;
        RECT 63.810 216.750 64.110 224.860 ;
        RECT 66.545 216.975 66.845 224.915 ;
        RECT 69.295 217.760 69.595 224.920 ;
        RECT 72.075 218.365 72.375 224.925 ;
        RECT 74.800 224.855 75.120 225.235 ;
        RECT 77.530 224.930 77.850 225.310 ;
        RECT 74.810 218.950 75.110 224.855 ;
        RECT 77.540 219.430 77.840 224.930 ;
        RECT 80.270 224.895 80.590 225.275 ;
        RECT 80.280 220.050 80.580 224.895 ;
        RECT 83.045 224.880 83.365 225.260 ;
        RECT 83.055 220.675 83.355 224.880 ;
        RECT 85.800 224.855 86.120 225.235 ;
        RECT 88.590 224.985 88.910 225.365 ;
        RECT 85.810 221.230 86.110 224.855 ;
        RECT 88.600 221.985 88.900 224.985 ;
        RECT 91.340 224.855 91.660 225.235 ;
        RECT 94.070 224.955 94.390 225.335 ;
        RECT 91.350 222.660 91.650 224.855 ;
        RECT 94.080 223.455 94.380 224.955 ;
        RECT 94.055 223.105 94.405 223.455 ;
        RECT 91.325 222.310 91.675 222.660 ;
        RECT 88.575 221.635 88.925 221.985 ;
        RECT 85.785 220.880 86.135 221.230 ;
        RECT 83.030 220.325 83.380 220.675 ;
        RECT 80.255 219.700 80.605 220.050 ;
        RECT 77.515 219.080 77.865 219.430 ;
        RECT 102.410 219.330 102.710 223.730 ;
        RECT 105.140 219.790 105.440 223.730 ;
        RECT 119.005 220.345 119.305 223.730 ;
        RECT 121.720 220.820 122.020 223.730 ;
        RECT 124.530 221.255 124.830 223.730 ;
        RECT 127.280 221.715 127.580 223.730 ;
        RECT 129.960 222.220 130.260 223.730 ;
        RECT 132.775 222.670 133.075 223.730 ;
        RECT 135.545 223.120 135.845 223.730 ;
        RECT 135.520 222.770 135.870 223.120 ;
        RECT 132.750 222.320 133.100 222.670 ;
        RECT 129.935 221.870 130.285 222.220 ;
        RECT 127.255 221.365 127.605 221.715 ;
        RECT 124.505 220.905 124.855 221.255 ;
        RECT 121.695 220.470 122.045 220.820 ;
        RECT 118.980 219.995 119.330 220.345 ;
        RECT 105.115 219.440 105.465 219.790 ;
        RECT 102.385 218.980 102.735 219.330 ;
        RECT 74.785 218.600 75.135 218.950 ;
        RECT 72.050 218.015 72.400 218.365 ;
        RECT 69.270 217.410 69.620 217.760 ;
        RECT 63.785 216.400 64.135 216.750 ;
        RECT 66.520 216.625 66.870 216.975 ;
        RECT 117.345 95.065 117.695 95.415 ;
        RECT 56.625 64.490 56.955 64.505 ;
        RECT 60.045 64.490 64.045 64.640 ;
        RECT 56.625 64.190 64.045 64.490 ;
        RECT 56.625 64.175 56.955 64.190 ;
        RECT 60.045 64.040 64.045 64.190 ;
        RECT 35.675 62.470 36.025 62.495 ;
        RECT 25.385 62.170 36.025 62.470 ;
        RECT 35.675 62.145 36.025 62.170 ;
        RECT 42.010 61.810 42.360 61.835 ;
        RECT 24.730 61.510 42.360 61.810 ;
        RECT 42.010 61.485 42.360 61.510 ;
        RECT 53.865 61.090 54.195 61.105 ;
        RECT 60.045 61.090 64.045 61.240 ;
        RECT 23.995 60.875 41.405 61.070 ;
        RECT 23.995 60.770 41.430 60.875 ;
        RECT 53.865 60.790 64.045 61.090 ;
        RECT 53.865 60.775 54.195 60.790 ;
        RECT 41.080 60.525 41.430 60.770 ;
        RECT 60.045 60.640 64.045 60.790 ;
        RECT 39.595 60.335 39.945 60.360 ;
        RECT 22.255 60.035 39.945 60.335 ;
        RECT 39.595 60.010 39.945 60.035 ;
        RECT 38.050 59.075 39.630 59.405 ;
        RECT 55.245 57.690 55.575 57.705 ;
        RECT 59.315 57.690 59.665 57.695 ;
        RECT 60.045 57.690 64.045 57.840 ;
        RECT 55.245 57.390 64.045 57.690 ;
        RECT 55.245 57.375 55.575 57.390 ;
        RECT 59.315 57.345 59.665 57.390 ;
        RECT 60.045 57.240 64.045 57.390 ;
        RECT 41.350 56.355 42.930 56.685 ;
        RECT 33.165 55.650 33.495 55.665 ;
        RECT 37.305 55.650 37.635 55.665 ;
        RECT 50.645 55.650 50.975 55.665 ;
        RECT 33.165 55.350 50.975 55.650 ;
        RECT 33.165 55.335 33.495 55.350 ;
        RECT 37.305 55.335 37.635 55.350 ;
        RECT 50.645 55.335 50.975 55.350 ;
        RECT 34.545 54.290 34.875 54.305 ;
        RECT 17.000 53.990 34.875 54.290 ;
        RECT 17.000 53.840 21.000 53.990 ;
        RECT 34.545 53.975 34.875 53.990 ;
        RECT 56.625 54.290 56.955 54.305 ;
        RECT 60.045 54.290 64.045 54.440 ;
        RECT 56.625 53.990 64.045 54.290 ;
        RECT 56.625 53.975 56.955 53.990 ;
        RECT 38.050 53.635 39.630 53.965 ;
        RECT 60.045 53.840 64.045 53.990 ;
        RECT 17.000 50.890 21.000 51.040 ;
        RECT 41.350 50.915 42.930 51.245 ;
        RECT 23.505 50.890 23.835 50.905 ;
        RECT 17.000 50.590 23.835 50.890 ;
        RECT 17.000 50.440 21.000 50.590 ;
        RECT 23.505 50.575 23.835 50.590 ;
        RECT 56.625 50.890 56.955 50.905 ;
        RECT 60.045 50.890 64.045 51.040 ;
        RECT 56.625 50.590 64.045 50.890 ;
        RECT 56.625 50.575 56.955 50.590 ;
        RECT 60.045 50.440 64.045 50.590 ;
        RECT 38.050 48.195 39.630 48.525 ;
        RECT 54.325 47.490 54.655 47.505 ;
        RECT 60.045 47.490 64.045 47.640 ;
        RECT 54.325 47.190 64.045 47.490 ;
        RECT 54.325 47.175 54.655 47.190 ;
        RECT 60.045 47.040 64.045 47.190 ;
        RECT 41.350 45.475 42.930 45.805 ;
        RECT 17.000 44.090 21.000 44.240 ;
        RECT 21.730 44.090 22.060 44.105 ;
        RECT 23.505 44.090 23.835 44.105 ;
        RECT 17.000 43.790 23.835 44.090 ;
        RECT 17.000 43.640 21.000 43.790 ;
        RECT 21.730 43.775 22.060 43.790 ;
        RECT 23.505 43.775 23.835 43.790 ;
        RECT 56.625 44.090 56.955 44.105 ;
        RECT 60.045 44.090 64.045 44.240 ;
        RECT 56.625 43.790 64.045 44.090 ;
        RECT 56.625 43.775 56.955 43.790 ;
        RECT 60.045 43.640 64.045 43.790 ;
        RECT 38.050 42.755 39.630 43.085 ;
        RECT 51.565 40.690 51.895 40.705 ;
        RECT 60.045 40.690 64.045 40.840 ;
        RECT 51.565 40.390 64.045 40.690 ;
        RECT 51.565 40.375 51.895 40.390 ;
        RECT 41.350 40.035 42.930 40.365 ;
        RECT 60.045 40.240 64.045 40.390 ;
        RECT 17.000 37.305 21.000 37.440 ;
        RECT 38.050 37.315 39.630 37.645 ;
        RECT 17.000 37.290 21.130 37.305 ;
        RECT 23.505 37.290 23.835 37.305 ;
        RECT 17.000 36.990 23.835 37.290 ;
        RECT 17.000 36.975 21.130 36.990 ;
        RECT 23.505 36.975 23.835 36.990 ;
        RECT 49.265 37.290 49.595 37.305 ;
        RECT 60.045 37.290 64.045 37.440 ;
        RECT 49.265 36.990 64.045 37.290 ;
        RECT 49.265 36.975 49.595 36.990 ;
        RECT 17.000 36.840 21.000 36.975 ;
        RECT 60.045 36.840 64.045 36.990 ;
        RECT 41.350 34.595 42.930 34.925 ;
        RECT 59.395 34.040 60.270 34.055 ;
        RECT 52.945 33.890 53.275 33.905 ;
        RECT 59.395 33.890 64.045 34.040 ;
        RECT 52.945 33.590 64.045 33.890 ;
        RECT 52.945 33.575 53.275 33.590 ;
        RECT 59.395 33.440 64.045 33.590 ;
        RECT 59.395 33.415 60.195 33.440 ;
        RECT 38.050 31.875 39.630 32.205 ;
        RECT 50.645 30.490 50.975 30.505 ;
        RECT 58.910 30.490 59.260 30.515 ;
        RECT 60.045 30.490 64.045 30.640 ;
        RECT 50.645 30.190 64.045 30.490 ;
        RECT 50.645 30.175 50.975 30.190 ;
        RECT 58.910 30.165 59.260 30.190 ;
        RECT 60.045 30.040 64.045 30.190 ;
        RECT 41.350 29.155 42.930 29.485 ;
        RECT 21.205 27.770 21.535 27.785 ;
        RECT 20.990 27.455 21.535 27.770 ;
        RECT 20.990 27.240 21.290 27.455 ;
        RECT 17.000 26.790 21.290 27.240 ;
        RECT 47.885 27.090 48.215 27.105 ;
        RECT 60.045 27.090 64.045 27.240 ;
        RECT 47.885 26.790 64.045 27.090 ;
        RECT 17.000 26.640 21.000 26.790 ;
        RECT 47.885 26.775 48.215 26.790 ;
        RECT 38.050 26.435 39.630 26.765 ;
        RECT 60.045 26.640 64.045 26.790 ;
        RECT 41.350 23.715 42.930 24.045 ;
        RECT 52.485 23.690 52.815 23.705 ;
        RECT 60.045 23.690 64.045 23.840 ;
        RECT 52.485 23.390 64.045 23.690 ;
        RECT 52.485 23.375 52.815 23.390 ;
        RECT 60.045 23.240 64.045 23.390 ;
        RECT 69.185 21.700 70.380 90.285 ;
        RECT 117.370 78.855 117.670 95.065 ;
        RECT 118.320 94.530 118.715 94.925 ;
        RECT 88.180 78.555 117.670 78.855 ;
        RECT 88.180 78.150 88.480 78.555 ;
        RECT 88.070 77.685 88.555 78.150 ;
        RECT 104.935 77.835 105.420 77.895 ;
        RECT 118.345 77.835 118.690 94.530 ;
        RECT 119.245 93.920 119.595 94.270 ;
        RECT 119.270 77.955 119.570 93.920 ;
        RECT 120.350 93.485 120.700 93.835 ;
        RECT 104.935 77.490 118.690 77.835 ;
        RECT 119.185 77.490 119.670 77.955 ;
        RECT 104.935 77.430 105.420 77.490 ;
        RECT 74.115 59.995 75.425 61.225 ;
        RECT 120.375 51.540 120.675 93.485 ;
        RECT 121.255 92.970 121.605 93.320 ;
        RECT 85.460 51.240 120.675 51.540 ;
        RECT 85.460 48.920 85.760 51.240 ;
        RECT 121.280 50.110 121.580 92.970 ;
        RECT 123.120 92.885 133.705 93.185 ;
        RECT 122.095 92.505 122.445 92.855 ;
        RECT 105.300 49.810 121.580 50.110 ;
        RECT 105.300 49.030 105.600 49.810 ;
        RECT 85.445 48.590 85.775 48.920 ;
        RECT 105.285 48.700 105.615 49.030 ;
        RECT 122.120 48.995 122.420 92.505 ;
        RECT 122.105 48.665 122.435 48.995 ;
        RECT 89.895 31.680 90.420 32.205 ;
        RECT 89.920 28.380 90.395 31.680 ;
        RECT 92.200 29.050 92.695 32.495 ;
        RECT 107.000 31.605 107.525 32.130 ;
        RECT 92.175 28.505 92.720 29.050 ;
        RECT 107.025 28.280 107.500 31.605 ;
        RECT 109.085 29.050 109.580 32.570 ;
        RECT 121.580 31.085 122.105 31.610 ;
        RECT 109.060 28.505 109.605 29.050 ;
        RECT 121.605 28.280 122.080 31.085 ;
        RECT 123.120 22.985 123.420 92.885 ;
        RECT 127.175 91.705 127.525 92.055 ;
        RECT 133.405 92.015 133.705 92.885 ;
        RECT 125.140 89.920 125.515 90.295 ;
        RECT 124.045 88.190 124.395 88.540 ;
        RECT 88.155 22.685 123.420 22.985 ;
        RECT 1.005 21.600 2.995 21.625 ;
        RECT 37.735 21.600 39.735 21.630 ;
        RECT 1.000 19.600 39.735 21.600 ;
        RECT 56.165 20.290 56.495 20.305 ;
        RECT 60.045 20.290 64.045 20.440 ;
        RECT 69.120 20.430 70.420 21.700 ;
        RECT 56.165 19.990 64.045 20.290 ;
        RECT 88.155 20.045 88.455 22.685 ;
        RECT 124.070 21.240 124.370 88.190 ;
        RECT 104.960 20.940 124.370 21.240 ;
        RECT 104.960 20.045 105.260 20.940 ;
        RECT 56.165 19.975 56.495 19.990 ;
        RECT 60.045 19.840 64.045 19.990 ;
        RECT 88.140 19.715 88.470 20.045 ;
        RECT 104.945 19.715 105.275 20.045 ;
        RECT 122.430 19.850 122.760 19.855 ;
        RECT 125.165 19.850 125.490 89.920 ;
        RECT 126.235 89.045 126.585 89.395 ;
        RECT 1.005 19.575 2.995 19.600 ;
        RECT 122.430 19.525 125.490 19.850 ;
        RECT 126.260 20.005 126.560 89.045 ;
        RECT 127.200 28.305 127.500 91.705 ;
        RECT 133.380 91.665 133.730 92.015 ;
        RECT 134.850 88.070 135.200 88.095 ;
        RECT 134.850 87.770 139.270 88.070 ;
        RECT 143.765 87.850 144.115 87.875 ;
        RECT 134.850 87.745 135.200 87.770 ;
        RECT 133.965 87.255 134.315 87.280 ;
        RECT 133.965 86.955 138.300 87.255 ;
        RECT 133.965 86.930 134.315 86.955 ;
        RECT 138.000 49.115 138.300 86.955 ;
        RECT 137.950 48.680 138.385 49.115 ;
        RECT 138.970 48.970 139.270 87.770 ;
        RECT 140.310 87.550 144.115 87.850 ;
        RECT 140.310 78.040 140.610 87.550 ;
        RECT 143.765 87.525 144.115 87.550 ;
        RECT 139.750 77.640 140.610 78.040 ;
        RECT 142.265 77.885 142.615 77.910 ;
        RECT 149.630 77.885 150.065 77.955 ;
        RECT 139.750 77.570 140.425 77.640 ;
        RECT 142.265 77.585 150.065 77.885 ;
        RECT 142.265 77.560 142.615 77.585 ;
        RECT 149.630 77.520 150.065 77.585 ;
        RECT 150.785 48.970 151.220 49.035 ;
        RECT 138.970 48.670 151.220 48.970 ;
        RECT 150.785 48.600 151.220 48.670 ;
        RECT 141.630 31.775 142.155 32.300 ;
        RECT 129.315 29.410 129.810 31.630 ;
        RECT 141.655 29.475 142.130 31.775 ;
        RECT 143.060 31.390 143.680 31.985 ;
        RECT 129.290 28.865 129.835 29.410 ;
        RECT 140.845 29.000 142.130 29.475 ;
        RECT 143.135 29.460 143.630 31.390 ;
        RECT 143.110 28.915 143.655 29.460 ;
        RECT 127.200 28.005 149.925 28.305 ;
        RECT 132.630 20.005 132.960 20.020 ;
        RECT 126.260 19.705 132.960 20.005 ;
        RECT 149.625 19.930 149.925 28.005 ;
        RECT 132.630 19.690 132.960 19.705 ;
        RECT 149.610 19.600 149.940 19.930 ;
        RECT 89.795 12.460 90.660 12.535 ;
        RECT 106.820 12.460 107.595 12.500 ;
        RECT 89.795 12.455 158.190 12.460 ;
        RECT 89.785 11.780 158.190 12.455 ;
        RECT 89.795 11.775 158.190 11.780 ;
        RECT 89.795 11.700 90.660 11.775 ;
        RECT 106.820 11.725 107.595 11.775 ;
        RECT 151.815 0.995 152.705 1.000 ;
        RECT 151.785 0.630 152.735 0.995 ;
        RECT 151.815 0.625 152.705 0.630 ;
      LAYER met4 ;
        RECT 64.090 225.055 64.145 225.385 ;
        RECT 64.090 224.885 64.125 225.055 ;
        RECT 66.455 224.965 66.550 225.295 ;
        RECT 69.305 225.275 69.310 225.465 ;
        RECT 66.530 224.940 66.550 224.965 ;
        RECT 66.850 224.940 66.860 225.270 ;
        RECT 69.280 224.945 69.310 225.275 ;
        RECT 69.610 225.135 69.635 225.465 ;
        RECT 72.060 225.225 72.070 225.280 ;
        RECT 71.995 224.895 72.070 225.225 ;
        RECT 72.370 224.950 72.390 225.280 ;
        RECT 74.785 224.945 74.830 225.275 ;
        RECT 77.525 225.085 77.590 225.285 ;
        RECT 80.295 225.250 80.350 225.255 ;
        RECT 74.795 224.880 74.830 224.945 ;
        RECT 77.515 224.760 77.590 225.085 ;
        RECT 80.265 224.920 80.350 225.250 ;
        RECT 88.585 225.245 88.630 225.340 ;
        RECT 83.040 225.085 83.110 225.235 ;
        RECT 83.025 224.760 83.110 225.085 ;
        RECT 85.795 224.880 85.870 225.245 ;
        RECT 88.535 224.915 88.630 225.245 ;
        RECT 91.335 224.880 91.390 225.210 ;
        RECT 94.065 224.980 94.150 225.310 ;
        RECT 91.350 224.835 91.390 224.880 ;
        RECT 94.125 224.815 94.150 224.980 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 102.395 225.110 102.430 225.440 ;
        RECT 105.125 225.110 105.190 225.440 ;
        RECT 119.290 225.090 119.320 225.420 ;
        RECT 121.705 225.025 121.750 225.355 ;
        RECT 124.810 225.040 124.845 225.370 ;
        RECT 127.265 225.050 127.270 225.380 ;
        RECT 127.570 225.050 127.595 225.380 ;
        RECT 129.945 225.105 130.030 225.435 ;
        RECT 132.760 224.970 132.790 225.300 ;
        RECT 135.530 225.000 135.550 225.330 ;
        RECT 135.850 225.000 135.860 225.330 ;
        RECT 138.235 225.010 138.310 225.340 ;
        RECT 144.130 224.790 144.160 225.120 ;
        RECT 77.515 224.755 77.845 224.760 ;
        RECT 83.025 224.755 83.355 224.760 ;
        RECT 8.880 61.445 14.220 61.450 ;
        RECT 6.000 59.840 76.035 61.445 ;
        RECT 8.880 59.770 14.220 59.840 ;
        RECT 38.040 23.640 39.640 59.480 ;
        RECT 41.340 58.675 42.945 59.840 ;
        RECT 41.340 23.640 42.940 58.675 ;
        RECT 38.140 22.860 39.335 23.640 ;
        RECT 38.140 21.780 39.330 22.860 ;
        RECT 38.140 21.655 39.335 21.780 ;
        RECT 69.120 21.655 70.420 21.700 ;
        RECT 38.140 21.605 90.750 21.655 ;
        RECT 37.730 20.460 90.750 21.605 ;
        RECT 37.730 20.400 39.740 20.460 ;
        RECT 69.120 20.430 70.420 20.460 ;
        RECT 89.810 11.775 90.495 20.460 ;
        RECT 16.570 1.000 17.470 1.020 ;
        RECT 35.890 1.000 36.790 1.020 ;
        RECT 55.210 1.000 56.110 1.020 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

