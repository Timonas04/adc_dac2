magic
tech sky130A
magscale 1 2
timestamp 1730800671
<< metal1 >>
rect 29536 44108 29588 44114
rect 29536 44050 29588 44056
rect 29448 44000 29500 44006
rect 29448 43942 29500 43948
rect 29368 43850 29374 43902
rect 29426 43850 29432 43902
rect 29262 43804 29314 43810
rect 29262 43746 29314 43752
rect 21670 41226 21722 41232
rect 21670 41168 21722 41174
rect 21682 40352 21710 41168
rect 21762 41116 21814 41122
rect 21762 41058 21814 41064
rect 21774 40466 21802 41058
rect 21858 41018 21910 41024
rect 21858 40960 21910 40966
rect 21870 40634 21898 40960
rect 21858 40628 21910 40634
rect 21858 40570 21910 40576
rect 21774 40438 21984 40466
rect 21682 40324 21874 40352
rect 21563 39775 21762 39781
rect 21563 34934 21762 39576
rect 21846 39302 21874 40324
rect 21956 39442 21984 40438
rect 29274 39994 29302 43746
rect 29256 39988 29320 39994
rect 29256 39936 29262 39988
rect 29314 39936 29320 39988
rect 29256 39930 29320 39936
rect 29386 39528 29414 43850
rect 29368 39476 29374 39528
rect 29426 39476 29432 39528
rect 21938 39436 22004 39442
rect 21938 39384 21944 39436
rect 21996 39384 22004 39436
rect 29460 39384 29488 43942
rect 29548 40822 29576 44050
rect 29530 40816 29594 40822
rect 29530 40764 29536 40816
rect 29588 40764 29594 40816
rect 29530 40758 29594 40764
rect 21938 39378 22004 39384
rect 29366 39356 29488 39384
rect 21846 39274 21908 39302
rect 21880 38246 21908 39274
rect 21880 38240 21986 38246
rect 29366 38240 29394 39356
rect 21880 38200 21934 38240
rect 29348 38188 29354 38240
rect 29406 38188 29412 38240
rect 21934 38182 21986 38188
rect 20054 34735 27899 34934
rect 20072 34470 20234 34735
rect 23890 34464 24026 34735
rect 27678 34416 27816 34735
<< via1 >>
rect 29536 44056 29588 44108
rect 29448 43948 29500 44000
rect 29374 43850 29426 43902
rect 29262 43752 29314 43804
rect 21670 41174 21722 41226
rect 21762 41064 21814 41116
rect 21858 40966 21910 41018
rect 21858 40576 21910 40628
rect 21563 39576 21762 39775
rect 29262 39936 29314 39988
rect 29374 39476 29426 39528
rect 21944 39384 21996 39436
rect 29536 40764 29588 40816
rect 21934 38188 21986 38240
rect 29354 38188 29406 38240
rect 23638 34324 23722 34596
rect 27440 34280 27524 34552
rect 31246 34306 31340 34576
<< metal2 >>
rect 13855 44240 13864 44300
rect 13924 44284 13933 44300
rect 13924 44256 14640 44284
rect 13924 44240 13933 44256
rect 14612 44248 14640 44256
rect 14612 44220 25026 44248
rect 14393 44148 14402 44208
rect 14462 44192 14471 44208
rect 14462 44164 24898 44192
rect 14462 44148 14471 44164
rect 14951 44064 14960 44124
rect 15020 44112 15029 44124
rect 24711 44112 24720 44122
rect 15020 44076 24720 44112
rect 15020 44064 15029 44076
rect 24711 44066 24720 44076
rect 24776 44066 24785 44122
rect 24870 44074 24898 44164
rect 24998 44130 25026 44220
rect 24998 44102 27780 44130
rect 27752 44096 27780 44102
rect 29530 44096 29536 44108
rect 24870 44046 27660 44074
rect 27752 44068 29536 44096
rect 29530 44056 29536 44068
rect 29588 44056 29594 44108
rect 16053 43948 16062 44008
rect 16122 43997 16131 44008
rect 27431 43997 27440 44006
rect 16122 43966 27440 43997
rect 16122 43959 16571 43966
rect 16705 43959 27440 43966
rect 16122 43948 16131 43959
rect 27431 43950 27440 43959
rect 27496 43950 27505 44006
rect 27632 43988 27660 44046
rect 29442 43988 29448 44000
rect 27632 43960 29448 43988
rect 29442 43948 29448 43960
rect 29500 43948 29506 44000
rect 16599 43878 16608 43938
rect 16668 43922 16677 43938
rect 16668 43894 23036 43922
rect 16668 43878 16677 43894
rect 23008 43890 23036 43894
rect 29374 43902 29426 43908
rect 23008 43862 29374 43890
rect 17153 43791 17162 43851
rect 17222 43844 17231 43851
rect 29374 43844 29426 43850
rect 17222 43798 22828 43844
rect 17222 43791 17231 43798
rect 29256 43792 29262 43804
rect 23000 43764 29262 43792
rect 18273 43697 18333 43706
rect 18819 43704 18828 43764
rect 18888 43748 18897 43764
rect 23000 43748 23028 43764
rect 29256 43752 29262 43764
rect 29314 43752 29320 43804
rect 18888 43720 23028 43748
rect 26070 43724 26146 43734
rect 18888 43704 18897 43720
rect 26070 43713 26080 43724
rect 23136 43683 26080 43713
rect 18333 43672 18792 43683
rect 18924 43680 26080 43683
rect 18924 43672 23169 43680
rect 18333 43650 23169 43672
rect 26070 43668 26080 43680
rect 26136 43668 26146 43724
rect 26070 43658 26146 43668
rect 28108 43714 28188 43724
rect 28108 43658 28120 43714
rect 28176 43702 28188 43714
rect 28773 43702 28782 43717
rect 28176 43671 28782 43702
rect 28176 43658 28188 43671
rect 28108 43650 28188 43658
rect 28773 43657 28782 43671
rect 28842 43657 28851 43717
rect 18768 43644 18950 43650
rect 18273 43628 18333 43637
rect 17701 43558 17710 43618
rect 17770 43602 17779 43618
rect 17770 43598 18242 43602
rect 18364 43598 22002 43602
rect 17770 43574 22002 43598
rect 17770 43558 17779 43574
rect 18196 43566 18396 43574
rect 15506 43548 15566 43557
rect 15566 43530 17673 43532
rect 17807 43530 21926 43532
rect 15566 43504 21926 43530
rect 17656 43502 17824 43504
rect 15506 43479 15566 43488
rect 13285 43408 13294 43468
rect 13354 43452 13363 43468
rect 13354 43450 15474 43452
rect 15596 43450 21802 43452
rect 13354 43424 21802 43450
rect 13354 43408 13363 43424
rect 15450 43422 15628 43424
rect 12757 43336 12766 43396
rect 12826 43380 12835 43396
rect 12826 43352 21710 43380
rect 12826 43336 12835 43352
rect 21682 41226 21710 43352
rect 21664 41174 21670 41226
rect 21722 41174 21728 41226
rect 21774 41116 21802 43424
rect 21756 41064 21762 41116
rect 21814 41064 21820 41116
rect 21898 41018 21926 43504
rect 21852 40966 21858 41018
rect 21910 40972 21926 41018
rect 21910 40966 21916 40972
rect 21974 40776 22002 43574
rect 29530 40816 29594 40822
rect 29530 40764 29536 40816
rect 29588 40764 29594 40816
rect 29530 40758 29594 40764
rect 21852 40576 21858 40628
rect 21910 40616 21916 40628
rect 21910 40576 21934 40616
rect 21898 40550 21934 40576
rect 21898 40252 21926 40550
rect 21062 40224 21926 40252
rect 21062 40132 21090 40224
rect 29256 39988 29320 39994
rect 29256 39936 29262 39988
rect 29314 39936 29320 39988
rect 29256 39930 29320 39936
rect 21260 39576 21269 39775
rect 21468 39576 21563 39775
rect 21762 39576 21768 39775
rect 29374 39528 29426 39534
rect 29374 39470 29426 39476
rect 21938 39436 22004 39442
rect 21938 39384 21944 39436
rect 21996 39384 22004 39436
rect 21938 39378 22004 39384
rect 29354 38240 29406 38246
rect 21928 38188 21934 38240
rect 21986 38228 21992 38240
rect 21986 38200 22002 38228
rect 21986 38188 21992 38200
rect 29354 38182 29406 38188
rect 23618 34596 23736 34614
rect 23618 34324 23638 34596
rect 23722 34324 23736 34596
rect 23618 34302 23736 34324
rect 27422 34552 27552 34580
rect 27422 34280 27440 34552
rect 27524 34280 27552 34552
rect 31226 34576 31356 34604
rect 31226 34306 31246 34576
rect 31340 34306 31356 34576
rect 31226 34282 31356 34306
rect 27422 34258 27552 34280
rect 25416 22879 25425 22939
rect 25540 22879 25549 22939
<< via2 >>
rect 13864 44240 13924 44300
rect 14402 44148 14462 44208
rect 14960 44064 15020 44124
rect 24720 44066 24776 44122
rect 16062 43948 16122 44008
rect 27440 43950 27496 44006
rect 16608 43878 16668 43938
rect 17162 43791 17222 43851
rect 18828 43704 18888 43764
rect 18273 43637 18333 43697
rect 26080 43668 26136 43724
rect 28120 43658 28176 43714
rect 28782 43657 28842 43717
rect 17710 43558 17770 43618
rect 15506 43488 15566 43548
rect 13294 43408 13354 43468
rect 12766 43336 12826 43396
rect 21269 39576 21468 39775
rect 23638 34324 23722 34596
rect 27440 34280 27524 34552
rect 31246 34306 31340 34576
rect 25425 22879 25540 22939
<< metal3 >>
rect 13862 45092 13926 45098
rect 12764 45076 12828 45082
rect 12764 45006 12828 45012
rect 13292 45058 13356 45064
rect 12766 43401 12826 45006
rect 28780 45088 28844 45094
rect 14958 45054 15022 45060
rect 13862 45022 13926 45028
rect 14400 45044 14464 45050
rect 13292 44988 13356 44994
rect 13294 43473 13354 44988
rect 13864 44305 13924 45022
rect 16060 45050 16124 45056
rect 14958 44984 15022 44990
rect 15504 45016 15568 45022
rect 14400 44974 14464 44980
rect 13859 44300 13929 44305
rect 13859 44240 13864 44300
rect 13924 44240 13929 44300
rect 13859 44235 13929 44240
rect 14402 44213 14462 44974
rect 14397 44208 14467 44213
rect 14397 44148 14402 44208
rect 14462 44148 14467 44208
rect 14397 44143 14467 44148
rect 14960 44129 15020 44984
rect 17160 45048 17224 45054
rect 16060 44980 16124 44986
rect 16606 45016 16670 45022
rect 15504 44946 15568 44952
rect 14955 44124 15025 44129
rect 14955 44064 14960 44124
rect 15020 44064 15025 44124
rect 14955 44059 15025 44064
rect 15506 43553 15566 44946
rect 16062 44013 16122 44980
rect 17160 44978 17224 44984
rect 17708 45048 17772 45054
rect 17708 44978 17772 44984
rect 18271 45032 18335 45038
rect 16606 44946 16670 44952
rect 16057 44008 16127 44013
rect 16057 43948 16062 44008
rect 16122 43948 16127 44008
rect 16057 43943 16127 43948
rect 16608 43943 16668 44946
rect 16603 43938 16673 43943
rect 16603 43878 16608 43938
rect 16668 43878 16673 43938
rect 16603 43873 16673 43878
rect 17162 43856 17222 44978
rect 17157 43851 17227 43856
rect 17157 43791 17162 43851
rect 17222 43791 17227 43851
rect 17157 43786 17227 43791
rect 17710 43623 17770 44978
rect 18271 44962 18335 44968
rect 18826 45028 18890 45034
rect 28780 45018 28844 45024
rect 18273 43702 18333 44962
rect 18826 44958 18890 44964
rect 18828 43769 18888 44958
rect 24715 44122 24781 44127
rect 24715 44066 24720 44122
rect 24776 44066 24781 44122
rect 24715 44061 24781 44066
rect 18823 43764 18893 43769
rect 18823 43704 18828 43764
rect 18888 43704 18893 43764
rect 24718 43708 24778 44061
rect 27435 44006 27501 44011
rect 27435 43950 27440 44006
rect 27496 43950 27501 44006
rect 27435 43945 27501 43950
rect 26070 43724 26146 43734
rect 18268 43697 18338 43702
rect 18823 43699 18893 43704
rect 18268 43637 18273 43697
rect 18333 43637 18338 43697
rect 26070 43668 26080 43724
rect 26136 43668 26146 43724
rect 26070 43658 26146 43668
rect 27438 43656 27498 43945
rect 28782 43722 28842 45018
rect 28115 43714 28181 43719
rect 28115 43658 28120 43714
rect 28176 43658 28181 43714
rect 28115 43653 28181 43658
rect 28777 43717 28847 43722
rect 28777 43657 28782 43717
rect 28842 43657 28847 43717
rect 28777 43652 28847 43657
rect 18268 43632 18338 43637
rect 17705 43618 17775 43623
rect 17705 43558 17710 43618
rect 17770 43558 17775 43618
rect 17705 43553 17775 43558
rect 15501 43548 15571 43553
rect 15501 43488 15506 43548
rect 15566 43488 15571 43548
rect 15501 43483 15571 43488
rect 13289 43468 13359 43473
rect 13289 43408 13294 43468
rect 13354 43408 13359 43468
rect 13289 43403 13359 43408
rect 12761 43396 12831 43401
rect 12761 43336 12766 43396
rect 12826 43336 12831 43396
rect 12761 43331 12831 43336
rect 1713 40492 2031 40497
rect 214 40172 220 40492
rect 540 40491 2032 40492
rect 540 40173 1713 40491
rect 2031 40173 2032 40491
rect 21702 40433 21905 40434
rect 21697 40232 21703 40433
rect 21904 40232 21910 40433
rect 540 40172 2032 40173
rect 1713 40167 2031 40172
rect 21256 39780 21482 39786
rect 21256 39571 21264 39780
rect 21473 39571 21482 39780
rect 21256 39562 21482 39571
rect 21702 34602 21905 40232
rect 23618 34602 23736 34614
rect 31226 34602 31356 34604
rect 21688 34596 31359 34602
rect 21688 34371 23638 34596
rect 23618 34324 23638 34371
rect 23722 34576 31359 34596
rect 23722 34552 31246 34576
rect 23722 34371 27440 34552
rect 23722 34324 23736 34371
rect 23618 34302 23736 34324
rect 27422 34280 27440 34371
rect 27524 34371 31246 34552
rect 27524 34280 27552 34371
rect 31226 34306 31246 34371
rect 31340 34371 31359 34576
rect 31340 34306 31356 34371
rect 31226 34282 31356 34306
rect 27422 34258 27552 34280
rect 25420 22939 25545 22944
rect 25420 22879 25425 22939
rect 25540 22879 25545 22939
rect 25420 22875 25545 22879
rect 25420 22752 25421 22875
rect 25544 22752 25545 22875
rect 25420 22751 25545 22752
rect 25421 22746 25544 22751
<< via3 >>
rect 12764 45012 12828 45076
rect 13292 44994 13356 45058
rect 13862 45028 13926 45092
rect 14400 44980 14464 45044
rect 14958 44990 15022 45054
rect 15504 44952 15568 45016
rect 16060 44986 16124 45050
rect 16606 44952 16670 45016
rect 17160 44984 17224 45048
rect 17708 44984 17772 45048
rect 18271 44968 18335 45032
rect 18826 44964 18890 45028
rect 28780 45024 28844 45088
rect 220 40172 540 40492
rect 1713 40173 2031 40491
rect 21703 40232 21904 40433
rect 21264 39775 21473 39780
rect 21264 39576 21269 39775
rect 21269 39576 21468 39775
rect 21468 39576 21473 39775
rect 21264 39571 21473 39576
rect 25421 22752 25544 22875
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 45077 12818 45152
rect 12758 45076 12829 45077
rect 12758 45012 12764 45076
rect 12828 45012 12829 45076
rect 13310 45059 13370 45152
rect 13862 45093 13922 45152
rect 12758 45011 12829 45012
rect 13291 45058 13370 45059
rect 12758 44952 12818 45011
rect 13291 44994 13292 45058
rect 13356 44994 13370 45058
rect 13861 45092 13927 45093
rect 13861 45028 13862 45092
rect 13926 45028 13927 45092
rect 14414 45045 14474 45152
rect 14966 45055 15026 45152
rect 13861 45027 13927 45028
rect 14399 45044 14474 45045
rect 13291 44993 13370 44994
rect 13310 44952 13370 44993
rect 13862 44952 13922 45027
rect 14399 44980 14400 45044
rect 14464 44980 14474 45044
rect 14957 45054 15026 45055
rect 14957 44990 14958 45054
rect 15022 44990 15026 45054
rect 15518 45017 15578 45152
rect 16070 45051 16130 45152
rect 14957 44989 15026 44990
rect 14399 44979 14474 44980
rect 14414 44952 14474 44979
rect 14966 44952 15026 44989
rect 15503 45016 15578 45017
rect 15503 44952 15504 45016
rect 15568 44952 15578 45016
rect 16059 45050 16130 45051
rect 16059 44986 16060 45050
rect 16124 44986 16130 45050
rect 16622 45017 16682 45152
rect 17174 45049 17234 45152
rect 17726 45049 17786 45152
rect 16059 44985 16130 44986
rect 16070 44952 16130 44985
rect 16605 45016 16682 45017
rect 16605 44952 16606 45016
rect 16670 44952 16682 45016
rect 17159 45048 17234 45049
rect 17159 44984 17160 45048
rect 17224 44984 17234 45048
rect 17159 44983 17234 44984
rect 17707 45048 17786 45049
rect 17707 44984 17708 45048
rect 17772 44984 17786 45048
rect 18278 45033 18338 45152
rect 17707 44983 17786 44984
rect 17174 44952 17234 44983
rect 17726 44952 17786 44983
rect 18270 45032 18338 45033
rect 18270 44968 18271 45032
rect 18335 44968 18338 45032
rect 18830 45029 18890 45152
rect 18270 44967 18338 44968
rect 18278 44952 18338 44967
rect 18825 45028 18891 45029
rect 18825 44964 18826 45028
rect 18890 44964 18891 45028
rect 18825 44963 18891 44964
rect 18830 44952 18890 44963
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 45089 28826 45152
rect 28766 45088 28845 45089
rect 28766 45024 28780 45088
rect 28844 45024 28845 45088
rect 28766 45023 28845 45024
rect 28766 44952 28826 45023
rect 29318 44952 29378 45152
rect 15503 44951 15569 44952
rect 16605 44951 16671 44952
rect 200 40492 600 44152
rect 200 40172 220 40492
rect 540 40172 600 40492
rect 200 1000 600 40172
rect 800 39832 1200 44152
rect 1712 40491 22656 40492
rect 1712 40173 1713 40491
rect 2031 40433 22656 40491
rect 2031 40232 21703 40433
rect 21904 40232 22656 40433
rect 2031 40173 22656 40232
rect 1712 40172 22656 40173
rect 800 39780 22606 39832
rect 800 39571 21264 39780
rect 21473 39571 22606 39780
rect 800 39512 22606 39571
rect 800 1000 1200 39512
rect 23618 34302 23736 34614
rect 25420 22875 30515 22876
rect 25420 22752 25421 22875
rect 25544 22752 30515 22875
rect 25420 22751 30515 22752
rect 30390 200 30515 22751
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use flash_adc  flash_adc_0
timestamp 1730795883
transform 0 1 18078 -1 0 22692
box -22008 1842 3604 13395
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
