VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  OBS
      LAYER nwell ;
        RECT 17.130 211.005 147.230 212.610 ;
      LAYER pwell ;
        RECT 17.325 209.805 18.695 210.615 ;
        RECT 18.705 209.805 24.215 210.615 ;
        RECT 24.225 209.805 29.735 210.615 ;
        RECT 30.215 209.890 30.645 210.675 ;
        RECT 30.665 209.805 36.175 210.615 ;
        RECT 36.185 209.805 41.695 210.615 ;
        RECT 41.705 209.805 43.075 210.615 ;
        RECT 43.095 209.890 43.525 210.675 ;
        RECT 43.545 209.805 49.055 210.615 ;
        RECT 49.065 209.805 54.575 210.615 ;
        RECT 54.585 209.805 55.955 210.615 ;
        RECT 55.975 209.890 56.405 210.675 ;
        RECT 56.425 209.805 60.095 210.615 ;
        RECT 60.565 209.805 63.175 210.715 ;
        RECT 63.325 209.805 68.835 210.615 ;
        RECT 68.855 209.890 69.285 210.675 ;
        RECT 69.305 209.805 74.815 210.615 ;
        RECT 74.825 209.805 78.495 210.615 ;
        RECT 78.505 209.805 79.875 210.615 ;
        RECT 79.885 210.485 81.230 210.715 ;
        RECT 79.885 209.805 81.715 210.485 ;
        RECT 81.735 209.890 82.165 210.675 ;
        RECT 85.605 210.625 86.555 210.715 ;
        RECT 83.105 209.805 84.475 210.585 ;
        RECT 85.605 209.805 87.535 210.625 ;
        RECT 87.705 209.805 89.075 210.585 ;
        RECT 89.085 209.805 90.455 210.615 ;
        RECT 90.475 209.805 91.825 210.715 ;
        RECT 91.845 209.805 94.595 210.615 ;
        RECT 94.615 209.890 95.045 210.675 ;
        RECT 95.985 210.485 97.330 210.715 ;
        RECT 95.985 209.805 97.815 210.485 ;
        RECT 97.825 209.805 103.335 210.615 ;
        RECT 103.345 209.805 107.015 210.615 ;
        RECT 107.495 209.890 107.925 210.675 ;
        RECT 107.945 209.805 113.455 210.615 ;
        RECT 113.465 209.805 118.975 210.615 ;
        RECT 118.985 209.805 120.355 210.615 ;
        RECT 120.375 209.890 120.805 210.675 ;
        RECT 120.825 209.805 126.335 210.615 ;
        RECT 126.345 209.805 131.855 210.615 ;
        RECT 131.865 209.805 133.235 210.615 ;
        RECT 133.255 209.890 133.685 210.675 ;
        RECT 133.705 209.805 139.215 210.615 ;
        RECT 139.225 209.805 144.735 210.615 ;
        RECT 145.665 209.805 147.035 210.615 ;
        RECT 17.465 209.595 17.635 209.805 ;
        RECT 18.845 209.595 19.015 209.805 ;
        RECT 24.365 209.595 24.535 209.805 ;
        RECT 29.885 209.755 30.055 209.785 ;
        RECT 29.880 209.645 30.055 209.755 ;
        RECT 29.885 209.595 30.055 209.645 ;
        RECT 30.805 209.615 30.975 209.805 ;
        RECT 35.405 209.595 35.575 209.785 ;
        RECT 36.325 209.615 36.495 209.805 ;
        RECT 40.925 209.595 41.095 209.785 ;
        RECT 41.845 209.615 42.015 209.805 ;
        RECT 42.760 209.645 42.880 209.755 ;
        RECT 43.685 209.595 43.855 209.805 ;
        RECT 49.205 209.595 49.375 209.805 ;
        RECT 51.960 209.645 52.080 209.755 ;
        RECT 53.800 209.595 53.970 209.785 ;
        RECT 54.725 209.615 54.895 209.805 ;
        RECT 55.640 209.595 55.810 209.785 ;
        RECT 56.115 209.640 56.275 209.750 ;
        RECT 56.565 209.615 56.735 209.805 ;
        RECT 57.025 209.595 57.195 209.785 ;
        RECT 60.240 209.645 60.360 209.755 ;
        RECT 60.710 209.595 60.880 209.805 ;
        RECT 62.085 209.595 62.255 209.785 ;
        RECT 63.465 209.615 63.635 209.805 ;
        RECT 69.445 209.785 69.615 209.805 ;
        RECT 65.765 209.595 65.935 209.785 ;
        RECT 68.525 209.595 68.695 209.785 ;
        RECT 69.445 209.615 69.620 209.785 ;
        RECT 69.450 209.595 69.620 209.615 ;
        RECT 70.825 209.595 70.995 209.785 ;
        RECT 74.965 209.615 75.135 209.805 ;
        RECT 76.345 209.595 76.515 209.785 ;
        RECT 78.645 209.615 78.815 209.805 ;
        RECT 80.035 209.640 80.195 209.750 ;
        RECT 80.945 209.595 81.115 209.785 ;
        RECT 81.405 209.615 81.575 209.805 ;
        RECT 82.335 209.650 82.495 209.760 ;
        RECT 83.255 209.615 83.425 209.805 ;
        RECT 87.385 209.785 87.535 209.805 ;
        RECT 84.625 209.595 84.795 209.785 ;
        RECT 86.005 209.595 86.175 209.785 ;
        RECT 87.385 209.615 87.555 209.785 ;
        RECT 87.855 209.615 88.025 209.805 ;
        RECT 89.225 209.615 89.395 209.805 ;
        RECT 89.690 209.595 89.860 209.785 ;
        RECT 90.605 209.615 90.775 209.805 ;
        RECT 91.985 209.615 92.155 209.805 ;
        RECT 92.900 209.645 93.020 209.755 ;
        RECT 93.360 209.595 93.530 209.785 ;
        RECT 17.325 208.785 18.695 209.595 ;
        RECT 18.705 208.785 24.215 209.595 ;
        RECT 24.225 208.785 29.735 209.595 ;
        RECT 29.745 208.785 35.255 209.595 ;
        RECT 35.265 208.785 40.775 209.595 ;
        RECT 40.785 208.785 42.615 209.595 ;
        RECT 43.095 208.725 43.525 209.510 ;
        RECT 43.545 208.785 49.055 209.595 ;
        RECT 49.065 208.785 51.815 209.595 ;
        RECT 52.345 208.685 54.115 209.595 ;
        RECT 54.185 208.685 55.955 209.595 ;
        RECT 56.995 208.915 60.460 209.595 ;
        RECT 59.540 208.685 60.460 208.915 ;
        RECT 60.565 208.685 61.915 209.595 ;
        RECT 61.945 208.785 65.615 209.595 ;
        RECT 65.625 208.785 66.995 209.595 ;
        RECT 67.005 208.685 68.820 209.595 ;
        RECT 68.855 208.725 69.285 209.510 ;
        RECT 69.305 208.685 70.655 209.595 ;
        RECT 70.685 208.785 76.195 209.595 ;
        RECT 76.205 208.785 79.875 209.595 ;
        RECT 80.915 208.915 84.380 209.595 ;
        RECT 83.460 208.685 84.380 208.915 ;
        RECT 84.485 208.785 85.855 209.595 ;
        RECT 85.975 208.915 89.440 209.595 ;
        RECT 88.520 208.685 89.440 208.915 ;
        RECT 89.545 208.685 92.465 209.595 ;
        RECT 93.245 208.685 94.595 209.595 ;
        RECT 95.210 209.565 95.380 209.785 ;
        RECT 97.505 209.615 97.675 209.805 ;
        RECT 97.965 209.615 98.135 209.805 ;
        RECT 98.435 209.640 98.595 209.750 ;
        RECT 99.345 209.595 99.515 209.785 ;
        RECT 102.565 209.615 102.735 209.785 ;
        RECT 103.485 209.615 103.655 209.805 ;
        RECT 102.570 209.595 102.735 209.615 ;
        RECT 104.865 209.595 105.035 209.785 ;
        RECT 107.160 209.645 107.280 209.755 ;
        RECT 108.085 209.615 108.255 209.805 ;
        RECT 110.385 209.595 110.555 209.785 ;
        RECT 113.605 209.615 113.775 209.805 ;
        RECT 115.905 209.595 116.075 209.785 ;
        RECT 119.125 209.615 119.295 209.805 ;
        RECT 119.595 209.640 119.755 209.750 ;
        RECT 120.965 209.595 121.135 209.805 ;
        RECT 126.485 209.595 126.655 209.805 ;
        RECT 132.005 209.595 132.175 209.805 ;
        RECT 133.845 209.615 134.015 209.805 ;
        RECT 137.525 209.595 137.695 209.785 ;
        RECT 139.365 209.615 139.535 209.805 ;
        RECT 143.045 209.595 143.215 209.785 ;
        RECT 144.895 209.650 145.055 209.760 ;
        RECT 146.725 209.595 146.895 209.805 ;
        RECT 97.340 209.565 98.275 209.595 ;
        RECT 94.615 208.725 95.045 209.510 ;
        RECT 95.210 209.365 98.275 209.565 ;
        RECT 95.065 208.885 98.275 209.365 ;
        RECT 95.065 208.685 95.995 208.885 ;
        RECT 97.325 208.685 98.275 208.885 ;
        RECT 99.305 208.685 102.415 209.595 ;
        RECT 102.570 208.915 104.405 209.595 ;
        RECT 103.475 208.685 104.405 208.915 ;
        RECT 104.725 208.785 110.235 209.595 ;
        RECT 110.245 208.785 115.755 209.595 ;
        RECT 115.765 208.785 119.435 209.595 ;
        RECT 120.375 208.725 120.805 209.510 ;
        RECT 120.825 208.785 126.335 209.595 ;
        RECT 126.345 208.785 131.855 209.595 ;
        RECT 131.865 208.785 137.375 209.595 ;
        RECT 137.385 208.785 142.895 209.595 ;
        RECT 142.905 208.785 145.655 209.595 ;
        RECT 145.665 208.785 147.035 209.595 ;
      LAYER nwell ;
        RECT 17.130 205.565 147.230 208.395 ;
      LAYER pwell ;
        RECT 17.325 204.365 18.695 205.175 ;
        RECT 18.705 204.365 24.215 205.175 ;
        RECT 24.225 204.365 29.735 205.175 ;
        RECT 30.215 204.450 30.645 205.235 ;
        RECT 30.665 204.365 36.175 205.175 ;
        RECT 36.185 204.365 41.695 205.175 ;
        RECT 41.705 204.365 47.215 205.175 ;
        RECT 47.225 204.365 49.055 205.175 ;
        RECT 49.160 205.045 50.080 205.275 ;
        RECT 49.160 204.365 52.625 205.045 ;
        RECT 52.745 204.365 55.855 205.275 ;
        RECT 55.975 204.450 56.405 205.235 ;
        RECT 56.465 205.045 57.815 205.275 ;
        RECT 59.350 205.045 60.260 205.265 ;
        RECT 64.285 205.045 65.635 205.275 ;
        RECT 67.170 205.045 68.080 205.265 ;
        RECT 56.465 204.365 63.775 205.045 ;
        RECT 64.285 204.365 71.595 205.045 ;
        RECT 71.605 204.365 77.115 205.175 ;
        RECT 77.125 204.365 80.795 205.175 ;
        RECT 81.735 204.450 82.165 205.235 ;
        RECT 82.685 205.045 84.035 205.275 ;
        RECT 85.570 205.045 86.480 205.265 ;
        RECT 93.520 205.045 94.430 205.265 ;
        RECT 95.965 205.045 97.315 205.275 ;
        RECT 100.880 205.045 101.790 205.265 ;
        RECT 103.325 205.045 104.675 205.275 ;
        RECT 82.685 204.365 89.995 205.045 ;
        RECT 90.005 204.365 97.315 205.045 ;
        RECT 97.365 204.365 104.675 205.045 ;
        RECT 104.735 204.365 107.475 205.045 ;
        RECT 107.495 204.450 107.925 205.235 ;
        RECT 107.945 204.365 113.455 205.175 ;
        RECT 113.465 204.365 118.975 205.175 ;
        RECT 118.985 204.365 124.495 205.175 ;
        RECT 124.505 204.365 130.015 205.175 ;
        RECT 130.025 204.365 132.775 205.175 ;
        RECT 133.255 204.450 133.685 205.235 ;
        RECT 133.705 204.365 139.215 205.175 ;
        RECT 139.225 204.365 144.735 205.175 ;
        RECT 145.665 204.365 147.035 205.175 ;
        RECT 17.465 204.155 17.635 204.365 ;
        RECT 18.845 204.155 19.015 204.365 ;
        RECT 24.365 204.155 24.535 204.365 ;
        RECT 29.885 204.315 30.055 204.345 ;
        RECT 29.880 204.205 30.055 204.315 ;
        RECT 29.885 204.155 30.055 204.205 ;
        RECT 30.805 204.175 30.975 204.365 ;
        RECT 35.405 204.155 35.575 204.345 ;
        RECT 36.325 204.175 36.495 204.365 ;
        RECT 40.925 204.155 41.095 204.345 ;
        RECT 41.845 204.175 42.015 204.365 ;
        RECT 42.760 204.205 42.880 204.315 ;
        RECT 43.685 204.155 43.855 204.345 ;
        RECT 45.980 204.155 46.150 204.345 ;
        RECT 46.445 204.155 46.615 204.345 ;
        RECT 47.365 204.175 47.535 204.365 ;
        RECT 52.425 204.175 52.595 204.365 ;
        RECT 53.805 204.155 53.975 204.345 ;
        RECT 55.645 204.175 55.815 204.365 ;
        RECT 63.465 204.175 63.635 204.365 ;
        RECT 63.920 204.205 64.040 204.315 ;
        RECT 64.385 204.155 64.555 204.345 ;
        RECT 64.840 204.205 64.960 204.315 ;
        RECT 65.305 204.155 65.475 204.345 ;
        RECT 71.285 204.175 71.455 204.365 ;
        RECT 71.745 204.175 71.915 204.365 ;
        RECT 72.665 204.155 72.835 204.345 ;
        RECT 73.125 204.155 73.295 204.345 ;
        RECT 77.265 204.175 77.435 204.365 ;
        RECT 80.485 204.155 80.655 204.345 ;
        RECT 80.955 204.210 81.115 204.320 ;
        RECT 82.320 204.205 82.440 204.315 ;
        RECT 87.855 204.200 88.015 204.310 ;
        RECT 88.770 204.155 88.940 204.345 ;
        RECT 89.685 204.175 89.855 204.365 ;
        RECT 90.145 204.175 90.315 204.365 ;
        RECT 97.505 204.345 97.675 204.365 ;
        RECT 93.365 204.155 93.535 204.345 ;
        RECT 93.835 204.200 93.995 204.310 ;
        RECT 17.325 203.345 18.695 204.155 ;
        RECT 18.705 203.345 24.215 204.155 ;
        RECT 24.225 203.345 29.735 204.155 ;
        RECT 29.745 203.345 35.255 204.155 ;
        RECT 35.265 203.345 40.775 204.155 ;
        RECT 40.785 203.345 42.615 204.155 ;
        RECT 43.095 203.285 43.525 204.070 ;
        RECT 43.545 203.345 44.915 204.155 ;
        RECT 44.945 203.245 46.295 204.155 ;
        RECT 46.305 203.475 53.615 204.155 ;
        RECT 53.665 203.475 60.975 204.155 ;
        RECT 49.820 203.255 50.730 203.475 ;
        RECT 52.265 203.245 53.615 203.475 ;
        RECT 57.180 203.255 58.090 203.475 ;
        RECT 59.625 203.245 60.975 203.475 ;
        RECT 61.120 203.475 64.585 204.155 ;
        RECT 65.275 203.475 68.740 204.155 ;
        RECT 61.120 203.245 62.040 203.475 ;
        RECT 67.820 203.245 68.740 203.475 ;
        RECT 68.855 203.285 69.285 204.070 ;
        RECT 69.445 203.245 72.895 204.155 ;
        RECT 72.985 203.475 80.295 204.155 ;
        RECT 80.345 203.475 87.655 204.155 ;
        RECT 76.500 203.255 77.410 203.475 ;
        RECT 78.945 203.245 80.295 203.475 ;
        RECT 83.860 203.255 84.770 203.475 ;
        RECT 86.305 203.245 87.655 203.475 ;
        RECT 88.625 203.245 92.280 204.155 ;
        RECT 92.315 203.245 93.665 204.155 ;
        RECT 95.200 204.125 95.370 204.345 ;
        RECT 97.505 204.175 97.680 204.345 ;
        RECT 107.165 204.175 107.335 204.365 ;
        RECT 97.510 204.155 97.680 204.175 ;
        RECT 108.085 204.155 108.255 204.365 ;
        RECT 108.545 204.155 108.715 204.345 ;
        RECT 113.605 204.175 113.775 204.365 ;
        RECT 114.065 204.155 114.235 204.345 ;
        RECT 119.125 204.175 119.295 204.365 ;
        RECT 119.595 204.200 119.755 204.310 ;
        RECT 120.965 204.155 121.135 204.345 ;
        RECT 124.645 204.175 124.815 204.365 ;
        RECT 126.485 204.155 126.655 204.345 ;
        RECT 130.165 204.175 130.335 204.365 ;
        RECT 132.005 204.155 132.175 204.345 ;
        RECT 132.920 204.205 133.040 204.315 ;
        RECT 133.845 204.175 134.015 204.365 ;
        RECT 137.525 204.155 137.695 204.345 ;
        RECT 139.365 204.175 139.535 204.365 ;
        RECT 143.045 204.155 143.215 204.345 ;
        RECT 144.895 204.210 145.055 204.320 ;
        RECT 146.725 204.155 146.895 204.365 ;
        RECT 96.400 204.125 97.355 204.155 ;
        RECT 94.615 203.285 95.045 204.070 ;
        RECT 95.075 203.445 97.355 204.125 ;
        RECT 96.400 203.245 97.355 203.445 ;
        RECT 97.365 203.475 100.950 204.155 ;
        RECT 101.085 203.475 108.395 204.155 ;
        RECT 97.365 203.245 98.285 203.475 ;
        RECT 101.085 203.245 102.435 203.475 ;
        RECT 103.970 203.255 104.880 203.475 ;
        RECT 108.405 203.345 113.915 204.155 ;
        RECT 113.925 203.345 119.435 204.155 ;
        RECT 120.375 203.285 120.805 204.070 ;
        RECT 120.825 203.345 126.335 204.155 ;
        RECT 126.345 203.345 131.855 204.155 ;
        RECT 131.865 203.345 137.375 204.155 ;
        RECT 137.385 203.345 142.895 204.155 ;
        RECT 142.905 203.345 145.655 204.155 ;
        RECT 145.665 203.345 147.035 204.155 ;
      LAYER nwell ;
        RECT 17.130 200.125 147.230 202.955 ;
      LAYER pwell ;
        RECT 17.325 198.925 18.695 199.735 ;
        RECT 18.705 198.925 24.215 199.735 ;
        RECT 24.225 198.925 29.735 199.735 ;
        RECT 30.215 199.010 30.645 199.795 ;
        RECT 30.665 198.925 36.175 199.735 ;
        RECT 36.185 198.925 41.695 199.735 ;
        RECT 41.705 198.925 45.375 199.735 ;
        RECT 49.360 199.605 50.270 199.825 ;
        RECT 51.805 199.605 53.155 199.835 ;
        RECT 45.845 198.925 53.155 199.605 ;
        RECT 54.125 198.925 55.940 199.835 ;
        RECT 55.975 199.010 56.405 199.795 ;
        RECT 58.500 199.605 59.635 199.835 ;
        RECT 56.425 198.925 59.635 199.605 ;
        RECT 60.105 199.605 61.025 199.835 ;
        RECT 60.105 198.925 62.395 199.605 ;
        RECT 62.505 198.925 65.615 199.835 ;
        RECT 69.140 199.605 70.050 199.825 ;
        RECT 71.585 199.605 72.935 199.835 ;
        RECT 74.320 199.635 75.275 199.835 ;
        RECT 65.625 198.925 72.935 199.605 ;
        RECT 72.995 198.955 75.275 199.635 ;
        RECT 17.465 198.715 17.635 198.925 ;
        RECT 18.845 198.715 19.015 198.925 ;
        RECT 24.365 198.715 24.535 198.925 ;
        RECT 29.885 198.875 30.055 198.905 ;
        RECT 29.880 198.765 30.055 198.875 ;
        RECT 29.885 198.715 30.055 198.765 ;
        RECT 30.805 198.735 30.975 198.925 ;
        RECT 35.405 198.715 35.575 198.905 ;
        RECT 36.325 198.735 36.495 198.925 ;
        RECT 40.925 198.715 41.095 198.905 ;
        RECT 41.845 198.735 42.015 198.925 ;
        RECT 42.760 198.765 42.880 198.875 ;
        RECT 43.685 198.715 43.855 198.905 ;
        RECT 45.520 198.765 45.640 198.875 ;
        RECT 45.985 198.735 46.155 198.925 ;
        RECT 49.205 198.715 49.375 198.905 ;
        RECT 50.590 198.715 50.760 198.905 ;
        RECT 51.965 198.715 52.135 198.905 ;
        RECT 53.355 198.770 53.515 198.880 ;
        RECT 54.720 198.765 54.840 198.875 ;
        RECT 55.645 198.735 55.815 198.925 ;
        RECT 56.105 198.715 56.275 198.905 ;
        RECT 56.565 198.715 56.735 198.925 ;
        RECT 59.780 198.765 59.900 198.875 ;
        RECT 62.085 198.715 62.255 198.925 ;
        RECT 62.545 198.735 62.715 198.925 ;
        RECT 65.300 198.715 65.470 198.905 ;
        RECT 65.765 198.735 65.935 198.925 ;
        RECT 68.525 198.715 68.695 198.905 ;
        RECT 70.825 198.715 70.995 198.905 ;
        RECT 71.285 198.715 71.455 198.905 ;
        RECT 73.120 198.735 73.290 198.955 ;
        RECT 74.320 198.925 75.275 198.955 ;
        RECT 75.285 198.925 80.795 199.735 ;
        RECT 81.735 199.010 82.165 199.795 ;
        RECT 82.645 199.605 85.470 199.835 ;
        RECT 86.420 199.605 87.340 199.835 ;
        RECT 90.005 199.635 90.950 199.835 ;
        RECT 92.285 199.635 93.215 199.835 ;
        RECT 82.645 198.925 86.175 199.605 ;
        RECT 86.420 198.925 89.885 199.605 ;
        RECT 90.005 199.155 93.215 199.635 ;
        RECT 94.275 199.605 95.205 199.835 ;
        RECT 90.005 198.955 93.075 199.155 ;
        RECT 90.005 198.925 90.950 198.955 ;
        RECT 75.425 198.735 75.595 198.925 ;
        RECT 85.975 198.905 86.175 198.925 ;
        RECT 76.805 198.715 76.975 198.905 ;
        RECT 80.955 198.770 81.115 198.880 ;
        RECT 82.325 198.875 82.495 198.905 ;
        RECT 82.320 198.765 82.495 198.875 ;
        RECT 85.080 198.765 85.200 198.875 ;
        RECT 82.325 198.715 82.495 198.765 ;
        RECT 85.545 198.715 85.715 198.905 ;
        RECT 86.005 198.735 86.175 198.905 ;
        RECT 88.305 198.715 88.475 198.905 ;
        RECT 89.685 198.735 89.855 198.925 ;
        RECT 92.905 198.735 93.075 198.955 ;
        RECT 93.370 198.925 95.205 199.605 ;
        RECT 95.525 198.925 97.355 199.735 ;
        RECT 97.365 198.925 101.025 199.835 ;
        RECT 101.045 198.925 106.555 199.735 ;
        RECT 107.495 199.010 107.925 199.795 ;
        RECT 107.945 198.925 113.455 199.735 ;
        RECT 113.465 198.925 118.975 199.735 ;
        RECT 118.985 198.925 124.495 199.735 ;
        RECT 124.505 198.925 130.015 199.735 ;
        RECT 130.025 198.925 132.775 199.735 ;
        RECT 133.255 199.010 133.685 199.795 ;
        RECT 133.705 198.925 139.215 199.735 ;
        RECT 139.225 198.925 144.735 199.735 ;
        RECT 145.665 198.925 147.035 199.735 ;
        RECT 93.370 198.905 93.535 198.925 ;
        RECT 93.365 198.735 93.535 198.905 ;
        RECT 93.835 198.760 93.995 198.870 ;
        RECT 95.210 198.715 95.380 198.905 ;
        RECT 95.665 198.735 95.835 198.925 ;
        RECT 96.585 198.715 96.755 198.905 ;
        RECT 100.730 198.735 100.900 198.925 ;
        RECT 101.185 198.735 101.355 198.925 ;
        RECT 102.105 198.715 102.275 198.905 ;
        RECT 106.715 198.770 106.875 198.880 ;
        RECT 107.625 198.715 107.795 198.905 ;
        RECT 108.085 198.735 108.255 198.925 ;
        RECT 110.380 198.765 110.500 198.875 ;
        RECT 110.845 198.715 111.015 198.905 ;
        RECT 113.605 198.735 113.775 198.925 ;
        RECT 114.525 198.715 114.695 198.905 ;
        RECT 119.125 198.735 119.295 198.925 ;
        RECT 120.040 198.765 120.160 198.875 ;
        RECT 120.965 198.715 121.135 198.905 ;
        RECT 124.645 198.735 124.815 198.925 ;
        RECT 126.485 198.715 126.655 198.905 ;
        RECT 130.165 198.735 130.335 198.925 ;
        RECT 132.005 198.715 132.175 198.905 ;
        RECT 132.920 198.765 133.040 198.875 ;
        RECT 133.845 198.735 134.015 198.925 ;
        RECT 137.525 198.715 137.695 198.905 ;
        RECT 139.365 198.735 139.535 198.925 ;
        RECT 143.045 198.715 143.215 198.905 ;
        RECT 144.895 198.770 145.055 198.880 ;
        RECT 146.725 198.715 146.895 198.925 ;
        RECT 17.325 197.905 18.695 198.715 ;
        RECT 18.705 197.905 24.215 198.715 ;
        RECT 24.225 197.905 29.735 198.715 ;
        RECT 29.745 197.905 35.255 198.715 ;
        RECT 35.265 197.905 40.775 198.715 ;
        RECT 40.785 197.905 42.615 198.715 ;
        RECT 43.095 197.845 43.525 198.630 ;
        RECT 43.545 197.905 49.055 198.715 ;
        RECT 49.065 197.905 50.435 198.715 ;
        RECT 50.445 197.805 51.795 198.715 ;
        RECT 51.825 197.905 54.575 198.715 ;
        RECT 55.055 197.805 56.405 198.715 ;
        RECT 56.425 197.905 61.935 198.715 ;
        RECT 61.945 197.905 63.775 198.715 ;
        RECT 63.845 197.805 65.615 198.715 ;
        RECT 66.545 198.035 68.835 198.715 ;
        RECT 66.545 197.805 67.465 198.035 ;
        RECT 68.855 197.845 69.285 198.630 ;
        RECT 69.305 198.035 71.135 198.715 ;
        RECT 69.305 197.805 70.650 198.035 ;
        RECT 71.145 197.905 76.655 198.715 ;
        RECT 76.665 197.905 82.175 198.715 ;
        RECT 82.185 197.905 84.935 198.715 ;
        RECT 85.405 197.805 88.155 198.715 ;
        RECT 88.165 197.905 93.675 198.715 ;
        RECT 94.615 197.845 95.045 198.630 ;
        RECT 95.065 197.805 96.415 198.715 ;
        RECT 96.445 197.905 101.955 198.715 ;
        RECT 101.965 197.905 107.475 198.715 ;
        RECT 107.485 197.905 110.235 198.715 ;
        RECT 110.815 198.035 114.280 198.715 ;
        RECT 113.360 197.805 114.280 198.035 ;
        RECT 114.385 197.905 119.895 198.715 ;
        RECT 120.375 197.845 120.805 198.630 ;
        RECT 120.825 197.905 126.335 198.715 ;
        RECT 126.345 197.905 131.855 198.715 ;
        RECT 131.865 197.905 137.375 198.715 ;
        RECT 137.385 197.905 142.895 198.715 ;
        RECT 142.905 197.905 145.655 198.715 ;
        RECT 145.665 197.905 147.035 198.715 ;
      LAYER nwell ;
        RECT 17.130 194.685 147.230 197.515 ;
      LAYER pwell ;
        RECT 17.325 193.485 18.695 194.295 ;
        RECT 18.705 193.485 24.215 194.295 ;
        RECT 24.225 193.485 26.055 194.295 ;
        RECT 26.065 193.485 27.895 194.395 ;
        RECT 27.905 193.485 29.735 194.295 ;
        RECT 30.215 193.570 30.645 194.355 ;
        RECT 30.665 193.485 36.175 194.295 ;
        RECT 36.185 193.485 38.935 194.295 ;
        RECT 38.945 193.485 40.775 194.165 ;
        RECT 40.785 193.485 46.295 194.295 ;
        RECT 46.305 193.485 51.815 194.295 ;
        RECT 51.825 193.485 53.655 194.295 ;
        RECT 54.715 194.165 55.645 194.395 ;
        RECT 53.810 193.485 55.645 194.165 ;
        RECT 55.975 193.570 56.405 194.355 ;
        RECT 56.425 193.485 59.175 194.395 ;
        RECT 59.200 193.485 61.015 194.395 ;
        RECT 61.025 193.485 66.535 194.295 ;
        RECT 66.545 193.485 72.055 194.295 ;
        RECT 72.065 193.485 77.575 194.295 ;
        RECT 77.585 193.485 79.415 194.295 ;
        RECT 79.885 193.485 81.715 194.395 ;
        RECT 81.735 193.570 82.165 194.355 ;
        RECT 85.700 194.165 86.610 194.385 ;
        RECT 88.145 194.165 89.495 194.395 ;
        RECT 82.185 193.485 89.495 194.165 ;
        RECT 89.640 194.165 90.560 194.395 ;
        RECT 93.225 194.195 94.170 194.395 ;
        RECT 95.505 194.195 96.435 194.395 ;
        RECT 89.640 193.485 93.105 194.165 ;
        RECT 93.225 193.715 96.435 194.195 ;
        RECT 99.960 194.165 100.870 194.385 ;
        RECT 102.405 194.165 103.755 194.395 ;
        RECT 93.225 193.515 96.295 193.715 ;
        RECT 93.225 193.485 94.170 193.515 ;
        RECT 17.465 193.275 17.635 193.485 ;
        RECT 18.845 193.275 19.015 193.485 ;
        RECT 20.225 193.275 20.395 193.465 ;
        RECT 21.605 193.275 21.775 193.465 ;
        RECT 24.365 193.295 24.535 193.485 ;
        RECT 25.285 193.275 25.455 193.465 ;
        RECT 27.580 193.295 27.750 193.485 ;
        RECT 28.045 193.295 28.215 193.485 ;
        RECT 29.880 193.325 30.000 193.435 ;
        RECT 30.805 193.295 30.975 193.485 ;
        RECT 32.645 193.275 32.815 193.465 ;
        RECT 36.325 193.295 36.495 193.485 ;
        RECT 39.085 193.295 39.255 193.485 ;
        RECT 40.010 193.275 40.180 193.465 ;
        RECT 40.925 193.295 41.095 193.485 ;
        RECT 42.765 193.275 42.935 193.465 ;
        RECT 46.445 193.295 46.615 193.485 ;
        RECT 49.205 193.275 49.375 193.465 ;
        RECT 49.665 193.275 49.835 193.465 ;
        RECT 51.045 193.275 51.215 193.465 ;
        RECT 51.965 193.295 52.135 193.485 ;
        RECT 53.810 193.465 53.975 193.485 ;
        RECT 53.805 193.275 53.975 193.465 ;
        RECT 17.325 192.465 18.695 193.275 ;
        RECT 18.705 192.495 20.075 193.275 ;
        RECT 20.085 192.465 21.455 193.275 ;
        RECT 21.465 192.595 24.215 193.275 ;
        RECT 25.145 192.595 32.455 193.275 ;
        RECT 32.505 192.595 39.815 193.275 ;
        RECT 23.285 192.365 24.215 192.595 ;
        RECT 28.660 192.375 29.570 192.595 ;
        RECT 31.105 192.365 32.455 192.595 ;
        RECT 36.020 192.375 36.930 192.595 ;
        RECT 38.465 192.365 39.815 192.595 ;
        RECT 39.865 192.365 41.215 193.275 ;
        RECT 41.245 192.595 43.075 193.275 ;
        RECT 41.245 192.365 42.590 192.595 ;
        RECT 43.095 192.405 43.525 193.190 ;
        RECT 43.695 192.365 49.515 193.275 ;
        RECT 49.525 192.465 50.895 193.275 ;
        RECT 50.905 192.365 53.310 193.275 ;
        RECT 53.665 192.595 56.875 193.275 ;
        RECT 57.030 193.245 57.200 193.465 ;
        RECT 58.865 193.295 59.035 193.485 ;
        RECT 59.325 193.295 59.495 193.485 ;
        RECT 60.705 193.275 60.875 193.465 ;
        RECT 61.165 193.295 61.335 193.485 ;
        RECT 64.385 193.275 64.555 193.465 ;
        RECT 64.845 193.275 65.015 193.465 ;
        RECT 66.685 193.295 66.855 193.485 ;
        RECT 68.520 193.325 68.640 193.435 ;
        RECT 69.440 193.325 69.560 193.435 ;
        RECT 72.205 193.295 72.375 193.485 ;
        RECT 73.125 193.275 73.295 193.465 ;
        RECT 75.425 193.295 75.595 193.465 ;
        RECT 75.880 193.325 76.000 193.435 ;
        RECT 77.725 193.295 77.895 193.485 ;
        RECT 79.560 193.325 79.680 193.435 ;
        RECT 80.030 193.295 80.200 193.485 ;
        RECT 75.425 193.275 75.575 193.295 ;
        RECT 80.945 193.275 81.115 193.465 ;
        RECT 82.325 193.275 82.495 193.485 ;
        RECT 82.785 193.275 82.955 193.465 ;
        RECT 86.475 193.320 86.635 193.430 ;
        RECT 87.385 193.275 87.555 193.465 ;
        RECT 92.905 193.295 93.075 193.485 ;
        RECT 95.480 193.275 95.650 193.465 ;
        RECT 96.125 193.295 96.295 193.515 ;
        RECT 96.445 193.485 103.755 194.165 ;
        RECT 103.900 194.165 104.820 194.395 ;
        RECT 103.900 193.485 107.365 194.165 ;
        RECT 107.495 193.570 107.925 194.355 ;
        RECT 108.445 194.165 109.795 194.395 ;
        RECT 111.330 194.165 112.240 194.385 ;
        RECT 108.445 193.485 115.755 194.165 ;
        RECT 115.765 193.485 121.275 194.295 ;
        RECT 121.285 193.485 126.795 194.295 ;
        RECT 126.805 193.485 132.315 194.295 ;
        RECT 133.255 193.570 133.685 194.355 ;
        RECT 133.705 193.485 139.215 194.295 ;
        RECT 139.225 193.485 144.735 194.295 ;
        RECT 145.665 193.485 147.035 194.295 ;
        RECT 96.585 193.295 96.755 193.485 ;
        RECT 99.340 193.295 99.510 193.465 ;
        RECT 99.375 193.275 99.510 193.295 ;
        RECT 103.030 193.275 103.200 193.465 ;
        RECT 106.245 193.275 106.415 193.465 ;
        RECT 107.165 193.295 107.335 193.485 ;
        RECT 107.625 193.275 107.795 193.465 ;
        RECT 108.080 193.325 108.200 193.435 ;
        RECT 114.710 193.275 114.880 193.465 ;
        RECT 115.445 193.275 115.615 193.485 ;
        RECT 115.905 193.295 116.075 193.485 ;
        RECT 119.125 193.275 119.295 193.465 ;
        RECT 120.965 193.275 121.135 193.465 ;
        RECT 121.425 193.295 121.595 193.485 ;
        RECT 126.485 193.275 126.655 193.465 ;
        RECT 126.945 193.295 127.115 193.485 ;
        RECT 132.005 193.275 132.175 193.465 ;
        RECT 132.475 193.330 132.635 193.440 ;
        RECT 133.845 193.295 134.015 193.485 ;
        RECT 137.525 193.275 137.695 193.465 ;
        RECT 139.365 193.295 139.535 193.485 ;
        RECT 143.045 193.275 143.215 193.465 ;
        RECT 144.895 193.330 145.055 193.440 ;
        RECT 146.725 193.275 146.895 193.485 ;
        RECT 59.605 193.245 60.555 193.275 ;
        RECT 55.740 192.365 56.875 192.595 ;
        RECT 56.885 192.565 60.555 193.245 ;
        RECT 59.605 192.365 60.555 192.565 ;
        RECT 60.565 192.365 63.315 193.275 ;
        RECT 63.335 192.365 64.685 193.275 ;
        RECT 64.705 192.465 68.375 193.275 ;
        RECT 68.855 192.405 69.285 193.190 ;
        RECT 69.860 192.595 73.325 193.275 ;
        RECT 69.860 192.365 70.780 192.595 ;
        RECT 73.645 192.455 75.575 193.275 ;
        RECT 76.440 192.595 81.255 193.275 ;
        RECT 73.645 192.365 74.595 192.455 ;
        RECT 81.275 192.365 82.625 193.275 ;
        RECT 82.755 192.595 86.220 193.275 ;
        RECT 87.245 192.595 94.555 193.275 ;
        RECT 85.300 192.365 86.220 192.595 ;
        RECT 90.760 192.375 91.670 192.595 ;
        RECT 93.205 192.365 94.555 192.595 ;
        RECT 94.615 192.405 95.045 193.190 ;
        RECT 95.065 192.595 98.965 193.275 ;
        RECT 95.065 192.365 95.995 192.595 ;
        RECT 99.375 192.365 102.875 193.275 ;
        RECT 102.885 192.365 105.805 193.275 ;
        RECT 106.115 192.365 107.465 193.275 ;
        RECT 107.485 192.465 111.155 193.275 ;
        RECT 111.395 192.595 115.295 193.275 ;
        RECT 114.365 192.365 115.295 192.595 ;
        RECT 115.305 192.465 118.975 193.275 ;
        RECT 118.985 192.465 120.355 193.275 ;
        RECT 120.375 192.405 120.805 193.190 ;
        RECT 120.825 192.465 126.335 193.275 ;
        RECT 126.345 192.465 131.855 193.275 ;
        RECT 131.865 192.465 137.375 193.275 ;
        RECT 137.385 192.465 142.895 193.275 ;
        RECT 142.905 192.465 145.655 193.275 ;
        RECT 145.665 192.465 147.035 193.275 ;
      LAYER nwell ;
        RECT 17.130 189.245 147.230 192.075 ;
      LAYER pwell ;
        RECT 17.325 188.045 18.695 188.855 ;
        RECT 18.705 188.045 21.455 188.855 ;
        RECT 24.980 188.725 25.890 188.945 ;
        RECT 27.425 188.725 28.775 188.955 ;
        RECT 21.465 188.045 28.775 188.725 ;
        RECT 28.845 188.045 30.195 188.955 ;
        RECT 30.215 188.130 30.645 188.915 ;
        RECT 30.675 188.045 33.405 188.955 ;
        RECT 34.475 188.725 35.405 188.955 ;
        RECT 33.570 188.045 35.405 188.725 ;
        RECT 35.725 188.725 36.645 188.955 ;
        RECT 35.725 188.045 38.015 188.725 ;
        RECT 38.945 188.045 41.555 188.955 ;
        RECT 42.165 188.275 45.365 188.955 ;
        RECT 46.435 188.725 47.365 188.955 ;
        RECT 42.310 188.045 45.365 188.275 ;
        RECT 45.530 188.045 47.365 188.725 ;
        RECT 48.620 188.045 50.435 188.955 ;
        RECT 51.585 188.865 52.535 188.955 ;
        RECT 50.605 188.045 52.535 188.865 ;
        RECT 53.035 188.045 55.955 188.955 ;
        RECT 55.975 188.130 56.405 188.915 ;
        RECT 56.435 188.045 57.785 188.955 ;
        RECT 59.385 188.725 62.385 188.955 ;
        RECT 57.805 188.635 62.385 188.725 ;
        RECT 62.405 188.755 63.350 188.955 ;
        RECT 64.685 188.755 65.615 188.955 ;
        RECT 57.805 188.275 62.395 188.635 ;
        RECT 57.805 188.045 59.375 188.275 ;
        RECT 61.465 188.085 62.395 188.275 ;
        RECT 62.405 188.275 65.615 188.755 ;
        RECT 61.465 188.045 62.385 188.085 ;
        RECT 62.405 188.075 65.475 188.275 ;
        RECT 62.405 188.045 63.350 188.075 ;
        RECT 17.465 187.835 17.635 188.045 ;
        RECT 18.845 187.995 19.015 188.045 ;
        RECT 18.840 187.885 19.015 187.995 ;
        RECT 18.845 187.855 19.015 187.885 ;
        RECT 21.605 187.855 21.775 188.045 ;
        RECT 26.205 187.835 26.375 188.025 ;
        RECT 28.960 187.855 29.130 188.045 ;
        RECT 29.425 187.835 29.595 188.025 ;
        RECT 29.890 187.835 30.060 188.025 ;
        RECT 30.805 187.855 30.975 188.045 ;
        RECT 33.570 188.025 33.735 188.045 ;
        RECT 33.100 187.885 33.220 187.995 ;
        RECT 33.560 187.855 33.735 188.025 ;
        RECT 37.705 187.855 37.875 188.045 ;
        RECT 39.090 188.025 39.260 188.045 ;
        RECT 38.175 187.890 38.335 188.000 ;
        RECT 17.325 187.025 18.695 187.835 ;
        RECT 19.205 187.155 26.515 187.835 ;
        RECT 26.525 187.155 29.735 187.835 ;
        RECT 19.205 186.925 20.555 187.155 ;
        RECT 22.090 186.935 23.000 187.155 ;
        RECT 26.525 186.925 27.660 187.155 ;
        RECT 29.745 186.925 32.665 187.835 ;
        RECT 33.560 187.805 33.730 187.855 ;
        RECT 38.625 187.835 38.795 188.025 ;
        RECT 39.085 187.855 39.260 188.025 ;
        RECT 41.840 187.885 41.960 187.995 ;
        RECT 42.310 187.855 42.480 188.045 ;
        RECT 45.530 188.025 45.695 188.045 ;
        RECT 39.085 187.835 39.255 187.855 ;
        RECT 43.690 187.835 43.860 188.025 ;
        RECT 45.525 187.855 45.695 188.025 ;
        RECT 47.365 187.835 47.535 188.025 ;
        RECT 47.825 187.835 47.995 188.025 ;
        RECT 48.745 187.855 48.915 188.045 ;
        RECT 50.605 188.025 50.755 188.045 ;
        RECT 50.585 187.995 50.755 188.025 ;
        RECT 50.580 187.885 50.755 187.995 ;
        RECT 50.585 187.855 50.755 187.885 ;
        RECT 51.040 187.835 51.210 188.025 ;
        RECT 34.760 187.805 35.715 187.835 ;
        RECT 33.435 187.125 35.715 187.805 ;
        RECT 34.760 186.925 35.715 187.125 ;
        RECT 35.725 186.925 38.935 187.835 ;
        RECT 38.945 186.925 42.155 187.835 ;
        RECT 43.095 186.965 43.525 187.750 ;
        RECT 43.690 187.605 45.380 187.835 ;
        RECT 43.545 186.925 45.380 187.605 ;
        RECT 45.845 187.155 47.675 187.835 ;
        RECT 47.685 187.025 50.435 187.835 ;
        RECT 50.925 186.925 52.275 187.835 ;
        RECT 52.420 187.805 52.590 188.025 ;
        RECT 54.725 187.835 54.895 188.025 ;
        RECT 55.640 187.855 55.810 188.045 ;
        RECT 57.485 187.855 57.655 188.045 ;
        RECT 57.945 187.855 58.115 188.045 ;
        RECT 61.160 187.835 61.330 188.025 ;
        RECT 63.925 187.835 64.095 188.025 ;
        RECT 64.385 187.835 64.555 188.025 ;
        RECT 65.305 187.855 65.475 188.075 ;
        RECT 65.625 188.045 67.455 188.955 ;
        RECT 67.465 188.045 68.835 188.855 ;
        RECT 68.845 188.045 70.195 188.955 ;
        RECT 73.740 188.725 74.650 188.945 ;
        RECT 76.185 188.725 77.535 188.955 ;
        RECT 70.225 188.045 77.535 188.725 ;
        RECT 78.050 188.045 79.415 188.725 ;
        RECT 79.425 188.045 81.255 188.855 ;
        RECT 81.735 188.130 82.165 188.915 ;
        RECT 82.185 188.045 84.015 188.855 ;
        RECT 84.035 188.045 86.765 188.955 ;
        RECT 86.785 188.045 88.615 188.855 ;
        RECT 89.085 188.045 90.435 188.955 ;
        RECT 90.485 188.045 91.835 188.955 ;
        RECT 91.855 188.045 93.205 188.955 ;
        RECT 93.235 188.045 95.965 188.955 ;
        RECT 95.985 188.045 99.655 188.955 ;
        RECT 99.975 188.725 100.905 188.955 ;
        RECT 99.975 188.045 101.810 188.725 ;
        RECT 101.980 188.045 105.635 188.955 ;
        RECT 105.655 188.045 107.005 188.955 ;
        RECT 107.495 188.130 107.925 188.915 ;
        RECT 107.945 188.045 109.295 188.955 ;
        RECT 110.245 188.725 111.175 188.955 ;
        RECT 114.480 188.725 115.400 188.955 ;
        RECT 110.245 188.045 114.145 188.725 ;
        RECT 114.480 188.045 117.945 188.725 ;
        RECT 118.065 188.045 121.735 188.855 ;
        RECT 122.205 188.045 125.415 188.955 ;
        RECT 125.425 188.045 130.935 188.855 ;
        RECT 130.945 188.045 132.775 188.855 ;
        RECT 133.255 188.130 133.685 188.915 ;
        RECT 133.705 188.045 139.215 188.855 ;
        RECT 139.225 188.045 144.735 188.855 ;
        RECT 145.665 188.045 147.035 188.855 ;
        RECT 65.770 187.855 65.940 188.045 ;
        RECT 67.605 187.855 67.775 188.045 ;
        RECT 68.075 187.880 68.235 187.990 ;
        RECT 68.990 187.855 69.160 188.045 ;
        RECT 69.445 187.835 69.615 188.025 ;
        RECT 70.365 187.855 70.535 188.045 ;
        RECT 71.290 187.835 71.460 188.025 ;
        RECT 77.725 187.855 77.895 188.025 ;
        RECT 79.565 187.855 79.735 188.045 ;
        RECT 80.025 187.835 80.195 188.025 ;
        RECT 80.480 187.885 80.600 187.995 ;
        RECT 80.945 187.835 81.115 188.025 ;
        RECT 81.400 187.885 81.520 187.995 ;
        RECT 82.325 187.855 82.495 188.045 ;
        RECT 84.165 187.855 84.335 188.045 ;
        RECT 86.925 187.855 87.095 188.045 ;
        RECT 88.305 187.835 88.475 188.025 ;
        RECT 88.760 187.885 88.880 187.995 ;
        RECT 90.150 187.855 90.320 188.045 ;
        RECT 91.520 187.855 91.690 188.045 ;
        RECT 92.905 187.855 93.075 188.045 ;
        RECT 93.835 187.880 93.995 187.990 ;
        RECT 95.205 187.835 95.375 188.025 ;
        RECT 95.665 187.855 95.835 188.045 ;
        RECT 96.125 187.855 96.295 188.045 ;
        RECT 101.645 188.025 101.810 188.045 ;
        RECT 97.965 187.835 98.135 188.025 ;
        RECT 101.180 187.885 101.300 187.995 ;
        RECT 101.645 187.855 101.815 188.025 ;
        RECT 104.400 187.835 104.570 188.025 ;
        RECT 104.865 187.835 105.035 188.025 ;
        RECT 105.320 187.855 105.490 188.045 ;
        RECT 105.785 187.855 105.955 188.045 ;
        RECT 106.245 187.835 106.415 188.025 ;
        RECT 107.160 187.885 107.280 187.995 ;
        RECT 107.625 187.835 107.795 188.025 ;
        RECT 108.090 187.855 108.260 188.045 ;
        RECT 109.475 187.890 109.635 188.000 ;
        RECT 110.660 187.855 110.830 188.045 ;
        RECT 114.985 187.835 115.155 188.025 ;
        RECT 117.745 187.855 117.915 188.045 ;
        RECT 118.205 187.855 118.375 188.045 ;
        RECT 121.240 187.835 121.410 188.025 ;
        RECT 121.880 187.885 122.000 187.995 ;
        RECT 125.105 187.855 125.275 188.045 ;
        RECT 125.565 187.855 125.735 188.045 ;
        RECT 131.085 187.855 131.255 188.045 ;
        RECT 132.925 187.995 133.095 188.025 ;
        RECT 132.920 187.885 133.095 187.995 ;
        RECT 132.925 187.835 133.095 187.885 ;
        RECT 133.845 187.855 134.015 188.045 ;
        RECT 134.765 187.835 134.935 188.025 ;
        RECT 135.225 187.835 135.395 188.025 ;
        RECT 139.365 187.855 139.535 188.045 ;
        RECT 140.745 187.835 140.915 188.025 ;
        RECT 144.425 187.835 144.595 188.025 ;
        RECT 144.895 187.890 145.055 188.000 ;
        RECT 146.725 187.835 146.895 188.045 ;
        RECT 53.620 187.805 54.575 187.835 ;
        RECT 52.295 187.125 54.575 187.805 ;
        RECT 53.620 186.925 54.575 187.125 ;
        RECT 54.585 186.925 57.795 187.835 ;
        RECT 58.000 186.925 61.475 187.835 ;
        RECT 61.495 186.925 64.225 187.835 ;
        RECT 64.245 187.025 67.915 187.835 ;
        RECT 68.855 186.965 69.285 187.750 ;
        RECT 69.305 187.025 71.135 187.835 ;
        RECT 71.145 186.925 72.915 187.835 ;
        RECT 73.025 187.155 80.335 187.835 ;
        RECT 80.805 187.155 88.115 187.835 ;
        RECT 73.025 186.925 74.375 187.155 ;
        RECT 75.910 186.935 76.820 187.155 ;
        RECT 84.320 186.935 85.230 187.155 ;
        RECT 86.765 186.925 88.115 187.155 ;
        RECT 88.165 187.025 93.675 187.835 ;
        RECT 94.615 186.965 95.045 187.750 ;
        RECT 95.065 187.025 97.815 187.835 ;
        RECT 97.825 186.925 101.035 187.835 ;
        RECT 101.795 186.925 104.715 187.835 ;
        RECT 104.735 186.925 106.085 187.835 ;
        RECT 106.105 187.025 107.475 187.835 ;
        RECT 107.485 187.155 114.795 187.835 ;
        RECT 111.000 186.935 111.910 187.155 ;
        RECT 113.445 186.925 114.795 187.155 ;
        RECT 114.845 187.025 120.355 187.835 ;
        RECT 120.375 186.965 120.805 187.750 ;
        RECT 120.825 187.155 124.725 187.835 ;
        RECT 125.925 187.155 133.235 187.835 ;
        RECT 133.245 187.155 135.075 187.835 ;
        RECT 120.825 186.925 121.755 187.155 ;
        RECT 125.925 186.925 127.275 187.155 ;
        RECT 128.810 186.935 129.720 187.155 ;
        RECT 135.085 187.025 140.595 187.835 ;
        RECT 140.605 187.025 144.275 187.835 ;
        RECT 144.285 187.025 145.655 187.835 ;
        RECT 145.665 187.025 147.035 187.835 ;
      LAYER nwell ;
        RECT 17.130 183.805 147.230 186.635 ;
      LAYER pwell ;
        RECT 17.325 182.605 18.695 183.415 ;
        RECT 18.705 182.605 22.375 183.415 ;
        RECT 22.845 183.285 23.765 183.515 ;
        RECT 26.065 183.285 26.985 183.515 ;
        RECT 22.845 182.605 25.135 183.285 ;
        RECT 26.065 182.605 28.355 183.285 ;
        RECT 28.375 182.605 29.725 183.515 ;
        RECT 30.215 182.690 30.645 183.475 ;
        RECT 30.665 182.605 36.175 183.415 ;
        RECT 36.185 182.605 37.555 183.415 ;
        RECT 37.565 182.605 40.315 183.515 ;
        RECT 40.345 182.605 41.695 183.515 ;
        RECT 41.905 183.425 42.855 183.515 ;
        RECT 41.905 182.605 43.835 183.425 ;
        RECT 44.060 182.605 54.080 183.515 ;
        RECT 54.125 182.605 55.955 183.415 ;
        RECT 55.975 182.690 56.405 183.475 ;
        RECT 56.425 182.605 59.635 183.515 ;
        RECT 59.845 183.425 60.795 183.515 ;
        RECT 59.845 182.605 61.775 183.425 ;
        RECT 61.945 182.605 67.455 183.415 ;
        RECT 67.465 182.605 71.135 183.415 ;
        RECT 71.145 182.605 72.515 183.415 ;
        RECT 72.625 182.605 75.735 183.515 ;
        RECT 76.900 182.605 81.715 183.285 ;
        RECT 81.735 182.690 82.165 183.475 ;
        RECT 82.185 182.605 87.695 183.415 ;
        RECT 87.705 182.605 91.375 183.415 ;
        RECT 91.480 183.285 92.400 183.515 ;
        RECT 98.580 183.285 99.490 183.505 ;
        RECT 101.025 183.285 102.375 183.515 ;
        RECT 91.480 182.605 94.945 183.285 ;
        RECT 95.065 182.605 102.375 183.285 ;
        RECT 102.425 183.285 103.355 183.515 ;
        RECT 102.425 182.605 106.325 183.285 ;
        RECT 107.495 182.690 107.925 183.475 ;
        RECT 111.460 183.285 112.370 183.505 ;
        RECT 113.905 183.285 115.255 183.515 ;
        RECT 107.945 182.605 115.255 183.285 ;
        RECT 115.305 182.605 118.055 183.415 ;
        RECT 118.065 183.285 118.995 183.515 ;
        RECT 124.860 183.285 125.780 183.515 ;
        RECT 118.065 182.605 121.965 183.285 ;
        RECT 122.315 182.605 125.780 183.285 ;
        RECT 125.885 182.605 127.255 183.415 ;
        RECT 129.920 183.285 130.840 183.515 ;
        RECT 131.430 183.285 132.775 183.515 ;
        RECT 127.375 182.605 130.840 183.285 ;
        RECT 130.945 182.605 132.775 183.285 ;
        RECT 133.255 182.690 133.685 183.475 ;
        RECT 133.705 182.605 136.915 183.515 ;
        RECT 136.925 182.605 142.435 183.415 ;
        RECT 142.445 182.605 145.195 183.415 ;
        RECT 145.665 182.605 147.035 183.415 ;
        RECT 17.465 182.395 17.635 182.605 ;
        RECT 18.845 182.395 19.015 182.605 ;
        RECT 24.825 182.585 24.995 182.605 ;
        RECT 22.520 182.445 22.640 182.555 ;
        RECT 24.360 182.445 24.480 182.555 ;
        RECT 24.820 182.415 24.995 182.585 ;
        RECT 25.295 182.450 25.455 182.560 ;
        RECT 24.820 182.395 24.990 182.415 ;
        RECT 26.205 182.395 26.375 182.585 ;
        RECT 28.045 182.415 28.215 182.605 ;
        RECT 28.505 182.415 28.675 182.605 ;
        RECT 29.880 182.445 30.000 182.555 ;
        RECT 30.805 182.415 30.975 182.605 ;
        RECT 31.725 182.395 31.895 182.585 ;
        RECT 36.325 182.415 36.495 182.605 ;
        RECT 37.710 182.415 37.880 182.605 ;
        RECT 38.620 182.395 38.790 182.585 ;
        RECT 40.460 182.415 40.630 182.605 ;
        RECT 43.685 182.585 43.835 182.605 ;
        RECT 42.300 182.395 42.470 182.585 ;
        RECT 42.760 182.445 42.880 182.555 ;
        RECT 43.685 182.395 43.855 182.585 ;
        RECT 44.145 182.415 44.315 182.605 ;
        RECT 48.745 182.395 48.915 182.585 ;
        RECT 54.265 182.395 54.435 182.605 ;
        RECT 54.725 182.395 54.895 182.585 ;
        RECT 56.565 182.395 56.735 182.605 ;
        RECT 61.625 182.585 61.775 182.605 ;
        RECT 59.780 182.395 59.950 182.585 ;
        RECT 60.240 182.445 60.360 182.555 ;
        RECT 17.325 181.585 18.695 182.395 ;
        RECT 18.705 181.585 24.215 182.395 ;
        RECT 24.705 181.485 26.055 182.395 ;
        RECT 26.065 181.585 31.575 182.395 ;
        RECT 31.585 181.585 35.255 182.395 ;
        RECT 35.460 181.485 38.935 182.395 ;
        RECT 39.140 181.485 42.615 182.395 ;
        RECT 43.095 181.525 43.525 182.310 ;
        RECT 43.545 181.715 48.360 182.395 ;
        RECT 48.655 181.485 51.815 182.395 ;
        RECT 52.485 181.585 54.575 182.395 ;
        RECT 54.585 181.585 56.415 182.395 ;
        RECT 56.435 181.485 57.785 182.395 ;
        RECT 57.820 181.715 60.095 182.395 ;
        RECT 60.710 182.365 60.880 182.585 ;
        RECT 61.625 182.415 61.795 182.585 ;
        RECT 62.085 182.415 62.255 182.605 ;
        RECT 63.465 182.395 63.635 182.585 ;
        RECT 66.685 182.415 66.855 182.585 ;
        RECT 67.605 182.415 67.775 182.605 ;
        RECT 66.690 182.395 66.855 182.415 ;
        RECT 70.825 182.395 70.995 182.585 ;
        RECT 71.285 182.395 71.455 182.605 ;
        RECT 72.665 182.415 72.835 182.605 ;
        RECT 75.895 182.450 76.055 182.560 ;
        RECT 76.805 182.395 76.975 182.585 ;
        RECT 77.260 182.445 77.380 182.555 ;
        RECT 77.725 182.415 77.895 182.585 ;
        RECT 80.950 182.395 81.120 182.585 ;
        RECT 81.405 182.415 81.575 182.605 ;
        RECT 82.325 182.395 82.495 182.605 ;
        RECT 87.845 182.415 88.015 182.605 ;
        RECT 89.040 182.395 89.210 182.585 ;
        RECT 92.905 182.395 93.075 182.585 ;
        RECT 94.745 182.415 94.915 182.605 ;
        RECT 95.205 182.555 95.375 182.605 ;
        RECT 95.200 182.445 95.375 182.555 ;
        RECT 95.205 182.415 95.375 182.445 ;
        RECT 95.940 182.395 96.110 182.585 ;
        RECT 99.805 182.395 99.975 182.585 ;
        RECT 102.840 182.415 103.010 182.605 ;
        RECT 103.485 182.395 103.655 182.585 ;
        RECT 106.715 182.450 106.875 182.560 ;
        RECT 107.165 182.395 107.335 182.585 ;
        RECT 108.085 182.415 108.255 182.605 ;
        RECT 108.820 182.395 108.990 182.585 ;
        RECT 115.445 182.415 115.615 182.605 ;
        RECT 115.905 182.395 116.075 182.585 ;
        RECT 116.640 182.395 116.810 182.585 ;
        RECT 118.480 182.415 118.650 182.605 ;
        RECT 120.965 182.395 121.135 182.585 ;
        RECT 122.345 182.415 122.515 182.605 ;
        RECT 126.025 182.415 126.195 182.605 ;
        RECT 127.405 182.415 127.575 182.605 ;
        RECT 131.085 182.415 131.255 182.605 ;
        RECT 131.545 182.395 131.715 182.585 ;
        RECT 132.005 182.415 132.175 182.585 ;
        RECT 132.920 182.445 133.040 182.555 ;
        RECT 136.605 182.415 136.775 182.605 ;
        RECT 137.065 182.415 137.235 182.605 ;
        RECT 132.010 182.395 132.175 182.415 ;
        RECT 141.205 182.395 141.375 182.585 ;
        RECT 141.665 182.395 141.835 182.585 ;
        RECT 142.585 182.415 142.755 182.605 ;
        RECT 145.340 182.445 145.460 182.555 ;
        RECT 146.725 182.395 146.895 182.605 ;
        RECT 62.370 182.365 63.315 182.395 ;
        RECT 57.820 181.485 59.190 181.715 ;
        RECT 60.565 181.685 63.315 182.365 ;
        RECT 62.370 181.485 63.315 181.685 ;
        RECT 63.325 181.485 66.535 182.395 ;
        RECT 66.690 181.715 68.525 182.395 ;
        RECT 67.595 181.485 68.525 181.715 ;
        RECT 68.855 181.525 69.285 182.310 ;
        RECT 69.305 181.485 71.120 182.395 ;
        RECT 71.145 181.715 73.435 182.395 ;
        RECT 72.515 181.485 73.435 181.715 ;
        RECT 73.540 181.715 77.005 182.395 ;
        RECT 77.990 181.715 80.415 182.395 ;
        RECT 73.540 181.485 74.460 181.715 ;
        RECT 80.805 181.485 82.155 182.395 ;
        RECT 82.185 181.585 87.695 182.395 ;
        RECT 88.625 181.715 92.525 182.395 ;
        RECT 88.625 181.485 89.555 181.715 ;
        RECT 92.765 181.585 94.595 182.395 ;
        RECT 94.615 181.525 95.045 182.310 ;
        RECT 95.525 181.715 99.425 182.395 ;
        RECT 99.775 181.715 103.240 182.395 ;
        RECT 103.455 181.715 106.920 182.395 ;
        RECT 95.525 181.485 96.455 181.715 ;
        RECT 102.320 181.485 103.240 181.715 ;
        RECT 106.000 181.485 106.920 181.715 ;
        RECT 107.025 181.585 108.395 182.395 ;
        RECT 108.405 181.715 112.305 182.395 ;
        RECT 112.640 181.715 116.105 182.395 ;
        RECT 116.225 181.715 120.125 182.395 ;
        RECT 108.405 181.485 109.335 181.715 ;
        RECT 112.640 181.485 113.560 181.715 ;
        RECT 116.225 181.485 117.155 181.715 ;
        RECT 120.375 181.525 120.805 182.310 ;
        RECT 120.825 181.715 128.135 182.395 ;
        RECT 124.340 181.495 125.250 181.715 ;
        RECT 126.785 181.485 128.135 181.715 ;
        RECT 128.280 181.715 131.745 182.395 ;
        RECT 132.010 181.715 133.845 182.395 ;
        RECT 128.280 181.485 129.200 181.715 ;
        RECT 132.915 181.485 133.845 181.715 ;
        RECT 134.205 181.715 141.515 182.395 ;
        RECT 134.205 181.485 135.555 181.715 ;
        RECT 137.090 181.495 138.000 181.715 ;
        RECT 141.525 181.585 145.195 182.395 ;
        RECT 145.665 181.585 147.035 182.395 ;
      LAYER nwell ;
        RECT 17.130 178.365 147.230 181.195 ;
      LAYER pwell ;
        RECT 17.325 177.165 18.695 177.975 ;
        RECT 18.705 177.165 22.375 177.975 ;
        RECT 22.385 177.845 23.305 178.075 ;
        RECT 25.735 177.845 26.665 178.075 ;
        RECT 22.385 177.165 24.675 177.845 ;
        RECT 24.830 177.165 26.665 177.845 ;
        RECT 26.995 177.165 28.345 178.075 ;
        RECT 28.365 177.165 29.715 178.075 ;
        RECT 30.215 177.250 30.645 178.035 ;
        RECT 30.665 177.165 34.335 177.975 ;
        RECT 35.000 177.165 38.475 178.075 ;
        RECT 38.505 177.165 39.855 178.075 ;
        RECT 39.865 177.875 40.795 178.075 ;
        RECT 42.130 177.875 43.075 178.075 ;
        RECT 39.865 177.395 43.075 177.875 ;
        RECT 40.005 177.195 43.075 177.395 ;
        RECT 17.465 176.955 17.635 177.165 ;
        RECT 18.845 176.975 19.015 177.165 ;
        RECT 19.765 176.955 19.935 177.145 ;
        RECT 24.365 176.975 24.535 177.165 ;
        RECT 24.830 177.145 24.995 177.165 ;
        RECT 24.825 176.975 24.995 177.145 ;
        RECT 27.125 176.955 27.295 177.165 ;
        RECT 29.430 176.975 29.600 177.165 ;
        RECT 29.880 177.005 30.000 177.115 ;
        RECT 30.805 176.975 30.975 177.165 ;
        RECT 31.265 176.955 31.435 177.145 ;
        RECT 31.725 176.955 31.895 177.145 ;
        RECT 33.105 176.955 33.275 177.145 ;
        RECT 34.480 177.005 34.600 177.115 ;
        RECT 36.780 177.005 36.900 177.115 ;
        RECT 37.245 176.975 37.415 177.145 ;
        RECT 38.160 176.975 38.330 177.165 ;
        RECT 38.620 176.975 38.790 177.165 ;
        RECT 40.005 176.975 40.175 177.195 ;
        RECT 42.130 177.165 43.075 177.195 ;
        RECT 43.320 177.165 48.135 177.845 ;
        RECT 48.145 177.165 53.655 177.975 ;
        RECT 53.665 177.165 55.495 177.975 ;
        RECT 55.975 177.250 56.405 178.035 ;
        RECT 56.885 177.165 58.715 178.075 ;
        RECT 58.725 177.165 61.130 178.075 ;
        RECT 61.485 177.165 65.145 178.075 ;
        RECT 65.165 177.165 70.675 177.975 ;
        RECT 70.685 177.165 72.055 177.975 ;
        RECT 72.065 177.165 73.835 178.075 ;
        RECT 73.945 177.845 75.295 178.075 ;
        RECT 76.830 177.845 77.740 178.065 ;
        RECT 73.945 177.165 81.255 177.845 ;
        RECT 81.735 177.250 82.165 178.035 ;
        RECT 82.185 177.165 84.015 177.975 ;
        RECT 88.000 177.845 88.910 178.065 ;
        RECT 90.445 177.845 91.795 178.075 ;
        RECT 84.485 177.165 91.795 177.845 ;
        RECT 92.805 177.845 94.155 178.075 ;
        RECT 95.690 177.845 96.600 178.065 ;
        RECT 100.125 177.845 101.055 178.075 ;
        RECT 92.805 177.165 100.115 177.845 ;
        RECT 100.125 177.165 104.025 177.845 ;
        RECT 104.265 177.165 107.015 177.975 ;
        RECT 107.495 177.250 107.925 178.035 ;
        RECT 107.945 177.165 111.155 178.075 ;
        RECT 111.165 177.165 116.675 177.975 ;
        RECT 116.725 177.845 118.075 178.075 ;
        RECT 119.610 177.845 120.520 178.065 ;
        RECT 116.725 177.165 124.035 177.845 ;
        RECT 124.045 177.165 127.255 178.075 ;
        RECT 127.265 177.875 128.220 178.075 ;
        RECT 127.265 177.195 129.545 177.875 ;
        RECT 127.265 177.165 128.220 177.195 ;
        RECT 37.255 176.955 37.415 176.975 ;
        RECT 41.390 176.955 41.560 177.145 ;
        RECT 42.760 177.005 42.880 177.115 ;
        RECT 43.685 176.955 43.855 177.145 ;
        RECT 46.905 176.955 47.075 177.145 ;
        RECT 47.825 176.975 47.995 177.165 ;
        RECT 48.285 176.975 48.455 177.165 ;
        RECT 52.425 176.955 52.595 177.145 ;
        RECT 53.805 176.975 53.975 177.165 ;
        RECT 55.640 177.005 55.760 177.115 ;
        RECT 56.560 177.005 56.680 177.115 ;
        RECT 57.030 176.975 57.200 177.165 ;
        RECT 57.945 176.955 58.115 177.145 ;
        RECT 58.865 176.975 59.035 177.165 ;
        RECT 60.700 177.005 60.820 177.115 ;
        RECT 61.170 176.955 61.340 177.145 ;
        RECT 62.540 177.005 62.660 177.115 ;
        RECT 62.995 176.955 63.165 177.145 ;
        RECT 64.850 176.975 65.020 177.165 ;
        RECT 65.305 176.975 65.475 177.165 ;
        RECT 66.225 176.955 66.395 177.145 ;
        RECT 69.445 176.955 69.615 177.145 ;
        RECT 70.825 176.975 70.995 177.165 ;
        RECT 72.210 176.975 72.380 177.165 ;
        RECT 73.125 176.955 73.295 177.145 ;
        RECT 74.505 176.955 74.675 177.145 ;
        RECT 78.190 176.955 78.360 177.145 ;
        RECT 79.565 176.955 79.735 177.145 ;
        RECT 80.945 176.975 81.115 177.165 ;
        RECT 81.400 177.005 81.520 177.115 ;
        RECT 82.325 176.975 82.495 177.165 ;
        RECT 84.160 177.005 84.280 177.115 ;
        RECT 84.625 176.975 84.795 177.165 ;
        RECT 85.085 176.955 85.255 177.145 ;
        RECT 86.920 177.005 87.040 177.115 ;
        RECT 87.385 176.955 87.555 177.145 ;
        RECT 91.995 177.010 92.155 177.120 ;
        RECT 98.425 176.955 98.595 177.145 ;
        RECT 99.805 176.975 99.975 177.165 ;
        RECT 100.540 176.975 100.710 177.165 ;
        RECT 102.105 176.955 102.275 177.145 ;
        RECT 104.405 176.975 104.575 177.165 ;
        RECT 105.785 176.955 105.955 177.145 ;
        RECT 106.245 176.975 106.415 177.145 ;
        RECT 107.160 177.005 107.280 177.115 ;
        RECT 110.845 176.975 111.015 177.165 ;
        RECT 111.305 176.975 111.475 177.165 ;
        RECT 112.225 176.955 112.395 177.145 ;
        RECT 112.685 176.955 112.855 177.145 ;
        RECT 118.205 176.955 118.375 177.145 ;
        RECT 120.040 177.005 120.160 177.115 ;
        RECT 120.965 176.955 121.135 177.145 ;
        RECT 123.725 177.115 123.895 177.165 ;
        RECT 123.720 177.005 123.895 177.115 ;
        RECT 123.725 176.975 123.895 177.005 ;
        RECT 126.025 176.975 126.195 177.145 ;
        RECT 126.025 176.955 126.190 176.975 ;
        RECT 126.485 176.955 126.655 177.145 ;
        RECT 126.945 176.975 127.115 177.165 ;
        RECT 129.250 176.975 129.420 177.195 ;
        RECT 129.565 177.165 133.235 178.075 ;
        RECT 133.255 177.250 133.685 178.035 ;
        RECT 137.220 177.845 138.130 178.065 ;
        RECT 139.665 177.845 141.015 178.075 ;
        RECT 133.705 177.165 141.015 177.845 ;
        RECT 141.065 177.165 144.275 178.075 ;
        RECT 144.285 177.165 145.655 177.975 ;
        RECT 145.665 177.165 147.035 177.975 ;
        RECT 129.700 176.955 129.870 177.145 ;
        RECT 130.175 177.000 130.335 177.110 ;
        RECT 131.080 176.955 131.250 177.145 ;
        RECT 132.920 176.975 133.090 177.165 ;
        RECT 133.845 176.975 134.015 177.165 ;
        RECT 135.220 176.955 135.390 177.145 ;
        RECT 137.065 176.955 137.235 177.145 ;
        RECT 137.525 176.955 137.695 177.145 ;
        RECT 143.965 176.975 144.135 177.165 ;
        RECT 144.425 176.975 144.595 177.165 ;
        RECT 144.895 177.000 145.055 177.110 ;
        RECT 146.725 176.955 146.895 177.165 ;
        RECT 17.325 176.145 18.695 176.955 ;
        RECT 19.625 176.275 26.935 176.955 ;
        RECT 26.985 176.275 29.275 176.955 ;
        RECT 23.140 176.055 24.050 176.275 ;
        RECT 25.585 176.045 26.935 176.275 ;
        RECT 28.355 176.045 29.275 176.275 ;
        RECT 29.285 176.275 31.575 176.955 ;
        RECT 29.285 176.045 30.205 176.275 ;
        RECT 31.595 176.045 32.945 176.955 ;
        RECT 32.965 176.145 36.635 176.955 ;
        RECT 37.255 176.045 40.910 176.955 ;
        RECT 41.245 176.045 42.595 176.955 ;
        RECT 43.095 176.085 43.525 176.870 ;
        RECT 43.625 176.045 46.625 176.955 ;
        RECT 46.765 176.145 52.275 176.955 ;
        RECT 52.285 176.145 57.795 176.955 ;
        RECT 57.805 176.145 60.555 176.955 ;
        RECT 61.025 176.045 62.375 176.955 ;
        RECT 62.865 176.045 66.075 176.955 ;
        RECT 66.085 176.145 68.835 176.955 ;
        RECT 68.855 176.085 69.285 176.870 ;
        RECT 69.305 176.145 72.975 176.955 ;
        RECT 72.985 176.145 74.355 176.955 ;
        RECT 74.475 176.275 77.940 176.955 ;
        RECT 77.020 176.045 77.940 176.275 ;
        RECT 78.045 176.045 79.395 176.955 ;
        RECT 79.425 176.145 84.935 176.955 ;
        RECT 84.945 176.145 86.775 176.955 ;
        RECT 87.245 176.275 94.555 176.955 ;
        RECT 90.760 176.055 91.670 176.275 ;
        RECT 93.205 176.045 94.555 176.275 ;
        RECT 94.615 176.085 95.045 176.870 ;
        RECT 95.160 176.275 98.625 176.955 ;
        RECT 98.840 176.275 102.305 176.955 ;
        RECT 102.520 176.275 105.985 176.955 ;
        RECT 106.510 176.275 108.935 176.955 ;
        RECT 109.325 176.275 112.535 176.955 ;
        RECT 95.160 176.045 96.080 176.275 ;
        RECT 98.840 176.045 99.760 176.275 ;
        RECT 102.520 176.045 103.440 176.275 ;
        RECT 109.325 176.045 110.460 176.275 ;
        RECT 112.545 176.145 118.055 176.955 ;
        RECT 118.065 176.145 119.895 176.955 ;
        RECT 120.375 176.085 120.805 176.870 ;
        RECT 120.825 176.145 123.575 176.955 ;
        RECT 124.355 176.275 126.190 176.955 ;
        RECT 126.345 176.275 128.635 176.955 ;
        RECT 124.355 176.045 125.285 176.275 ;
        RECT 127.715 176.045 128.635 176.275 ;
        RECT 128.665 176.045 130.015 176.955 ;
        RECT 130.965 176.045 132.315 176.955 ;
        RECT 132.615 176.045 135.535 176.955 ;
        RECT 135.545 176.275 137.375 176.955 ;
        RECT 137.385 176.275 144.695 176.955 ;
        RECT 140.900 176.055 141.810 176.275 ;
        RECT 143.345 176.045 144.695 176.275 ;
        RECT 145.665 176.145 147.035 176.955 ;
      LAYER nwell ;
        RECT 17.130 172.925 147.230 175.755 ;
      LAYER pwell ;
        RECT 17.325 171.725 18.695 172.535 ;
        RECT 18.705 171.725 21.455 172.535 ;
        RECT 21.965 172.405 23.315 172.635 ;
        RECT 24.850 172.405 25.760 172.625 ;
        RECT 21.965 171.725 29.275 172.405 ;
        RECT 30.215 171.810 30.645 172.595 ;
        RECT 30.665 171.725 36.175 172.535 ;
        RECT 36.185 171.725 37.555 172.535 ;
        RECT 37.695 171.725 40.695 172.635 ;
        RECT 40.785 172.405 41.705 172.635 ;
        RECT 40.785 171.725 44.370 172.405 ;
        RECT 44.485 171.725 45.835 172.635 ;
        RECT 46.345 172.405 47.695 172.635 ;
        RECT 49.230 172.405 50.140 172.625 ;
        RECT 46.345 171.725 53.655 172.405 ;
        RECT 53.665 171.725 55.495 172.535 ;
        RECT 55.975 171.810 56.405 172.595 ;
        RECT 56.425 171.725 61.935 172.535 ;
        RECT 61.945 171.725 63.775 172.535 ;
        RECT 64.245 172.405 65.165 172.635 ;
        RECT 64.245 171.725 66.535 172.405 ;
        RECT 66.545 171.725 68.360 172.635 ;
        RECT 68.385 171.725 69.735 172.635 ;
        RECT 71.825 172.545 72.775 172.635 ;
        RECT 70.845 171.725 72.775 172.545 ;
        RECT 73.025 172.405 74.375 172.635 ;
        RECT 75.910 172.405 76.820 172.625 ;
        RECT 73.025 171.725 80.335 172.405 ;
        RECT 80.345 171.725 81.715 172.535 ;
        RECT 81.735 171.810 82.165 172.595 ;
        RECT 82.185 171.725 85.855 172.535 ;
        RECT 89.840 172.405 90.750 172.625 ;
        RECT 92.285 172.405 93.635 172.635 ;
        RECT 86.325 171.725 93.635 172.405 ;
        RECT 93.685 172.405 94.615 172.635 ;
        RECT 93.685 171.725 97.585 172.405 ;
        RECT 97.825 171.725 100.575 172.535 ;
        RECT 100.585 172.405 101.515 172.635 ;
        RECT 100.585 171.725 104.485 172.405 ;
        RECT 105.665 171.725 107.015 172.635 ;
        RECT 107.495 171.810 107.925 172.595 ;
        RECT 111.460 172.405 112.370 172.625 ;
        RECT 113.905 172.405 115.255 172.635 ;
        RECT 107.945 171.725 115.255 172.405 ;
        RECT 115.305 171.725 120.815 172.535 ;
        RECT 120.825 171.725 122.655 172.535 ;
        RECT 123.145 171.725 124.495 172.635 ;
        RECT 124.505 171.725 130.015 172.535 ;
        RECT 130.505 171.725 131.855 172.635 ;
        RECT 131.885 171.725 133.235 172.635 ;
        RECT 133.255 171.810 133.685 172.595 ;
        RECT 133.705 171.725 135.055 172.635 ;
        RECT 136.005 171.725 139.215 172.635 ;
        RECT 139.235 171.725 140.585 172.635 ;
        RECT 140.605 171.725 141.955 172.635 ;
        RECT 141.985 171.725 145.655 172.535 ;
        RECT 145.665 171.725 147.035 172.535 ;
        RECT 17.465 171.515 17.635 171.725 ;
        RECT 18.845 171.515 19.015 171.725 ;
        RECT 21.600 171.565 21.720 171.675 ;
        RECT 24.365 171.515 24.535 171.705 ;
        RECT 28.965 171.535 29.135 171.725 ;
        RECT 29.435 171.570 29.595 171.680 ;
        RECT 29.885 171.515 30.055 171.705 ;
        RECT 30.805 171.535 30.975 171.725 ;
        RECT 33.565 171.515 33.735 171.705 ;
        RECT 36.325 171.535 36.495 171.725 ;
        RECT 38.160 171.515 38.330 171.705 ;
        RECT 38.625 171.535 38.795 171.705 ;
        RECT 40.465 171.535 40.635 171.725 ;
        RECT 40.930 171.705 41.100 171.725 ;
        RECT 40.925 171.535 41.100 171.705 ;
        RECT 42.760 171.565 42.880 171.675 ;
        RECT 38.630 171.515 38.795 171.535 ;
        RECT 40.925 171.515 41.095 171.535 ;
        RECT 43.690 171.515 43.860 171.705 ;
        RECT 44.600 171.535 44.770 171.725 ;
        RECT 45.980 171.565 46.100 171.675 ;
        RECT 47.365 171.515 47.535 171.705 ;
        RECT 50.585 171.535 50.755 171.705 ;
        RECT 50.605 171.515 50.755 171.535 ;
        RECT 52.885 171.515 53.055 171.705 ;
        RECT 53.345 171.535 53.515 171.725 ;
        RECT 53.805 171.535 53.975 171.725 ;
        RECT 56.565 171.675 56.735 171.725 ;
        RECT 55.640 171.565 55.760 171.675 ;
        RECT 56.560 171.565 56.735 171.675 ;
        RECT 56.565 171.535 56.735 171.565 ;
        RECT 58.400 171.515 58.570 171.705 ;
        RECT 61.625 171.515 61.795 171.705 ;
        RECT 62.085 171.515 62.255 171.725 ;
        RECT 63.920 171.565 64.040 171.675 ;
        RECT 66.225 171.535 66.395 171.725 ;
        RECT 68.065 171.535 68.235 171.725 ;
        RECT 68.530 171.705 68.700 171.725 ;
        RECT 70.845 171.705 70.995 171.725 ;
        RECT 68.525 171.535 68.700 171.705 ;
        RECT 69.915 171.570 70.075 171.680 ;
        RECT 70.825 171.535 70.995 171.705 ;
        RECT 68.525 171.515 68.695 171.535 ;
        RECT 72.665 171.515 72.835 171.705 ;
        RECT 74.500 171.515 74.670 171.705 ;
        RECT 74.965 171.515 75.135 171.705 ;
        RECT 77.725 171.515 77.895 171.705 ;
        RECT 80.025 171.535 80.195 171.725 ;
        RECT 80.485 171.535 80.655 171.725 ;
        RECT 82.325 171.535 82.495 171.725 ;
        RECT 85.085 171.515 85.255 171.705 ;
        RECT 86.000 171.565 86.120 171.675 ;
        RECT 86.465 171.535 86.635 171.725 ;
        RECT 90.605 171.515 90.775 171.705 ;
        RECT 94.100 171.535 94.270 171.725 ;
        RECT 94.280 171.565 94.400 171.675 ;
        RECT 95.480 171.515 95.650 171.705 ;
        RECT 97.965 171.535 98.135 171.725 ;
        RECT 99.345 171.515 99.515 171.705 ;
        RECT 101.000 171.535 101.170 171.725 ;
        RECT 101.185 171.515 101.355 171.705 ;
        RECT 104.875 171.570 105.035 171.680 ;
        RECT 106.245 171.515 106.415 171.705 ;
        RECT 106.700 171.535 106.870 171.725 ;
        RECT 107.160 171.565 107.280 171.675 ;
        RECT 108.085 171.515 108.255 171.725 ;
        RECT 115.445 171.535 115.615 171.725 ;
        RECT 116.365 171.535 116.535 171.705 ;
        RECT 120.040 171.565 120.160 171.675 ;
        RECT 116.365 171.515 116.565 171.535 ;
        RECT 120.965 171.515 121.135 171.725 ;
        RECT 122.800 171.565 122.920 171.675 ;
        RECT 123.260 171.535 123.430 171.725 ;
        RECT 124.645 171.535 124.815 171.725 ;
        RECT 126.485 171.515 126.655 171.705 ;
        RECT 128.330 171.515 128.500 171.705 ;
        RECT 129.705 171.515 129.875 171.705 ;
        RECT 130.160 171.565 130.280 171.675 ;
        RECT 131.540 171.535 131.710 171.725 ;
        RECT 132.920 171.535 133.090 171.725 ;
        RECT 133.850 171.535 134.020 171.725 ;
        RECT 135.235 171.570 135.395 171.680 ;
        RECT 135.690 171.515 135.860 171.705 ;
        RECT 136.145 171.535 136.315 171.725 ;
        RECT 137.985 171.535 138.155 171.705 ;
        RECT 137.985 171.515 138.135 171.535 ;
        RECT 138.450 171.515 138.620 171.705 ;
        RECT 139.825 171.515 139.995 171.705 ;
        RECT 140.285 171.535 140.455 171.725 ;
        RECT 141.670 171.535 141.840 171.725 ;
        RECT 142.125 171.535 142.295 171.725 ;
        RECT 145.340 171.565 145.460 171.675 ;
        RECT 146.725 171.515 146.895 171.725 ;
        RECT 17.325 170.705 18.695 171.515 ;
        RECT 18.705 170.705 24.215 171.515 ;
        RECT 24.225 170.705 29.735 171.515 ;
        RECT 29.745 170.705 33.415 171.515 ;
        RECT 33.425 170.705 34.795 171.515 ;
        RECT 34.805 170.835 38.475 171.515 ;
        RECT 38.630 170.835 40.465 171.515 ;
        RECT 37.550 170.605 38.475 170.835 ;
        RECT 39.535 170.605 40.465 170.835 ;
        RECT 40.785 170.705 42.615 171.515 ;
        RECT 43.095 170.645 43.525 171.430 ;
        RECT 43.545 170.835 47.130 171.515 ;
        RECT 43.545 170.605 44.465 170.835 ;
        RECT 47.265 170.605 50.435 171.515 ;
        RECT 50.605 170.695 52.535 171.515 ;
        RECT 52.745 170.705 56.415 171.515 ;
        RECT 51.585 170.605 52.535 170.695 ;
        RECT 56.945 170.605 58.715 171.515 ;
        RECT 58.725 170.605 61.835 171.515 ;
        RECT 62.045 170.605 65.155 171.515 ;
        RECT 65.260 170.835 68.725 171.515 ;
        RECT 65.260 170.605 66.180 170.835 ;
        RECT 68.855 170.645 69.285 171.430 ;
        RECT 69.400 170.835 72.865 171.515 ;
        RECT 69.400 170.605 70.320 170.835 ;
        RECT 73.045 170.605 74.815 171.515 ;
        RECT 74.825 170.705 77.575 171.515 ;
        RECT 77.585 170.835 84.895 171.515 ;
        RECT 81.100 170.615 82.010 170.835 ;
        RECT 83.545 170.605 84.895 170.835 ;
        RECT 84.945 170.705 90.455 171.515 ;
        RECT 90.465 170.705 94.135 171.515 ;
        RECT 94.615 170.645 95.045 171.430 ;
        RECT 95.065 170.835 98.965 171.515 ;
        RECT 95.065 170.605 95.995 170.835 ;
        RECT 99.205 170.705 101.035 171.515 ;
        RECT 101.045 170.835 105.860 171.515 ;
        RECT 106.105 170.705 107.935 171.515 ;
        RECT 107.945 170.835 115.255 171.515 ;
        RECT 116.365 170.835 119.895 171.515 ;
        RECT 111.460 170.615 112.370 170.835 ;
        RECT 113.905 170.605 115.255 170.835 ;
        RECT 117.070 170.605 119.895 170.835 ;
        RECT 120.375 170.645 120.805 171.430 ;
        RECT 120.825 170.705 126.335 171.515 ;
        RECT 126.360 170.605 128.175 171.515 ;
        RECT 128.185 170.605 129.535 171.515 ;
        RECT 129.565 170.705 132.315 171.515 ;
        RECT 132.325 170.605 135.985 171.515 ;
        RECT 136.205 170.695 138.135 171.515 ;
        RECT 136.205 170.605 137.155 170.695 ;
        RECT 138.305 170.605 139.655 171.515 ;
        RECT 139.685 170.705 145.195 171.515 ;
        RECT 145.665 170.705 147.035 171.515 ;
      LAYER nwell ;
        RECT 17.130 167.485 147.230 170.315 ;
      LAYER pwell ;
        RECT 17.325 166.285 18.695 167.095 ;
        RECT 18.705 166.285 22.375 167.095 ;
        RECT 22.385 166.285 23.755 167.095 ;
        RECT 23.775 166.285 25.125 167.195 ;
        RECT 25.805 167.105 26.755 167.195 ;
        RECT 25.805 166.285 27.735 167.105 ;
        RECT 27.905 166.285 29.735 167.095 ;
        RECT 30.215 166.370 30.645 167.155 ;
        RECT 30.665 166.285 33.875 167.195 ;
        RECT 33.885 166.285 36.175 167.195 ;
        RECT 36.185 166.285 37.535 167.195 ;
        RECT 37.565 166.285 43.075 167.095 ;
        RECT 45.350 166.995 46.295 167.195 ;
        RECT 43.545 166.315 46.295 166.995 ;
        RECT 47.675 166.965 48.595 167.195 ;
        RECT 17.465 166.075 17.635 166.285 ;
        RECT 18.845 166.075 19.015 166.285 ;
        RECT 22.525 166.095 22.695 166.285 ;
        RECT 22.525 166.075 22.690 166.095 ;
        RECT 24.825 166.075 24.995 166.285 ;
        RECT 27.585 166.265 27.735 166.285 ;
        RECT 25.280 166.125 25.400 166.235 ;
        RECT 27.125 166.095 27.295 166.265 ;
        RECT 27.585 166.235 27.755 166.265 ;
        RECT 27.580 166.125 27.755 166.235 ;
        RECT 27.585 166.095 27.755 166.125 ;
        RECT 28.045 166.095 28.215 166.285 ;
        RECT 30.805 166.265 30.975 166.285 ;
        RECT 29.880 166.125 30.000 166.235 ;
        RECT 30.800 166.095 30.975 166.265 ;
        RECT 27.125 166.075 27.290 166.095 ;
        RECT 30.800 166.075 30.970 166.095 ;
        RECT 32.185 166.075 32.355 166.265 ;
        RECT 32.645 166.075 32.815 166.265 ;
        RECT 35.865 166.095 36.035 166.285 ;
        RECT 36.320 166.125 36.440 166.235 ;
        RECT 37.250 166.095 37.420 166.285 ;
        RECT 37.705 166.095 37.875 166.285 ;
        RECT 38.625 166.095 38.795 166.265 ;
        RECT 38.625 166.075 38.790 166.095 ;
        RECT 40.005 166.075 40.175 166.265 ;
        RECT 40.465 166.075 40.635 166.265 ;
        RECT 42.760 166.075 42.930 166.265 ;
        RECT 43.220 166.125 43.340 166.235 ;
        RECT 43.690 166.095 43.860 166.315 ;
        RECT 45.350 166.285 46.295 166.315 ;
        RECT 46.305 166.285 48.595 166.965 ;
        RECT 48.615 166.285 49.965 167.195 ;
        RECT 49.985 166.285 52.735 167.095 ;
        RECT 53.215 166.285 54.565 167.195 ;
        RECT 54.585 166.285 55.955 167.095 ;
        RECT 55.975 166.370 56.405 167.155 ;
        RECT 56.905 166.285 58.255 167.195 ;
        RECT 61.780 166.965 62.690 167.185 ;
        RECT 64.225 166.965 65.575 167.195 ;
        RECT 58.265 166.285 65.575 166.965 ;
        RECT 65.665 166.965 67.015 167.195 ;
        RECT 68.550 166.965 69.460 167.185 ;
        RECT 65.665 166.285 72.975 166.965 ;
        RECT 72.985 166.285 78.495 167.095 ;
        RECT 78.505 166.285 81.255 167.095 ;
        RECT 81.735 166.370 82.165 167.155 ;
        RECT 82.185 166.285 84.015 167.095 ;
        RECT 87.140 166.965 88.060 167.195 ;
        RECT 84.595 166.285 88.060 166.965 ;
        RECT 88.165 166.285 91.835 167.095 ;
        RECT 91.845 166.285 93.215 167.095 ;
        RECT 96.740 166.965 97.650 167.185 ;
        RECT 99.185 166.965 100.535 167.195 ;
        RECT 93.225 166.285 100.535 166.965 ;
        RECT 100.585 166.965 101.515 167.195 ;
        RECT 100.585 166.285 104.485 166.965 ;
        RECT 105.645 166.285 107.460 167.195 ;
        RECT 107.495 166.370 107.925 167.155 ;
        RECT 107.955 166.285 109.305 167.195 ;
        RECT 109.325 166.965 113.255 167.195 ;
        RECT 113.925 166.995 114.875 167.195 ;
        RECT 118.745 167.105 119.695 167.195 ;
        RECT 109.325 166.285 113.740 166.965 ;
        RECT 113.925 166.315 117.595 166.995 ;
        RECT 113.925 166.285 114.875 166.315 ;
        RECT 46.445 166.075 46.615 166.285 ;
        RECT 47.830 166.075 48.000 166.265 ;
        RECT 48.280 166.125 48.400 166.235 ;
        RECT 48.745 166.095 48.915 166.285 ;
        RECT 50.125 166.095 50.295 166.285 ;
        RECT 52.880 166.125 53.000 166.235 ;
        RECT 53.345 166.095 53.515 166.285 ;
        RECT 54.725 166.095 54.895 166.285 ;
        RECT 55.645 166.075 55.815 166.265 ;
        RECT 56.105 166.075 56.275 166.265 ;
        RECT 56.560 166.125 56.680 166.235 ;
        RECT 57.940 166.095 58.110 166.285 ;
        RECT 58.405 166.095 58.575 166.285 ;
        RECT 61.625 166.075 61.795 166.265 ;
        RECT 69.445 166.075 69.615 166.265 ;
        RECT 72.665 166.095 72.835 166.285 ;
        RECT 73.125 166.095 73.295 166.285 ;
        RECT 74.965 166.075 75.135 166.265 ;
        RECT 78.645 166.095 78.815 166.285 ;
        RECT 81.400 166.125 81.520 166.235 ;
        RECT 82.325 166.095 82.495 166.285 ;
        RECT 83.705 166.075 83.875 166.265 ;
        RECT 84.170 166.235 84.340 166.265 ;
        RECT 84.160 166.125 84.340 166.235 ;
        RECT 84.170 166.075 84.340 166.125 ;
        RECT 84.625 166.095 84.795 166.285 ;
        RECT 87.850 166.075 88.020 166.265 ;
        RECT 88.305 166.095 88.475 166.285 ;
        RECT 91.065 166.075 91.235 166.265 ;
        RECT 91.985 166.095 92.155 166.285 ;
        RECT 93.365 166.095 93.535 166.285 ;
        RECT 95.205 166.075 95.375 166.265 ;
        RECT 98.880 166.075 99.050 166.265 ;
        RECT 101.000 166.095 101.170 166.285 ;
        RECT 104.875 166.130 105.035 166.240 ;
        RECT 107.165 166.075 107.335 166.285 ;
        RECT 108.085 166.095 108.255 166.285 ;
        RECT 113.630 166.265 113.740 166.285 ;
        RECT 110.845 166.075 111.015 166.265 ;
        RECT 111.305 166.095 111.475 166.265 ;
        RECT 113.630 166.095 113.800 166.265 ;
        RECT 111.305 166.075 111.505 166.095 ;
        RECT 17.325 165.265 18.695 166.075 ;
        RECT 18.705 165.265 20.535 166.075 ;
        RECT 20.855 165.395 22.690 166.075 ;
        RECT 22.845 165.395 25.135 166.075 ;
        RECT 25.455 165.395 27.290 166.075 ;
        RECT 20.855 165.165 21.785 165.395 ;
        RECT 22.845 165.165 23.765 165.395 ;
        RECT 25.455 165.165 26.385 165.395 ;
        RECT 28.195 165.165 31.115 166.075 ;
        RECT 31.135 165.165 32.485 166.075 ;
        RECT 32.505 165.265 36.175 166.075 ;
        RECT 36.955 165.395 38.790 166.075 ;
        RECT 36.955 165.165 37.885 165.395 ;
        RECT 38.955 165.165 40.305 166.075 ;
        RECT 40.325 165.265 41.695 166.075 ;
        RECT 41.725 165.165 43.075 166.075 ;
        RECT 43.095 165.205 43.525 165.990 ;
        RECT 43.545 165.165 46.755 166.075 ;
        RECT 46.765 165.165 48.115 166.075 ;
        RECT 48.645 165.395 55.955 166.075 ;
        RECT 48.645 165.165 49.995 165.395 ;
        RECT 51.530 165.175 52.440 165.395 ;
        RECT 55.965 165.265 61.475 166.075 ;
        RECT 61.485 165.395 68.795 166.075 ;
        RECT 65.000 165.175 65.910 165.395 ;
        RECT 67.445 165.165 68.795 165.395 ;
        RECT 68.855 165.205 69.285 165.990 ;
        RECT 69.305 165.265 74.815 166.075 ;
        RECT 74.825 165.265 76.655 166.075 ;
        RECT 76.705 165.395 84.015 166.075 ;
        RECT 84.025 165.395 87.610 166.075 ;
        RECT 76.705 165.165 78.055 165.395 ;
        RECT 79.590 165.175 80.500 165.395 ;
        RECT 84.025 165.165 84.945 165.395 ;
        RECT 87.705 165.165 90.820 166.075 ;
        RECT 90.925 165.265 94.595 166.075 ;
        RECT 94.615 165.205 95.045 165.990 ;
        RECT 95.065 165.265 98.735 166.075 ;
        RECT 98.765 165.165 100.115 166.075 ;
        RECT 100.165 165.395 107.475 166.075 ;
        RECT 107.580 165.395 111.045 166.075 ;
        RECT 111.305 165.395 114.835 166.075 ;
        RECT 114.990 166.045 115.160 166.265 ;
        RECT 117.280 166.095 117.450 166.315 ;
        RECT 117.765 166.285 119.695 167.105 ;
        RECT 119.925 166.285 121.275 167.195 ;
        RECT 121.285 166.285 122.655 167.095 ;
        RECT 122.665 166.995 123.610 167.195 ;
        RECT 124.945 166.995 125.875 167.195 ;
        RECT 122.665 166.515 125.875 166.995 ;
        RECT 127.705 166.965 128.635 167.195 ;
        RECT 122.665 166.315 125.735 166.515 ;
        RECT 122.665 166.285 123.610 166.315 ;
        RECT 117.765 166.265 117.915 166.285 ;
        RECT 117.745 166.095 117.915 166.265 ;
        RECT 118.665 166.075 118.835 166.265 ;
        RECT 120.040 166.095 120.210 166.285 ;
        RECT 121.425 166.095 121.595 166.285 ;
        RECT 122.805 166.075 122.975 166.265 ;
        RECT 123.265 166.075 123.435 166.265 ;
        RECT 125.565 166.095 125.735 166.315 ;
        RECT 125.885 166.285 128.635 166.965 ;
        RECT 128.645 166.285 130.460 167.195 ;
        RECT 130.505 166.285 131.855 167.195 ;
        RECT 131.865 166.285 133.235 167.095 ;
        RECT 133.255 166.370 133.685 167.155 ;
        RECT 135.040 166.995 135.995 167.195 ;
        RECT 133.715 166.315 135.995 166.995 ;
        RECT 126.025 166.095 126.195 166.285 ;
        RECT 128.335 166.120 128.495 166.230 ;
        RECT 129.245 166.095 129.415 166.265 ;
        RECT 130.165 166.095 130.335 166.285 ;
        RECT 131.540 166.095 131.710 166.285 ;
        RECT 132.005 166.095 132.175 166.285 ;
        RECT 133.380 166.125 133.500 166.235 ;
        RECT 133.840 166.095 134.010 166.315 ;
        RECT 135.040 166.285 135.995 166.315 ;
        RECT 136.005 166.285 137.355 167.195 ;
        RECT 137.385 166.285 142.895 167.095 ;
        RECT 143.825 166.965 145.170 167.195 ;
        RECT 143.825 166.285 145.655 166.965 ;
        RECT 145.665 166.285 147.035 167.095 ;
        RECT 135.685 166.095 135.855 166.265 ;
        RECT 136.140 166.125 136.260 166.235 ;
        RECT 129.255 166.075 129.415 166.095 ;
        RECT 135.685 166.075 135.850 166.095 ;
        RECT 136.605 166.075 136.775 166.265 ;
        RECT 137.070 166.095 137.240 166.285 ;
        RECT 137.525 166.095 137.695 166.285 ;
        RECT 143.055 166.130 143.215 166.240 ;
        RECT 143.965 166.075 144.135 166.265 ;
        RECT 145.345 166.095 145.515 166.285 ;
        RECT 146.725 166.075 146.895 166.285 ;
        RECT 117.565 166.045 118.515 166.075 ;
        RECT 100.165 165.165 101.515 165.395 ;
        RECT 103.050 165.175 103.960 165.395 ;
        RECT 107.580 165.165 108.500 165.395 ;
        RECT 112.010 165.165 114.835 165.395 ;
        RECT 114.845 165.365 118.515 166.045 ;
        RECT 117.565 165.165 118.515 165.365 ;
        RECT 118.525 165.265 120.355 166.075 ;
        RECT 120.375 165.205 120.805 165.990 ;
        RECT 120.825 165.395 123.115 166.075 ;
        RECT 123.125 165.395 127.940 166.075 ;
        RECT 120.825 165.165 121.745 165.395 ;
        RECT 129.255 165.165 132.910 166.075 ;
        RECT 134.015 165.395 135.850 166.075 ;
        RECT 136.465 165.395 143.775 166.075 ;
        RECT 143.825 165.395 145.655 166.075 ;
        RECT 134.015 165.165 134.945 165.395 ;
        RECT 139.980 165.175 140.890 165.395 ;
        RECT 142.425 165.165 143.775 165.395 ;
        RECT 144.310 165.165 145.655 165.395 ;
        RECT 145.665 165.265 147.035 166.075 ;
      LAYER nwell ;
        RECT 17.130 162.045 147.230 164.875 ;
      LAYER pwell ;
        RECT 17.325 160.845 18.695 161.655 ;
        RECT 22.680 161.525 23.590 161.745 ;
        RECT 25.125 161.525 26.475 161.755 ;
        RECT 19.165 160.845 26.475 161.525 ;
        RECT 26.525 160.845 27.875 161.755 ;
        RECT 29.275 161.525 30.195 161.755 ;
        RECT 27.905 160.845 30.195 161.525 ;
        RECT 30.215 160.930 30.645 161.715 ;
        RECT 34.180 161.525 35.090 161.745 ;
        RECT 36.625 161.525 37.975 161.755 ;
        RECT 39.165 161.665 40.115 161.755 ;
        RECT 30.665 160.845 37.975 161.525 ;
        RECT 38.185 160.845 40.115 161.665 ;
        RECT 43.215 161.525 44.145 161.755 ;
        RECT 45.835 161.525 46.755 161.755 ;
        RECT 40.325 160.845 42.155 161.525 ;
        RECT 42.310 160.845 44.145 161.525 ;
        RECT 44.465 160.845 46.755 161.525 ;
        RECT 46.865 160.845 49.975 161.755 ;
        RECT 51.125 161.665 52.075 161.755 ;
        RECT 50.145 160.845 52.075 161.665 ;
        RECT 52.285 160.845 55.955 161.655 ;
        RECT 55.975 160.930 56.405 161.715 ;
        RECT 56.425 160.845 61.935 161.655 ;
        RECT 61.945 160.845 67.455 161.655 ;
        RECT 67.465 160.845 72.975 161.655 ;
        RECT 72.985 160.845 78.495 161.655 ;
        RECT 78.505 160.845 81.255 161.655 ;
        RECT 81.735 160.930 82.165 161.715 ;
        RECT 82.645 161.075 85.395 161.755 ;
        RECT 85.405 161.555 86.335 161.755 ;
        RECT 87.665 161.555 88.615 161.755 ;
        RECT 85.405 161.075 88.615 161.555 ;
        RECT 82.785 160.845 85.395 161.075 ;
        RECT 85.550 160.875 88.615 161.075 ;
        RECT 17.465 160.635 17.635 160.845 ;
        RECT 18.845 160.795 19.015 160.825 ;
        RECT 18.840 160.685 19.015 160.795 ;
        RECT 18.845 160.635 19.015 160.685 ;
        RECT 19.305 160.655 19.475 160.845 ;
        RECT 22.065 160.635 22.235 160.825 ;
        RECT 22.525 160.635 22.695 160.825 ;
        RECT 27.590 160.655 27.760 160.845 ;
        RECT 28.045 160.655 28.215 160.845 ;
        RECT 29.885 160.635 30.055 160.825 ;
        RECT 30.805 160.655 30.975 160.845 ;
        RECT 38.185 160.825 38.335 160.845 ;
        RECT 32.185 160.635 32.355 160.825 ;
        RECT 34.940 160.685 35.060 160.795 ;
        RECT 35.405 160.635 35.575 160.825 ;
        RECT 38.165 160.655 38.335 160.825 ;
        RECT 41.845 160.655 42.015 160.845 ;
        RECT 42.310 160.825 42.475 160.845 ;
        RECT 42.305 160.655 42.475 160.825 ;
        RECT 42.760 160.685 42.880 160.795 ;
        RECT 43.685 160.635 43.855 160.825 ;
        RECT 44.605 160.655 44.775 160.845 ;
        RECT 46.905 160.655 47.075 160.845 ;
        RECT 50.145 160.825 50.295 160.845 ;
        RECT 50.125 160.655 50.295 160.825 ;
        RECT 51.965 160.635 52.135 160.825 ;
        RECT 52.425 160.635 52.595 160.845 ;
        RECT 56.565 160.655 56.735 160.845 ;
        RECT 57.945 160.635 58.115 160.825 ;
        RECT 61.620 160.685 61.740 160.795 ;
        RECT 62.085 160.655 62.255 160.845 ;
        RECT 63.005 160.635 63.175 160.825 ;
        RECT 63.475 160.680 63.635 160.790 ;
        RECT 67.605 160.635 67.775 160.845 ;
        RECT 68.075 160.680 68.235 160.790 ;
        RECT 69.445 160.635 69.615 160.825 ;
        RECT 73.125 160.655 73.295 160.845 ;
        RECT 74.965 160.635 75.135 160.825 ;
        RECT 78.645 160.655 78.815 160.845 ;
        RECT 79.565 160.635 79.735 160.825 ;
        RECT 81.400 160.685 81.520 160.795 ;
        RECT 82.320 160.685 82.440 160.795 ;
        RECT 82.785 160.655 82.955 160.845 ;
        RECT 83.245 160.635 83.415 160.825 ;
        RECT 85.550 160.655 85.720 160.875 ;
        RECT 87.680 160.845 88.615 160.875 ;
        RECT 88.625 160.845 89.975 161.755 ;
        RECT 93.980 161.525 94.890 161.745 ;
        RECT 96.425 161.525 97.775 161.755 ;
        RECT 102.980 161.525 103.900 161.755 ;
        RECT 90.465 160.845 97.775 161.525 ;
        RECT 98.060 160.845 102.875 161.525 ;
        RECT 102.980 160.845 106.445 161.525 ;
        RECT 107.495 160.930 107.925 161.715 ;
        RECT 107.995 160.845 111.155 161.755 ;
        RECT 111.165 161.555 112.095 161.755 ;
        RECT 113.425 161.555 114.375 161.755 ;
        RECT 111.165 161.075 114.375 161.555 ;
        RECT 111.310 160.875 114.375 161.075 ;
        RECT 89.690 160.825 89.860 160.845 ;
        RECT 89.685 160.655 89.860 160.825 ;
        RECT 90.605 160.825 90.775 160.845 ;
        RECT 90.140 160.685 90.260 160.795 ;
        RECT 90.605 160.655 90.780 160.825 ;
        RECT 95.205 160.655 95.375 160.825 ;
        RECT 97.500 160.685 97.620 160.795 ;
        RECT 89.685 160.635 89.855 160.655 ;
        RECT 90.610 160.635 90.780 160.655 ;
        RECT 95.210 160.635 95.375 160.655 ;
        RECT 101.645 160.635 101.815 160.825 ;
        RECT 102.565 160.655 102.735 160.845 ;
        RECT 105.325 160.635 105.495 160.825 ;
        RECT 106.245 160.655 106.415 160.845 ;
        RECT 106.715 160.690 106.875 160.800 ;
        RECT 108.085 160.655 108.255 160.845 ;
        RECT 108.545 160.635 108.715 160.825 ;
        RECT 109.015 160.680 109.175 160.790 ;
        RECT 111.310 160.655 111.480 160.875 ;
        RECT 113.440 160.845 114.375 160.875 ;
        RECT 114.465 160.845 116.675 161.755 ;
        RECT 117.615 160.845 120.345 161.755 ;
        RECT 120.835 160.845 123.565 161.755 ;
        RECT 124.245 160.845 126.335 161.655 ;
        RECT 126.495 160.845 130.150 161.755 ;
        RECT 130.795 161.525 131.725 161.755 ;
        RECT 130.795 160.845 132.630 161.525 ;
        RECT 133.255 160.930 133.685 161.715 ;
        RECT 135.040 161.555 135.995 161.755 ;
        RECT 133.715 160.875 135.995 161.555 ;
        RECT 115.440 160.635 115.610 160.825 ;
        RECT 115.905 160.635 116.075 160.825 ;
        RECT 116.360 160.655 116.530 160.845 ;
        RECT 116.835 160.690 116.995 160.800 ;
        RECT 117.745 160.655 117.915 160.845 ;
        RECT 120.965 160.825 121.135 160.845 ;
        RECT 118.210 160.635 118.380 160.825 ;
        RECT 118.660 160.685 118.780 160.795 ;
        RECT 119.120 160.635 119.290 160.825 ;
        RECT 120.500 160.685 120.620 160.795 ;
        RECT 120.960 160.655 121.135 160.825 ;
        RECT 17.325 159.825 18.695 160.635 ;
        RECT 18.705 159.825 20.075 160.635 ;
        RECT 20.085 159.955 22.375 160.635 ;
        RECT 22.385 159.955 29.695 160.635 ;
        RECT 29.745 159.955 32.035 160.635 ;
        RECT 20.085 159.725 21.005 159.955 ;
        RECT 25.900 159.735 26.810 159.955 ;
        RECT 28.345 159.725 29.695 159.955 ;
        RECT 31.115 159.725 32.035 159.955 ;
        RECT 32.045 159.825 34.795 160.635 ;
        RECT 35.265 159.955 42.575 160.635 ;
        RECT 38.780 159.735 39.690 159.955 ;
        RECT 41.225 159.725 42.575 159.955 ;
        RECT 43.095 159.765 43.525 160.550 ;
        RECT 43.545 159.825 44.915 160.635 ;
        RECT 44.965 159.955 52.275 160.635 ;
        RECT 44.965 159.725 46.315 159.955 ;
        RECT 47.850 159.735 48.760 159.955 ;
        RECT 52.285 159.825 57.795 160.635 ;
        RECT 57.805 159.825 61.475 160.635 ;
        RECT 61.955 159.725 63.305 160.635 ;
        RECT 64.340 159.955 67.805 160.635 ;
        RECT 64.340 159.725 65.260 159.955 ;
        RECT 68.855 159.765 69.285 160.550 ;
        RECT 69.305 159.825 74.815 160.635 ;
        RECT 74.825 159.825 78.495 160.635 ;
        RECT 79.535 159.955 83.000 160.635 ;
        RECT 82.080 159.725 83.000 159.955 ;
        RECT 83.105 159.825 86.775 160.635 ;
        RECT 88.155 160.605 89.995 160.635 ;
        RECT 86.830 159.955 89.995 160.605 ;
        RECT 86.830 159.925 89.510 159.955 ;
        RECT 88.155 159.725 89.510 159.925 ;
        RECT 90.465 159.725 94.355 160.635 ;
        RECT 94.615 159.765 95.045 160.550 ;
        RECT 95.210 159.955 97.045 160.635 ;
        RECT 96.115 159.725 97.045 159.955 ;
        RECT 97.825 159.725 101.955 160.635 ;
        RECT 102.060 159.955 105.525 160.635 ;
        RECT 102.060 159.725 102.980 159.955 ;
        RECT 105.645 159.725 108.855 160.635 ;
        RECT 110.045 159.725 115.755 160.635 ;
        RECT 115.775 159.725 117.125 160.635 ;
        RECT 117.145 159.725 118.495 160.635 ;
        RECT 119.005 159.725 120.355 160.635 ;
        RECT 120.960 160.605 121.130 160.655 ;
        RECT 123.265 160.635 123.435 160.825 ;
        RECT 126.025 160.655 126.195 160.845 ;
        RECT 126.495 160.825 126.655 160.845 ;
        RECT 132.465 160.825 132.630 160.845 ;
        RECT 126.485 160.655 126.655 160.825 ;
        RECT 131.540 160.635 131.710 160.825 ;
        RECT 132.005 160.635 132.175 160.825 ;
        RECT 132.465 160.655 132.635 160.825 ;
        RECT 132.920 160.685 133.040 160.795 ;
        RECT 133.840 160.655 134.010 160.875 ;
        RECT 135.040 160.845 135.995 160.875 ;
        RECT 136.005 160.845 137.375 161.655 ;
        RECT 137.385 161.525 138.315 161.755 ;
        RECT 141.620 161.525 142.540 161.755 ;
        RECT 137.385 160.845 141.285 161.525 ;
        RECT 141.620 160.845 145.085 161.525 ;
        RECT 145.665 160.845 147.035 161.655 ;
        RECT 135.220 160.685 135.340 160.795 ;
        RECT 135.685 160.635 135.855 160.825 ;
        RECT 136.145 160.655 136.315 160.845 ;
        RECT 137.800 160.655 137.970 160.845 ;
        RECT 143.055 160.680 143.215 160.790 ;
        RECT 143.965 160.635 144.135 160.825 ;
        RECT 144.885 160.655 145.055 160.845 ;
        RECT 145.340 160.685 145.460 160.795 ;
        RECT 146.725 160.635 146.895 160.845 ;
        RECT 122.160 160.605 123.115 160.635 ;
        RECT 120.375 159.765 120.805 160.550 ;
        RECT 120.835 159.925 123.115 160.605 ;
        RECT 123.125 159.955 127.940 160.635 ;
        RECT 122.160 159.725 123.115 159.925 ;
        RECT 128.380 159.725 131.855 160.635 ;
        RECT 131.865 159.725 135.075 160.635 ;
        RECT 135.545 159.955 142.855 160.635 ;
        RECT 143.825 159.955 145.655 160.635 ;
        RECT 139.060 159.735 139.970 159.955 ;
        RECT 141.505 159.725 142.855 159.955 ;
        RECT 144.310 159.725 145.655 159.955 ;
        RECT 145.665 159.825 147.035 160.635 ;
      LAYER nwell ;
        RECT 17.130 156.605 147.230 159.435 ;
      LAYER pwell ;
        RECT 17.325 155.405 18.695 156.215 ;
        RECT 18.705 155.405 24.215 156.215 ;
        RECT 24.225 155.405 29.735 156.215 ;
        RECT 30.215 155.490 30.645 156.275 ;
        RECT 30.665 155.405 36.175 156.215 ;
        RECT 36.645 156.085 37.565 156.315 ;
        RECT 36.645 155.405 38.935 156.085 ;
        RECT 38.945 155.405 44.455 156.215 ;
        RECT 44.465 155.405 49.975 156.215 ;
        RECT 49.985 155.405 55.495 156.215 ;
        RECT 55.975 155.490 56.405 156.275 ;
        RECT 56.425 155.405 58.255 156.215 ;
        RECT 61.380 156.085 62.300 156.315 ;
        RECT 58.835 155.405 62.300 156.085 ;
        RECT 62.415 155.405 65.145 156.315 ;
        RECT 66.395 156.085 67.325 156.315 ;
        RECT 66.395 155.405 68.230 156.085 ;
        RECT 68.385 155.405 70.215 156.085 ;
        RECT 70.225 155.405 71.575 156.315 ;
        RECT 75.120 156.085 76.030 156.305 ;
        RECT 77.565 156.085 78.915 156.315 ;
        RECT 71.605 155.405 78.915 156.085 ;
        RECT 78.965 156.085 79.885 156.315 ;
        RECT 78.965 155.405 81.255 156.085 ;
        RECT 81.735 155.490 82.165 156.275 ;
        RECT 82.185 155.405 87.695 156.215 ;
        RECT 87.705 155.405 93.215 156.215 ;
        RECT 93.225 155.405 96.895 156.215 ;
        RECT 97.365 155.405 98.715 156.315 ;
        RECT 98.745 155.405 104.255 156.215 ;
        RECT 104.265 155.405 107.015 156.215 ;
        RECT 107.495 155.490 107.925 156.275 ;
        RECT 107.945 155.405 111.615 156.215 ;
        RECT 114.740 156.085 115.660 156.315 ;
        RECT 112.195 155.405 115.660 156.085 ;
        RECT 115.765 155.405 119.265 156.315 ;
        RECT 119.445 155.405 121.275 156.215 ;
        RECT 121.765 155.405 123.115 156.315 ;
        RECT 127.855 156.085 128.785 156.315 ;
        RECT 123.530 155.405 125.955 156.085 ;
        RECT 126.950 155.405 128.785 156.085 ;
        RECT 129.105 155.405 131.855 156.315 ;
        RECT 131.865 155.405 133.235 156.215 ;
        RECT 133.255 155.490 133.685 156.275 ;
        RECT 133.705 155.405 135.535 156.315 ;
        RECT 135.545 155.405 136.915 156.185 ;
        RECT 136.925 156.085 137.855 156.315 ;
        RECT 141.160 156.085 142.080 156.315 ;
        RECT 136.925 155.405 140.825 156.085 ;
        RECT 141.160 155.405 144.625 156.085 ;
        RECT 145.665 155.405 147.035 156.215 ;
        RECT 17.465 155.195 17.635 155.405 ;
        RECT 18.845 155.195 19.015 155.405 ;
        RECT 20.685 155.195 20.855 155.385 ;
        RECT 24.365 155.215 24.535 155.405 ;
        RECT 26.205 155.195 26.375 155.385 ;
        RECT 29.880 155.245 30.000 155.355 ;
        RECT 30.805 155.215 30.975 155.405 ;
        RECT 31.725 155.195 31.895 155.385 ;
        RECT 36.320 155.245 36.440 155.355 ;
        RECT 37.245 155.195 37.415 155.385 ;
        RECT 38.625 155.215 38.795 155.405 ;
        RECT 39.085 155.215 39.255 155.405 ;
        RECT 42.760 155.245 42.880 155.355 ;
        RECT 43.685 155.195 43.855 155.385 ;
        RECT 44.605 155.215 44.775 155.405 ;
        RECT 49.205 155.195 49.375 155.385 ;
        RECT 50.125 155.215 50.295 155.405 ;
        RECT 54.725 155.195 54.895 155.385 ;
        RECT 55.640 155.245 55.760 155.355 ;
        RECT 56.105 155.215 56.275 155.385 ;
        RECT 56.565 155.215 56.735 155.405 ;
        RECT 58.400 155.245 58.520 155.355 ;
        RECT 56.255 155.195 56.275 155.215 ;
        RECT 58.865 155.195 59.035 155.405 ;
        RECT 62.545 155.215 62.715 155.405 ;
        RECT 68.065 155.385 68.230 155.405 ;
        RECT 65.315 155.250 65.475 155.360 ;
        RECT 66.225 155.195 66.395 155.385 ;
        RECT 68.065 155.215 68.235 155.385 ;
        RECT 69.905 155.215 70.075 155.405 ;
        RECT 70.370 155.215 70.540 155.405 ;
        RECT 71.745 155.195 71.915 155.405 ;
        RECT 72.205 155.195 72.375 155.385 ;
        RECT 75.885 155.195 76.055 155.385 ;
        RECT 80.945 155.215 81.115 155.405 ;
        RECT 81.400 155.245 81.520 155.355 ;
        RECT 82.325 155.215 82.495 155.405 ;
        RECT 86.465 155.195 86.635 155.385 ;
        RECT 86.930 155.195 87.100 155.385 ;
        RECT 87.845 155.215 88.015 155.405 ;
        RECT 89.235 155.240 89.395 155.350 ;
        RECT 90.145 155.215 90.315 155.385 ;
        RECT 93.365 155.195 93.535 155.405 ;
        RECT 95.205 155.195 95.375 155.385 ;
        RECT 97.040 155.245 97.160 155.355 ;
        RECT 97.510 155.215 97.680 155.405 ;
        RECT 98.885 155.215 99.055 155.405 ;
        RECT 100.725 155.195 100.895 155.385 ;
        RECT 102.560 155.245 102.680 155.355 ;
        RECT 103.025 155.195 103.195 155.385 ;
        RECT 104.405 155.215 104.575 155.405 ;
        RECT 107.160 155.245 107.280 155.355 ;
        RECT 108.085 155.215 108.255 155.405 ;
        RECT 110.395 155.240 110.555 155.350 ;
        RECT 111.760 155.245 111.880 155.355 ;
        RECT 112.225 155.215 112.395 155.405 ;
        RECT 119.130 155.385 119.265 155.405 ;
        RECT 114.065 155.195 114.235 155.385 ;
        RECT 17.325 154.385 18.695 155.195 ;
        RECT 18.705 154.515 20.535 155.195 ;
        RECT 19.190 154.285 20.535 154.515 ;
        RECT 20.545 154.385 26.055 155.195 ;
        RECT 26.065 154.385 31.575 155.195 ;
        RECT 31.585 154.385 37.095 155.195 ;
        RECT 37.105 154.385 42.615 155.195 ;
        RECT 43.095 154.325 43.525 155.110 ;
        RECT 43.545 154.385 49.055 155.195 ;
        RECT 49.065 154.385 54.575 155.195 ;
        RECT 54.585 154.385 55.955 155.195 ;
        RECT 56.255 154.515 58.705 155.195 ;
        RECT 58.725 154.515 66.035 155.195 ;
        RECT 66.085 154.515 68.835 155.195 ;
        RECT 56.745 154.285 58.705 154.515 ;
        RECT 62.240 154.295 63.150 154.515 ;
        RECT 64.685 154.285 66.035 154.515 ;
        RECT 67.905 154.285 68.835 154.515 ;
        RECT 68.855 154.325 69.285 155.110 ;
        RECT 69.305 154.285 72.055 155.195 ;
        RECT 72.175 154.515 75.640 155.195 ;
        RECT 75.745 154.515 83.055 155.195 ;
        RECT 74.720 154.285 75.640 154.515 ;
        RECT 79.260 154.295 80.170 154.515 ;
        RECT 81.705 154.285 83.055 154.515 ;
        RECT 83.200 154.515 86.665 155.195 ;
        RECT 86.785 154.515 89.060 155.195 ;
        RECT 90.410 154.515 92.835 155.195 ;
        RECT 83.200 154.285 84.120 154.515 ;
        RECT 87.690 154.285 89.060 154.515 ;
        RECT 93.225 154.385 94.595 155.195 ;
        RECT 94.615 154.325 95.045 155.110 ;
        RECT 95.065 154.385 100.575 155.195 ;
        RECT 100.585 154.385 102.415 155.195 ;
        RECT 102.885 154.515 110.195 155.195 ;
        RECT 106.400 154.295 107.310 154.515 ;
        RECT 108.845 154.285 110.195 154.515 ;
        RECT 111.165 154.285 114.375 155.195 ;
        RECT 114.385 155.165 115.340 155.195 ;
        RECT 116.370 155.165 116.540 155.385 ;
        RECT 116.825 155.195 116.995 155.385 ;
        RECT 118.205 155.215 118.375 155.385 ;
        RECT 119.130 155.215 119.300 155.385 ;
        RECT 119.585 155.215 119.755 155.405 ;
        RECT 118.210 155.195 118.375 155.215 ;
        RECT 120.965 155.195 121.135 155.385 ;
        RECT 121.420 155.245 121.540 155.355 ;
        RECT 122.800 155.215 122.970 155.405 ;
        RECT 126.950 155.385 127.115 155.405 ;
        RECT 123.265 155.215 123.435 155.385 ;
        RECT 124.185 155.195 124.355 155.385 ;
        RECT 126.480 155.245 126.600 155.355 ;
        RECT 126.945 155.215 127.115 155.385 ;
        RECT 129.705 155.195 129.875 155.385 ;
        RECT 131.545 155.215 131.715 155.405 ;
        RECT 132.005 155.215 132.175 155.405 ;
        RECT 132.465 155.195 132.635 155.385 ;
        RECT 134.305 155.195 134.475 155.385 ;
        RECT 135.040 155.195 135.210 155.385 ;
        RECT 135.220 155.215 135.390 155.405 ;
        RECT 135.685 155.215 135.855 155.405 ;
        RECT 137.340 155.215 137.510 155.405 ;
        RECT 142.125 155.195 142.295 155.385 ;
        RECT 142.585 155.195 142.755 155.385 ;
        RECT 143.965 155.195 144.135 155.385 ;
        RECT 144.425 155.215 144.595 155.405 ;
        RECT 144.895 155.250 145.055 155.360 ;
        RECT 146.725 155.195 146.895 155.405 ;
        RECT 114.385 154.485 116.665 155.165 ;
        RECT 114.385 154.285 115.340 154.485 ;
        RECT 116.695 154.285 118.045 155.195 ;
        RECT 118.210 154.515 120.045 155.195 ;
        RECT 119.115 154.285 120.045 154.515 ;
        RECT 120.375 154.325 120.805 155.110 ;
        RECT 120.825 154.285 124.035 155.195 ;
        RECT 124.045 154.385 129.555 155.195 ;
        RECT 129.565 154.415 130.935 155.195 ;
        RECT 130.945 154.515 132.775 155.195 ;
        RECT 132.785 154.515 134.615 155.195 ;
        RECT 134.625 154.515 138.525 155.195 ;
        RECT 138.860 154.515 142.325 155.195 ;
        RECT 130.945 154.285 132.290 154.515 ;
        RECT 132.785 154.285 134.130 154.515 ;
        RECT 134.625 154.285 135.555 154.515 ;
        RECT 138.860 154.285 139.780 154.515 ;
        RECT 142.445 154.415 143.815 155.195 ;
        RECT 143.825 154.515 145.655 155.195 ;
        RECT 144.310 154.285 145.655 154.515 ;
        RECT 145.665 154.385 147.035 155.195 ;
      LAYER nwell ;
        RECT 17.130 151.165 147.230 153.995 ;
      LAYER pwell ;
        RECT 17.325 149.965 18.695 150.775 ;
        RECT 18.705 149.965 24.215 150.775 ;
        RECT 24.225 149.965 29.735 150.775 ;
        RECT 30.215 150.050 30.645 150.835 ;
        RECT 30.665 149.965 33.415 150.775 ;
        RECT 34.195 150.645 35.125 150.875 ;
        RECT 36.185 150.645 37.105 150.875 ;
        RECT 34.195 149.965 36.030 150.645 ;
        RECT 36.185 149.965 38.475 150.645 ;
        RECT 38.485 149.965 40.315 150.875 ;
        RECT 40.325 149.965 43.075 150.875 ;
        RECT 43.085 149.965 46.755 150.775 ;
        RECT 48.135 150.645 49.055 150.875 ;
        RECT 46.765 149.965 49.055 150.645 ;
        RECT 49.065 149.965 54.575 150.775 ;
        RECT 54.585 149.965 55.935 150.875 ;
        RECT 55.975 150.050 56.405 150.835 ;
        RECT 57.795 150.645 58.715 150.875 ;
        RECT 62.240 150.645 63.150 150.865 ;
        RECT 64.685 150.645 66.035 150.875 ;
        RECT 56.425 149.965 58.715 150.645 ;
        RECT 58.725 149.965 66.035 150.645 ;
        RECT 66.095 149.965 68.825 150.875 ;
        RECT 68.845 149.965 70.195 150.875 ;
        RECT 70.780 150.645 71.700 150.875 ;
        RECT 77.880 150.645 78.790 150.865 ;
        RECT 80.325 150.645 81.675 150.875 ;
        RECT 70.780 149.965 74.245 150.645 ;
        RECT 74.365 149.965 81.675 150.645 ;
        RECT 81.735 150.050 82.165 150.835 ;
        RECT 82.185 149.965 83.535 150.875 ;
        RECT 83.565 149.965 85.395 150.775 ;
        RECT 85.420 149.965 87.235 150.875 ;
        RECT 87.735 150.675 89.115 150.875 ;
        RECT 87.735 149.995 90.440 150.675 ;
        RECT 93.980 150.645 94.890 150.865 ;
        RECT 96.425 150.645 97.775 150.875 ;
        RECT 87.735 149.965 89.115 149.995 ;
        RECT 17.465 149.755 17.635 149.965 ;
        RECT 18.845 149.755 19.015 149.965 ;
        RECT 24.365 149.755 24.535 149.965 ;
        RECT 29.880 149.910 30.000 149.915 ;
        RECT 29.880 149.805 30.055 149.910 ;
        RECT 29.895 149.800 30.055 149.805 ;
        RECT 30.805 149.775 30.975 149.965 ;
        RECT 35.865 149.945 36.030 149.965 ;
        RECT 31.730 149.755 31.900 149.945 ;
        RECT 32.185 149.755 32.355 149.945 ;
        RECT 33.560 149.805 33.680 149.915 ;
        RECT 34.485 149.755 34.655 149.945 ;
        RECT 35.865 149.775 36.035 149.945 ;
        RECT 38.165 149.775 38.335 149.965 ;
        RECT 40.000 149.775 40.170 149.965 ;
        RECT 41.845 149.755 42.015 149.945 ;
        RECT 42.765 149.775 42.935 149.965 ;
        RECT 43.225 149.775 43.395 149.965 ;
        RECT 43.685 149.755 43.855 149.945 ;
        RECT 45.525 149.755 45.695 149.945 ;
        RECT 46.905 149.775 47.075 149.965 ;
        RECT 48.745 149.755 48.915 149.945 ;
        RECT 49.205 149.775 49.375 149.965 ;
        RECT 50.130 149.755 50.300 149.945 ;
        RECT 54.730 149.775 54.900 149.965 ;
        RECT 56.565 149.945 56.735 149.965 ;
        RECT 55.185 149.755 55.355 149.945 ;
        RECT 55.655 149.800 55.815 149.910 ;
        RECT 56.565 149.775 56.740 149.945 ;
        RECT 58.865 149.775 59.035 149.965 ;
        RECT 60.255 149.800 60.415 149.910 ;
        RECT 56.570 149.755 56.740 149.775 ;
        RECT 61.165 149.755 61.335 149.945 ;
        RECT 66.225 149.775 66.395 149.965 ;
        RECT 69.910 149.945 70.080 149.965 ;
        RECT 66.225 149.755 66.390 149.775 ;
        RECT 66.685 149.755 66.855 149.945 ;
        RECT 68.520 149.805 68.640 149.915 ;
        RECT 69.440 149.805 69.560 149.915 ;
        RECT 69.905 149.775 70.080 149.945 ;
        RECT 70.360 149.805 70.480 149.915 ;
        RECT 74.045 149.775 74.215 149.965 ;
        RECT 74.505 149.775 74.675 149.965 ;
        RECT 69.905 149.755 70.075 149.775 ;
        RECT 77.265 149.755 77.435 149.945 ;
        RECT 80.020 149.805 80.140 149.915 ;
        RECT 80.485 149.755 80.655 149.945 ;
        RECT 82.330 149.775 82.500 149.965 ;
        RECT 83.705 149.775 83.875 149.965 ;
        RECT 85.545 149.775 85.715 149.965 ;
        RECT 87.380 149.805 87.500 149.915 ;
        RECT 89.685 149.755 89.855 149.945 ;
        RECT 90.145 149.775 90.315 149.995 ;
        RECT 90.465 149.965 97.775 150.645 ;
        RECT 98.785 150.645 100.135 150.875 ;
        RECT 101.670 150.645 102.580 150.865 ;
        RECT 98.785 149.965 106.095 150.645 ;
        RECT 106.105 149.965 107.475 150.775 ;
        RECT 107.495 150.050 107.925 150.835 ;
        RECT 107.945 150.645 108.875 150.875 ;
        RECT 107.945 149.965 111.845 150.645 ;
        RECT 112.085 149.965 113.435 150.875 ;
        RECT 113.465 149.965 118.975 150.775 ;
        RECT 119.005 149.965 120.355 150.875 ;
        RECT 120.365 149.965 122.195 150.775 ;
        RECT 122.675 149.965 124.025 150.875 ;
        RECT 125.255 149.965 128.175 150.875 ;
        RECT 128.185 149.965 129.535 150.875 ;
        RECT 129.565 149.965 133.235 150.775 ;
        RECT 133.255 150.050 133.685 150.835 ;
        RECT 137.220 150.645 138.130 150.865 ;
        RECT 139.665 150.645 141.015 150.875 ;
        RECT 133.705 149.965 141.015 150.645 ;
        RECT 141.065 150.645 141.995 150.875 ;
        RECT 141.065 149.965 144.965 150.645 ;
        RECT 145.665 149.965 147.035 150.775 ;
        RECT 90.605 149.775 90.775 149.965 ;
        RECT 93.365 149.755 93.535 149.945 ;
        RECT 95.480 149.755 95.650 149.945 ;
        RECT 97.975 149.810 98.135 149.920 ;
        RECT 99.620 149.755 99.790 149.945 ;
        RECT 104.405 149.755 104.575 149.945 ;
        RECT 105.140 149.755 105.310 149.945 ;
        RECT 105.785 149.775 105.955 149.965 ;
        RECT 106.245 149.775 106.415 149.965 ;
        RECT 108.360 149.775 108.530 149.965 ;
        RECT 109.005 149.755 109.175 149.945 ;
        RECT 110.845 149.755 111.015 149.945 ;
        RECT 112.230 149.775 112.400 149.965 ;
        RECT 113.605 149.775 113.775 149.965 ;
        RECT 114.530 149.755 114.700 149.945 ;
        RECT 117.740 149.755 117.910 149.945 ;
        RECT 118.210 149.755 118.380 149.945 ;
        RECT 119.120 149.775 119.290 149.965 ;
        RECT 120.040 149.805 120.160 149.915 ;
        RECT 120.505 149.775 120.675 149.965 ;
        RECT 120.960 149.805 121.080 149.915 ;
        RECT 122.340 149.805 122.460 149.915 ;
        RECT 122.805 149.775 122.975 149.965 ;
        RECT 124.180 149.920 124.350 149.945 ;
        RECT 124.180 149.810 124.355 149.920 ;
        RECT 124.180 149.755 124.350 149.810 ;
        RECT 124.640 149.755 124.810 149.945 ;
        RECT 126.035 149.800 126.195 149.910 ;
        RECT 126.945 149.775 127.115 149.945 ;
        RECT 127.860 149.775 128.030 149.965 ;
        RECT 129.250 149.945 129.420 149.965 ;
        RECT 129.245 149.775 129.420 149.945 ;
        RECT 129.705 149.775 129.875 149.965 ;
        RECT 126.950 149.755 127.115 149.775 ;
        RECT 129.245 149.755 129.415 149.775 ;
        RECT 132.465 149.755 132.635 149.945 ;
        RECT 133.845 149.775 134.015 149.965 ;
        RECT 134.305 149.755 134.475 149.945 ;
        RECT 141.480 149.775 141.650 149.965 ;
        RECT 141.940 149.755 142.110 149.945 ;
        RECT 145.340 149.805 145.460 149.915 ;
        RECT 146.725 149.755 146.895 149.965 ;
        RECT 17.325 148.945 18.695 149.755 ;
        RECT 18.705 148.945 24.215 149.755 ;
        RECT 24.225 148.945 29.735 149.755 ;
        RECT 30.665 148.845 32.015 149.755 ;
        RECT 32.045 149.075 34.335 149.755 ;
        RECT 34.345 149.075 41.655 149.755 ;
        RECT 33.415 148.845 34.335 149.075 ;
        RECT 37.860 148.855 38.770 149.075 ;
        RECT 40.305 148.845 41.655 149.075 ;
        RECT 41.705 148.945 43.075 149.755 ;
        RECT 43.095 148.885 43.525 149.670 ;
        RECT 43.545 148.945 45.375 149.755 ;
        RECT 45.385 148.845 48.595 149.755 ;
        RECT 48.605 148.945 49.975 149.755 ;
        RECT 49.985 148.845 53.640 149.755 ;
        RECT 53.665 148.845 55.480 149.755 ;
        RECT 56.425 148.845 60.080 149.755 ;
        RECT 61.025 148.845 64.235 149.755 ;
        RECT 64.555 149.075 66.390 149.755 ;
        RECT 64.555 148.845 65.485 149.075 ;
        RECT 66.545 148.945 68.375 149.755 ;
        RECT 68.855 148.885 69.285 149.670 ;
        RECT 69.765 149.075 77.075 149.755 ;
        RECT 73.280 148.855 74.190 149.075 ;
        RECT 75.725 148.845 77.075 149.075 ;
        RECT 77.125 148.945 79.875 149.755 ;
        RECT 80.345 149.075 89.450 149.755 ;
        RECT 89.655 149.075 93.120 149.755 ;
        RECT 92.200 148.845 93.120 149.075 ;
        RECT 93.225 148.945 94.595 149.755 ;
        RECT 94.615 148.885 95.045 149.670 ;
        RECT 95.065 149.075 98.965 149.755 ;
        RECT 99.205 149.075 103.105 149.755 ;
        RECT 95.065 148.845 95.995 149.075 ;
        RECT 99.205 148.845 100.135 149.075 ;
        RECT 103.355 148.845 104.705 149.755 ;
        RECT 104.725 149.075 108.625 149.755 ;
        RECT 104.725 148.845 105.655 149.075 ;
        RECT 108.865 148.945 110.695 149.755 ;
        RECT 110.815 149.075 114.280 149.755 ;
        RECT 113.360 148.845 114.280 149.075 ;
        RECT 114.385 148.845 116.215 149.755 ;
        RECT 116.225 148.845 118.055 149.755 ;
        RECT 118.065 148.845 119.895 149.755 ;
        RECT 120.375 148.885 120.805 149.670 ;
        RECT 121.575 148.845 124.495 149.755 ;
        RECT 124.525 148.845 125.875 149.755 ;
        RECT 126.950 149.075 128.785 149.755 ;
        RECT 127.855 148.845 128.785 149.075 ;
        RECT 129.105 148.845 132.315 149.755 ;
        RECT 132.325 148.945 134.155 149.755 ;
        RECT 134.165 149.075 141.475 149.755 ;
        RECT 137.680 148.855 138.590 149.075 ;
        RECT 140.125 148.845 141.475 149.075 ;
        RECT 141.525 149.075 145.425 149.755 ;
        RECT 141.525 148.845 142.455 149.075 ;
        RECT 145.665 148.945 147.035 149.755 ;
      LAYER nwell ;
        RECT 17.130 145.725 147.230 148.555 ;
      LAYER pwell ;
        RECT 17.325 144.525 18.695 145.335 ;
        RECT 18.705 144.525 24.215 145.335 ;
        RECT 24.225 144.525 29.735 145.335 ;
        RECT 30.215 144.610 30.645 145.395 ;
        RECT 31.165 145.205 32.515 145.435 ;
        RECT 34.050 145.205 34.960 145.425 ;
        RECT 31.165 144.525 38.475 145.205 ;
        RECT 38.485 144.525 41.405 145.435 ;
        RECT 42.165 144.525 45.375 145.435 ;
        RECT 45.395 144.525 48.125 145.435 ;
        RECT 48.145 144.525 53.655 145.335 ;
        RECT 53.665 144.525 55.495 145.335 ;
        RECT 55.975 144.610 56.405 145.395 ;
        RECT 58.485 145.345 59.435 145.435 ;
        RECT 57.505 144.525 59.435 145.345 ;
        RECT 59.645 145.235 60.575 145.435 ;
        RECT 61.905 145.235 62.855 145.435 ;
        RECT 59.645 144.755 62.855 145.235 ;
        RECT 59.790 144.555 62.855 144.755 ;
        RECT 17.465 144.315 17.635 144.525 ;
        RECT 18.845 144.315 19.015 144.525 ;
        RECT 24.365 144.315 24.535 144.525 ;
        RECT 29.885 144.475 30.055 144.505 ;
        RECT 29.880 144.365 30.055 144.475 ;
        RECT 30.800 144.365 30.920 144.475 ;
        RECT 31.720 144.365 31.840 144.475 ;
        RECT 29.885 144.315 30.055 144.365 ;
        RECT 32.185 144.315 32.355 144.505 ;
        RECT 34.955 144.360 35.115 144.470 ;
        RECT 38.165 144.315 38.335 144.525 ;
        RECT 38.630 144.335 38.800 144.525 ;
        RECT 41.385 144.315 41.555 144.505 ;
        RECT 41.845 144.475 42.015 144.505 ;
        RECT 41.840 144.365 42.015 144.475 ;
        RECT 41.845 144.315 42.015 144.365 ;
        RECT 43.685 144.315 43.855 144.505 ;
        RECT 45.075 144.335 45.245 144.525 ;
        RECT 47.825 144.335 47.995 144.525 ;
        RECT 48.285 144.335 48.455 144.525 ;
        RECT 49.205 144.315 49.375 144.505 ;
        RECT 53.805 144.335 53.975 144.525 ;
        RECT 57.505 144.505 57.655 144.525 ;
        RECT 55.650 144.475 55.820 144.505 ;
        RECT 55.640 144.365 55.820 144.475 ;
        RECT 56.100 144.365 56.220 144.475 ;
        RECT 55.650 144.315 55.820 144.365 ;
        RECT 17.325 143.505 18.695 144.315 ;
        RECT 18.705 143.505 24.215 144.315 ;
        RECT 24.225 143.505 29.735 144.315 ;
        RECT 29.745 143.505 31.575 144.315 ;
        RECT 32.045 143.635 34.795 144.315 ;
        RECT 33.865 143.405 34.795 143.635 ;
        RECT 35.735 143.405 38.465 144.315 ;
        RECT 38.485 143.635 41.695 144.315 ;
        RECT 38.485 143.405 39.620 143.635 ;
        RECT 41.705 143.505 43.075 144.315 ;
        RECT 43.095 143.445 43.525 144.230 ;
        RECT 43.545 143.505 49.055 144.315 ;
        RECT 49.065 143.505 54.575 144.315 ;
        RECT 54.585 143.405 55.935 144.315 ;
        RECT 56.570 144.285 56.740 144.505 ;
        RECT 57.485 144.335 57.655 144.505 ;
        RECT 59.790 144.475 59.960 144.555 ;
        RECT 61.920 144.525 62.855 144.555 ;
        RECT 63.175 145.205 64.105 145.435 ;
        RECT 63.175 144.525 65.010 145.205 ;
        RECT 65.165 144.525 70.675 145.335 ;
        RECT 70.685 144.525 76.195 145.335 ;
        RECT 76.975 145.205 77.905 145.435 ;
        RECT 76.975 144.525 78.810 145.205 ;
        RECT 78.975 144.525 80.325 145.435 ;
        RECT 80.345 144.525 81.715 145.335 ;
        RECT 81.735 144.610 82.165 145.395 ;
        RECT 82.185 144.525 85.855 145.335 ;
        RECT 85.865 144.525 87.235 145.335 ;
        RECT 87.285 145.205 88.635 145.435 ;
        RECT 90.170 145.205 91.080 145.425 ;
        RECT 98.120 145.205 99.030 145.425 ;
        RECT 100.565 145.205 101.915 145.435 ;
        RECT 105.540 145.205 106.460 145.435 ;
        RECT 87.285 144.525 94.595 145.205 ;
        RECT 94.605 144.525 101.915 145.205 ;
        RECT 102.995 144.525 106.460 145.205 ;
        RECT 107.495 144.610 107.925 145.395 ;
        RECT 107.985 145.205 109.335 145.435 ;
        RECT 110.870 145.205 111.780 145.425 ;
        RECT 115.305 145.205 116.235 145.435 ;
        RECT 122.100 145.205 123.020 145.435 ;
        RECT 107.985 144.525 115.295 145.205 ;
        RECT 115.305 144.525 119.205 145.205 ;
        RECT 119.555 144.525 123.020 145.205 ;
        RECT 123.125 144.525 124.955 145.435 ;
        RECT 124.965 145.205 125.895 145.435 ;
        RECT 129.200 145.205 130.120 145.435 ;
        RECT 124.965 144.525 128.865 145.205 ;
        RECT 129.200 144.525 132.665 145.205 ;
        RECT 133.255 144.610 133.685 145.395 ;
        RECT 137.680 145.205 138.590 145.425 ;
        RECT 140.125 145.205 141.475 145.435 ;
        RECT 144.640 145.205 145.560 145.435 ;
        RECT 134.165 144.525 141.475 145.205 ;
        RECT 142.095 144.525 145.560 145.205 ;
        RECT 145.665 144.525 147.035 145.335 ;
        RECT 64.845 144.505 65.010 144.525 ;
        RECT 59.780 144.365 59.960 144.475 ;
        RECT 59.790 144.335 59.960 144.365 ;
        RECT 60.245 144.315 60.415 144.505 ;
        RECT 64.845 144.335 65.015 144.505 ;
        RECT 65.305 144.335 65.475 144.525 ;
        RECT 67.605 144.315 67.775 144.505 ;
        RECT 69.445 144.315 69.615 144.505 ;
        RECT 70.825 144.335 70.995 144.525 ;
        RECT 78.645 144.505 78.810 144.525 ;
        RECT 72.200 144.315 72.370 144.505 ;
        RECT 73.585 144.315 73.755 144.505 ;
        RECT 76.340 144.365 76.460 144.475 ;
        RECT 77.080 144.315 77.250 144.505 ;
        RECT 78.645 144.335 78.815 144.505 ;
        RECT 80.025 144.335 80.195 144.525 ;
        RECT 80.485 144.335 80.655 144.525 ;
        RECT 80.940 144.365 81.060 144.475 ;
        RECT 82.325 144.335 82.495 144.525 ;
        RECT 86.005 144.335 86.175 144.525 ;
        RECT 88.765 144.315 88.935 144.505 ;
        RECT 89.225 144.315 89.395 144.505 ;
        RECT 91.985 144.315 92.155 144.505 ;
        RECT 94.285 144.335 94.455 144.525 ;
        RECT 94.745 144.335 94.915 144.525 ;
        RECT 98.425 144.315 98.595 144.505 ;
        RECT 98.885 144.315 99.055 144.505 ;
        RECT 100.265 144.315 100.435 144.505 ;
        RECT 102.115 144.370 102.275 144.480 ;
        RECT 103.025 144.335 103.195 144.525 ;
        RECT 103.945 144.315 104.115 144.505 ;
        RECT 106.705 144.315 106.875 144.505 ;
        RECT 112.225 144.315 112.395 144.505 ;
        RECT 114.985 144.335 115.155 144.525 ;
        RECT 115.720 144.335 115.890 144.525 ;
        RECT 119.585 144.335 119.755 144.525 ;
        RECT 120.965 144.315 121.135 144.505 ;
        RECT 124.185 144.315 124.355 144.505 ;
        RECT 124.640 144.335 124.810 144.525 ;
        RECT 125.380 144.335 125.550 144.525 ;
        RECT 131.545 144.315 131.715 144.505 ;
        RECT 132.465 144.335 132.635 144.525 ;
        RECT 132.920 144.365 133.040 144.475 ;
        RECT 133.840 144.365 133.960 144.475 ;
        RECT 134.305 144.335 134.475 144.525 ;
        RECT 137.060 144.365 137.180 144.475 ;
        RECT 137.525 144.315 137.695 144.505 ;
        RECT 139.825 144.315 139.995 144.505 ;
        RECT 140.285 144.315 140.455 144.505 ;
        RECT 141.660 144.365 141.780 144.475 ;
        RECT 142.125 144.315 142.295 144.525 ;
        RECT 146.725 144.315 146.895 144.525 ;
        RECT 58.700 144.285 59.635 144.315 ;
        RECT 56.570 144.085 59.635 144.285 ;
        RECT 56.425 143.605 59.635 144.085 ;
        RECT 60.105 143.635 67.415 144.315 ;
        RECT 56.425 143.405 57.355 143.605 ;
        RECT 58.685 143.405 59.635 143.605 ;
        RECT 63.620 143.415 64.530 143.635 ;
        RECT 66.065 143.405 67.415 143.635 ;
        RECT 67.465 143.505 68.835 144.315 ;
        RECT 68.855 143.445 69.285 144.230 ;
        RECT 69.305 143.505 72.055 144.315 ;
        RECT 72.085 143.405 73.435 144.315 ;
        RECT 73.445 143.405 76.195 144.315 ;
        RECT 76.665 143.635 80.565 144.315 ;
        RECT 81.345 143.635 89.075 144.315 ;
        RECT 76.665 143.405 77.595 143.635 ;
        RECT 81.345 143.405 83.115 143.635 ;
        RECT 84.650 143.415 85.560 143.635 ;
        RECT 89.085 143.505 91.835 144.315 ;
        RECT 91.845 143.405 94.595 144.315 ;
        RECT 94.615 143.445 95.045 144.230 ;
        RECT 95.160 143.635 98.625 144.315 ;
        RECT 95.160 143.405 96.080 143.635 ;
        RECT 98.745 143.505 100.115 144.315 ;
        RECT 100.235 143.635 103.700 144.315 ;
        RECT 102.780 143.405 103.700 143.635 ;
        RECT 103.805 143.405 106.555 144.315 ;
        RECT 106.565 143.505 112.075 144.315 ;
        RECT 112.085 143.635 119.395 144.315 ;
        RECT 115.600 143.415 116.510 143.635 ;
        RECT 118.045 143.405 119.395 143.635 ;
        RECT 120.375 143.445 120.805 144.230 ;
        RECT 120.825 143.405 124.035 144.315 ;
        RECT 124.045 143.635 131.355 144.315 ;
        RECT 127.560 143.415 128.470 143.635 ;
        RECT 130.005 143.405 131.355 143.635 ;
        RECT 131.405 143.505 136.915 144.315 ;
        RECT 137.385 143.535 138.755 144.315 ;
        RECT 138.765 143.535 140.135 144.315 ;
        RECT 140.145 143.635 141.975 144.315 ;
        RECT 142.095 143.635 145.560 144.315 ;
        RECT 140.630 143.405 141.975 143.635 ;
        RECT 144.640 143.405 145.560 143.635 ;
        RECT 145.665 143.505 147.035 144.315 ;
      LAYER nwell ;
        RECT 17.130 140.285 147.230 143.115 ;
      LAYER pwell ;
        RECT 17.325 139.085 18.695 139.895 ;
        RECT 18.705 139.085 24.215 139.895 ;
        RECT 24.225 139.085 29.735 139.895 ;
        RECT 30.215 139.170 30.645 139.955 ;
        RECT 30.665 139.085 32.495 139.895 ;
        RECT 32.505 139.795 33.435 139.995 ;
        RECT 34.765 139.795 35.715 139.995 ;
        RECT 32.505 139.315 35.715 139.795 ;
        RECT 39.240 139.765 40.150 139.985 ;
        RECT 41.685 139.765 43.035 139.995 ;
        RECT 32.650 139.115 35.715 139.315 ;
        RECT 17.465 138.875 17.635 139.085 ;
        RECT 18.845 138.895 19.015 139.085 ;
        RECT 20.225 138.875 20.395 139.065 ;
        RECT 20.685 138.875 20.855 139.065 ;
        RECT 24.365 138.895 24.535 139.085 ;
        RECT 26.205 138.875 26.375 139.065 ;
        RECT 28.960 138.925 29.080 139.035 ;
        RECT 29.880 138.925 30.000 139.035 ;
        RECT 30.805 138.895 30.975 139.085 ;
        RECT 32.650 138.895 32.820 139.115 ;
        RECT 34.780 139.085 35.715 139.115 ;
        RECT 35.725 139.085 43.035 139.765 ;
        RECT 43.085 139.085 44.455 139.895 ;
        RECT 44.700 139.085 49.515 139.765 ;
        RECT 49.525 139.085 52.275 139.895 ;
        RECT 52.745 139.085 55.665 139.995 ;
        RECT 55.975 139.170 56.405 139.955 ;
        RECT 56.425 139.085 57.795 139.895 ;
        RECT 57.805 139.085 62.620 139.765 ;
        RECT 62.960 139.085 66.830 139.995 ;
        RECT 67.005 139.765 67.925 139.995 ;
        RECT 67.005 139.085 69.295 139.765 ;
        RECT 69.305 139.085 71.135 139.995 ;
        RECT 74.660 139.765 75.570 139.985 ;
        RECT 77.105 139.765 78.455 139.995 ;
        RECT 80.580 139.765 81.715 139.995 ;
        RECT 71.145 139.085 78.455 139.765 ;
        RECT 78.505 139.085 81.715 139.765 ;
        RECT 81.735 139.170 82.165 139.955 ;
        RECT 85.385 139.765 86.315 139.995 ;
        RECT 82.415 139.085 86.315 139.765 ;
        RECT 86.335 139.085 89.065 139.995 ;
        RECT 89.085 139.085 90.455 139.895 ;
        RECT 93.980 139.765 94.890 139.985 ;
        RECT 96.425 139.765 97.775 139.995 ;
        RECT 101.505 139.765 102.435 139.995 ;
        RECT 106.085 139.765 107.015 139.995 ;
        RECT 90.465 139.085 97.775 139.765 ;
        RECT 97.825 139.085 100.565 139.765 ;
        RECT 101.505 139.085 104.255 139.765 ;
        RECT 104.265 139.085 107.015 139.765 ;
        RECT 107.495 139.170 107.925 139.955 ;
        RECT 107.945 139.085 113.455 139.895 ;
        RECT 113.465 139.085 118.975 139.895 ;
        RECT 118.985 139.085 120.355 139.895 ;
        RECT 120.365 139.085 123.575 139.995 ;
        RECT 123.605 139.085 124.955 139.995 ;
        RECT 124.965 139.085 128.635 139.895 ;
        RECT 128.645 139.085 130.015 139.895 ;
        RECT 130.025 139.085 133.235 139.995 ;
        RECT 133.255 139.170 133.685 139.955 ;
        RECT 134.625 139.765 135.555 139.995 ;
        RECT 138.860 139.765 139.780 139.995 ;
        RECT 134.625 139.085 138.525 139.765 ;
        RECT 138.860 139.085 142.325 139.765 ;
        RECT 142.445 139.085 143.815 139.865 ;
        RECT 144.310 139.765 145.655 139.995 ;
        RECT 143.825 139.085 145.655 139.765 ;
        RECT 145.665 139.085 147.035 139.895 ;
        RECT 35.865 138.895 36.035 139.085 ;
        RECT 36.325 138.875 36.495 139.065 ;
        RECT 36.785 138.875 36.955 139.065 ;
        RECT 40.005 138.895 40.175 139.065 ;
        RECT 40.005 138.875 40.170 138.895 ;
        RECT 40.465 138.875 40.635 139.065 ;
        RECT 43.225 138.895 43.395 139.085 ;
        RECT 43.695 138.920 43.855 139.030 ;
        RECT 44.605 138.895 44.775 139.065 ;
        RECT 48.740 138.925 48.860 139.035 ;
        RECT 49.205 138.895 49.375 139.085 ;
        RECT 49.665 138.895 49.835 139.085 ;
        RECT 44.630 138.875 44.775 138.895 ;
        RECT 49.225 138.875 49.375 138.895 ;
        RECT 17.325 138.065 18.695 138.875 ;
        RECT 18.705 138.195 20.535 138.875 ;
        RECT 18.705 137.965 20.050 138.195 ;
        RECT 20.545 138.065 26.055 138.875 ;
        RECT 26.065 138.065 28.815 138.875 ;
        RECT 29.325 138.195 36.635 138.875 ;
        RECT 29.325 137.965 30.675 138.195 ;
        RECT 32.210 137.975 33.120 138.195 ;
        RECT 36.645 138.065 38.015 138.875 ;
        RECT 38.335 138.195 40.170 138.875 ;
        RECT 38.335 137.965 39.265 138.195 ;
        RECT 40.335 137.965 43.065 138.875 ;
        RECT 43.095 138.005 43.525 138.790 ;
        RECT 44.630 137.965 48.500 138.875 ;
        RECT 49.225 138.055 51.155 138.875 ;
        RECT 51.510 138.845 51.680 139.065 ;
        RECT 52.420 138.925 52.540 139.035 ;
        RECT 52.890 138.895 53.060 139.085 ;
        RECT 54.735 138.920 54.895 139.030 ;
        RECT 56.565 138.895 56.735 139.085 ;
        RECT 57.945 138.895 58.115 139.085 ;
        RECT 66.685 139.065 66.830 139.085 ;
        RECT 62.545 138.875 62.715 139.065 ;
        RECT 64.845 138.895 65.015 139.065 ;
        RECT 64.845 138.875 65.010 138.895 ;
        RECT 65.305 138.875 65.475 139.065 ;
        RECT 66.685 138.895 66.855 139.065 ;
        RECT 68.985 138.895 69.155 139.085 ;
        RECT 69.450 138.895 69.620 139.085 ;
        RECT 70.365 138.875 70.535 139.065 ;
        RECT 71.285 138.895 71.455 139.085 ;
        RECT 77.735 138.920 77.895 139.030 ;
        RECT 78.645 138.875 78.815 139.085 ;
        RECT 82.325 138.875 82.495 139.065 ;
        RECT 85.730 138.895 85.900 139.085 ;
        RECT 53.640 138.845 54.575 138.875 ;
        RECT 51.510 138.645 54.575 138.845 ;
        RECT 50.205 137.965 51.155 138.055 ;
        RECT 51.365 138.165 54.575 138.645 ;
        RECT 51.365 137.965 52.295 138.165 ;
        RECT 53.625 137.965 54.575 138.165 ;
        RECT 55.545 138.195 62.855 138.875 ;
        RECT 63.175 138.195 65.010 138.875 ;
        RECT 55.545 137.965 56.895 138.195 ;
        RECT 58.430 137.975 59.340 138.195 ;
        RECT 63.175 137.965 64.105 138.195 ;
        RECT 65.165 138.065 68.835 138.875 ;
        RECT 68.855 138.005 69.285 138.790 ;
        RECT 70.225 138.195 77.535 138.875 ;
        RECT 78.615 138.195 82.080 138.875 ;
        RECT 82.295 138.195 85.760 138.875 ;
        RECT 86.005 138.845 86.175 139.065 ;
        RECT 88.765 138.875 88.935 139.085 ;
        RECT 89.225 138.895 89.395 139.085 ;
        RECT 90.605 138.895 90.775 139.085 ;
        RECT 94.280 138.925 94.400 139.035 ;
        RECT 95.205 138.875 95.375 139.065 ;
        RECT 97.965 138.895 98.135 139.085 ;
        RECT 100.735 138.875 100.905 139.065 ;
        RECT 101.195 138.920 101.355 139.030 ;
        RECT 102.105 138.875 102.275 139.065 ;
        RECT 103.945 138.895 104.115 139.085 ;
        RECT 104.405 138.895 104.575 139.085 ;
        RECT 107.160 138.925 107.280 139.035 ;
        RECT 108.085 138.895 108.255 139.085 ;
        RECT 109.465 138.875 109.635 139.065 ;
        RECT 113.605 138.895 113.775 139.085 ;
        RECT 116.825 138.875 116.995 139.065 ;
        RECT 119.125 138.895 119.295 139.085 ;
        RECT 120.505 138.895 120.675 139.085 ;
        RECT 123.720 138.895 123.890 139.085 ;
        RECT 124.185 138.875 124.355 139.065 ;
        RECT 124.645 138.875 124.815 139.065 ;
        RECT 125.105 138.895 125.275 139.085 ;
        RECT 128.325 138.875 128.495 139.065 ;
        RECT 128.785 138.895 128.955 139.085 ;
        RECT 129.705 138.875 129.875 139.065 ;
        RECT 130.165 138.895 130.335 139.085 ;
        RECT 132.920 138.925 133.040 139.035 ;
        RECT 133.385 138.875 133.555 139.065 ;
        RECT 133.855 138.930 134.015 139.040 ;
        RECT 135.040 138.895 135.210 139.085 ;
        RECT 140.745 138.875 140.915 139.065 ;
        RECT 142.125 138.875 142.295 139.085 ;
        RECT 143.505 138.895 143.675 139.085 ;
        RECT 143.965 138.875 144.135 139.085 ;
        RECT 146.725 138.875 146.895 139.085 ;
        RECT 87.205 138.845 88.585 138.875 ;
        RECT 73.740 137.975 74.650 138.195 ;
        RECT 76.185 137.965 77.535 138.195 ;
        RECT 81.160 137.965 82.080 138.195 ;
        RECT 84.840 137.965 85.760 138.195 ;
        RECT 85.880 138.165 88.585 138.845 ;
        RECT 87.205 137.965 88.585 138.165 ;
        RECT 88.625 138.065 94.135 138.875 ;
        RECT 94.615 138.005 95.045 138.790 ;
        RECT 95.065 138.065 97.815 138.875 ;
        RECT 97.825 137.965 101.035 138.875 ;
        RECT 101.965 138.195 109.275 138.875 ;
        RECT 109.325 138.195 116.635 138.875 ;
        RECT 105.480 137.975 106.390 138.195 ;
        RECT 107.925 137.965 109.275 138.195 ;
        RECT 112.840 137.975 113.750 138.195 ;
        RECT 115.285 137.965 116.635 138.195 ;
        RECT 116.685 138.065 120.355 138.875 ;
        RECT 120.375 138.005 120.805 138.790 ;
        RECT 120.920 138.195 124.385 138.875 ;
        RECT 120.920 137.965 121.840 138.195 ;
        RECT 124.505 138.065 128.175 138.875 ;
        RECT 128.185 138.065 129.555 138.875 ;
        RECT 129.565 137.965 132.775 138.875 ;
        RECT 133.245 138.195 140.555 138.875 ;
        RECT 136.760 137.975 137.670 138.195 ;
        RECT 139.205 137.965 140.555 138.195 ;
        RECT 140.605 138.095 141.975 138.875 ;
        RECT 141.985 138.195 143.815 138.875 ;
        RECT 143.825 138.195 145.655 138.875 ;
        RECT 142.470 137.965 143.815 138.195 ;
        RECT 144.310 137.965 145.655 138.195 ;
        RECT 145.665 138.065 147.035 138.875 ;
      LAYER nwell ;
        RECT 17.130 134.845 147.230 137.675 ;
      LAYER pwell ;
        RECT 17.325 133.645 18.695 134.455 ;
        RECT 18.705 134.325 20.050 134.555 ;
        RECT 18.705 133.645 20.535 134.325 ;
        RECT 20.545 133.645 26.055 134.455 ;
        RECT 26.065 133.645 29.735 134.455 ;
        RECT 30.215 133.730 30.645 134.515 ;
        RECT 30.665 133.645 34.335 134.455 ;
        RECT 36.635 134.325 37.555 134.555 ;
        RECT 35.265 133.645 37.555 134.325 ;
        RECT 37.565 134.355 38.495 134.555 ;
        RECT 39.825 134.355 40.775 134.555 ;
        RECT 37.565 133.875 40.775 134.355 ;
        RECT 44.300 134.325 45.210 134.545 ;
        RECT 46.745 134.325 48.095 134.555 ;
        RECT 49.515 134.325 50.435 134.555 ;
        RECT 52.415 134.325 53.345 134.555 ;
        RECT 55.035 134.325 55.955 134.555 ;
        RECT 37.710 133.675 40.775 133.875 ;
        RECT 17.465 133.435 17.635 133.645 ;
        RECT 18.840 133.485 18.960 133.595 ;
        RECT 19.305 133.435 19.475 133.625 ;
        RECT 20.225 133.455 20.395 133.645 ;
        RECT 20.685 133.455 20.855 133.645 ;
        RECT 26.205 133.455 26.375 133.645 ;
        RECT 26.675 133.480 26.835 133.590 ;
        RECT 27.585 133.455 27.755 133.625 ;
        RECT 29.885 133.595 30.055 133.625 ;
        RECT 29.880 133.485 30.055 133.595 ;
        RECT 27.590 133.435 27.755 133.455 ;
        RECT 29.885 133.435 30.055 133.485 ;
        RECT 30.805 133.455 30.975 133.645 ;
        RECT 34.495 133.490 34.655 133.600 ;
        RECT 35.405 133.595 35.575 133.645 ;
        RECT 35.400 133.485 35.575 133.595 ;
        RECT 35.405 133.455 35.575 133.485 ;
        RECT 35.865 133.435 36.035 133.625 ;
        RECT 37.710 133.455 37.880 133.675 ;
        RECT 39.840 133.645 40.775 133.675 ;
        RECT 40.785 133.645 48.095 134.325 ;
        RECT 48.145 133.645 50.435 134.325 ;
        RECT 51.510 133.645 53.345 134.325 ;
        RECT 53.665 133.645 55.955 134.325 ;
        RECT 55.975 133.730 56.405 134.515 ;
        RECT 59.940 134.325 60.850 134.545 ;
        RECT 62.385 134.325 63.735 134.555 ;
        RECT 56.425 133.645 63.735 134.325 ;
        RECT 63.785 133.645 69.295 134.455 ;
        RECT 69.305 133.645 72.055 134.455 ;
        RECT 75.580 134.325 76.490 134.545 ;
        RECT 78.025 134.325 79.375 134.555 ;
        RECT 72.065 133.645 79.375 134.325 ;
        RECT 79.425 133.645 81.255 134.555 ;
        RECT 81.735 133.730 82.165 134.515 ;
        RECT 82.280 134.325 83.200 134.555 ;
        RECT 82.280 133.645 85.745 134.325 ;
        RECT 85.885 133.645 87.235 134.555 ;
        RECT 91.680 134.325 92.590 134.545 ;
        RECT 94.125 134.325 95.475 134.555 ;
        RECT 88.165 133.645 95.475 134.325 ;
        RECT 95.525 133.645 96.895 134.455 ;
        RECT 96.905 133.645 100.115 134.555 ;
        RECT 100.125 133.645 102.875 134.455 ;
        RECT 103.345 134.325 104.275 134.555 ;
        RECT 103.345 133.645 107.245 134.325 ;
        RECT 107.495 133.730 107.925 134.515 ;
        RECT 107.945 134.325 108.875 134.555 ;
        RECT 107.945 133.645 111.845 134.325 ;
        RECT 112.085 133.645 117.595 134.455 ;
        RECT 118.565 134.325 119.915 134.555 ;
        RECT 121.450 134.325 122.360 134.545 ;
        RECT 128.540 134.325 129.460 134.555 ;
        RECT 118.565 133.645 125.875 134.325 ;
        RECT 125.995 133.645 129.460 134.325 ;
        RECT 129.565 133.645 133.235 134.455 ;
        RECT 133.255 133.730 133.685 134.515 ;
        RECT 137.220 134.325 138.130 134.545 ;
        RECT 139.665 134.325 141.015 134.555 ;
        RECT 133.705 133.645 141.015 134.325 ;
        RECT 141.160 134.325 142.080 134.555 ;
        RECT 141.160 133.645 144.625 134.325 ;
        RECT 145.665 133.645 147.035 134.455 ;
        RECT 40.925 133.455 41.095 133.645 ;
        RECT 44.610 133.435 44.780 133.625 ;
        RECT 45.065 133.435 45.235 133.625 ;
        RECT 48.285 133.455 48.455 133.645 ;
        RECT 51.510 133.625 51.675 133.645 ;
        RECT 50.595 133.480 50.755 133.600 ;
        RECT 51.505 133.455 51.675 133.625 ;
        RECT 53.805 133.455 53.975 133.645 ;
        RECT 56.565 133.455 56.735 133.645 ;
        RECT 58.405 133.435 58.575 133.625 ;
        RECT 58.865 133.435 59.035 133.625 ;
        RECT 63.925 133.455 64.095 133.645 ;
        RECT 64.385 133.435 64.555 133.625 ;
        RECT 65.765 133.435 65.935 133.625 ;
        RECT 69.445 133.435 69.615 133.645 ;
        RECT 72.205 133.455 72.375 133.645 ;
        RECT 74.505 133.435 74.675 133.625 ;
        RECT 77.270 133.435 77.440 133.625 ;
        RECT 79.105 133.435 79.275 133.625 ;
        RECT 79.570 133.455 79.740 133.645 ;
        RECT 81.400 133.485 81.520 133.595 ;
        RECT 84.620 133.485 84.740 133.595 ;
        RECT 85.085 133.435 85.255 133.625 ;
        RECT 85.545 133.455 85.715 133.645 ;
        RECT 86.000 133.455 86.170 133.645 ;
        RECT 86.465 133.435 86.635 133.625 ;
        RECT 87.395 133.490 87.555 133.600 ;
        RECT 88.305 133.455 88.475 133.645 ;
        RECT 88.760 133.485 88.880 133.595 ;
        RECT 89.500 133.435 89.670 133.625 ;
        RECT 93.365 133.435 93.535 133.625 ;
        RECT 95.205 133.435 95.375 133.625 ;
        RECT 95.665 133.455 95.835 133.645 ;
        RECT 97.035 133.455 97.205 133.645 ;
        RECT 100.265 133.455 100.435 133.645 ;
        RECT 100.725 133.435 100.895 133.625 ;
        RECT 102.565 133.435 102.735 133.625 ;
        RECT 103.020 133.485 103.140 133.595 ;
        RECT 103.760 133.455 103.930 133.645 ;
        RECT 106.245 133.435 106.415 133.625 ;
        RECT 108.085 133.435 108.255 133.625 ;
        RECT 108.360 133.455 108.530 133.645 ;
        RECT 112.225 133.455 112.395 133.645 ;
        RECT 113.145 133.435 113.315 133.625 ;
        RECT 113.605 133.435 113.775 133.625 ;
        RECT 117.280 133.485 117.400 133.595 ;
        RECT 117.755 133.490 117.915 133.600 ;
        RECT 120.045 133.435 120.215 133.625 ;
        RECT 125.565 133.455 125.735 133.645 ;
        RECT 126.025 133.455 126.195 133.645 ;
        RECT 127.865 133.435 128.035 133.625 ;
        RECT 128.325 133.435 128.495 133.625 ;
        RECT 129.705 133.455 129.875 133.645 ;
        RECT 131.085 133.435 131.255 133.625 ;
        RECT 133.845 133.455 134.015 133.645 ;
        RECT 134.120 133.435 134.290 133.625 ;
        RECT 138.260 133.435 138.430 133.625 ;
        RECT 142.125 133.435 142.295 133.625 ;
        RECT 143.500 133.485 143.620 133.595 ;
        RECT 143.965 133.435 144.135 133.625 ;
        RECT 144.425 133.455 144.595 133.645 ;
        RECT 144.895 133.490 145.055 133.600 ;
        RECT 146.725 133.435 146.895 133.645 ;
        RECT 17.325 132.625 18.695 133.435 ;
        RECT 19.165 132.755 26.475 133.435 ;
        RECT 27.590 132.755 29.425 133.435 ;
        RECT 22.680 132.535 23.590 132.755 ;
        RECT 25.125 132.525 26.475 132.755 ;
        RECT 28.495 132.525 29.425 132.755 ;
        RECT 29.745 132.625 35.255 133.435 ;
        RECT 35.725 132.755 43.035 133.435 ;
        RECT 39.240 132.535 40.150 132.755 ;
        RECT 41.685 132.525 43.035 132.755 ;
        RECT 43.095 132.565 43.525 133.350 ;
        RECT 43.545 132.525 44.895 133.435 ;
        RECT 44.925 132.625 50.435 133.435 ;
        RECT 51.405 132.755 58.715 133.435 ;
        RECT 51.405 132.525 52.755 132.755 ;
        RECT 54.290 132.535 55.200 132.755 ;
        RECT 58.725 132.625 64.235 133.435 ;
        RECT 64.245 132.625 65.615 133.435 ;
        RECT 65.675 132.525 68.835 133.435 ;
        RECT 68.855 132.565 69.285 133.350 ;
        RECT 69.305 132.755 74.120 133.435 ;
        RECT 74.365 132.625 77.115 133.435 ;
        RECT 77.125 132.525 78.955 133.435 ;
        RECT 78.965 132.625 84.475 133.435 ;
        RECT 84.955 132.525 86.305 133.435 ;
        RECT 86.325 132.755 88.615 133.435 ;
        RECT 87.695 132.525 88.615 132.755 ;
        RECT 89.085 132.755 92.985 133.435 ;
        RECT 89.085 132.525 90.015 132.755 ;
        RECT 93.225 132.625 94.595 133.435 ;
        RECT 94.615 132.565 95.045 133.350 ;
        RECT 95.065 132.625 100.575 133.435 ;
        RECT 100.585 132.625 102.415 133.435 ;
        RECT 102.535 132.755 106.000 133.435 ;
        RECT 105.080 132.525 106.000 132.755 ;
        RECT 106.105 132.625 107.935 133.435 ;
        RECT 107.945 132.525 110.695 133.435 ;
        RECT 110.715 132.755 113.455 133.435 ;
        RECT 113.465 132.625 117.135 133.435 ;
        RECT 117.605 132.525 120.355 133.435 ;
        RECT 120.375 132.565 120.805 133.350 ;
        RECT 120.865 132.755 128.175 133.435 ;
        RECT 120.865 132.525 122.215 132.755 ;
        RECT 123.750 132.535 124.660 132.755 ;
        RECT 128.185 132.525 130.935 133.435 ;
        RECT 130.945 132.625 133.695 133.435 ;
        RECT 133.705 132.755 137.605 133.435 ;
        RECT 137.845 132.755 141.745 133.435 ;
        RECT 133.705 132.525 134.635 132.755 ;
        RECT 137.845 132.525 138.775 132.755 ;
        RECT 141.985 132.655 143.355 133.435 ;
        RECT 143.825 132.755 145.655 133.435 ;
        RECT 144.310 132.525 145.655 132.755 ;
        RECT 145.665 132.625 147.035 133.435 ;
      LAYER nwell ;
        RECT 17.130 129.405 147.230 132.235 ;
      LAYER pwell ;
        RECT 17.325 128.205 18.695 129.015 ;
        RECT 18.705 128.885 19.635 129.115 ;
        RECT 22.885 128.885 24.235 129.115 ;
        RECT 25.770 128.885 26.680 129.105 ;
        RECT 18.705 128.205 22.605 128.885 ;
        RECT 22.885 128.205 30.195 128.885 ;
        RECT 30.215 128.290 30.645 129.075 ;
        RECT 30.745 128.205 33.745 129.115 ;
        RECT 33.885 128.205 39.395 129.015 ;
        RECT 39.405 128.205 44.915 129.015 ;
        RECT 44.925 128.205 50.435 129.015 ;
        RECT 50.445 128.205 55.955 129.015 ;
        RECT 55.975 128.290 56.405 129.075 ;
        RECT 56.425 128.205 61.935 129.015 ;
        RECT 61.945 128.205 67.455 129.015 ;
        RECT 67.465 128.205 68.835 129.015 ;
        RECT 68.885 128.205 72.055 129.115 ;
        RECT 72.065 128.915 73.015 129.115 ;
        RECT 74.345 128.915 75.275 129.115 ;
        RECT 72.065 128.435 75.275 128.915 ;
        RECT 72.065 128.235 75.130 128.435 ;
        RECT 72.065 128.205 73.000 128.235 ;
        RECT 17.465 127.995 17.635 128.205 ;
        RECT 19.120 128.015 19.290 128.205 ;
        RECT 20.225 127.995 20.395 128.185 ;
        RECT 20.695 127.995 20.865 128.185 ;
        RECT 22.065 127.995 22.235 128.185 ;
        RECT 24.825 127.995 24.995 128.185 ;
        RECT 29.885 128.015 30.055 128.205 ;
        RECT 30.805 128.015 30.975 128.205 ;
        RECT 32.185 127.995 32.355 128.185 ;
        RECT 33.565 127.995 33.735 128.185 ;
        RECT 34.025 128.015 34.195 128.205 ;
        RECT 39.085 127.995 39.255 128.185 ;
        RECT 39.545 128.015 39.715 128.205 ;
        RECT 42.760 128.045 42.880 128.155 ;
        RECT 43.685 127.995 43.855 128.185 ;
        RECT 45.065 128.015 45.235 128.205 ;
        RECT 49.205 127.995 49.375 128.185 ;
        RECT 50.585 128.015 50.755 128.205 ;
        RECT 54.725 127.995 54.895 128.185 ;
        RECT 56.565 128.015 56.735 128.205 ;
        RECT 60.245 127.995 60.415 128.185 ;
        RECT 62.085 128.015 62.255 128.205 ;
        RECT 63.925 127.995 64.095 128.185 ;
        RECT 66.220 127.995 66.390 128.185 ;
        RECT 67.605 128.015 67.775 128.205 ;
        RECT 68.525 128.015 68.695 128.185 ;
        RECT 68.985 128.015 69.155 128.205 ;
        RECT 68.525 127.995 68.690 128.015 ;
        RECT 69.445 127.995 69.615 128.185 ;
        RECT 74.960 128.015 75.130 128.235 ;
        RECT 75.285 128.205 80.795 129.015 ;
        RECT 81.735 128.290 82.165 129.075 ;
        RECT 83.980 128.915 84.935 129.115 ;
        RECT 82.655 128.235 84.935 128.915 ;
        RECT 84.945 128.915 85.875 129.115 ;
        RECT 87.210 128.915 88.155 129.115 ;
        RECT 84.945 128.435 88.155 128.915 ;
        RECT 75.425 128.015 75.595 128.205 ;
        RECT 82.780 128.185 82.950 128.235 ;
        RECT 83.980 128.205 84.935 128.235 ;
        RECT 85.085 128.235 88.155 128.435 ;
        RECT 77.730 127.995 77.900 128.185 ;
        RECT 78.185 127.995 78.355 128.185 ;
        RECT 17.325 127.185 18.695 127.995 ;
        RECT 18.705 127.315 20.535 127.995 ;
        RECT 18.705 127.085 20.050 127.315 ;
        RECT 20.545 127.215 21.915 127.995 ;
        RECT 21.925 127.185 24.675 127.995 ;
        RECT 24.685 127.315 31.995 127.995 ;
        RECT 28.200 127.095 29.110 127.315 ;
        RECT 30.645 127.085 31.995 127.315 ;
        RECT 32.055 127.085 33.405 127.995 ;
        RECT 33.425 127.185 38.935 127.995 ;
        RECT 38.945 127.185 42.615 127.995 ;
        RECT 43.095 127.125 43.525 127.910 ;
        RECT 43.545 127.185 49.055 127.995 ;
        RECT 49.065 127.185 54.575 127.995 ;
        RECT 54.585 127.185 60.095 127.995 ;
        RECT 60.105 127.185 63.775 127.995 ;
        RECT 63.785 127.185 65.155 127.995 ;
        RECT 65.185 127.085 66.535 127.995 ;
        RECT 66.855 127.315 68.690 127.995 ;
        RECT 66.855 127.085 67.785 127.315 ;
        RECT 68.855 127.125 69.285 127.910 ;
        RECT 69.305 127.315 76.615 127.995 ;
        RECT 72.820 127.095 73.730 127.315 ;
        RECT 75.265 127.085 76.615 127.315 ;
        RECT 76.665 127.085 78.015 127.995 ;
        RECT 78.045 127.185 79.415 127.995 ;
        RECT 79.565 127.965 79.735 128.185 ;
        RECT 80.955 128.050 81.115 128.160 ;
        RECT 82.320 128.045 82.440 128.155 ;
        RECT 82.780 128.015 82.955 128.185 ;
        RECT 85.085 128.015 85.255 128.235 ;
        RECT 87.210 128.205 88.155 128.235 ;
        RECT 88.165 128.885 89.095 129.115 ;
        RECT 92.305 128.885 93.235 129.115 ;
        RECT 88.165 128.205 92.065 128.885 ;
        RECT 92.305 128.205 96.205 128.885 ;
        RECT 96.445 128.205 100.115 129.015 ;
        RECT 100.585 128.205 104.455 129.115 ;
        RECT 104.725 128.205 107.475 129.115 ;
        RECT 107.495 128.290 107.925 129.075 ;
        RECT 107.945 128.205 109.775 129.015 ;
        RECT 110.340 128.885 111.260 129.115 ;
        RECT 117.440 128.885 118.350 129.105 ;
        RECT 119.885 128.885 121.235 129.115 ;
        RECT 124.800 128.885 125.710 129.105 ;
        RECT 127.245 128.885 128.595 129.115 ;
        RECT 110.340 128.205 113.805 128.885 ;
        RECT 113.925 128.205 121.235 128.885 ;
        RECT 121.285 128.205 128.595 128.885 ;
        RECT 128.645 128.205 130.475 129.015 ;
        RECT 132.305 128.885 133.235 129.115 ;
        RECT 130.485 128.205 133.235 128.885 ;
        RECT 133.255 128.290 133.685 129.075 ;
        RECT 133.705 128.205 136.915 129.115 ;
        RECT 140.900 128.885 141.810 129.105 ;
        RECT 143.345 128.885 144.695 129.115 ;
        RECT 137.385 128.205 144.695 128.885 ;
        RECT 145.665 128.205 147.035 129.015 ;
        RECT 86.015 128.040 86.175 128.150 ;
        RECT 81.690 127.965 82.635 127.995 ;
        RECT 79.565 127.765 82.635 127.965 ;
        RECT 82.785 127.965 82.955 128.015 ;
        RECT 86.925 127.995 87.095 128.185 ;
        RECT 88.580 128.015 88.750 128.205 ;
        RECT 92.720 128.015 92.890 128.205 ;
        RECT 95.205 127.995 95.375 128.185 ;
        RECT 96.585 128.015 96.755 128.205 ;
        RECT 98.895 128.040 99.055 128.150 ;
        RECT 100.260 128.045 100.380 128.155 ;
        RECT 100.730 128.015 100.900 128.205 ;
        RECT 104.865 128.015 105.035 128.205 ;
        RECT 106.705 127.995 106.875 128.185 ;
        RECT 107.165 127.995 107.335 128.185 ;
        RECT 108.085 128.015 108.255 128.205 ;
        RECT 109.920 128.045 110.040 128.155 ;
        RECT 113.605 128.015 113.775 128.205 ;
        RECT 114.065 128.015 114.235 128.205 ;
        RECT 114.525 127.995 114.695 128.185 ;
        RECT 116.360 128.045 116.480 128.155 ;
        RECT 116.825 127.995 116.995 128.185 ;
        RECT 119.595 128.040 119.755 128.150 ;
        RECT 121.425 128.015 121.595 128.205 ;
        RECT 128.785 128.185 128.955 128.205 ;
        RECT 124.185 127.995 124.355 128.185 ;
        RECT 127.865 127.995 128.035 128.185 ;
        RECT 128.320 128.045 128.440 128.155 ;
        RECT 128.775 128.015 128.955 128.185 ;
        RECT 130.625 128.015 130.795 128.205 ;
        RECT 133.835 128.015 134.005 128.205 ;
        RECT 128.775 127.995 128.945 128.015 ;
        RECT 135.410 127.995 135.580 128.185 ;
        RECT 136.145 127.995 136.315 128.185 ;
        RECT 137.060 128.045 137.180 128.155 ;
        RECT 137.525 128.015 137.695 128.205 ;
        RECT 143.500 128.045 143.620 128.155 ;
        RECT 143.965 127.995 144.135 128.185 ;
        RECT 144.895 128.050 145.055 128.160 ;
        RECT 146.725 127.995 146.895 128.205 ;
        RECT 84.910 127.965 85.855 127.995 ;
        RECT 82.785 127.765 85.855 127.965 ;
        RECT 79.425 127.285 82.635 127.765 ;
        RECT 79.425 127.085 80.355 127.285 ;
        RECT 81.690 127.085 82.635 127.285 ;
        RECT 82.645 127.285 85.855 127.765 ;
        RECT 86.785 127.315 94.515 127.995 ;
        RECT 82.645 127.085 83.575 127.285 ;
        RECT 84.910 127.085 85.855 127.285 ;
        RECT 90.300 127.095 91.210 127.315 ;
        RECT 92.745 127.085 94.515 127.315 ;
        RECT 94.615 127.125 95.045 127.910 ;
        RECT 95.065 127.185 98.735 127.995 ;
        RECT 99.705 127.315 107.015 127.995 ;
        RECT 107.025 127.315 114.335 127.995 ;
        RECT 99.705 127.085 101.055 127.315 ;
        RECT 102.590 127.095 103.500 127.315 ;
        RECT 110.540 127.095 111.450 127.315 ;
        RECT 112.985 127.085 114.335 127.315 ;
        RECT 114.385 127.185 116.215 127.995 ;
        RECT 116.685 127.085 119.435 127.995 ;
        RECT 120.375 127.125 120.805 127.910 ;
        RECT 120.920 127.315 124.385 127.995 ;
        RECT 124.600 127.315 128.065 127.995 ;
        RECT 120.920 127.085 121.840 127.315 ;
        RECT 124.600 127.085 125.520 127.315 ;
        RECT 128.645 127.085 131.855 127.995 ;
        RECT 132.095 127.315 135.995 127.995 ;
        RECT 136.005 127.315 143.315 127.995 ;
        RECT 143.825 127.315 145.655 127.995 ;
        RECT 135.065 127.085 135.995 127.315 ;
        RECT 139.520 127.095 140.430 127.315 ;
        RECT 141.965 127.085 143.315 127.315 ;
        RECT 144.310 127.085 145.655 127.315 ;
        RECT 145.665 127.185 147.035 127.995 ;
      LAYER nwell ;
        RECT 17.130 123.965 147.230 126.795 ;
      LAYER pwell ;
        RECT 17.325 122.765 18.695 123.575 ;
        RECT 22.680 123.445 23.590 123.665 ;
        RECT 25.125 123.445 26.475 123.675 ;
        RECT 19.165 122.765 26.475 123.445 ;
        RECT 27.065 122.765 30.065 123.675 ;
        RECT 30.215 122.850 30.645 123.635 ;
        RECT 30.975 123.445 31.905 123.675 ;
        RECT 30.975 122.765 32.810 123.445 ;
        RECT 32.975 122.765 34.325 123.675 ;
        RECT 34.345 122.765 39.855 123.575 ;
        RECT 39.865 122.765 45.375 123.575 ;
        RECT 45.385 122.765 50.895 123.575 ;
        RECT 50.905 122.765 54.575 123.575 ;
        RECT 54.585 122.765 55.955 123.575 ;
        RECT 55.975 122.850 56.405 123.635 ;
        RECT 56.425 122.765 61.935 123.575 ;
        RECT 65.460 123.445 66.370 123.665 ;
        RECT 67.905 123.445 69.675 123.675 ;
        RECT 61.945 122.765 69.675 123.445 ;
        RECT 69.965 123.585 70.915 123.675 ;
        RECT 69.965 122.765 71.895 123.585 ;
        RECT 76.040 123.445 76.950 123.665 ;
        RECT 78.485 123.445 79.835 123.675 ;
        RECT 72.525 122.765 79.835 123.445 ;
        RECT 79.885 122.765 81.715 123.575 ;
        RECT 81.735 122.850 82.165 123.635 ;
        RECT 82.185 122.765 83.555 123.575 ;
        RECT 86.765 123.445 87.695 123.675 ;
        RECT 91.220 123.445 92.130 123.665 ;
        RECT 93.665 123.445 95.435 123.675 ;
        RECT 83.795 122.765 87.695 123.445 ;
        RECT 87.705 122.765 95.435 123.445 ;
        RECT 95.620 123.445 96.540 123.675 ;
        RECT 102.320 123.445 103.240 123.675 ;
        RECT 106.545 123.445 107.475 123.675 ;
        RECT 95.620 122.765 99.085 123.445 ;
        RECT 99.775 122.765 103.240 123.445 ;
        RECT 103.575 122.765 107.475 123.445 ;
        RECT 107.495 122.850 107.925 123.635 ;
        RECT 111.460 123.445 112.370 123.665 ;
        RECT 113.905 123.445 115.255 123.675 ;
        RECT 107.945 122.765 115.255 123.445 ;
        RECT 115.305 122.765 120.815 123.575 ;
        RECT 120.825 122.765 123.575 123.675 ;
        RECT 123.585 122.765 129.095 123.575 ;
        RECT 129.105 122.765 132.775 123.575 ;
        RECT 133.255 122.850 133.685 123.635 ;
        RECT 135.525 123.445 136.455 123.675 ;
        RECT 133.705 122.765 136.455 123.445 ;
        RECT 136.465 122.765 141.975 123.575 ;
        RECT 142.470 123.445 143.815 123.675 ;
        RECT 144.310 123.445 145.655 123.675 ;
        RECT 141.985 122.765 143.815 123.445 ;
        RECT 143.825 122.765 145.655 123.445 ;
        RECT 145.665 122.765 147.035 123.575 ;
        RECT 17.465 122.555 17.635 122.765 ;
        RECT 18.840 122.605 18.960 122.715 ;
        RECT 19.305 122.575 19.475 122.765 ;
        RECT 20.225 122.555 20.395 122.745 ;
        RECT 20.685 122.555 20.855 122.745 ;
        RECT 22.340 122.555 22.510 122.745 ;
        RECT 26.205 122.555 26.375 122.745 ;
        RECT 26.660 122.605 26.780 122.715 ;
        RECT 27.125 122.575 27.295 122.765 ;
        RECT 32.645 122.745 32.810 122.765 ;
        RECT 31.725 122.555 31.895 122.745 ;
        RECT 32.645 122.575 32.815 122.745 ;
        RECT 34.025 122.575 34.195 122.765 ;
        RECT 34.485 122.575 34.655 122.765 ;
        RECT 37.245 122.555 37.415 122.745 ;
        RECT 40.005 122.575 40.175 122.765 ;
        RECT 42.760 122.605 42.880 122.715 ;
        RECT 43.685 122.555 43.855 122.745 ;
        RECT 45.525 122.575 45.695 122.765 ;
        RECT 49.205 122.555 49.375 122.745 ;
        RECT 51.045 122.575 51.215 122.765 ;
        RECT 54.725 122.555 54.895 122.765 ;
        RECT 56.565 122.575 56.735 122.765 ;
        RECT 60.240 122.605 60.360 122.715 ;
        RECT 60.705 122.555 60.875 122.745 ;
        RECT 62.085 122.575 62.255 122.765 ;
        RECT 71.745 122.745 71.895 122.765 ;
        RECT 63.925 122.555 64.095 122.745 ;
        RECT 69.445 122.555 69.615 122.745 ;
        RECT 71.745 122.575 71.915 122.745 ;
        RECT 72.200 122.605 72.320 122.715 ;
        RECT 72.665 122.575 72.835 122.765 ;
        RECT 80.025 122.575 80.195 122.765 ;
        RECT 82.325 122.575 82.495 122.765 ;
        RECT 84.165 122.555 84.335 122.745 ;
        RECT 84.635 122.600 84.795 122.710 ;
        RECT 85.545 122.555 85.715 122.745 ;
        RECT 87.110 122.575 87.280 122.765 ;
        RECT 87.845 122.575 88.015 122.765 ;
        RECT 93.365 122.555 93.535 122.745 ;
        RECT 95.205 122.555 95.375 122.745 ;
        RECT 97.965 122.555 98.135 122.745 ;
        RECT 98.885 122.575 99.055 122.765 ;
        RECT 99.340 122.605 99.460 122.715 ;
        RECT 99.805 122.575 99.975 122.765 ;
        RECT 101.645 122.555 101.815 122.745 ;
        RECT 105.325 122.555 105.495 122.745 ;
        RECT 106.890 122.575 107.060 122.765 ;
        RECT 108.085 122.575 108.255 122.765 ;
        RECT 109.475 122.555 109.645 122.745 ;
        RECT 109.925 122.555 110.095 122.745 ;
        RECT 111.765 122.555 111.935 122.745 ;
        RECT 115.445 122.575 115.615 122.765 ;
        RECT 119.125 122.555 119.295 122.745 ;
        RECT 120.965 122.575 121.135 122.765 ;
        RECT 123.265 122.555 123.435 122.745 ;
        RECT 123.725 122.555 123.895 122.765 ;
        RECT 129.245 122.715 129.415 122.765 ;
        RECT 129.240 122.605 129.415 122.715 ;
        RECT 129.245 122.575 129.415 122.605 ;
        RECT 129.705 122.555 129.875 122.745 ;
        RECT 132.465 122.555 132.635 122.745 ;
        RECT 132.920 122.605 133.040 122.715 ;
        RECT 133.845 122.575 134.015 122.765 ;
        RECT 135.220 122.605 135.340 122.715 ;
        RECT 135.960 122.555 136.130 122.745 ;
        RECT 136.605 122.575 136.775 122.765 ;
        RECT 139.825 122.555 139.995 122.745 ;
        RECT 142.125 122.575 142.295 122.765 ;
        RECT 143.965 122.575 144.135 122.765 ;
        RECT 145.340 122.605 145.460 122.715 ;
        RECT 146.725 122.555 146.895 122.765 ;
        RECT 17.325 121.745 18.695 122.555 ;
        RECT 18.705 121.875 20.535 122.555 ;
        RECT 18.705 121.645 20.050 121.875 ;
        RECT 20.545 121.745 21.915 122.555 ;
        RECT 21.925 121.875 25.825 122.555 ;
        RECT 21.925 121.645 22.855 121.875 ;
        RECT 26.065 121.745 31.575 122.555 ;
        RECT 31.585 121.745 37.095 122.555 ;
        RECT 37.105 121.745 42.615 122.555 ;
        RECT 43.095 121.685 43.525 122.470 ;
        RECT 43.545 121.745 49.055 122.555 ;
        RECT 49.065 121.745 54.575 122.555 ;
        RECT 54.585 121.745 60.095 122.555 ;
        RECT 60.615 121.645 63.775 122.555 ;
        RECT 63.785 121.875 68.600 122.555 ;
        RECT 68.855 121.685 69.285 122.470 ;
        RECT 69.305 121.875 77.035 122.555 ;
        RECT 72.820 121.655 73.730 121.875 ;
        RECT 75.265 121.645 77.035 121.875 ;
        RECT 77.165 121.875 84.475 122.555 ;
        RECT 85.405 121.875 93.135 122.555 ;
        RECT 77.165 121.645 78.515 121.875 ;
        RECT 80.050 121.655 80.960 121.875 ;
        RECT 88.920 121.655 89.830 121.875 ;
        RECT 91.365 121.645 93.135 121.875 ;
        RECT 93.225 121.745 94.595 122.555 ;
        RECT 94.615 121.685 95.045 122.470 ;
        RECT 95.065 121.745 97.815 122.555 ;
        RECT 97.935 121.875 101.400 122.555 ;
        RECT 100.480 121.645 101.400 121.875 ;
        RECT 101.505 121.745 105.175 122.555 ;
        RECT 105.185 121.745 106.555 122.555 ;
        RECT 106.565 121.645 109.775 122.555 ;
        RECT 109.785 121.745 111.615 122.555 ;
        RECT 111.625 121.875 118.935 122.555 ;
        RECT 115.140 121.655 116.050 121.875 ;
        RECT 117.585 121.645 118.935 121.875 ;
        RECT 118.985 121.745 120.355 122.555 ;
        RECT 120.375 121.685 120.805 122.470 ;
        RECT 120.825 121.875 123.575 122.555 ;
        RECT 120.825 121.645 121.755 121.875 ;
        RECT 123.585 121.745 129.095 122.555 ;
        RECT 129.565 121.875 132.315 122.555 ;
        RECT 131.385 121.645 132.315 121.875 ;
        RECT 132.325 121.745 135.075 122.555 ;
        RECT 135.545 121.875 139.445 122.555 ;
        RECT 135.545 121.645 136.475 121.875 ;
        RECT 139.685 121.745 145.195 122.555 ;
        RECT 145.665 121.745 147.035 122.555 ;
      LAYER nwell ;
        RECT 17.130 118.525 147.230 121.355 ;
      LAYER pwell ;
        RECT 17.325 117.325 18.695 118.135 ;
        RECT 18.705 118.005 20.050 118.235 ;
        RECT 20.545 118.005 21.890 118.235 ;
        RECT 18.705 117.325 20.535 118.005 ;
        RECT 20.545 117.325 22.375 118.005 ;
        RECT 22.385 117.325 26.055 118.135 ;
        RECT 27.115 118.005 28.045 118.235 ;
        RECT 26.210 117.325 28.045 118.005 ;
        RECT 28.365 117.325 30.195 118.135 ;
        RECT 30.215 117.410 30.645 118.195 ;
        RECT 30.665 117.325 36.175 118.135 ;
        RECT 36.185 117.325 41.695 118.135 ;
        RECT 41.705 117.325 47.215 118.135 ;
        RECT 47.225 117.325 52.735 118.135 ;
        RECT 52.745 117.325 55.495 118.135 ;
        RECT 55.975 117.410 56.405 118.195 ;
        RECT 56.425 117.325 61.935 118.135 ;
        RECT 61.945 117.325 64.695 118.135 ;
        RECT 64.705 118.005 65.635 118.235 ;
        RECT 64.705 117.325 68.605 118.005 ;
        RECT 68.845 117.325 71.595 118.135 ;
        RECT 71.605 118.005 72.535 118.235 ;
        RECT 71.605 117.325 75.505 118.005 ;
        RECT 75.745 117.325 81.255 118.135 ;
        RECT 81.735 117.410 82.165 118.195 ;
        RECT 82.185 118.005 83.115 118.235 ;
        RECT 82.185 117.325 86.085 118.005 ;
        RECT 86.325 117.325 89.995 118.135 ;
        RECT 90.005 117.325 91.375 118.135 ;
        RECT 96.445 118.005 97.375 118.235 ;
        RECT 100.585 118.005 101.515 118.235 ;
        RECT 91.620 117.325 96.435 118.005 ;
        RECT 96.445 117.325 100.345 118.005 ;
        RECT 100.585 117.325 104.485 118.005 ;
        RECT 104.725 117.325 107.475 118.135 ;
        RECT 107.495 117.410 107.925 118.195 ;
        RECT 110.685 118.005 111.615 118.235 ;
        RECT 108.865 117.325 111.615 118.005 ;
        RECT 111.625 118.005 112.555 118.235 ;
        RECT 111.625 117.325 115.525 118.005 ;
        RECT 115.765 117.325 117.595 118.135 ;
        RECT 117.605 117.325 120.815 118.235 ;
        RECT 124.340 118.005 125.250 118.225 ;
        RECT 126.785 118.005 128.135 118.235 ;
        RECT 120.825 117.325 128.135 118.005 ;
        RECT 128.185 117.325 130.015 118.135 ;
        RECT 132.305 118.005 133.235 118.235 ;
        RECT 130.485 117.325 133.235 118.005 ;
        RECT 133.255 117.410 133.685 118.195 ;
        RECT 133.705 117.325 136.915 118.235 ;
        RECT 140.900 118.005 141.810 118.225 ;
        RECT 143.345 118.005 144.695 118.235 ;
        RECT 137.385 117.325 144.695 118.005 ;
        RECT 145.665 117.325 147.035 118.135 ;
        RECT 17.465 117.115 17.635 117.325 ;
        RECT 18.855 117.160 19.015 117.270 ;
        RECT 19.765 117.115 19.935 117.305 ;
        RECT 20.225 117.135 20.395 117.325 ;
        RECT 21.605 117.115 21.775 117.305 ;
        RECT 22.065 117.135 22.235 117.325 ;
        RECT 22.525 117.135 22.695 117.325 ;
        RECT 26.210 117.305 26.375 117.325 ;
        RECT 26.205 117.135 26.375 117.305 ;
        RECT 28.505 117.135 28.675 117.325 ;
        RECT 29.885 117.115 30.055 117.305 ;
        RECT 30.345 117.115 30.515 117.305 ;
        RECT 30.805 117.135 30.975 117.325 ;
        RECT 34.485 117.115 34.655 117.305 ;
        RECT 36.325 117.135 36.495 117.325 ;
        RECT 40.005 117.115 40.175 117.305 ;
        RECT 41.845 117.135 42.015 117.325 ;
        RECT 42.760 117.165 42.880 117.275 ;
        RECT 43.685 117.115 43.855 117.305 ;
        RECT 47.365 117.135 47.535 117.325 ;
        RECT 49.205 117.115 49.375 117.305 ;
        RECT 52.885 117.135 53.055 117.325 ;
        RECT 54.725 117.115 54.895 117.305 ;
        RECT 55.640 117.165 55.760 117.275 ;
        RECT 56.565 117.135 56.735 117.325 ;
        RECT 60.245 117.115 60.415 117.305 ;
        RECT 62.085 117.135 62.255 117.325 ;
        RECT 65.120 117.135 65.290 117.325 ;
        RECT 65.765 117.115 65.935 117.305 ;
        RECT 68.520 117.165 68.640 117.275 ;
        RECT 68.985 117.135 69.155 117.325 ;
        RECT 69.445 117.115 69.615 117.305 ;
        RECT 72.020 117.135 72.190 117.325 ;
        RECT 74.965 117.115 75.135 117.305 ;
        RECT 75.885 117.135 76.055 117.325 ;
        RECT 80.485 117.115 80.655 117.305 ;
        RECT 81.400 117.165 81.520 117.275 ;
        RECT 82.600 117.135 82.770 117.325 ;
        RECT 86.015 117.160 86.175 117.270 ;
        RECT 86.465 117.135 86.635 117.325 ;
        RECT 86.925 117.115 87.095 117.305 ;
        RECT 89.685 117.115 89.855 117.305 ;
        RECT 90.145 117.135 90.315 117.325 ;
        RECT 95.205 117.115 95.375 117.305 ;
        RECT 96.125 117.135 96.295 117.325 ;
        RECT 96.860 117.135 97.030 117.325 ;
        RECT 101.000 117.135 101.170 117.325 ;
        RECT 103.940 117.115 104.110 117.305 ;
        RECT 104.405 117.115 104.575 117.305 ;
        RECT 104.865 117.135 105.035 117.325 ;
        RECT 108.095 117.170 108.255 117.280 ;
        RECT 109.005 117.135 109.175 117.325 ;
        RECT 109.925 117.115 110.095 117.305 ;
        RECT 112.040 117.135 112.210 117.325 ;
        RECT 113.600 117.165 113.720 117.275 ;
        RECT 114.340 117.115 114.510 117.305 ;
        RECT 115.905 117.135 116.075 117.325 ;
        RECT 117.735 117.135 117.905 117.325 ;
        RECT 118.205 117.115 118.375 117.305 ;
        RECT 120.040 117.165 120.160 117.275 ;
        RECT 120.965 117.135 121.135 117.325 ;
        RECT 121.885 117.115 122.055 117.305 ;
        RECT 127.220 117.115 127.390 117.305 ;
        RECT 128.325 117.135 128.495 117.325 ;
        RECT 130.160 117.165 130.280 117.275 ;
        RECT 130.625 117.135 130.795 117.325 ;
        RECT 131.085 117.115 131.255 117.305 ;
        RECT 132.465 117.115 132.635 117.305 ;
        RECT 133.835 117.135 134.005 117.325 ;
        RECT 137.060 117.165 137.180 117.275 ;
        RECT 137.525 117.135 137.695 117.325 ;
        RECT 139.825 117.115 139.995 117.305 ;
        RECT 141.660 117.165 141.780 117.275 ;
        RECT 142.125 117.115 142.295 117.305 ;
        RECT 143.965 117.115 144.135 117.305 ;
        RECT 144.895 117.170 145.055 117.280 ;
        RECT 146.725 117.115 146.895 117.325 ;
        RECT 17.325 116.305 18.695 117.115 ;
        RECT 19.625 116.435 21.455 117.115 ;
        RECT 21.465 116.305 22.835 117.115 ;
        RECT 22.885 116.435 30.195 117.115 ;
        RECT 22.885 116.205 24.235 116.435 ;
        RECT 25.770 116.215 26.680 116.435 ;
        RECT 30.205 116.205 34.265 117.115 ;
        RECT 34.345 116.305 39.855 117.115 ;
        RECT 39.865 116.305 42.615 117.115 ;
        RECT 43.095 116.245 43.525 117.030 ;
        RECT 43.545 116.305 49.055 117.115 ;
        RECT 49.065 116.305 54.575 117.115 ;
        RECT 54.585 116.305 60.095 117.115 ;
        RECT 60.105 116.305 65.615 117.115 ;
        RECT 65.625 116.305 68.375 117.115 ;
        RECT 68.855 116.245 69.285 117.030 ;
        RECT 69.305 116.305 74.815 117.115 ;
        RECT 74.825 116.305 80.335 117.115 ;
        RECT 80.345 116.305 85.855 117.115 ;
        RECT 86.785 116.305 88.875 117.115 ;
        RECT 89.545 116.435 94.360 117.115 ;
        RECT 94.615 116.245 95.045 117.030 ;
        RECT 95.065 116.435 102.375 117.115 ;
        RECT 98.580 116.215 99.490 116.435 ;
        RECT 101.025 116.205 102.375 116.435 ;
        RECT 102.485 116.205 104.255 117.115 ;
        RECT 104.265 116.305 109.775 117.115 ;
        RECT 109.785 116.305 113.455 117.115 ;
        RECT 113.925 116.435 117.825 117.115 ;
        RECT 113.925 116.205 114.855 116.435 ;
        RECT 118.065 116.305 119.895 117.115 ;
        RECT 120.375 116.245 120.805 117.030 ;
        RECT 121.745 116.435 126.560 117.115 ;
        RECT 126.805 116.435 130.705 117.115 ;
        RECT 126.805 116.205 127.735 116.435 ;
        RECT 130.945 116.305 132.315 117.115 ;
        RECT 132.325 116.435 139.635 117.115 ;
        RECT 135.840 116.215 136.750 116.435 ;
        RECT 138.285 116.205 139.635 116.435 ;
        RECT 139.685 116.305 141.515 117.115 ;
        RECT 141.985 116.435 143.815 117.115 ;
        RECT 143.825 116.435 145.655 117.115 ;
        RECT 142.470 116.205 143.815 116.435 ;
        RECT 144.310 116.205 145.655 116.435 ;
        RECT 145.665 116.305 147.035 117.115 ;
      LAYER nwell ;
        RECT 17.130 113.085 147.230 115.915 ;
      LAYER pwell ;
        RECT 17.325 111.885 18.695 112.695 ;
        RECT 22.680 112.565 23.590 112.785 ;
        RECT 25.125 112.565 26.475 112.795 ;
        RECT 19.165 111.885 26.475 112.565 ;
        RECT 26.985 112.565 28.350 112.795 ;
        RECT 26.985 111.885 30.195 112.565 ;
        RECT 30.215 111.970 30.645 112.755 ;
        RECT 34.180 112.565 35.090 112.785 ;
        RECT 36.625 112.565 37.975 112.795 ;
        RECT 30.665 111.885 37.975 112.565 ;
        RECT 38.025 111.885 43.535 112.695 ;
        RECT 43.545 111.885 49.055 112.695 ;
        RECT 49.065 111.885 54.575 112.695 ;
        RECT 54.585 111.885 55.955 112.695 ;
        RECT 55.975 111.970 56.405 112.755 ;
        RECT 56.425 111.885 61.935 112.695 ;
        RECT 61.945 111.885 67.455 112.695 ;
        RECT 67.465 111.885 72.975 112.695 ;
        RECT 72.985 111.885 78.495 112.695 ;
        RECT 78.505 111.885 81.255 112.695 ;
        RECT 81.735 111.970 82.165 112.755 ;
        RECT 82.185 111.885 85.855 112.695 ;
        RECT 88.605 112.565 89.535 112.795 ;
        RECT 86.785 111.885 89.535 112.565 ;
        RECT 90.665 111.885 92.755 112.695 ;
        RECT 96.740 112.565 97.650 112.785 ;
        RECT 99.185 112.565 100.535 112.795 ;
        RECT 93.225 111.885 100.535 112.565 ;
        RECT 100.585 112.115 105.175 112.795 ;
        RECT 101.545 111.885 105.175 112.115 ;
        RECT 105.185 111.885 107.015 112.565 ;
        RECT 107.495 111.970 107.925 112.755 ;
        RECT 107.945 111.885 111.155 112.795 ;
        RECT 111.165 111.885 112.995 112.695 ;
        RECT 116.980 112.565 117.890 112.785 ;
        RECT 119.425 112.565 120.775 112.795 ;
        RECT 113.465 111.885 120.775 112.565 ;
        RECT 120.825 111.885 125.640 112.565 ;
        RECT 125.885 111.885 129.555 112.695 ;
        RECT 129.565 111.885 133.220 112.795 ;
        RECT 133.255 111.970 133.685 112.755 ;
        RECT 133.705 112.565 134.635 112.795 ;
        RECT 133.705 111.885 137.605 112.565 ;
        RECT 137.845 111.885 141.515 112.695 ;
        RECT 142.470 112.565 143.815 112.795 ;
        RECT 144.310 112.565 145.655 112.795 ;
        RECT 141.985 111.885 143.815 112.565 ;
        RECT 143.825 111.885 145.655 112.565 ;
        RECT 145.665 111.885 147.035 112.695 ;
        RECT 17.465 111.675 17.635 111.885 ;
        RECT 18.855 111.835 19.025 111.865 ;
        RECT 18.840 111.725 19.025 111.835 ;
        RECT 18.855 111.675 19.025 111.725 ;
        RECT 19.305 111.695 19.475 111.885 ;
        RECT 20.235 111.675 20.405 111.865 ;
        RECT 21.880 111.675 22.050 111.865 ;
        RECT 25.740 111.725 25.860 111.835 ;
        RECT 26.205 111.675 26.375 111.865 ;
        RECT 26.660 111.725 26.780 111.835 ;
        RECT 29.880 111.695 30.050 111.885 ;
        RECT 30.805 111.695 30.975 111.885 ;
        RECT 33.570 111.675 33.740 111.865 ;
        RECT 36.785 111.675 36.955 111.865 ;
        RECT 38.165 111.695 38.335 111.885 ;
        RECT 42.315 111.720 42.475 111.830 ;
        RECT 43.685 111.675 43.855 111.885 ;
        RECT 49.205 111.675 49.375 111.885 ;
        RECT 54.725 111.675 54.895 111.885 ;
        RECT 56.565 111.695 56.735 111.885 ;
        RECT 60.245 111.675 60.415 111.865 ;
        RECT 62.085 111.695 62.255 111.885 ;
        RECT 65.765 111.675 65.935 111.865 ;
        RECT 67.605 111.695 67.775 111.885 ;
        RECT 68.520 111.725 68.640 111.835 ;
        RECT 69.445 111.675 69.615 111.865 ;
        RECT 73.125 111.695 73.295 111.885 ;
        RECT 74.045 111.675 74.215 111.865 ;
        RECT 76.805 111.675 76.975 111.865 ;
        RECT 78.460 111.675 78.630 111.865 ;
        RECT 78.645 111.695 78.815 111.885 ;
        RECT 81.400 111.725 81.520 111.835 ;
        RECT 82.325 111.675 82.495 111.885 ;
        RECT 84.160 111.725 84.280 111.835 ;
        RECT 84.900 111.675 85.070 111.865 ;
        RECT 86.015 111.730 86.175 111.840 ;
        RECT 86.925 111.695 87.095 111.885 ;
        RECT 88.765 111.675 88.935 111.865 ;
        RECT 89.680 111.725 89.800 111.835 ;
        RECT 90.610 111.675 90.780 111.865 ;
        RECT 92.445 111.695 92.615 111.885 ;
        RECT 92.900 111.725 93.020 111.835 ;
        RECT 93.365 111.695 93.535 111.885 ;
        RECT 95.215 111.720 95.375 111.830 ;
        RECT 97.505 111.675 97.675 111.865 ;
        RECT 97.970 111.675 98.140 111.865 ;
        RECT 102.565 111.695 102.735 111.865 ;
        RECT 104.860 111.695 105.030 111.885 ;
        RECT 106.705 111.695 106.875 111.885 ;
        RECT 107.160 111.725 107.280 111.835 ;
        RECT 108.075 111.695 108.245 111.885 ;
        RECT 102.595 111.675 102.735 111.695 ;
        RECT 111.030 111.675 111.200 111.865 ;
        RECT 111.305 111.695 111.475 111.885 ;
        RECT 111.775 111.720 111.935 111.830 ;
        RECT 112.685 111.675 112.855 111.865 ;
        RECT 113.140 111.725 113.260 111.835 ;
        RECT 113.605 111.695 113.775 111.885 ;
        RECT 115.445 111.675 115.615 111.865 ;
        RECT 119.125 111.675 119.295 111.865 ;
        RECT 120.965 111.835 121.135 111.885 ;
        RECT 120.960 111.725 121.135 111.835 ;
        RECT 120.965 111.695 121.135 111.725 ;
        RECT 121.425 111.675 121.595 111.865 ;
        RECT 126.025 111.695 126.195 111.885 ;
        RECT 129.060 111.675 129.230 111.865 ;
        RECT 129.710 111.695 129.880 111.885 ;
        RECT 132.925 111.675 133.095 111.865 ;
        RECT 134.120 111.695 134.290 111.885 ;
        RECT 134.765 111.675 134.935 111.865 ;
        RECT 137.525 111.675 137.695 111.865 ;
        RECT 137.985 111.695 138.155 111.885 ;
        RECT 141.660 111.725 141.780 111.835 ;
        RECT 142.125 111.695 142.295 111.885 ;
        RECT 143.965 111.695 144.135 111.885 ;
        RECT 144.895 111.720 145.055 111.830 ;
        RECT 146.725 111.675 146.895 111.885 ;
        RECT 17.325 110.865 18.695 111.675 ;
        RECT 18.705 110.895 20.075 111.675 ;
        RECT 20.085 110.895 21.455 111.675 ;
        RECT 21.465 110.995 25.365 111.675 ;
        RECT 26.065 110.995 33.375 111.675 ;
        RECT 33.425 110.995 36.635 111.675 ;
        RECT 21.465 110.765 22.395 110.995 ;
        RECT 29.580 110.775 30.490 110.995 ;
        RECT 32.025 110.765 33.375 110.995 ;
        RECT 35.270 110.765 36.635 110.995 ;
        RECT 36.645 110.865 42.155 111.675 ;
        RECT 43.095 110.805 43.525 111.590 ;
        RECT 43.545 110.865 49.055 111.675 ;
        RECT 49.065 110.865 54.575 111.675 ;
        RECT 54.585 110.865 60.095 111.675 ;
        RECT 60.105 110.865 65.615 111.675 ;
        RECT 65.625 110.865 68.375 111.675 ;
        RECT 68.855 110.805 69.285 111.590 ;
        RECT 69.305 110.865 72.975 111.675 ;
        RECT 73.905 110.995 76.655 111.675 ;
        RECT 75.725 110.765 76.655 110.995 ;
        RECT 76.665 110.865 78.035 111.675 ;
        RECT 78.045 110.995 81.945 111.675 ;
        RECT 78.045 110.765 78.975 110.995 ;
        RECT 82.185 110.865 84.015 111.675 ;
        RECT 84.485 110.995 88.385 111.675 ;
        RECT 84.485 110.765 85.415 110.995 ;
        RECT 88.625 110.865 90.455 111.675 ;
        RECT 90.465 110.765 94.335 111.675 ;
        RECT 94.615 110.805 95.045 111.590 ;
        RECT 95.985 110.995 97.815 111.675 ;
        RECT 97.825 111.445 101.455 111.675 ;
        RECT 102.595 111.445 106.365 111.675 ;
        RECT 95.985 110.765 97.330 110.995 ;
        RECT 97.825 110.765 102.415 111.445 ;
        RECT 102.595 110.765 106.945 111.445 ;
        RECT 107.715 110.995 111.615 111.675 ;
        RECT 112.545 110.995 115.295 111.675 ;
        RECT 110.685 110.765 111.615 110.995 ;
        RECT 114.365 110.765 115.295 110.995 ;
        RECT 115.305 110.865 118.975 111.675 ;
        RECT 118.985 110.865 120.355 111.675 ;
        RECT 120.375 110.805 120.805 111.590 ;
        RECT 121.285 110.995 128.595 111.675 ;
        RECT 124.800 110.775 125.710 110.995 ;
        RECT 127.245 110.765 128.595 110.995 ;
        RECT 128.645 110.995 132.545 111.675 ;
        RECT 128.645 110.765 129.575 110.995 ;
        RECT 132.785 110.865 134.615 111.675 ;
        RECT 134.625 110.995 137.375 111.675 ;
        RECT 137.385 110.995 144.695 111.675 ;
        RECT 136.445 110.765 137.375 110.995 ;
        RECT 140.900 110.775 141.810 110.995 ;
        RECT 143.345 110.765 144.695 110.995 ;
        RECT 145.665 110.865 147.035 111.675 ;
      LAYER nwell ;
        RECT 17.130 107.645 147.230 110.475 ;
      LAYER pwell ;
        RECT 17.325 106.445 18.695 107.255 ;
        RECT 18.705 106.445 24.215 107.255 ;
        RECT 24.225 106.445 27.895 107.255 ;
        RECT 28.845 106.445 30.195 107.355 ;
        RECT 30.215 106.530 30.645 107.315 ;
        RECT 30.665 106.445 36.175 107.255 ;
        RECT 36.185 106.445 41.695 107.255 ;
        RECT 41.705 106.445 47.215 107.255 ;
        RECT 47.225 106.445 52.735 107.255 ;
        RECT 52.745 106.445 55.495 107.255 ;
        RECT 55.975 106.530 56.405 107.315 ;
        RECT 56.425 106.445 61.935 107.255 ;
        RECT 61.945 106.445 67.455 107.255 ;
        RECT 67.465 106.445 71.135 107.255 ;
        RECT 72.965 107.125 73.895 107.355 ;
        RECT 77.420 107.125 78.330 107.345 ;
        RECT 79.865 107.125 81.215 107.355 ;
        RECT 71.145 106.445 73.895 107.125 ;
        RECT 73.905 106.445 81.215 107.125 ;
        RECT 81.735 106.530 82.165 107.315 ;
        RECT 85.700 107.125 86.610 107.345 ;
        RECT 88.145 107.125 89.495 107.355 ;
        RECT 82.185 106.445 89.495 107.125 ;
        RECT 90.465 107.125 91.395 107.355 ;
        RECT 90.465 106.445 94.365 107.125 ;
        RECT 94.605 106.445 98.475 107.355 ;
        RECT 99.005 106.445 102.875 107.355 ;
        RECT 103.345 107.125 104.275 107.355 ;
        RECT 103.345 106.445 107.245 107.125 ;
        RECT 107.495 106.530 107.925 107.315 ;
        RECT 107.985 107.125 109.335 107.355 ;
        RECT 110.870 107.125 111.780 107.345 ;
        RECT 107.985 106.445 115.295 107.125 ;
        RECT 115.305 106.445 120.815 107.255 ;
        RECT 123.105 107.125 124.035 107.355 ;
        RECT 121.285 106.445 124.035 107.125 ;
        RECT 124.045 107.125 124.975 107.355 ;
        RECT 124.045 106.445 126.795 107.125 ;
        RECT 126.805 106.445 132.315 107.255 ;
        RECT 133.255 106.530 133.685 107.315 ;
        RECT 133.705 106.445 136.455 107.255 ;
        RECT 136.465 107.125 137.395 107.355 ;
        RECT 136.465 106.445 140.365 107.125 ;
        RECT 140.620 106.445 144.275 107.355 ;
        RECT 144.285 106.445 145.655 107.255 ;
        RECT 145.665 106.445 147.035 107.255 ;
        RECT 17.465 106.235 17.635 106.445 ;
        RECT 18.845 106.255 19.015 106.445 ;
        RECT 20.225 106.235 20.395 106.425 ;
        RECT 20.685 106.235 20.855 106.425 ;
        RECT 24.365 106.255 24.535 106.445 ;
        RECT 25.930 106.235 26.100 106.425 ;
        RECT 26.660 106.285 26.780 106.395 ;
        RECT 27.125 106.235 27.295 106.425 ;
        RECT 28.055 106.290 28.215 106.400 ;
        RECT 29.880 106.255 30.050 106.445 ;
        RECT 30.805 106.255 30.975 106.445 ;
        RECT 34.485 106.235 34.655 106.425 ;
        RECT 36.325 106.255 36.495 106.445 ;
        RECT 40.005 106.235 40.175 106.425 ;
        RECT 41.845 106.255 42.015 106.445 ;
        RECT 42.760 106.285 42.880 106.395 ;
        RECT 43.685 106.235 43.855 106.425 ;
        RECT 47.365 106.255 47.535 106.445 ;
        RECT 49.205 106.235 49.375 106.425 ;
        RECT 52.885 106.255 53.055 106.445 ;
        RECT 54.725 106.235 54.895 106.425 ;
        RECT 55.640 106.285 55.760 106.395 ;
        RECT 56.565 106.255 56.735 106.445 ;
        RECT 60.245 106.235 60.415 106.425 ;
        RECT 62.085 106.255 62.255 106.445 ;
        RECT 65.765 106.235 65.935 106.425 ;
        RECT 67.605 106.255 67.775 106.445 ;
        RECT 68.520 106.285 68.640 106.395 ;
        RECT 69.445 106.235 69.615 106.425 ;
        RECT 71.285 106.235 71.455 106.445 ;
        RECT 74.045 106.255 74.215 106.445 ;
        RECT 78.920 106.235 79.090 106.425 ;
        RECT 81.400 106.285 81.520 106.395 ;
        RECT 82.325 106.255 82.495 106.445 ;
        RECT 82.790 106.235 82.960 106.425 ;
        RECT 86.460 106.285 86.580 106.395 ;
        RECT 86.925 106.235 87.095 106.425 ;
        RECT 89.695 106.290 89.855 106.400 ;
        RECT 90.880 106.255 91.050 106.445 ;
        RECT 94.280 106.285 94.400 106.395 ;
        RECT 94.750 106.255 94.920 106.445 ;
        RECT 102.560 106.425 102.730 106.445 ;
        RECT 98.880 106.235 99.050 106.425 ;
        RECT 99.345 106.235 99.515 106.425 ;
        RECT 102.105 106.235 102.275 106.425 ;
        RECT 102.560 106.255 102.735 106.425 ;
        RECT 103.020 106.285 103.140 106.395 ;
        RECT 103.760 106.255 103.930 106.445 ;
        RECT 102.565 106.235 102.735 106.255 ;
        RECT 109.925 106.235 110.095 106.425 ;
        RECT 113.145 106.235 113.315 106.425 ;
        RECT 114.985 106.255 115.155 106.445 ;
        RECT 115.445 106.255 115.615 106.445 ;
        RECT 118.665 106.235 118.835 106.425 ;
        RECT 120.965 106.395 121.135 106.425 ;
        RECT 120.960 106.285 121.135 106.395 ;
        RECT 120.965 106.235 121.135 106.285 ;
        RECT 121.425 106.255 121.595 106.445 ;
        RECT 122.345 106.235 122.515 106.425 ;
        RECT 126.485 106.255 126.655 106.445 ;
        RECT 126.945 106.255 127.115 106.445 ;
        RECT 129.980 106.235 130.150 106.425 ;
        RECT 132.475 106.290 132.635 106.400 ;
        RECT 133.845 106.235 134.015 106.445 ;
        RECT 135.960 106.235 136.130 106.425 ;
        RECT 136.880 106.255 137.050 106.445 ;
        RECT 143.960 106.425 144.130 106.445 ;
        RECT 140.100 106.235 140.270 106.425 ;
        RECT 143.960 106.255 144.135 106.425 ;
        RECT 144.425 106.255 144.595 106.445 ;
        RECT 143.965 106.235 144.135 106.255 ;
        RECT 146.725 106.235 146.895 106.445 ;
        RECT 17.325 105.425 18.695 106.235 ;
        RECT 18.705 105.555 20.535 106.235 ;
        RECT 18.705 105.325 20.050 105.555 ;
        RECT 20.545 105.425 22.375 106.235 ;
        RECT 22.615 105.555 26.515 106.235 ;
        RECT 26.985 105.555 34.295 106.235 ;
        RECT 25.585 105.325 26.515 105.555 ;
        RECT 30.500 105.335 31.410 105.555 ;
        RECT 32.945 105.325 34.295 105.555 ;
        RECT 34.345 105.425 39.855 106.235 ;
        RECT 39.865 105.425 42.615 106.235 ;
        RECT 43.095 105.365 43.525 106.150 ;
        RECT 43.545 105.425 49.055 106.235 ;
        RECT 49.065 105.425 54.575 106.235 ;
        RECT 54.585 105.425 60.095 106.235 ;
        RECT 60.105 105.425 65.615 106.235 ;
        RECT 65.625 105.425 68.375 106.235 ;
        RECT 68.855 105.365 69.285 106.150 ;
        RECT 69.305 105.425 71.135 106.235 ;
        RECT 71.145 105.555 78.455 106.235 ;
        RECT 74.660 105.335 75.570 105.555 ;
        RECT 77.105 105.325 78.455 105.555 ;
        RECT 78.505 105.555 82.405 106.235 ;
        RECT 78.505 105.325 79.435 105.555 ;
        RECT 82.645 105.325 86.300 106.235 ;
        RECT 86.785 105.555 94.095 106.235 ;
        RECT 90.300 105.335 91.210 105.555 ;
        RECT 92.745 105.325 94.095 105.555 ;
        RECT 94.615 105.365 95.045 106.150 ;
        RECT 95.325 105.325 99.195 106.235 ;
        RECT 99.205 105.425 100.575 106.235 ;
        RECT 100.585 105.555 102.415 106.235 ;
        RECT 102.425 105.555 109.735 106.235 ;
        RECT 105.940 105.335 106.850 105.555 ;
        RECT 108.385 105.325 109.735 105.555 ;
        RECT 109.785 105.325 112.995 106.235 ;
        RECT 113.005 105.425 118.515 106.235 ;
        RECT 118.525 105.425 120.355 106.235 ;
        RECT 120.375 105.365 120.805 106.150 ;
        RECT 120.825 105.425 122.195 106.235 ;
        RECT 122.205 105.555 129.515 106.235 ;
        RECT 125.720 105.335 126.630 105.555 ;
        RECT 128.165 105.325 129.515 105.555 ;
        RECT 129.565 105.555 133.465 106.235 ;
        RECT 129.565 105.325 130.495 105.555 ;
        RECT 133.705 105.425 135.535 106.235 ;
        RECT 135.545 105.555 139.445 106.235 ;
        RECT 139.685 105.555 143.585 106.235 ;
        RECT 143.825 105.555 145.655 106.235 ;
        RECT 135.545 105.325 136.475 105.555 ;
        RECT 139.685 105.325 140.615 105.555 ;
        RECT 144.310 105.325 145.655 105.555 ;
        RECT 145.665 105.425 147.035 106.235 ;
      LAYER nwell ;
        RECT 17.130 102.205 147.230 105.035 ;
      LAYER pwell ;
        RECT 17.325 101.005 18.695 101.815 ;
        RECT 19.205 101.685 20.555 101.915 ;
        RECT 22.090 101.685 23.000 101.905 ;
        RECT 19.205 101.005 26.515 101.685 ;
        RECT 26.525 101.005 30.195 101.815 ;
        RECT 30.215 101.090 30.645 101.875 ;
        RECT 30.665 101.685 31.595 101.915 ;
        RECT 30.665 101.005 34.565 101.685 ;
        RECT 34.805 101.005 40.315 101.815 ;
        RECT 40.325 101.005 45.835 101.815 ;
        RECT 45.845 101.005 51.355 101.815 ;
        RECT 51.365 101.005 55.035 101.815 ;
        RECT 55.975 101.090 56.405 101.875 ;
        RECT 56.425 101.005 61.935 101.815 ;
        RECT 61.945 101.005 63.315 101.815 ;
        RECT 66.840 101.685 67.750 101.905 ;
        RECT 69.285 101.685 70.635 101.915 ;
        RECT 63.325 101.005 70.635 101.685 ;
        RECT 70.685 101.685 71.615 101.915 ;
        RECT 70.685 101.005 74.585 101.685 ;
        RECT 74.825 101.005 80.335 101.815 ;
        RECT 80.345 101.005 81.715 101.815 ;
        RECT 81.735 101.090 82.165 101.875 ;
        RECT 84.005 101.685 84.935 101.915 ;
        RECT 82.185 101.005 84.935 101.685 ;
        RECT 84.945 101.005 88.615 101.815 ;
        RECT 88.625 101.005 91.835 101.915 ;
        RECT 91.845 101.005 97.355 101.815 ;
        RECT 97.365 101.005 102.875 101.815 ;
        RECT 102.885 101.685 103.815 101.915 ;
        RECT 102.885 101.005 105.635 101.685 ;
        RECT 105.645 101.005 107.475 101.815 ;
        RECT 107.495 101.090 107.925 101.875 ;
        RECT 109.765 101.685 110.695 101.915 ;
        RECT 107.945 101.005 110.695 101.685 ;
        RECT 110.705 101.005 112.535 101.815 ;
        RECT 116.205 101.685 117.135 101.915 ;
        RECT 120.660 101.685 121.570 101.905 ;
        RECT 123.105 101.685 124.455 101.915 ;
        RECT 113.235 101.005 117.135 101.685 ;
        RECT 117.145 101.005 124.455 101.685 ;
        RECT 124.505 101.005 130.015 101.815 ;
        RECT 132.305 101.685 133.235 101.915 ;
        RECT 130.485 101.005 133.235 101.685 ;
        RECT 133.255 101.090 133.685 101.875 ;
        RECT 133.705 101.005 135.535 101.815 ;
        RECT 139.520 101.685 140.430 101.905 ;
        RECT 141.965 101.685 143.315 101.915 ;
        RECT 144.310 101.685 145.655 101.915 ;
        RECT 136.005 101.005 143.315 101.685 ;
        RECT 143.825 101.005 145.655 101.685 ;
        RECT 145.665 101.005 147.035 101.815 ;
        RECT 17.465 100.795 17.635 101.005 ;
        RECT 18.840 100.845 18.960 100.955 ;
        RECT 20.225 100.795 20.395 100.985 ;
        RECT 20.680 100.845 20.800 100.955 ;
        RECT 26.205 100.815 26.375 101.005 ;
        RECT 26.665 100.815 26.835 101.005 ;
        RECT 28.045 100.795 28.215 100.985 ;
        RECT 28.780 100.795 28.950 100.985 ;
        RECT 31.080 100.815 31.250 101.005 ;
        RECT 32.645 100.795 32.815 100.985 ;
        RECT 34.945 100.815 35.115 101.005 ;
        RECT 38.165 100.795 38.335 100.985 ;
        RECT 40.465 100.815 40.635 101.005 ;
        RECT 41.845 100.795 42.015 100.985 ;
        RECT 43.685 100.795 43.855 100.985 ;
        RECT 45.985 100.815 46.155 101.005 ;
        RECT 49.205 100.795 49.375 100.985 ;
        RECT 51.505 100.815 51.675 101.005 ;
        RECT 54.725 100.795 54.895 100.985 ;
        RECT 55.195 100.850 55.355 100.960 ;
        RECT 56.565 100.815 56.735 101.005 ;
        RECT 60.245 100.795 60.415 100.985 ;
        RECT 62.085 100.815 62.255 101.005 ;
        RECT 63.465 100.815 63.635 101.005 ;
        RECT 63.920 100.845 64.040 100.955 ;
        RECT 66.685 100.795 66.855 100.985 ;
        RECT 67.145 100.795 67.315 100.985 ;
        RECT 69.445 100.795 69.615 100.985 ;
        RECT 71.100 100.815 71.270 101.005 ;
        RECT 74.965 100.795 75.135 101.005 ;
        RECT 80.485 100.795 80.655 101.005 ;
        RECT 82.325 100.815 82.495 101.005 ;
        RECT 85.085 100.815 85.255 101.005 ;
        RECT 86.005 100.795 86.175 100.985 ;
        RECT 91.525 100.795 91.695 101.005 ;
        RECT 91.985 100.815 92.155 101.005 ;
        RECT 94.280 100.845 94.400 100.955 ;
        RECT 95.205 100.795 95.375 100.985 ;
        RECT 97.505 100.815 97.675 101.005 ;
        RECT 100.725 100.795 100.895 100.985 ;
        RECT 105.325 100.815 105.495 101.005 ;
        RECT 105.785 100.815 105.955 101.005 ;
        RECT 106.255 100.840 106.415 100.950 ;
        RECT 107.165 100.795 107.335 100.985 ;
        RECT 108.085 100.815 108.255 101.005 ;
        RECT 109.925 100.795 110.095 100.985 ;
        RECT 110.845 100.815 111.015 101.005 ;
        RECT 112.680 100.845 112.800 100.955 ;
        RECT 115.455 100.840 115.615 100.950 ;
        RECT 116.365 100.795 116.535 100.985 ;
        RECT 116.550 100.815 116.720 101.005 ;
        RECT 117.285 100.815 117.455 101.005 ;
        RECT 119.125 100.795 119.295 100.985 ;
        RECT 120.965 100.795 121.135 100.985 ;
        RECT 124.645 100.815 124.815 101.005 ;
        RECT 126.485 100.795 126.655 100.985 ;
        RECT 130.160 100.845 130.280 100.955 ;
        RECT 130.625 100.815 130.795 101.005 ;
        RECT 132.005 100.795 132.175 100.985 ;
        RECT 133.845 100.795 134.015 101.005 ;
        RECT 135.680 100.845 135.800 100.955 ;
        RECT 136.145 100.815 136.315 101.005 ;
        RECT 136.605 100.795 136.775 100.985 ;
        RECT 143.500 100.845 143.620 100.955 ;
        RECT 143.965 100.795 144.135 101.005 ;
        RECT 146.725 100.795 146.895 101.005 ;
        RECT 17.325 99.985 18.695 100.795 ;
        RECT 18.705 100.115 20.535 100.795 ;
        RECT 21.045 100.115 28.355 100.795 ;
        RECT 28.365 100.115 32.265 100.795 ;
        RECT 18.705 99.885 20.050 100.115 ;
        RECT 21.045 99.885 22.395 100.115 ;
        RECT 23.930 99.895 24.840 100.115 ;
        RECT 28.365 99.885 29.295 100.115 ;
        RECT 32.505 99.985 38.015 100.795 ;
        RECT 38.025 99.985 41.695 100.795 ;
        RECT 41.705 99.985 43.075 100.795 ;
        RECT 43.095 99.925 43.525 100.710 ;
        RECT 43.545 99.985 49.055 100.795 ;
        RECT 49.065 99.985 54.575 100.795 ;
        RECT 54.585 99.985 60.095 100.795 ;
        RECT 60.105 99.985 63.775 100.795 ;
        RECT 64.245 100.115 66.995 100.795 ;
        RECT 64.245 99.885 65.175 100.115 ;
        RECT 67.005 99.985 68.835 100.795 ;
        RECT 68.855 99.925 69.285 100.710 ;
        RECT 69.305 99.985 74.815 100.795 ;
        RECT 74.825 99.985 80.335 100.795 ;
        RECT 80.345 99.985 85.855 100.795 ;
        RECT 85.865 99.985 91.375 100.795 ;
        RECT 91.385 99.985 94.135 100.795 ;
        RECT 94.615 99.925 95.045 100.710 ;
        RECT 95.065 99.985 100.575 100.795 ;
        RECT 100.585 99.985 106.095 100.795 ;
        RECT 107.025 100.115 109.775 100.795 ;
        RECT 108.845 99.885 109.775 100.115 ;
        RECT 109.785 99.985 115.295 100.795 ;
        RECT 116.225 100.115 118.975 100.795 ;
        RECT 118.045 99.885 118.975 100.115 ;
        RECT 118.985 99.985 120.355 100.795 ;
        RECT 120.375 99.925 120.805 100.710 ;
        RECT 120.825 99.985 126.335 100.795 ;
        RECT 126.345 99.985 131.855 100.795 ;
        RECT 131.865 99.985 133.695 100.795 ;
        RECT 133.705 100.115 136.455 100.795 ;
        RECT 136.465 100.115 143.775 100.795 ;
        RECT 143.825 100.115 145.655 100.795 ;
        RECT 135.525 99.885 136.455 100.115 ;
        RECT 139.980 99.895 140.890 100.115 ;
        RECT 142.425 99.885 143.775 100.115 ;
        RECT 144.310 99.885 145.655 100.115 ;
        RECT 145.665 99.985 147.035 100.795 ;
      LAYER nwell ;
        RECT 17.130 96.765 147.230 99.595 ;
      LAYER pwell ;
        RECT 17.325 95.565 18.695 96.375 ;
        RECT 19.205 96.245 20.555 96.475 ;
        RECT 22.090 96.245 23.000 96.465 ;
        RECT 19.205 95.565 26.515 96.245 ;
        RECT 26.525 95.565 27.895 96.375 ;
        RECT 27.905 96.275 28.860 96.475 ;
        RECT 27.905 95.595 30.185 96.275 ;
        RECT 30.215 95.650 30.645 96.435 ;
        RECT 27.905 95.565 28.860 95.595 ;
        RECT 17.465 95.355 17.635 95.565 ;
        RECT 18.840 95.405 18.960 95.515 ;
        RECT 20.225 95.355 20.395 95.545 ;
        RECT 22.065 95.355 22.235 95.545 ;
        RECT 25.930 95.355 26.100 95.545 ;
        RECT 26.205 95.375 26.375 95.565 ;
        RECT 26.665 95.375 26.835 95.565 ;
        RECT 26.940 95.355 27.110 95.545 ;
        RECT 29.890 95.375 30.060 95.595 ;
        RECT 30.745 95.565 34.195 96.475 ;
        RECT 36.150 96.275 37.095 96.475 ;
        RECT 34.345 95.595 37.095 96.275 ;
        RECT 30.805 95.515 30.975 95.565 ;
        RECT 30.800 95.405 30.975 95.515 ;
        RECT 30.805 95.375 30.975 95.405 ;
        RECT 31.270 95.355 31.440 95.545 ;
        RECT 34.490 95.375 34.660 95.595 ;
        RECT 36.150 95.565 37.095 95.595 ;
        RECT 37.105 95.565 42.615 96.375 ;
        RECT 42.625 95.565 48.135 96.375 ;
        RECT 48.145 95.565 53.655 96.375 ;
        RECT 53.665 95.565 55.495 96.375 ;
        RECT 55.975 95.650 56.405 96.435 ;
        RECT 56.425 95.565 61.935 96.375 ;
        RECT 63.765 96.245 64.695 96.475 ;
        RECT 61.945 95.565 64.695 96.245 ;
        RECT 64.705 95.565 67.455 96.375 ;
        RECT 67.465 96.245 68.395 96.475 ;
        RECT 67.465 95.565 71.365 96.245 ;
        RECT 71.605 95.565 74.815 96.475 ;
        RECT 74.825 95.565 78.495 96.375 ;
        RECT 80.785 96.245 81.715 96.475 ;
        RECT 78.965 95.565 81.715 96.245 ;
        RECT 81.735 95.650 82.165 96.435 ;
        RECT 82.185 95.565 84.015 96.375 ;
        RECT 84.025 96.245 84.955 96.475 ;
        RECT 84.025 95.565 87.925 96.245 ;
        RECT 88.165 95.565 89.995 96.375 ;
        RECT 90.465 95.565 94.120 96.475 ;
        RECT 94.145 95.565 95.515 96.375 ;
        RECT 97.365 96.245 101.295 96.475 ;
        RECT 101.965 96.245 102.895 96.475 ;
        RECT 95.525 95.565 97.355 96.245 ;
        RECT 97.365 95.565 101.780 96.245 ;
        RECT 101.965 95.565 105.865 96.245 ;
        RECT 106.105 95.565 107.475 96.375 ;
        RECT 107.495 95.650 107.925 96.435 ;
        RECT 108.405 96.245 109.335 96.475 ;
        RECT 108.405 95.565 112.305 96.245 ;
        RECT 112.545 95.565 114.375 96.375 ;
        RECT 114.385 95.565 118.040 96.475 ;
        RECT 118.065 95.565 123.575 96.375 ;
        RECT 123.585 95.565 126.335 96.375 ;
        RECT 128.165 96.245 129.095 96.475 ;
        RECT 126.345 95.565 129.095 96.245 ;
        RECT 129.105 95.565 130.935 96.245 ;
        RECT 130.945 95.565 132.775 96.245 ;
        RECT 133.255 95.650 133.685 96.435 ;
        RECT 135.525 96.245 136.455 96.475 ;
        RECT 133.705 95.565 136.455 96.245 ;
        RECT 136.465 95.565 139.675 96.475 ;
        RECT 139.685 95.565 141.515 96.375 ;
        RECT 142.470 96.245 143.815 96.475 ;
        RECT 144.310 96.245 145.655 96.475 ;
        RECT 141.985 95.565 143.815 96.245 ;
        RECT 143.825 95.565 145.655 96.245 ;
        RECT 145.665 95.565 147.035 96.375 ;
        RECT 17.325 94.545 18.695 95.355 ;
        RECT 18.705 94.675 20.535 95.355 ;
        RECT 20.545 94.675 22.375 95.355 ;
        RECT 22.615 94.675 26.515 95.355 ;
        RECT 18.705 94.445 20.050 94.675 ;
        RECT 20.545 94.445 21.890 94.675 ;
        RECT 25.585 94.445 26.515 94.675 ;
        RECT 26.525 94.675 30.425 95.355 ;
        RECT 26.525 94.445 27.455 94.675 ;
        RECT 31.125 94.445 32.475 95.355 ;
        RECT 32.505 95.325 33.455 95.355 ;
        RECT 35.860 95.325 36.030 95.545 ;
        RECT 36.320 95.405 36.440 95.515 ;
        RECT 36.785 95.355 36.955 95.545 ;
        RECT 37.245 95.375 37.415 95.565 ;
        RECT 40.000 95.405 40.120 95.515 ;
        RECT 41.380 95.355 41.550 95.545 ;
        RECT 41.845 95.355 42.015 95.545 ;
        RECT 42.765 95.375 42.935 95.565 ;
        RECT 43.685 95.355 43.855 95.545 ;
        RECT 48.285 95.375 48.455 95.565 ;
        RECT 49.205 95.355 49.375 95.545 ;
        RECT 53.805 95.375 53.975 95.565 ;
        RECT 54.725 95.355 54.895 95.545 ;
        RECT 55.640 95.405 55.760 95.515 ;
        RECT 56.565 95.375 56.735 95.565 ;
        RECT 58.400 95.405 58.520 95.515 ;
        RECT 61.165 95.355 61.335 95.545 ;
        RECT 61.625 95.355 61.795 95.545 ;
        RECT 62.085 95.375 62.255 95.565 ;
        RECT 64.845 95.375 65.015 95.565 ;
        RECT 67.880 95.375 68.050 95.565 ;
        RECT 69.720 95.355 69.890 95.545 ;
        RECT 71.745 95.375 71.915 95.565 ;
        RECT 73.585 95.355 73.755 95.545 ;
        RECT 74.965 95.375 75.135 95.565 ;
        RECT 76.620 95.355 76.790 95.545 ;
        RECT 78.640 95.405 78.760 95.515 ;
        RECT 79.105 95.375 79.275 95.565 ;
        RECT 80.485 95.355 80.655 95.545 ;
        RECT 82.325 95.375 82.495 95.565 ;
        RECT 84.440 95.375 84.610 95.565 ;
        RECT 88.120 95.355 88.290 95.545 ;
        RECT 88.305 95.375 88.475 95.565 ;
        RECT 90.140 95.405 90.260 95.515 ;
        RECT 90.610 95.375 90.780 95.565 ;
        RECT 91.985 95.355 92.155 95.545 ;
        RECT 94.285 95.375 94.455 95.565 ;
        RECT 95.205 95.355 95.375 95.545 ;
        RECT 95.665 95.375 95.835 95.565 ;
        RECT 101.670 95.545 101.780 95.565 ;
        RECT 101.670 95.375 101.840 95.545 ;
        RECT 102.380 95.375 102.550 95.565 ;
        RECT 102.840 95.355 103.010 95.545 ;
        RECT 106.245 95.375 106.415 95.565 ;
        RECT 106.700 95.405 106.820 95.515 ;
        RECT 107.165 95.355 107.335 95.545 ;
        RECT 108.080 95.405 108.200 95.515 ;
        RECT 108.820 95.375 108.990 95.565 ;
        RECT 112.685 95.375 112.855 95.565 ;
        RECT 114.530 95.375 114.700 95.565 ;
        RECT 114.800 95.355 114.970 95.545 ;
        RECT 118.205 95.375 118.375 95.565 ;
        RECT 118.665 95.355 118.835 95.545 ;
        RECT 121.240 95.355 121.410 95.545 ;
        RECT 123.725 95.375 123.895 95.565 ;
        RECT 125.105 95.355 125.275 95.545 ;
        RECT 126.485 95.355 126.655 95.565 ;
        RECT 129.245 95.375 129.415 95.565 ;
        RECT 132.465 95.375 132.635 95.565 ;
        RECT 132.920 95.405 133.040 95.515 ;
        RECT 133.845 95.355 134.015 95.565 ;
        RECT 135.680 95.405 135.800 95.515 ;
        RECT 136.420 95.355 136.590 95.545 ;
        RECT 139.365 95.375 139.535 95.565 ;
        RECT 139.825 95.375 139.995 95.565 ;
        RECT 141.660 95.405 141.780 95.515 ;
        RECT 142.125 95.375 142.295 95.565 ;
        RECT 143.045 95.355 143.215 95.545 ;
        RECT 143.500 95.405 143.620 95.515 ;
        RECT 143.965 95.355 144.135 95.565 ;
        RECT 146.725 95.355 146.895 95.565 ;
        RECT 32.505 94.645 36.175 95.325 ;
        RECT 32.505 94.445 33.455 94.645 ;
        RECT 36.725 94.445 39.725 95.355 ;
        RECT 40.345 94.445 41.695 95.355 ;
        RECT 41.705 94.545 43.075 95.355 ;
        RECT 43.095 94.485 43.525 95.270 ;
        RECT 43.545 94.545 49.055 95.355 ;
        RECT 49.065 94.545 54.575 95.355 ;
        RECT 54.585 94.545 58.255 95.355 ;
        RECT 58.725 94.675 61.475 95.355 ;
        RECT 61.485 94.675 68.795 95.355 ;
        RECT 58.725 94.445 59.655 94.675 ;
        RECT 65.000 94.455 65.910 94.675 ;
        RECT 67.445 94.445 68.795 94.675 ;
        RECT 68.855 94.485 69.285 95.270 ;
        RECT 69.305 94.675 73.205 95.355 ;
        RECT 73.445 94.675 76.195 95.355 ;
        RECT 69.305 94.445 70.235 94.675 ;
        RECT 75.265 94.445 76.195 94.675 ;
        RECT 76.205 94.675 80.105 95.355 ;
        RECT 80.345 94.675 87.655 95.355 ;
        RECT 76.205 94.445 77.135 94.675 ;
        RECT 83.860 94.455 84.770 94.675 ;
        RECT 86.305 94.445 87.655 94.675 ;
        RECT 87.705 94.675 91.605 95.355 ;
        RECT 91.845 94.675 94.595 95.355 ;
        RECT 87.705 94.445 88.635 94.675 ;
        RECT 93.665 94.445 94.595 94.675 ;
        RECT 94.615 94.485 95.045 95.270 ;
        RECT 95.065 94.675 102.375 95.355 ;
        RECT 98.580 94.455 99.490 94.675 ;
        RECT 101.025 94.445 102.375 94.675 ;
        RECT 102.425 94.675 106.325 95.355 ;
        RECT 107.025 94.675 114.335 95.355 ;
        RECT 102.425 94.445 103.355 94.675 ;
        RECT 110.540 94.455 111.450 94.675 ;
        RECT 112.985 94.445 114.335 94.675 ;
        RECT 114.385 94.675 118.285 95.355 ;
        RECT 114.385 94.445 115.315 94.675 ;
        RECT 118.525 94.545 120.355 95.355 ;
        RECT 120.375 94.485 120.805 95.270 ;
        RECT 120.825 94.675 124.725 95.355 ;
        RECT 120.825 94.445 121.755 94.675 ;
        RECT 124.965 94.545 126.335 95.355 ;
        RECT 126.345 94.675 133.655 95.355 ;
        RECT 133.705 94.675 135.535 95.355 ;
        RECT 136.005 94.675 139.905 95.355 ;
        RECT 129.860 94.455 130.770 94.675 ;
        RECT 132.305 94.445 133.655 94.675 ;
        RECT 136.005 94.445 136.935 94.675 ;
        RECT 140.145 94.445 143.355 95.355 ;
        RECT 143.825 94.675 145.655 95.355 ;
        RECT 144.310 94.445 145.655 94.675 ;
        RECT 145.665 94.545 147.035 95.355 ;
      LAYER nwell ;
        RECT 17.130 91.325 147.230 94.155 ;
      LAYER pwell ;
        RECT 17.325 90.125 18.695 90.935 ;
        RECT 18.705 90.125 21.455 90.935 ;
        RECT 24.980 90.805 25.890 91.025 ;
        RECT 27.425 90.805 28.775 91.035 ;
        RECT 21.465 90.125 28.775 90.805 ;
        RECT 28.845 90.125 30.195 91.035 ;
        RECT 30.215 90.210 30.645 90.995 ;
        RECT 31.665 90.125 35.115 91.035 ;
        RECT 35.345 90.125 38.795 91.035 ;
        RECT 39.025 90.125 42.475 91.035 ;
        RECT 42.705 90.125 46.155 91.035 ;
        RECT 48.125 90.805 49.055 91.035 ;
        RECT 46.305 90.125 49.055 90.805 ;
        RECT 49.065 90.125 54.575 90.935 ;
        RECT 54.585 90.125 55.955 90.935 ;
        RECT 55.975 90.210 56.405 90.995 ;
        RECT 56.425 90.125 57.795 90.935 ;
        RECT 61.320 90.805 62.230 91.025 ;
        RECT 63.765 90.805 65.115 91.035 ;
        RECT 68.680 90.805 69.590 91.025 ;
        RECT 71.125 90.805 72.475 91.035 ;
        RECT 73.010 90.805 74.355 91.035 ;
        RECT 77.880 90.805 78.790 91.025 ;
        RECT 80.325 90.805 81.675 91.035 ;
        RECT 57.805 90.125 65.115 90.805 ;
        RECT 65.165 90.125 72.475 90.805 ;
        RECT 72.525 90.125 74.355 90.805 ;
        RECT 74.365 90.125 81.675 90.805 ;
        RECT 81.735 90.210 82.165 90.995 ;
        RECT 82.185 90.125 85.395 91.035 ;
        RECT 85.405 90.125 87.235 90.935 ;
        RECT 90.760 90.805 91.670 91.025 ;
        RECT 93.205 90.805 94.555 91.035 ;
        RECT 87.245 90.125 94.555 90.805 ;
        RECT 94.605 90.125 95.975 90.905 ;
        RECT 99.500 90.805 100.410 91.025 ;
        RECT 101.945 90.805 103.295 91.035 ;
        RECT 95.985 90.125 103.295 90.805 ;
        RECT 103.345 90.125 107.000 91.035 ;
        RECT 107.495 90.210 107.925 90.995 ;
        RECT 111.460 90.805 112.370 91.025 ;
        RECT 113.905 90.805 115.255 91.035 ;
        RECT 118.820 90.805 119.730 91.025 ;
        RECT 121.265 90.805 122.615 91.035 ;
        RECT 126.180 90.805 127.090 91.025 ;
        RECT 128.625 90.805 129.975 91.035 ;
        RECT 107.945 90.125 115.255 90.805 ;
        RECT 115.305 90.125 122.615 90.805 ;
        RECT 122.665 90.125 129.975 90.805 ;
        RECT 130.025 90.805 130.955 91.035 ;
        RECT 130.025 90.125 132.775 90.805 ;
        RECT 133.255 90.210 133.685 90.995 ;
        RECT 137.680 90.805 138.590 91.025 ;
        RECT 140.125 90.805 141.475 91.035 ;
        RECT 134.165 90.125 141.475 90.805 ;
        RECT 141.525 90.805 142.455 91.035 ;
        RECT 141.525 90.125 145.425 90.805 ;
        RECT 145.665 90.125 147.035 90.935 ;
        RECT 17.465 89.915 17.635 90.125 ;
        RECT 18.845 90.075 19.015 90.125 ;
        RECT 18.840 89.965 19.015 90.075 ;
        RECT 18.845 89.935 19.015 89.965 ;
        RECT 21.605 89.935 21.775 90.125 ;
        RECT 26.205 89.915 26.375 90.105 ;
        RECT 26.940 89.915 27.110 90.105 ;
        RECT 29.880 89.935 30.050 90.125 ;
        RECT 31.725 90.105 31.895 90.125 ;
        RECT 30.815 89.960 30.975 90.080 ;
        RECT 31.725 89.935 31.900 90.105 ;
        RECT 31.730 89.915 31.900 89.935 ;
        RECT 34.945 89.915 35.115 90.105 ;
        RECT 35.405 89.935 35.575 90.125 ;
        RECT 39.085 89.935 39.255 90.125 ;
        RECT 17.325 89.105 18.695 89.915 ;
        RECT 19.205 89.235 26.515 89.915 ;
        RECT 26.525 89.235 30.425 89.915 ;
        RECT 19.205 89.005 20.555 89.235 ;
        RECT 22.090 89.015 23.000 89.235 ;
        RECT 26.525 89.005 27.455 89.235 ;
        RECT 31.585 89.005 34.505 89.915 ;
        RECT 34.885 89.005 38.335 89.915 ;
        RECT 38.485 89.885 39.430 89.915 ;
        RECT 40.920 89.885 41.090 90.105 ;
        RECT 41.390 89.915 41.560 90.105 ;
        RECT 42.765 90.075 42.935 90.125 ;
        RECT 42.760 89.965 42.935 90.075 ;
        RECT 42.765 89.935 42.935 89.965 ;
        RECT 43.685 89.915 43.855 90.105 ;
        RECT 46.445 89.915 46.615 90.125 ;
        RECT 49.205 89.935 49.375 90.125 ;
        RECT 51.965 89.915 52.135 90.105 ;
        RECT 54.725 89.935 54.895 90.125 ;
        RECT 56.565 89.935 56.735 90.125 ;
        RECT 57.945 89.935 58.115 90.125 ;
        RECT 58.405 89.915 58.575 90.105 ;
        RECT 58.865 89.915 59.035 90.105 ;
        RECT 60.705 89.915 60.875 90.105 ;
        RECT 65.305 89.935 65.475 90.125 ;
        RECT 68.075 89.960 68.235 90.070 ;
        RECT 69.720 89.915 69.890 90.105 ;
        RECT 72.665 89.935 72.835 90.125 ;
        RECT 73.585 89.915 73.755 90.105 ;
        RECT 74.505 89.935 74.675 90.125 ;
        RECT 76.805 89.915 76.975 90.105 ;
        RECT 82.325 89.915 82.495 90.125 ;
        RECT 83.705 89.915 83.875 90.105 ;
        RECT 85.545 89.935 85.715 90.125 ;
        RECT 87.385 89.935 87.555 90.125 ;
        RECT 91.070 89.915 91.240 90.105 ;
        RECT 95.480 89.915 95.650 90.105 ;
        RECT 95.655 89.935 95.825 90.125 ;
        RECT 96.125 89.935 96.295 90.125 ;
        RECT 99.345 89.915 99.515 90.105 ;
        RECT 102.105 89.915 102.275 90.105 ;
        RECT 103.490 89.935 103.660 90.125 ;
        RECT 104.865 89.915 105.035 90.105 ;
        RECT 107.160 89.965 107.280 90.075 ;
        RECT 107.625 89.915 107.795 90.105 ;
        RECT 108.085 89.935 108.255 90.125 ;
        RECT 111.305 89.915 111.475 90.105 ;
        RECT 112.685 89.915 112.855 90.105 ;
        RECT 115.445 90.075 115.615 90.125 ;
        RECT 115.440 89.965 115.615 90.075 ;
        RECT 115.445 89.935 115.615 89.965 ;
        RECT 116.180 89.915 116.350 90.105 ;
        RECT 120.040 89.965 120.160 90.075 ;
        RECT 120.965 89.915 121.135 90.105 ;
        RECT 122.805 89.935 122.975 90.125 ;
        RECT 123.725 89.915 123.895 90.105 ;
        RECT 131.360 89.915 131.530 90.105 ;
        RECT 132.465 89.935 132.635 90.125 ;
        RECT 132.920 89.965 133.040 90.075 ;
        RECT 133.840 89.965 133.960 90.075 ;
        RECT 134.305 89.935 134.475 90.125 ;
        RECT 136.135 89.915 136.305 90.105 ;
        RECT 136.605 89.915 136.775 90.105 ;
        RECT 141.940 89.935 142.110 90.125 ;
        RECT 143.965 89.915 144.135 90.105 ;
        RECT 146.725 89.915 146.895 90.125 ;
        RECT 38.485 89.205 41.235 89.885 ;
        RECT 38.485 89.005 39.430 89.205 ;
        RECT 41.245 89.005 42.595 89.915 ;
        RECT 43.095 89.045 43.525 89.830 ;
        RECT 43.545 89.005 46.295 89.915 ;
        RECT 46.305 89.105 51.815 89.915 ;
        RECT 51.825 89.105 57.335 89.915 ;
        RECT 57.345 89.135 58.715 89.915 ;
        RECT 58.725 89.105 60.555 89.915 ;
        RECT 60.565 89.235 67.875 89.915 ;
        RECT 64.080 89.015 64.990 89.235 ;
        RECT 66.525 89.005 67.875 89.235 ;
        RECT 68.855 89.045 69.285 89.830 ;
        RECT 69.305 89.235 73.205 89.915 ;
        RECT 69.305 89.005 70.235 89.235 ;
        RECT 73.445 89.005 76.655 89.915 ;
        RECT 76.665 89.105 82.175 89.915 ;
        RECT 82.185 89.105 83.555 89.915 ;
        RECT 83.565 89.235 90.875 89.915 ;
        RECT 87.080 89.015 87.990 89.235 ;
        RECT 89.525 89.005 90.875 89.235 ;
        RECT 90.925 89.005 94.580 89.915 ;
        RECT 94.615 89.045 95.045 89.830 ;
        RECT 95.065 89.235 98.965 89.915 ;
        RECT 99.205 89.235 101.955 89.915 ;
        RECT 95.065 89.005 95.995 89.235 ;
        RECT 101.025 89.005 101.955 89.235 ;
        RECT 101.965 89.105 104.715 89.915 ;
        RECT 104.725 89.235 107.475 89.915 ;
        RECT 106.545 89.005 107.475 89.235 ;
        RECT 107.485 89.105 111.155 89.915 ;
        RECT 111.165 89.105 112.535 89.915 ;
        RECT 112.545 89.235 115.295 89.915 ;
        RECT 114.365 89.005 115.295 89.235 ;
        RECT 115.765 89.235 119.665 89.915 ;
        RECT 115.765 89.005 116.695 89.235 ;
        RECT 120.375 89.045 120.805 89.830 ;
        RECT 120.825 89.105 123.575 89.915 ;
        RECT 123.585 89.235 130.895 89.915 ;
        RECT 127.100 89.015 128.010 89.235 ;
        RECT 129.545 89.005 130.895 89.235 ;
        RECT 130.945 89.235 134.845 89.915 ;
        RECT 130.945 89.005 131.875 89.235 ;
        RECT 135.085 89.135 136.455 89.915 ;
        RECT 136.465 89.235 143.775 89.915 ;
        RECT 143.825 89.235 145.655 89.915 ;
        RECT 139.980 89.015 140.890 89.235 ;
        RECT 142.425 89.005 143.775 89.235 ;
        RECT 144.310 89.005 145.655 89.235 ;
        RECT 145.665 89.105 147.035 89.915 ;
      LAYER nwell ;
        RECT 17.130 85.885 147.230 88.715 ;
      LAYER pwell ;
        RECT 17.325 84.685 18.695 85.495 ;
        RECT 18.705 84.685 20.075 85.465 ;
        RECT 20.085 84.685 21.455 85.465 ;
        RECT 21.925 85.365 23.270 85.595 ;
        RECT 21.925 84.685 23.755 85.365 ;
        RECT 23.765 84.685 25.135 85.465 ;
        RECT 25.145 84.685 26.515 85.465 ;
        RECT 26.525 84.685 28.355 85.495 ;
        RECT 28.850 85.365 30.195 85.595 ;
        RECT 28.365 84.685 30.195 85.365 ;
        RECT 30.215 84.770 30.645 85.555 ;
        RECT 30.665 84.685 32.035 85.465 ;
        RECT 32.125 84.685 35.125 85.595 ;
        RECT 35.265 84.685 36.635 85.465 ;
        RECT 36.645 84.685 38.015 85.495 ;
        RECT 38.025 84.685 39.395 85.465 ;
        RECT 39.405 84.685 41.235 85.495 ;
        RECT 41.245 84.685 42.615 85.465 ;
        RECT 43.095 84.770 43.525 85.555 ;
        RECT 44.465 84.685 45.835 85.465 ;
        RECT 45.845 84.685 47.675 85.495 ;
        RECT 47.685 84.685 49.055 85.465 ;
        RECT 49.065 84.685 50.895 85.495 ;
        RECT 50.905 84.685 52.275 85.465 ;
        RECT 52.285 84.685 54.115 85.495 ;
        RECT 54.125 84.685 55.495 85.465 ;
        RECT 55.975 84.770 56.405 85.555 ;
        RECT 56.425 85.365 57.770 85.595 ;
        RECT 58.265 85.365 59.610 85.595 ;
        RECT 60.105 85.365 61.450 85.595 ;
        RECT 61.945 85.365 62.875 85.595 ;
        RECT 67.445 85.365 68.375 85.595 ;
        RECT 56.425 84.685 58.255 85.365 ;
        RECT 58.265 84.685 60.095 85.365 ;
        RECT 60.105 84.685 61.935 85.365 ;
        RECT 61.945 84.685 64.695 85.365 ;
        RECT 65.625 84.685 68.375 85.365 ;
        RECT 68.855 84.770 69.285 85.555 ;
        RECT 69.305 85.365 70.235 85.595 ;
        RECT 73.930 85.365 75.275 85.595 ;
        RECT 69.305 84.685 73.205 85.365 ;
        RECT 73.445 84.685 75.275 85.365 ;
        RECT 76.205 85.365 77.550 85.595 ;
        RECT 78.530 85.365 79.875 85.595 ;
        RECT 80.370 85.365 81.715 85.595 ;
        RECT 76.205 84.685 78.035 85.365 ;
        RECT 78.045 84.685 79.875 85.365 ;
        RECT 79.885 84.685 81.715 85.365 ;
        RECT 81.735 84.770 82.165 85.555 ;
        RECT 82.185 84.685 83.555 85.495 ;
        RECT 85.385 85.365 86.315 85.595 ;
        RECT 89.065 85.365 89.995 85.595 ;
        RECT 83.565 84.685 86.315 85.365 ;
        RECT 87.245 84.685 89.995 85.365 ;
        RECT 90.005 85.365 91.350 85.595 ;
        RECT 92.330 85.365 93.675 85.595 ;
        RECT 90.005 84.685 91.835 85.365 ;
        RECT 91.845 84.685 93.675 85.365 ;
        RECT 94.615 84.770 95.045 85.555 ;
        RECT 95.550 85.365 96.895 85.595 ;
        RECT 97.390 85.365 98.735 85.595 ;
        RECT 95.065 84.685 96.895 85.365 ;
        RECT 96.905 84.685 98.735 85.365 ;
        RECT 99.205 85.365 100.550 85.595 ;
        RECT 99.205 84.685 101.035 85.365 ;
        RECT 101.045 84.685 102.415 85.495 ;
        RECT 102.425 85.365 103.770 85.595 ;
        RECT 102.425 84.685 104.255 85.365 ;
        RECT 104.265 84.685 105.635 85.495 ;
        RECT 105.645 85.365 106.990 85.595 ;
        RECT 105.645 84.685 107.475 85.365 ;
        RECT 107.495 84.770 107.925 85.555 ;
        RECT 108.865 85.365 110.210 85.595 ;
        RECT 108.865 84.685 110.695 85.365 ;
        RECT 110.705 84.685 112.075 85.495 ;
        RECT 112.085 85.365 113.430 85.595 ;
        RECT 115.745 85.365 116.675 85.595 ;
        RECT 112.085 84.685 113.915 85.365 ;
        RECT 113.925 84.685 116.675 85.365 ;
        RECT 117.145 84.685 120.355 85.595 ;
        RECT 120.375 84.770 120.805 85.555 ;
        RECT 121.310 85.365 122.655 85.595 ;
        RECT 123.150 85.365 124.495 85.595 ;
        RECT 120.825 84.685 122.655 85.365 ;
        RECT 122.665 84.685 124.495 85.365 ;
        RECT 124.505 85.365 125.850 85.595 ;
        RECT 129.545 85.365 130.475 85.595 ;
        RECT 130.970 85.365 132.315 85.595 ;
        RECT 124.505 84.685 126.335 85.365 ;
        RECT 126.575 84.685 130.475 85.365 ;
        RECT 130.485 84.685 132.315 85.365 ;
        RECT 133.255 84.770 133.685 85.555 ;
        RECT 133.720 84.685 137.375 85.595 ;
        RECT 139.205 85.365 140.135 85.595 ;
        RECT 140.630 85.365 141.975 85.595 ;
        RECT 142.470 85.365 143.815 85.595 ;
        RECT 144.310 85.365 145.655 85.595 ;
        RECT 137.385 84.685 140.135 85.365 ;
        RECT 140.145 84.685 141.975 85.365 ;
        RECT 141.985 84.685 143.815 85.365 ;
        RECT 143.825 84.685 145.655 85.365 ;
        RECT 145.665 84.685 147.035 85.495 ;
        RECT 17.465 84.495 17.635 84.685 ;
        RECT 18.855 84.495 19.025 84.685 ;
        RECT 20.225 84.495 20.395 84.685 ;
        RECT 21.600 84.525 21.720 84.635 ;
        RECT 23.445 84.495 23.615 84.685 ;
        RECT 23.915 84.495 24.085 84.685 ;
        RECT 25.295 84.495 25.465 84.685 ;
        RECT 26.665 84.495 26.835 84.685 ;
        RECT 28.505 84.495 28.675 84.685 ;
        RECT 30.815 84.495 30.985 84.685 ;
        RECT 32.185 84.495 32.355 84.685 ;
        RECT 35.405 84.495 35.575 84.685 ;
        RECT 36.785 84.495 36.955 84.685 ;
        RECT 38.165 84.495 38.335 84.685 ;
        RECT 39.545 84.495 39.715 84.685 ;
        RECT 42.295 84.495 42.465 84.685 ;
        RECT 42.760 84.525 42.880 84.635 ;
        RECT 43.695 84.530 43.855 84.640 ;
        RECT 45.515 84.495 45.685 84.685 ;
        RECT 45.985 84.495 46.155 84.685 ;
        RECT 48.735 84.495 48.905 84.685 ;
        RECT 49.205 84.495 49.375 84.685 ;
        RECT 51.965 84.495 52.135 84.685 ;
        RECT 52.425 84.495 52.595 84.685 ;
        RECT 55.185 84.495 55.355 84.685 ;
        RECT 55.640 84.525 55.760 84.635 ;
        RECT 57.945 84.495 58.115 84.685 ;
        RECT 59.785 84.495 59.955 84.685 ;
        RECT 61.625 84.495 61.795 84.685 ;
        RECT 64.385 84.495 64.555 84.685 ;
        RECT 64.855 84.530 65.015 84.640 ;
        RECT 65.765 84.495 65.935 84.685 ;
        RECT 68.520 84.525 68.640 84.635 ;
        RECT 69.720 84.495 69.890 84.685 ;
        RECT 73.585 84.495 73.755 84.685 ;
        RECT 75.435 84.530 75.595 84.640 ;
        RECT 77.725 84.495 77.895 84.685 ;
        RECT 78.185 84.495 78.355 84.685 ;
        RECT 80.025 84.495 80.195 84.685 ;
        RECT 82.325 84.495 82.495 84.685 ;
        RECT 83.705 84.495 83.875 84.685 ;
        RECT 86.475 84.530 86.635 84.640 ;
        RECT 87.385 84.495 87.555 84.685 ;
        RECT 91.525 84.495 91.695 84.685 ;
        RECT 91.985 84.495 92.155 84.685 ;
        RECT 93.835 84.530 93.995 84.640 ;
        RECT 95.205 84.495 95.375 84.685 ;
        RECT 97.045 84.495 97.215 84.685 ;
        RECT 98.880 84.525 99.000 84.635 ;
        RECT 100.725 84.495 100.895 84.685 ;
        RECT 101.185 84.495 101.355 84.685 ;
        RECT 103.945 84.495 104.115 84.685 ;
        RECT 104.405 84.495 104.575 84.685 ;
        RECT 107.165 84.495 107.335 84.685 ;
        RECT 108.095 84.530 108.255 84.640 ;
        RECT 110.385 84.495 110.555 84.685 ;
        RECT 110.845 84.495 111.015 84.685 ;
        RECT 113.605 84.495 113.775 84.685 ;
        RECT 114.065 84.495 114.235 84.685 ;
        RECT 116.820 84.525 116.940 84.635 ;
        RECT 120.045 84.495 120.215 84.685 ;
        RECT 120.965 84.495 121.135 84.685 ;
        RECT 122.805 84.495 122.975 84.685 ;
        RECT 126.025 84.495 126.195 84.685 ;
        RECT 129.890 84.495 130.060 84.685 ;
        RECT 130.625 84.495 130.795 84.685 ;
        RECT 132.475 84.530 132.635 84.640 ;
        RECT 137.060 84.495 137.230 84.685 ;
        RECT 137.525 84.495 137.695 84.685 ;
        RECT 140.285 84.495 140.455 84.685 ;
        RECT 142.125 84.495 142.295 84.685 ;
        RECT 143.965 84.495 144.135 84.685 ;
        RECT 146.725 84.495 146.895 84.685 ;
      LAYER li1 ;
        RECT 17.320 212.335 147.040 212.505 ;
        RECT 17.405 211.245 18.615 212.335 ;
        RECT 18.785 211.900 24.130 212.335 ;
        RECT 24.305 211.900 29.650 212.335 ;
        RECT 17.405 210.535 17.925 211.075 ;
        RECT 18.095 210.705 18.615 211.245 ;
        RECT 17.405 209.785 18.615 210.535 ;
        RECT 20.370 210.330 20.710 211.160 ;
        RECT 22.190 210.650 22.540 211.900 ;
        RECT 25.890 210.330 26.230 211.160 ;
        RECT 27.710 210.650 28.060 211.900 ;
        RECT 30.285 211.170 30.575 212.335 ;
        RECT 30.745 211.900 36.090 212.335 ;
        RECT 36.265 211.900 41.610 212.335 ;
        RECT 18.785 209.785 24.130 210.330 ;
        RECT 24.305 209.785 29.650 210.330 ;
        RECT 30.285 209.785 30.575 210.510 ;
        RECT 32.330 210.330 32.670 211.160 ;
        RECT 34.150 210.650 34.500 211.900 ;
        RECT 37.850 210.330 38.190 211.160 ;
        RECT 39.670 210.650 40.020 211.900 ;
        RECT 41.785 211.245 42.995 212.335 ;
        RECT 41.785 210.535 42.305 211.075 ;
        RECT 42.475 210.705 42.995 211.245 ;
        RECT 43.165 211.170 43.455 212.335 ;
        RECT 43.625 211.900 48.970 212.335 ;
        RECT 49.145 211.900 54.490 212.335 ;
        RECT 30.745 209.785 36.090 210.330 ;
        RECT 36.265 209.785 41.610 210.330 ;
        RECT 41.785 209.785 42.995 210.535 ;
        RECT 43.165 209.785 43.455 210.510 ;
        RECT 45.210 210.330 45.550 211.160 ;
        RECT 47.030 210.650 47.380 211.900 ;
        RECT 50.730 210.330 51.070 211.160 ;
        RECT 52.550 210.650 52.900 211.900 ;
        RECT 54.665 211.245 55.875 212.335 ;
        RECT 54.665 210.535 55.185 211.075 ;
        RECT 55.355 210.705 55.875 211.245 ;
        RECT 56.045 211.170 56.335 212.335 ;
        RECT 56.505 211.245 60.015 212.335 ;
        RECT 56.505 210.555 58.155 211.075 ;
        RECT 58.325 210.725 60.015 211.245 ;
        RECT 60.655 211.355 60.985 212.165 ;
        RECT 61.155 211.535 61.395 212.335 ;
        RECT 60.655 211.185 61.370 211.355 ;
        RECT 60.650 210.775 61.030 211.015 ;
        RECT 61.200 210.945 61.370 211.185 ;
        RECT 61.575 211.315 61.745 212.165 ;
        RECT 61.915 211.535 62.245 212.335 ;
        RECT 62.415 211.315 62.585 212.165 ;
        RECT 61.575 211.145 62.585 211.315 ;
        RECT 62.755 211.185 63.085 212.335 ;
        RECT 63.405 211.900 68.750 212.335 ;
        RECT 61.200 210.775 61.700 210.945 ;
        RECT 61.200 210.605 61.370 210.775 ;
        RECT 62.090 210.635 62.585 211.145 ;
        RECT 62.085 210.605 62.585 210.635 ;
        RECT 43.625 209.785 48.970 210.330 ;
        RECT 49.145 209.785 54.490 210.330 ;
        RECT 54.665 209.785 55.875 210.535 ;
        RECT 56.045 209.785 56.335 210.510 ;
        RECT 56.505 209.785 60.015 210.555 ;
        RECT 60.735 210.435 61.370 210.605 ;
        RECT 61.575 210.435 62.585 210.605 ;
        RECT 60.735 209.955 60.905 210.435 ;
        RECT 61.085 209.785 61.325 210.265 ;
        RECT 61.575 209.955 61.745 210.435 ;
        RECT 61.915 209.785 62.245 210.265 ;
        RECT 62.415 209.955 62.585 210.435 ;
        RECT 62.755 209.785 63.085 210.585 ;
        RECT 64.990 210.330 65.330 211.160 ;
        RECT 66.810 210.650 67.160 211.900 ;
        RECT 68.925 211.170 69.215 212.335 ;
        RECT 69.385 211.900 74.730 212.335 ;
        RECT 63.405 209.785 68.750 210.330 ;
        RECT 68.925 209.785 69.215 210.510 ;
        RECT 70.970 210.330 71.310 211.160 ;
        RECT 72.790 210.650 73.140 211.900 ;
        RECT 74.905 211.245 78.415 212.335 ;
        RECT 78.585 211.245 79.795 212.335 ;
        RECT 74.905 210.555 76.555 211.075 ;
        RECT 76.725 210.725 78.415 211.245 ;
        RECT 69.385 209.785 74.730 210.330 ;
        RECT 74.905 209.785 78.415 210.555 ;
        RECT 78.585 210.535 79.105 211.075 ;
        RECT 79.275 210.705 79.795 211.245 ;
        RECT 79.970 211.185 80.230 212.335 ;
        RECT 80.405 211.260 80.660 212.165 ;
        RECT 80.830 211.575 81.160 212.335 ;
        RECT 81.375 211.405 81.545 212.165 ;
        RECT 78.585 209.785 79.795 210.535 ;
        RECT 79.970 209.785 80.230 210.625 ;
        RECT 80.405 210.530 80.575 211.260 ;
        RECT 80.830 211.235 81.545 211.405 ;
        RECT 80.830 211.025 81.000 211.235 ;
        RECT 81.805 211.170 82.095 212.335 ;
        RECT 83.265 211.405 83.445 212.165 ;
        RECT 83.625 211.575 83.955 212.335 ;
        RECT 83.265 211.235 83.940 211.405 ;
        RECT 84.125 211.260 84.395 212.165 ;
        RECT 83.770 211.090 83.940 211.235 ;
        RECT 80.745 210.695 81.000 211.025 ;
        RECT 80.405 209.955 80.660 210.530 ;
        RECT 80.830 210.505 81.000 210.695 ;
        RECT 81.280 210.685 81.635 211.055 ;
        RECT 83.205 210.685 83.545 211.055 ;
        RECT 83.770 210.760 84.045 211.090 ;
        RECT 80.830 210.335 81.545 210.505 ;
        RECT 80.830 209.785 81.160 210.165 ;
        RECT 81.375 209.955 81.545 210.335 ;
        RECT 81.805 209.785 82.095 210.510 ;
        RECT 83.770 210.505 83.940 210.760 ;
        RECT 83.275 210.335 83.940 210.505 ;
        RECT 84.215 210.460 84.395 211.260 ;
        RECT 83.275 209.955 83.445 210.335 ;
        RECT 83.625 209.785 83.955 210.165 ;
        RECT 84.135 209.955 84.395 210.460 ;
        RECT 85.485 211.615 85.945 212.165 ;
        RECT 86.135 211.615 86.465 212.335 ;
        RECT 85.485 210.245 85.735 211.615 ;
        RECT 86.665 211.445 86.965 211.995 ;
        RECT 87.135 211.665 87.415 212.335 ;
        RECT 86.025 211.275 86.965 211.445 ;
        RECT 87.865 211.405 88.045 212.165 ;
        RECT 88.225 211.575 88.555 212.335 ;
        RECT 86.025 211.025 86.195 211.275 ;
        RECT 87.335 211.025 87.600 211.385 ;
        RECT 87.865 211.235 88.540 211.405 ;
        RECT 88.725 211.260 88.995 212.165 ;
        RECT 88.370 211.090 88.540 211.235 ;
        RECT 85.905 210.695 86.195 211.025 ;
        RECT 86.365 210.775 86.705 211.025 ;
        RECT 86.925 210.775 87.600 211.025 ;
        RECT 86.025 210.605 86.195 210.695 ;
        RECT 87.805 210.685 88.145 211.055 ;
        RECT 88.370 210.760 88.645 211.090 ;
        RECT 86.025 210.415 87.415 210.605 ;
        RECT 88.370 210.505 88.540 210.760 ;
        RECT 85.485 209.955 86.045 210.245 ;
        RECT 86.215 209.785 86.465 210.245 ;
        RECT 87.085 210.055 87.415 210.415 ;
        RECT 87.875 210.335 88.540 210.505 ;
        RECT 88.815 210.460 88.995 211.260 ;
        RECT 89.165 211.245 90.375 212.335 ;
        RECT 87.875 209.955 88.045 210.335 ;
        RECT 88.225 209.785 88.555 210.165 ;
        RECT 88.735 209.955 88.995 210.460 ;
        RECT 89.165 210.535 89.685 211.075 ;
        RECT 89.855 210.705 90.375 211.245 ;
        RECT 90.585 211.195 90.815 212.335 ;
        RECT 90.985 211.185 91.315 212.165 ;
        RECT 91.485 211.195 91.695 212.335 ;
        RECT 91.925 211.245 94.515 212.335 ;
        RECT 90.565 210.775 90.895 211.025 ;
        RECT 89.165 209.785 90.375 210.535 ;
        RECT 90.585 209.785 90.815 210.605 ;
        RECT 91.065 210.585 91.315 211.185 ;
        RECT 90.985 209.955 91.315 210.585 ;
        RECT 91.485 209.785 91.695 210.605 ;
        RECT 91.925 210.555 93.135 211.075 ;
        RECT 93.305 210.725 94.515 211.245 ;
        RECT 94.685 211.170 94.975 212.335 ;
        RECT 96.070 211.185 96.330 212.335 ;
        RECT 96.505 211.260 96.760 212.165 ;
        RECT 96.930 211.575 97.260 212.335 ;
        RECT 97.475 211.405 97.645 212.165 ;
        RECT 97.905 211.900 103.250 212.335 ;
        RECT 91.925 209.785 94.515 210.555 ;
        RECT 94.685 209.785 94.975 210.510 ;
        RECT 96.070 209.785 96.330 210.625 ;
        RECT 96.505 210.530 96.675 211.260 ;
        RECT 96.930 211.235 97.645 211.405 ;
        RECT 96.930 211.025 97.100 211.235 ;
        RECT 96.845 210.695 97.100 211.025 ;
        RECT 96.505 209.955 96.760 210.530 ;
        RECT 96.930 210.505 97.100 210.695 ;
        RECT 97.380 210.685 97.735 211.055 ;
        RECT 96.930 210.335 97.645 210.505 ;
        RECT 96.930 209.785 97.260 210.165 ;
        RECT 97.475 209.955 97.645 210.335 ;
        RECT 99.490 210.330 99.830 211.160 ;
        RECT 101.310 210.650 101.660 211.900 ;
        RECT 103.425 211.245 106.935 212.335 ;
        RECT 103.425 210.555 105.075 211.075 ;
        RECT 105.245 210.725 106.935 211.245 ;
        RECT 107.565 211.170 107.855 212.335 ;
        RECT 108.025 211.900 113.370 212.335 ;
        RECT 113.545 211.900 118.890 212.335 ;
        RECT 97.905 209.785 103.250 210.330 ;
        RECT 103.425 209.785 106.935 210.555 ;
        RECT 107.565 209.785 107.855 210.510 ;
        RECT 109.610 210.330 109.950 211.160 ;
        RECT 111.430 210.650 111.780 211.900 ;
        RECT 115.130 210.330 115.470 211.160 ;
        RECT 116.950 210.650 117.300 211.900 ;
        RECT 119.065 211.245 120.275 212.335 ;
        RECT 119.065 210.535 119.585 211.075 ;
        RECT 119.755 210.705 120.275 211.245 ;
        RECT 120.445 211.170 120.735 212.335 ;
        RECT 120.905 211.900 126.250 212.335 ;
        RECT 126.425 211.900 131.770 212.335 ;
        RECT 108.025 209.785 113.370 210.330 ;
        RECT 113.545 209.785 118.890 210.330 ;
        RECT 119.065 209.785 120.275 210.535 ;
        RECT 120.445 209.785 120.735 210.510 ;
        RECT 122.490 210.330 122.830 211.160 ;
        RECT 124.310 210.650 124.660 211.900 ;
        RECT 128.010 210.330 128.350 211.160 ;
        RECT 129.830 210.650 130.180 211.900 ;
        RECT 131.945 211.245 133.155 212.335 ;
        RECT 131.945 210.535 132.465 211.075 ;
        RECT 132.635 210.705 133.155 211.245 ;
        RECT 133.325 211.170 133.615 212.335 ;
        RECT 133.785 211.900 139.130 212.335 ;
        RECT 139.305 211.900 144.650 212.335 ;
        RECT 120.905 209.785 126.250 210.330 ;
        RECT 126.425 209.785 131.770 210.330 ;
        RECT 131.945 209.785 133.155 210.535 ;
        RECT 133.325 209.785 133.615 210.510 ;
        RECT 135.370 210.330 135.710 211.160 ;
        RECT 137.190 210.650 137.540 211.900 ;
        RECT 140.890 210.330 141.230 211.160 ;
        RECT 142.710 210.650 143.060 211.900 ;
        RECT 145.745 211.245 146.955 212.335 ;
        RECT 145.745 210.705 146.265 211.245 ;
        RECT 146.435 210.535 146.955 211.075 ;
        RECT 133.785 209.785 139.130 210.330 ;
        RECT 139.305 209.785 144.650 210.330 ;
        RECT 145.745 209.785 146.955 210.535 ;
        RECT 17.320 209.615 147.040 209.785 ;
        RECT 17.405 208.865 18.615 209.615 ;
        RECT 18.785 209.070 24.130 209.615 ;
        RECT 24.305 209.070 29.650 209.615 ;
        RECT 29.825 209.070 35.170 209.615 ;
        RECT 35.345 209.070 40.690 209.615 ;
        RECT 17.405 208.325 17.925 208.865 ;
        RECT 18.095 208.155 18.615 208.695 ;
        RECT 20.370 208.240 20.710 209.070 ;
        RECT 17.405 207.065 18.615 208.155 ;
        RECT 22.190 207.500 22.540 208.750 ;
        RECT 25.890 208.240 26.230 209.070 ;
        RECT 27.710 207.500 28.060 208.750 ;
        RECT 31.410 208.240 31.750 209.070 ;
        RECT 33.230 207.500 33.580 208.750 ;
        RECT 36.930 208.240 37.270 209.070 ;
        RECT 40.865 208.845 42.535 209.615 ;
        RECT 43.165 208.890 43.455 209.615 ;
        RECT 43.625 209.070 48.970 209.615 ;
        RECT 38.750 207.500 39.100 208.750 ;
        RECT 40.865 208.325 41.615 208.845 ;
        RECT 41.785 208.155 42.535 208.675 ;
        RECT 45.210 208.240 45.550 209.070 ;
        RECT 49.145 208.845 51.735 209.615 ;
        RECT 52.435 209.215 52.765 209.615 ;
        RECT 52.935 209.045 53.105 209.315 ;
        RECT 53.275 209.215 53.605 209.615 ;
        RECT 53.775 209.045 54.030 209.315 ;
        RECT 54.275 209.215 54.605 209.615 ;
        RECT 54.775 209.045 54.945 209.315 ;
        RECT 55.115 209.215 55.445 209.615 ;
        RECT 55.615 209.045 55.870 209.315 ;
        RECT 18.785 207.065 24.130 207.500 ;
        RECT 24.305 207.065 29.650 207.500 ;
        RECT 29.825 207.065 35.170 207.500 ;
        RECT 35.345 207.065 40.690 207.500 ;
        RECT 40.865 207.065 42.535 208.155 ;
        RECT 43.165 207.065 43.455 208.230 ;
        RECT 47.030 207.500 47.380 208.750 ;
        RECT 49.145 208.325 50.355 208.845 ;
        RECT 50.525 208.155 51.735 208.675 ;
        RECT 43.625 207.065 48.970 207.500 ;
        RECT 49.145 207.065 51.735 208.155 ;
        RECT 52.365 208.035 52.635 209.045 ;
        RECT 52.805 208.875 54.030 209.045 ;
        RECT 52.805 208.205 52.975 208.875 ;
        RECT 53.145 208.375 53.525 208.705 ;
        RECT 53.695 208.375 54.030 208.705 ;
        RECT 52.805 208.035 53.120 208.205 ;
        RECT 52.370 207.065 52.685 207.865 ;
        RECT 52.950 207.420 53.120 208.035 ;
        RECT 53.290 207.695 53.525 208.375 ;
        RECT 53.695 207.420 54.030 208.205 ;
        RECT 54.205 208.035 54.475 209.045 ;
        RECT 54.645 208.875 55.870 209.045 ;
        RECT 57.080 208.985 57.365 209.445 ;
        RECT 57.535 209.155 57.805 209.615 ;
        RECT 54.645 208.205 54.815 208.875 ;
        RECT 57.080 208.815 58.035 208.985 ;
        RECT 54.985 208.375 55.365 208.705 ;
        RECT 55.535 208.375 55.870 208.705 ;
        RECT 54.645 208.035 54.960 208.205 ;
        RECT 52.950 207.250 54.030 207.420 ;
        RECT 54.210 207.065 54.525 207.865 ;
        RECT 54.790 207.420 54.960 208.035 ;
        RECT 55.130 207.695 55.365 208.375 ;
        RECT 55.535 207.420 55.870 208.205 ;
        RECT 56.965 208.085 57.655 208.645 ;
        RECT 57.825 207.915 58.035 208.815 ;
        RECT 54.790 207.250 55.870 207.420 ;
        RECT 57.080 207.695 58.035 207.915 ;
        RECT 58.205 208.645 58.605 209.445 ;
        RECT 58.795 208.985 59.075 209.445 ;
        RECT 59.595 209.155 59.920 209.615 ;
        RECT 58.795 208.815 59.920 208.985 ;
        RECT 60.090 208.875 60.475 209.445 ;
        RECT 59.470 208.705 59.920 208.815 ;
        RECT 58.205 208.085 59.300 208.645 ;
        RECT 59.470 208.375 60.025 208.705 ;
        RECT 57.080 207.235 57.365 207.695 ;
        RECT 57.535 207.065 57.805 207.525 ;
        RECT 58.205 207.235 58.605 208.085 ;
        RECT 59.470 207.915 59.920 208.375 ;
        RECT 60.195 208.205 60.475 208.875 ;
        RECT 60.665 208.805 60.905 209.615 ;
        RECT 61.075 208.805 61.405 209.445 ;
        RECT 61.575 208.805 61.845 209.615 ;
        RECT 62.025 208.845 65.535 209.615 ;
        RECT 65.705 208.865 66.915 209.615 ;
        RECT 67.095 208.885 67.395 209.615 ;
        RECT 60.645 208.375 60.995 208.625 ;
        RECT 61.165 208.205 61.335 208.805 ;
        RECT 61.505 208.375 61.855 208.625 ;
        RECT 62.025 208.325 63.675 208.845 ;
        RECT 58.795 207.695 59.920 207.915 ;
        RECT 58.795 207.235 59.075 207.695 ;
        RECT 59.595 207.065 59.920 207.525 ;
        RECT 60.090 207.235 60.475 208.205 ;
        RECT 60.655 208.035 61.335 208.205 ;
        RECT 60.655 207.250 60.985 208.035 ;
        RECT 61.515 207.065 61.845 208.205 ;
        RECT 63.845 208.155 65.535 208.675 ;
        RECT 65.705 208.325 66.225 208.865 ;
        RECT 67.575 208.705 67.805 209.325 ;
        RECT 68.005 209.055 68.230 209.435 ;
        RECT 68.400 209.225 68.730 209.615 ;
        RECT 68.005 208.875 68.335 209.055 ;
        RECT 66.395 208.155 66.915 208.695 ;
        RECT 67.100 208.375 67.395 208.705 ;
        RECT 67.575 208.375 67.990 208.705 ;
        RECT 68.160 208.205 68.335 208.875 ;
        RECT 68.505 208.375 68.745 209.025 ;
        RECT 68.925 208.890 69.215 209.615 ;
        RECT 69.405 208.805 69.645 209.615 ;
        RECT 69.815 208.805 70.145 209.445 ;
        RECT 70.315 208.805 70.585 209.615 ;
        RECT 70.765 209.070 76.110 209.615 ;
        RECT 69.385 208.375 69.735 208.625 ;
        RECT 62.025 207.065 65.535 208.155 ;
        RECT 65.705 207.065 66.915 208.155 ;
        RECT 67.095 207.845 67.990 208.175 ;
        RECT 68.160 208.015 68.745 208.205 ;
        RECT 67.095 207.675 68.300 207.845 ;
        RECT 67.095 207.245 67.425 207.675 ;
        RECT 67.605 207.065 67.800 207.505 ;
        RECT 67.970 207.245 68.300 207.675 ;
        RECT 68.470 207.245 68.745 208.015 ;
        RECT 68.925 207.065 69.215 208.230 ;
        RECT 69.905 208.205 70.075 208.805 ;
        RECT 70.245 208.375 70.595 208.625 ;
        RECT 72.350 208.240 72.690 209.070 ;
        RECT 76.285 208.845 79.795 209.615 ;
        RECT 81.000 208.985 81.285 209.445 ;
        RECT 81.455 209.155 81.725 209.615 ;
        RECT 69.395 208.035 70.075 208.205 ;
        RECT 69.395 207.250 69.725 208.035 ;
        RECT 70.255 207.065 70.585 208.205 ;
        RECT 74.170 207.500 74.520 208.750 ;
        RECT 76.285 208.325 77.935 208.845 ;
        RECT 81.000 208.815 81.955 208.985 ;
        RECT 78.105 208.155 79.795 208.675 ;
        RECT 70.765 207.065 76.110 207.500 ;
        RECT 76.285 207.065 79.795 208.155 ;
        RECT 80.885 208.085 81.575 208.645 ;
        RECT 81.745 207.915 81.955 208.815 ;
        RECT 81.000 207.695 81.955 207.915 ;
        RECT 82.125 208.645 82.525 209.445 ;
        RECT 82.715 208.985 82.995 209.445 ;
        RECT 83.515 209.155 83.840 209.615 ;
        RECT 82.715 208.815 83.840 208.985 ;
        RECT 84.010 208.875 84.395 209.445 ;
        RECT 83.390 208.705 83.840 208.815 ;
        RECT 82.125 208.085 83.220 208.645 ;
        RECT 83.390 208.375 83.945 208.705 ;
        RECT 81.000 207.235 81.285 207.695 ;
        RECT 81.455 207.065 81.725 207.525 ;
        RECT 82.125 207.235 82.525 208.085 ;
        RECT 83.390 207.915 83.840 208.375 ;
        RECT 84.115 208.205 84.395 208.875 ;
        RECT 84.565 208.865 85.775 209.615 ;
        RECT 86.060 208.985 86.345 209.445 ;
        RECT 86.515 209.155 86.785 209.615 ;
        RECT 84.565 208.325 85.085 208.865 ;
        RECT 86.060 208.815 87.015 208.985 ;
        RECT 82.715 207.695 83.840 207.915 ;
        RECT 82.715 207.235 82.995 207.695 ;
        RECT 83.515 207.065 83.840 207.525 ;
        RECT 84.010 207.235 84.395 208.205 ;
        RECT 85.255 208.155 85.775 208.695 ;
        RECT 84.565 207.065 85.775 208.155 ;
        RECT 85.945 208.085 86.635 208.645 ;
        RECT 86.805 207.915 87.015 208.815 ;
        RECT 86.060 207.695 87.015 207.915 ;
        RECT 87.185 208.645 87.585 209.445 ;
        RECT 87.775 208.985 88.055 209.445 ;
        RECT 88.575 209.155 88.900 209.615 ;
        RECT 87.775 208.815 88.900 208.985 ;
        RECT 89.070 208.875 89.455 209.445 ;
        RECT 88.450 208.705 88.900 208.815 ;
        RECT 87.185 208.085 88.280 208.645 ;
        RECT 88.450 208.375 89.005 208.705 ;
        RECT 86.060 207.235 86.345 207.695 ;
        RECT 86.515 207.065 86.785 207.525 ;
        RECT 87.185 207.235 87.585 208.085 ;
        RECT 88.450 207.915 88.900 208.375 ;
        RECT 89.175 208.205 89.455 208.875 ;
        RECT 87.775 207.695 88.900 207.915 ;
        RECT 87.775 207.235 88.055 207.695 ;
        RECT 88.575 207.065 88.900 207.525 ;
        RECT 89.070 207.235 89.455 208.205 ;
        RECT 89.635 208.890 89.965 209.400 ;
        RECT 90.135 209.215 90.465 209.615 ;
        RECT 91.515 209.045 91.845 209.385 ;
        RECT 92.015 209.215 92.345 209.615 ;
        RECT 89.635 208.125 89.825 208.890 ;
        RECT 90.135 208.875 92.500 209.045 ;
        RECT 90.135 208.705 90.305 208.875 ;
        RECT 89.995 208.375 90.305 208.705 ;
        RECT 90.475 208.375 90.780 208.705 ;
        RECT 89.635 207.275 89.965 208.125 ;
        RECT 90.135 207.065 90.385 208.205 ;
        RECT 90.565 208.045 90.780 208.375 ;
        RECT 90.955 208.045 91.240 208.705 ;
        RECT 91.435 208.045 91.700 208.705 ;
        RECT 91.915 208.045 92.160 208.705 ;
        RECT 92.330 207.875 92.500 208.875 ;
        RECT 93.305 208.815 93.615 209.615 ;
        RECT 93.820 208.815 94.515 209.445 ;
        RECT 94.685 208.890 94.975 209.615 ;
        RECT 93.315 208.375 93.650 208.645 ;
        RECT 93.820 208.255 93.990 208.815 ;
        RECT 95.145 208.795 95.405 209.615 ;
        RECT 95.575 208.795 95.905 209.215 ;
        RECT 96.085 209.130 96.875 209.395 ;
        RECT 95.655 208.705 95.905 208.795 ;
        RECT 94.160 208.375 94.495 208.625 ;
        RECT 93.820 208.215 93.995 208.255 ;
        RECT 90.575 207.705 91.865 207.875 ;
        RECT 90.575 207.285 90.825 207.705 ;
        RECT 91.055 207.065 91.385 207.535 ;
        RECT 91.615 207.285 91.865 207.705 ;
        RECT 92.045 207.705 92.500 207.875 ;
        RECT 92.045 207.275 92.375 207.705 ;
        RECT 93.305 207.065 93.585 208.205 ;
        RECT 93.755 207.235 94.085 208.215 ;
        RECT 94.255 207.065 94.515 208.205 ;
        RECT 94.685 207.065 94.975 208.230 ;
        RECT 95.145 207.745 95.485 208.625 ;
        RECT 95.655 208.455 96.450 208.705 ;
        RECT 95.145 207.065 95.405 207.575 ;
        RECT 95.655 207.235 95.825 208.455 ;
        RECT 96.620 208.275 96.875 209.130 ;
        RECT 97.045 208.975 97.245 209.395 ;
        RECT 97.435 209.155 97.765 209.615 ;
        RECT 97.045 208.455 97.455 208.975 ;
        RECT 97.935 208.965 98.195 209.445 ;
        RECT 97.625 208.275 97.855 208.705 ;
        RECT 96.065 208.105 97.855 208.275 ;
        RECT 96.065 207.740 96.315 208.105 ;
        RECT 96.485 207.745 96.815 207.935 ;
        RECT 97.035 207.810 97.750 208.105 ;
        RECT 98.025 207.935 98.195 208.965 ;
        RECT 96.485 207.570 96.680 207.745 ;
        RECT 96.065 207.065 96.680 207.570 ;
        RECT 96.850 207.235 97.325 207.575 ;
        RECT 97.495 207.065 97.710 207.610 ;
        RECT 97.920 207.235 98.195 207.935 ;
        RECT 99.285 208.875 99.750 209.420 ;
        RECT 99.285 207.915 99.455 208.875 ;
        RECT 100.255 208.795 100.425 209.615 ;
        RECT 100.595 208.965 100.925 209.445 ;
        RECT 101.095 209.225 101.445 209.615 ;
        RECT 101.615 209.045 101.845 209.445 ;
        RECT 101.335 208.965 101.845 209.045 ;
        RECT 100.595 208.875 101.845 208.965 ;
        RECT 102.015 208.875 102.335 209.355 ;
        RECT 102.670 209.105 102.910 209.615 ;
        RECT 103.090 209.105 103.370 209.435 ;
        RECT 103.600 209.105 103.815 209.615 ;
        RECT 100.595 208.795 101.505 208.875 ;
        RECT 99.625 208.255 99.870 208.705 ;
        RECT 100.130 208.425 100.825 208.625 ;
        RECT 100.995 208.455 101.595 208.625 ;
        RECT 100.995 208.255 101.165 208.455 ;
        RECT 101.825 208.285 101.995 208.705 ;
        RECT 99.625 208.085 101.165 208.255 ;
        RECT 101.335 208.115 101.995 208.285 ;
        RECT 101.335 207.915 101.505 208.115 ;
        RECT 102.165 207.945 102.335 208.875 ;
        RECT 102.565 208.375 102.920 208.935 ;
        RECT 103.090 208.205 103.260 209.105 ;
        RECT 103.430 208.375 103.695 208.935 ;
        RECT 103.985 208.875 104.600 209.445 ;
        RECT 104.805 209.070 110.150 209.615 ;
        RECT 110.325 209.070 115.670 209.615 ;
        RECT 103.945 208.205 104.115 208.705 ;
        RECT 99.285 207.745 101.505 207.915 ;
        RECT 101.675 207.745 102.335 207.945 ;
        RECT 102.690 208.035 104.115 208.205 ;
        RECT 102.690 207.860 103.080 208.035 ;
        RECT 99.285 207.065 99.585 207.575 ;
        RECT 99.755 207.235 100.085 207.745 ;
        RECT 101.675 207.575 101.845 207.745 ;
        RECT 100.255 207.065 100.885 207.575 ;
        RECT 101.465 207.405 101.845 207.575 ;
        RECT 102.015 207.065 102.315 207.575 ;
        RECT 103.565 207.065 103.895 207.865 ;
        RECT 104.285 207.855 104.600 208.875 ;
        RECT 106.390 208.240 106.730 209.070 ;
        RECT 104.065 207.235 104.600 207.855 ;
        RECT 108.210 207.500 108.560 208.750 ;
        RECT 111.910 208.240 112.250 209.070 ;
        RECT 115.845 208.845 119.355 209.615 ;
        RECT 120.445 208.890 120.735 209.615 ;
        RECT 120.905 209.070 126.250 209.615 ;
        RECT 126.425 209.070 131.770 209.615 ;
        RECT 131.945 209.070 137.290 209.615 ;
        RECT 137.465 209.070 142.810 209.615 ;
        RECT 113.730 207.500 114.080 208.750 ;
        RECT 115.845 208.325 117.495 208.845 ;
        RECT 117.665 208.155 119.355 208.675 ;
        RECT 122.490 208.240 122.830 209.070 ;
        RECT 104.805 207.065 110.150 207.500 ;
        RECT 110.325 207.065 115.670 207.500 ;
        RECT 115.845 207.065 119.355 208.155 ;
        RECT 120.445 207.065 120.735 208.230 ;
        RECT 124.310 207.500 124.660 208.750 ;
        RECT 128.010 208.240 128.350 209.070 ;
        RECT 129.830 207.500 130.180 208.750 ;
        RECT 133.530 208.240 133.870 209.070 ;
        RECT 135.350 207.500 135.700 208.750 ;
        RECT 139.050 208.240 139.390 209.070 ;
        RECT 142.985 208.845 145.575 209.615 ;
        RECT 145.745 208.865 146.955 209.615 ;
        RECT 140.870 207.500 141.220 208.750 ;
        RECT 142.985 208.325 144.195 208.845 ;
        RECT 144.365 208.155 145.575 208.675 ;
        RECT 120.905 207.065 126.250 207.500 ;
        RECT 126.425 207.065 131.770 207.500 ;
        RECT 131.945 207.065 137.290 207.500 ;
        RECT 137.465 207.065 142.810 207.500 ;
        RECT 142.985 207.065 145.575 208.155 ;
        RECT 145.745 208.155 146.265 208.695 ;
        RECT 146.435 208.325 146.955 208.865 ;
        RECT 145.745 207.065 146.955 208.155 ;
        RECT 17.320 206.895 147.040 207.065 ;
        RECT 17.405 205.805 18.615 206.895 ;
        RECT 18.785 206.460 24.130 206.895 ;
        RECT 24.305 206.460 29.650 206.895 ;
        RECT 17.405 205.095 17.925 205.635 ;
        RECT 18.095 205.265 18.615 205.805 ;
        RECT 17.405 204.345 18.615 205.095 ;
        RECT 20.370 204.890 20.710 205.720 ;
        RECT 22.190 205.210 22.540 206.460 ;
        RECT 25.890 204.890 26.230 205.720 ;
        RECT 27.710 205.210 28.060 206.460 ;
        RECT 30.285 205.730 30.575 206.895 ;
        RECT 30.745 206.460 36.090 206.895 ;
        RECT 36.265 206.460 41.610 206.895 ;
        RECT 41.785 206.460 47.130 206.895 ;
        RECT 18.785 204.345 24.130 204.890 ;
        RECT 24.305 204.345 29.650 204.890 ;
        RECT 30.285 204.345 30.575 205.070 ;
        RECT 32.330 204.890 32.670 205.720 ;
        RECT 34.150 205.210 34.500 206.460 ;
        RECT 37.850 204.890 38.190 205.720 ;
        RECT 39.670 205.210 40.020 206.460 ;
        RECT 43.370 204.890 43.710 205.720 ;
        RECT 45.190 205.210 45.540 206.460 ;
        RECT 47.305 205.805 48.975 206.895 ;
        RECT 47.305 205.115 48.055 205.635 ;
        RECT 48.225 205.285 48.975 205.805 ;
        RECT 49.145 205.755 49.530 206.725 ;
        RECT 49.700 206.435 50.025 206.895 ;
        RECT 50.545 206.265 50.825 206.725 ;
        RECT 49.700 206.045 50.825 206.265 ;
        RECT 30.745 204.345 36.090 204.890 ;
        RECT 36.265 204.345 41.610 204.890 ;
        RECT 41.785 204.345 47.130 204.890 ;
        RECT 47.305 204.345 48.975 205.115 ;
        RECT 49.145 205.085 49.425 205.755 ;
        RECT 49.700 205.585 50.150 206.045 ;
        RECT 51.015 205.875 51.415 206.725 ;
        RECT 51.815 206.435 52.085 206.895 ;
        RECT 52.255 206.265 52.540 206.725 ;
        RECT 52.845 206.385 53.145 206.895 ;
        RECT 53.315 206.385 53.695 206.555 ;
        RECT 54.275 206.385 54.905 206.895 ;
        RECT 49.595 205.255 50.150 205.585 ;
        RECT 50.320 205.315 51.415 205.875 ;
        RECT 49.700 205.145 50.150 205.255 ;
        RECT 49.145 204.515 49.530 205.085 ;
        RECT 49.700 204.975 50.825 205.145 ;
        RECT 49.700 204.345 50.025 204.805 ;
        RECT 50.545 204.515 50.825 204.975 ;
        RECT 51.015 204.515 51.415 205.315 ;
        RECT 51.585 206.045 52.540 206.265 ;
        RECT 53.315 206.215 53.485 206.385 ;
        RECT 55.075 206.215 55.405 206.725 ;
        RECT 55.575 206.385 55.875 206.895 ;
        RECT 51.585 205.145 51.795 206.045 ;
        RECT 52.825 206.015 53.485 206.215 ;
        RECT 53.655 206.045 55.875 206.215 ;
        RECT 51.965 205.315 52.655 205.875 ;
        RECT 51.585 204.975 52.540 205.145 ;
        RECT 51.815 204.345 52.085 204.805 ;
        RECT 52.255 204.515 52.540 204.975 ;
        RECT 52.825 205.085 52.995 206.015 ;
        RECT 53.655 205.845 53.825 206.045 ;
        RECT 53.165 205.675 53.825 205.845 ;
        RECT 53.995 205.705 55.535 205.875 ;
        RECT 53.165 205.255 53.335 205.675 ;
        RECT 53.995 205.505 54.165 205.705 ;
        RECT 53.565 205.335 54.165 205.505 ;
        RECT 54.335 205.335 55.030 205.535 ;
        RECT 55.290 205.255 55.535 205.705 ;
        RECT 53.655 205.085 54.565 205.165 ;
        RECT 52.825 204.605 53.145 205.085 ;
        RECT 53.315 204.995 54.565 205.085 ;
        RECT 53.315 204.915 53.825 204.995 ;
        RECT 53.315 204.515 53.545 204.915 ;
        RECT 53.715 204.345 54.065 204.735 ;
        RECT 54.235 204.515 54.565 204.995 ;
        RECT 54.735 204.345 54.905 205.165 ;
        RECT 55.705 205.085 55.875 206.045 ;
        RECT 56.045 205.730 56.335 206.895 ;
        RECT 56.565 205.835 56.895 206.680 ;
        RECT 57.065 205.885 57.235 206.895 ;
        RECT 57.405 206.165 57.745 206.725 ;
        RECT 57.975 206.395 58.290 206.895 ;
        RECT 58.470 206.425 59.355 206.595 ;
        RECT 56.505 205.755 56.895 205.835 ;
        RECT 57.405 205.790 58.300 206.165 ;
        RECT 55.410 204.540 55.875 205.085 ;
        RECT 56.505 205.705 56.720 205.755 ;
        RECT 56.505 205.125 56.675 205.705 ;
        RECT 57.405 205.585 57.595 205.790 ;
        RECT 58.470 205.585 58.640 206.425 ;
        RECT 59.580 206.395 59.830 206.725 ;
        RECT 56.845 205.255 57.595 205.585 ;
        RECT 57.765 205.255 58.640 205.585 ;
        RECT 56.505 205.085 56.730 205.125 ;
        RECT 57.395 205.085 57.595 205.255 ;
        RECT 56.045 204.345 56.335 205.070 ;
        RECT 56.505 205.000 56.885 205.085 ;
        RECT 56.555 204.565 56.885 205.000 ;
        RECT 57.055 204.345 57.225 204.955 ;
        RECT 57.395 204.560 57.725 205.085 ;
        RECT 57.985 204.345 58.195 204.875 ;
        RECT 58.470 204.795 58.640 205.255 ;
        RECT 58.810 205.295 59.130 206.255 ;
        RECT 59.300 205.505 59.490 206.225 ;
        RECT 59.660 205.325 59.830 206.395 ;
        RECT 60.000 206.095 60.170 206.895 ;
        RECT 60.340 206.450 61.445 206.620 ;
        RECT 60.340 205.835 60.510 206.450 ;
        RECT 61.655 206.300 61.905 206.725 ;
        RECT 62.075 206.435 62.340 206.895 ;
        RECT 60.680 205.915 61.210 206.280 ;
        RECT 61.655 206.170 61.960 206.300 ;
        RECT 60.000 205.745 60.510 205.835 ;
        RECT 60.000 205.575 60.870 205.745 ;
        RECT 60.000 205.505 60.170 205.575 ;
        RECT 60.290 205.325 60.490 205.355 ;
        RECT 58.810 204.965 59.275 205.295 ;
        RECT 59.660 205.025 60.490 205.325 ;
        RECT 59.660 204.795 59.830 205.025 ;
        RECT 58.470 204.625 59.255 204.795 ;
        RECT 59.425 204.625 59.830 204.795 ;
        RECT 60.010 204.345 60.380 204.845 ;
        RECT 60.700 204.795 60.870 205.575 ;
        RECT 61.040 205.215 61.210 205.915 ;
        RECT 61.380 205.385 61.620 205.980 ;
        RECT 61.040 204.995 61.565 205.215 ;
        RECT 61.790 205.065 61.960 206.170 ;
        RECT 61.735 204.935 61.960 205.065 ;
        RECT 62.130 204.975 62.410 205.925 ;
        RECT 61.735 204.795 61.905 204.935 ;
        RECT 60.700 204.625 61.375 204.795 ;
        RECT 61.570 204.625 61.905 204.795 ;
        RECT 62.075 204.345 62.325 204.805 ;
        RECT 62.580 204.605 62.765 206.725 ;
        RECT 62.935 206.395 63.265 206.895 ;
        RECT 63.435 206.225 63.605 206.725 ;
        RECT 62.940 206.055 63.605 206.225 ;
        RECT 62.940 205.065 63.170 206.055 ;
        RECT 63.340 205.235 63.690 205.885 ;
        RECT 64.385 205.835 64.715 206.680 ;
        RECT 64.885 205.885 65.055 206.895 ;
        RECT 65.225 206.165 65.565 206.725 ;
        RECT 65.795 206.395 66.110 206.895 ;
        RECT 66.290 206.425 67.175 206.595 ;
        RECT 64.325 205.755 64.715 205.835 ;
        RECT 65.225 205.790 66.120 206.165 ;
        RECT 64.325 205.705 64.540 205.755 ;
        RECT 64.325 205.125 64.495 205.705 ;
        RECT 65.225 205.585 65.415 205.790 ;
        RECT 66.290 205.585 66.460 206.425 ;
        RECT 67.400 206.395 67.650 206.725 ;
        RECT 64.665 205.255 65.415 205.585 ;
        RECT 65.585 205.255 66.460 205.585 ;
        RECT 64.325 205.085 64.550 205.125 ;
        RECT 65.215 205.085 65.415 205.255 ;
        RECT 62.940 204.895 63.605 205.065 ;
        RECT 64.325 205.000 64.705 205.085 ;
        RECT 62.935 204.345 63.265 204.725 ;
        RECT 63.435 204.605 63.605 204.895 ;
        RECT 64.375 204.565 64.705 205.000 ;
        RECT 64.875 204.345 65.045 204.955 ;
        RECT 65.215 204.560 65.545 205.085 ;
        RECT 65.805 204.345 66.015 204.875 ;
        RECT 66.290 204.795 66.460 205.255 ;
        RECT 66.630 205.295 66.950 206.255 ;
        RECT 67.120 205.505 67.310 206.225 ;
        RECT 67.480 205.325 67.650 206.395 ;
        RECT 67.820 206.095 67.990 206.895 ;
        RECT 68.160 206.450 69.265 206.620 ;
        RECT 68.160 205.835 68.330 206.450 ;
        RECT 69.475 206.300 69.725 206.725 ;
        RECT 69.895 206.435 70.160 206.895 ;
        RECT 68.500 205.915 69.030 206.280 ;
        RECT 69.475 206.170 69.780 206.300 ;
        RECT 67.820 205.745 68.330 205.835 ;
        RECT 67.820 205.575 68.690 205.745 ;
        RECT 67.820 205.505 67.990 205.575 ;
        RECT 68.110 205.325 68.310 205.355 ;
        RECT 66.630 204.965 67.095 205.295 ;
        RECT 67.480 205.025 68.310 205.325 ;
        RECT 67.480 204.795 67.650 205.025 ;
        RECT 66.290 204.625 67.075 204.795 ;
        RECT 67.245 204.625 67.650 204.795 ;
        RECT 67.830 204.345 68.200 204.845 ;
        RECT 68.520 204.795 68.690 205.575 ;
        RECT 68.860 205.215 69.030 205.915 ;
        RECT 69.200 205.385 69.440 205.980 ;
        RECT 68.860 204.995 69.385 205.215 ;
        RECT 69.610 205.065 69.780 206.170 ;
        RECT 69.555 204.935 69.780 205.065 ;
        RECT 69.950 204.975 70.230 205.925 ;
        RECT 69.555 204.795 69.725 204.935 ;
        RECT 68.520 204.625 69.195 204.795 ;
        RECT 69.390 204.625 69.725 204.795 ;
        RECT 69.895 204.345 70.145 204.805 ;
        RECT 70.400 204.605 70.585 206.725 ;
        RECT 70.755 206.395 71.085 206.895 ;
        RECT 71.255 206.225 71.425 206.725 ;
        RECT 71.685 206.460 77.030 206.895 ;
        RECT 70.760 206.055 71.425 206.225 ;
        RECT 70.760 205.065 70.990 206.055 ;
        RECT 71.160 205.235 71.510 205.885 ;
        RECT 70.760 204.895 71.425 205.065 ;
        RECT 70.755 204.345 71.085 204.725 ;
        RECT 71.255 204.605 71.425 204.895 ;
        RECT 73.270 204.890 73.610 205.720 ;
        RECT 75.090 205.210 75.440 206.460 ;
        RECT 77.205 205.805 80.715 206.895 ;
        RECT 77.205 205.115 78.855 205.635 ;
        RECT 79.025 205.285 80.715 205.805 ;
        RECT 81.805 205.730 82.095 206.895 ;
        RECT 82.785 205.835 83.115 206.680 ;
        RECT 83.285 205.885 83.455 206.895 ;
        RECT 83.625 206.165 83.965 206.725 ;
        RECT 84.195 206.395 84.510 206.895 ;
        RECT 84.690 206.425 85.575 206.595 ;
        RECT 82.725 205.755 83.115 205.835 ;
        RECT 83.625 205.790 84.520 206.165 ;
        RECT 82.725 205.705 82.940 205.755 ;
        RECT 82.725 205.125 82.895 205.705 ;
        RECT 83.625 205.585 83.815 205.790 ;
        RECT 84.690 205.585 84.860 206.425 ;
        RECT 85.800 206.395 86.050 206.725 ;
        RECT 83.065 205.255 83.815 205.585 ;
        RECT 83.985 205.255 84.860 205.585 ;
        RECT 71.685 204.345 77.030 204.890 ;
        RECT 77.205 204.345 80.715 205.115 ;
        RECT 82.725 205.085 82.950 205.125 ;
        RECT 83.615 205.085 83.815 205.255 ;
        RECT 81.805 204.345 82.095 205.070 ;
        RECT 82.725 205.000 83.105 205.085 ;
        RECT 82.775 204.565 83.105 205.000 ;
        RECT 83.275 204.345 83.445 204.955 ;
        RECT 83.615 204.560 83.945 205.085 ;
        RECT 84.205 204.345 84.415 204.875 ;
        RECT 84.690 204.795 84.860 205.255 ;
        RECT 85.030 205.295 85.350 206.255 ;
        RECT 85.520 205.505 85.710 206.225 ;
        RECT 85.880 205.325 86.050 206.395 ;
        RECT 86.220 206.095 86.390 206.895 ;
        RECT 86.560 206.450 87.665 206.620 ;
        RECT 86.560 205.835 86.730 206.450 ;
        RECT 87.875 206.300 88.125 206.725 ;
        RECT 88.295 206.435 88.560 206.895 ;
        RECT 86.900 205.915 87.430 206.280 ;
        RECT 87.875 206.170 88.180 206.300 ;
        RECT 86.220 205.745 86.730 205.835 ;
        RECT 86.220 205.575 87.090 205.745 ;
        RECT 86.220 205.505 86.390 205.575 ;
        RECT 86.510 205.325 86.710 205.355 ;
        RECT 85.030 204.965 85.495 205.295 ;
        RECT 85.880 205.025 86.710 205.325 ;
        RECT 85.880 204.795 86.050 205.025 ;
        RECT 84.690 204.625 85.475 204.795 ;
        RECT 85.645 204.625 86.050 204.795 ;
        RECT 86.230 204.345 86.600 204.845 ;
        RECT 86.920 204.795 87.090 205.575 ;
        RECT 87.260 205.215 87.430 205.915 ;
        RECT 87.600 205.385 87.840 205.980 ;
        RECT 87.260 204.995 87.785 205.215 ;
        RECT 88.010 205.065 88.180 206.170 ;
        RECT 87.955 204.935 88.180 205.065 ;
        RECT 88.350 204.975 88.630 205.925 ;
        RECT 87.955 204.795 88.125 204.935 ;
        RECT 86.920 204.625 87.595 204.795 ;
        RECT 87.790 204.625 88.125 204.795 ;
        RECT 88.295 204.345 88.545 204.805 ;
        RECT 88.800 204.605 88.985 206.725 ;
        RECT 89.155 206.395 89.485 206.895 ;
        RECT 89.655 206.225 89.825 206.725 ;
        RECT 89.160 206.055 89.825 206.225 ;
        RECT 90.175 206.225 90.345 206.725 ;
        RECT 90.515 206.395 90.845 206.895 ;
        RECT 90.175 206.055 90.840 206.225 ;
        RECT 89.160 205.065 89.390 206.055 ;
        RECT 89.560 205.235 89.910 205.885 ;
        RECT 90.090 205.235 90.440 205.885 ;
        RECT 90.610 205.065 90.840 206.055 ;
        RECT 89.160 204.895 89.825 205.065 ;
        RECT 89.155 204.345 89.485 204.725 ;
        RECT 89.655 204.605 89.825 204.895 ;
        RECT 90.175 204.895 90.840 205.065 ;
        RECT 90.175 204.605 90.345 204.895 ;
        RECT 90.515 204.345 90.845 204.725 ;
        RECT 91.015 204.605 91.200 206.725 ;
        RECT 91.440 206.435 91.705 206.895 ;
        RECT 91.875 206.300 92.125 206.725 ;
        RECT 92.335 206.450 93.440 206.620 ;
        RECT 91.820 206.170 92.125 206.300 ;
        RECT 91.370 204.975 91.650 205.925 ;
        RECT 91.820 205.065 91.990 206.170 ;
        RECT 92.160 205.385 92.400 205.980 ;
        RECT 92.570 205.915 93.100 206.280 ;
        RECT 92.570 205.215 92.740 205.915 ;
        RECT 93.270 205.835 93.440 206.450 ;
        RECT 93.610 206.095 93.780 206.895 ;
        RECT 93.950 206.395 94.200 206.725 ;
        RECT 94.425 206.425 95.310 206.595 ;
        RECT 93.270 205.745 93.780 205.835 ;
        RECT 91.820 204.935 92.045 205.065 ;
        RECT 92.215 204.995 92.740 205.215 ;
        RECT 92.910 205.575 93.780 205.745 ;
        RECT 91.455 204.345 91.705 204.805 ;
        RECT 91.875 204.795 92.045 204.935 ;
        RECT 92.910 204.795 93.080 205.575 ;
        RECT 93.610 205.505 93.780 205.575 ;
        RECT 93.290 205.325 93.490 205.355 ;
        RECT 93.950 205.325 94.120 206.395 ;
        RECT 94.290 205.505 94.480 206.225 ;
        RECT 93.290 205.025 94.120 205.325 ;
        RECT 94.650 205.295 94.970 206.255 ;
        RECT 91.875 204.625 92.210 204.795 ;
        RECT 92.405 204.625 93.080 204.795 ;
        RECT 93.400 204.345 93.770 204.845 ;
        RECT 93.950 204.795 94.120 205.025 ;
        RECT 94.505 204.965 94.970 205.295 ;
        RECT 95.140 205.585 95.310 206.425 ;
        RECT 95.490 206.395 95.805 206.895 ;
        RECT 96.035 206.165 96.375 206.725 ;
        RECT 95.480 205.790 96.375 206.165 ;
        RECT 96.545 205.885 96.715 206.895 ;
        RECT 96.185 205.585 96.375 205.790 ;
        RECT 96.885 205.835 97.215 206.680 ;
        RECT 97.535 206.225 97.705 206.725 ;
        RECT 97.875 206.395 98.205 206.895 ;
        RECT 97.535 206.055 98.200 206.225 ;
        RECT 96.885 205.755 97.275 205.835 ;
        RECT 97.060 205.705 97.275 205.755 ;
        RECT 95.140 205.255 96.015 205.585 ;
        RECT 96.185 205.255 96.935 205.585 ;
        RECT 95.140 204.795 95.310 205.255 ;
        RECT 96.185 205.085 96.385 205.255 ;
        RECT 97.105 205.125 97.275 205.705 ;
        RECT 97.450 205.235 97.800 205.885 ;
        RECT 97.050 205.085 97.275 205.125 ;
        RECT 93.950 204.625 94.355 204.795 ;
        RECT 94.525 204.625 95.310 204.795 ;
        RECT 95.585 204.345 95.795 204.875 ;
        RECT 96.055 204.560 96.385 205.085 ;
        RECT 96.895 205.000 97.275 205.085 ;
        RECT 97.970 205.065 98.200 206.055 ;
        RECT 96.555 204.345 96.725 204.955 ;
        RECT 96.895 204.565 97.225 205.000 ;
        RECT 97.535 204.895 98.200 205.065 ;
        RECT 97.535 204.605 97.705 204.895 ;
        RECT 97.875 204.345 98.205 204.725 ;
        RECT 98.375 204.605 98.560 206.725 ;
        RECT 98.800 206.435 99.065 206.895 ;
        RECT 99.235 206.300 99.485 206.725 ;
        RECT 99.695 206.450 100.800 206.620 ;
        RECT 99.180 206.170 99.485 206.300 ;
        RECT 98.730 204.975 99.010 205.925 ;
        RECT 99.180 205.065 99.350 206.170 ;
        RECT 99.520 205.385 99.760 205.980 ;
        RECT 99.930 205.915 100.460 206.280 ;
        RECT 99.930 205.215 100.100 205.915 ;
        RECT 100.630 205.835 100.800 206.450 ;
        RECT 100.970 206.095 101.140 206.895 ;
        RECT 101.310 206.395 101.560 206.725 ;
        RECT 101.785 206.425 102.670 206.595 ;
        RECT 100.630 205.745 101.140 205.835 ;
        RECT 99.180 204.935 99.405 205.065 ;
        RECT 99.575 204.995 100.100 205.215 ;
        RECT 100.270 205.575 101.140 205.745 ;
        RECT 98.815 204.345 99.065 204.805 ;
        RECT 99.235 204.795 99.405 204.935 ;
        RECT 100.270 204.795 100.440 205.575 ;
        RECT 100.970 205.505 101.140 205.575 ;
        RECT 100.650 205.325 100.850 205.355 ;
        RECT 101.310 205.325 101.480 206.395 ;
        RECT 101.650 205.505 101.840 206.225 ;
        RECT 100.650 205.025 101.480 205.325 ;
        RECT 102.010 205.295 102.330 206.255 ;
        RECT 99.235 204.625 99.570 204.795 ;
        RECT 99.765 204.625 100.440 204.795 ;
        RECT 100.760 204.345 101.130 204.845 ;
        RECT 101.310 204.795 101.480 205.025 ;
        RECT 101.865 204.965 102.330 205.295 ;
        RECT 102.500 205.585 102.670 206.425 ;
        RECT 102.850 206.395 103.165 206.895 ;
        RECT 103.395 206.165 103.735 206.725 ;
        RECT 102.840 205.790 103.735 206.165 ;
        RECT 103.905 205.885 104.075 206.895 ;
        RECT 103.545 205.585 103.735 205.790 ;
        RECT 104.245 205.835 104.575 206.680 ;
        RECT 104.860 206.025 105.145 206.895 ;
        RECT 105.315 206.265 105.575 206.725 ;
        RECT 105.750 206.435 106.005 206.895 ;
        RECT 106.175 206.265 106.435 206.725 ;
        RECT 105.315 206.095 106.435 206.265 ;
        RECT 106.605 206.095 106.915 206.895 ;
        RECT 105.315 205.845 105.575 206.095 ;
        RECT 107.085 205.925 107.395 206.725 ;
        RECT 104.245 205.755 104.635 205.835 ;
        RECT 104.420 205.705 104.635 205.755 ;
        RECT 102.500 205.255 103.375 205.585 ;
        RECT 103.545 205.255 104.295 205.585 ;
        RECT 102.500 204.795 102.670 205.255 ;
        RECT 103.545 205.085 103.745 205.255 ;
        RECT 104.465 205.125 104.635 205.705 ;
        RECT 104.410 205.085 104.635 205.125 ;
        RECT 101.310 204.625 101.715 204.795 ;
        RECT 101.885 204.625 102.670 204.795 ;
        RECT 102.945 204.345 103.155 204.875 ;
        RECT 103.415 204.560 103.745 205.085 ;
        RECT 104.255 205.000 104.635 205.085 ;
        RECT 104.820 205.675 105.575 205.845 ;
        RECT 106.365 205.755 107.395 205.925 ;
        RECT 104.820 205.165 105.225 205.675 ;
        RECT 106.365 205.505 106.535 205.755 ;
        RECT 105.395 205.335 106.535 205.505 ;
        RECT 103.915 204.345 104.085 204.955 ;
        RECT 104.255 204.565 104.585 205.000 ;
        RECT 104.820 204.995 106.470 205.165 ;
        RECT 106.705 205.015 107.055 205.585 ;
        RECT 104.865 204.345 105.145 204.825 ;
        RECT 105.315 204.605 105.575 204.995 ;
        RECT 105.750 204.345 106.005 204.825 ;
        RECT 106.175 204.605 106.470 204.995 ;
        RECT 107.225 204.845 107.395 205.755 ;
        RECT 107.565 205.730 107.855 206.895 ;
        RECT 108.025 206.460 113.370 206.895 ;
        RECT 113.545 206.460 118.890 206.895 ;
        RECT 119.065 206.460 124.410 206.895 ;
        RECT 124.585 206.460 129.930 206.895 ;
        RECT 106.650 204.345 106.925 204.825 ;
        RECT 107.095 204.515 107.395 204.845 ;
        RECT 107.565 204.345 107.855 205.070 ;
        RECT 109.610 204.890 109.950 205.720 ;
        RECT 111.430 205.210 111.780 206.460 ;
        RECT 115.130 204.890 115.470 205.720 ;
        RECT 116.950 205.210 117.300 206.460 ;
        RECT 120.650 204.890 120.990 205.720 ;
        RECT 122.470 205.210 122.820 206.460 ;
        RECT 126.170 204.890 126.510 205.720 ;
        RECT 127.990 205.210 128.340 206.460 ;
        RECT 130.105 205.805 132.695 206.895 ;
        RECT 130.105 205.115 131.315 205.635 ;
        RECT 131.485 205.285 132.695 205.805 ;
        RECT 133.325 205.730 133.615 206.895 ;
        RECT 133.785 206.460 139.130 206.895 ;
        RECT 139.305 206.460 144.650 206.895 ;
        RECT 108.025 204.345 113.370 204.890 ;
        RECT 113.545 204.345 118.890 204.890 ;
        RECT 119.065 204.345 124.410 204.890 ;
        RECT 124.585 204.345 129.930 204.890 ;
        RECT 130.105 204.345 132.695 205.115 ;
        RECT 133.325 204.345 133.615 205.070 ;
        RECT 135.370 204.890 135.710 205.720 ;
        RECT 137.190 205.210 137.540 206.460 ;
        RECT 140.890 204.890 141.230 205.720 ;
        RECT 142.710 205.210 143.060 206.460 ;
        RECT 145.745 205.805 146.955 206.895 ;
        RECT 145.745 205.265 146.265 205.805 ;
        RECT 146.435 205.095 146.955 205.635 ;
        RECT 133.785 204.345 139.130 204.890 ;
        RECT 139.305 204.345 144.650 204.890 ;
        RECT 145.745 204.345 146.955 205.095 ;
        RECT 17.320 204.175 147.040 204.345 ;
        RECT 17.405 203.425 18.615 204.175 ;
        RECT 18.785 203.630 24.130 204.175 ;
        RECT 24.305 203.630 29.650 204.175 ;
        RECT 29.825 203.630 35.170 204.175 ;
        RECT 35.345 203.630 40.690 204.175 ;
        RECT 17.405 202.885 17.925 203.425 ;
        RECT 18.095 202.715 18.615 203.255 ;
        RECT 20.370 202.800 20.710 203.630 ;
        RECT 17.405 201.625 18.615 202.715 ;
        RECT 22.190 202.060 22.540 203.310 ;
        RECT 25.890 202.800 26.230 203.630 ;
        RECT 27.710 202.060 28.060 203.310 ;
        RECT 31.410 202.800 31.750 203.630 ;
        RECT 33.230 202.060 33.580 203.310 ;
        RECT 36.930 202.800 37.270 203.630 ;
        RECT 40.865 203.405 42.535 204.175 ;
        RECT 43.165 203.450 43.455 204.175 ;
        RECT 43.625 203.425 44.835 204.175 ;
        RECT 38.750 202.060 39.100 203.310 ;
        RECT 40.865 202.885 41.615 203.405 ;
        RECT 41.785 202.715 42.535 203.235 ;
        RECT 43.625 202.885 44.145 203.425 ;
        RECT 45.015 203.365 45.285 204.175 ;
        RECT 45.455 203.365 45.785 204.005 ;
        RECT 45.955 203.365 46.195 204.175 ;
        RECT 46.475 203.625 46.645 203.915 ;
        RECT 46.815 203.795 47.145 204.175 ;
        RECT 46.475 203.455 47.140 203.625 ;
        RECT 18.785 201.625 24.130 202.060 ;
        RECT 24.305 201.625 29.650 202.060 ;
        RECT 29.825 201.625 35.170 202.060 ;
        RECT 35.345 201.625 40.690 202.060 ;
        RECT 40.865 201.625 42.535 202.715 ;
        RECT 43.165 201.625 43.455 202.790 ;
        RECT 44.315 202.715 44.835 203.255 ;
        RECT 45.005 202.935 45.355 203.185 ;
        RECT 45.525 202.765 45.695 203.365 ;
        RECT 45.865 202.935 46.215 203.185 ;
        RECT 43.625 201.625 44.835 202.715 ;
        RECT 45.015 201.625 45.345 202.765 ;
        RECT 45.525 202.595 46.205 202.765 ;
        RECT 46.390 202.635 46.740 203.285 ;
        RECT 45.875 201.810 46.205 202.595 ;
        RECT 46.910 202.465 47.140 203.455 ;
        RECT 46.475 202.295 47.140 202.465 ;
        RECT 46.475 201.795 46.645 202.295 ;
        RECT 46.815 201.625 47.145 202.125 ;
        RECT 47.315 201.795 47.500 203.915 ;
        RECT 47.755 203.715 48.005 204.175 ;
        RECT 48.175 203.725 48.510 203.895 ;
        RECT 48.705 203.725 49.380 203.895 ;
        RECT 48.175 203.585 48.345 203.725 ;
        RECT 47.670 202.595 47.950 203.545 ;
        RECT 48.120 203.455 48.345 203.585 ;
        RECT 48.120 202.350 48.290 203.455 ;
        RECT 48.515 203.305 49.040 203.525 ;
        RECT 48.460 202.540 48.700 203.135 ;
        RECT 48.870 202.605 49.040 203.305 ;
        RECT 49.210 202.945 49.380 203.725 ;
        RECT 49.700 203.675 50.070 204.175 ;
        RECT 50.250 203.725 50.655 203.895 ;
        RECT 50.825 203.725 51.610 203.895 ;
        RECT 50.250 203.495 50.420 203.725 ;
        RECT 49.590 203.195 50.420 203.495 ;
        RECT 50.805 203.225 51.270 203.555 ;
        RECT 49.590 203.165 49.790 203.195 ;
        RECT 49.910 202.945 50.080 203.015 ;
        RECT 49.210 202.775 50.080 202.945 ;
        RECT 49.570 202.685 50.080 202.775 ;
        RECT 48.120 202.220 48.425 202.350 ;
        RECT 48.870 202.240 49.400 202.605 ;
        RECT 47.740 201.625 48.005 202.085 ;
        RECT 48.175 201.795 48.425 202.220 ;
        RECT 49.570 202.070 49.740 202.685 ;
        RECT 48.635 201.900 49.740 202.070 ;
        RECT 49.910 201.625 50.080 202.425 ;
        RECT 50.250 202.125 50.420 203.195 ;
        RECT 50.590 202.295 50.780 203.015 ;
        RECT 50.950 202.265 51.270 203.225 ;
        RECT 51.440 203.265 51.610 203.725 ;
        RECT 51.885 203.645 52.095 204.175 ;
        RECT 52.355 203.435 52.685 203.960 ;
        RECT 52.855 203.565 53.025 204.175 ;
        RECT 53.195 203.520 53.525 203.955 ;
        RECT 53.835 203.625 54.005 203.915 ;
        RECT 54.175 203.795 54.505 204.175 ;
        RECT 53.195 203.435 53.575 203.520 ;
        RECT 53.835 203.455 54.500 203.625 ;
        RECT 52.485 203.265 52.685 203.435 ;
        RECT 53.350 203.395 53.575 203.435 ;
        RECT 51.440 202.935 52.315 203.265 ;
        RECT 52.485 202.935 53.235 203.265 ;
        RECT 50.250 201.795 50.500 202.125 ;
        RECT 51.440 202.095 51.610 202.935 ;
        RECT 52.485 202.730 52.675 202.935 ;
        RECT 53.405 202.815 53.575 203.395 ;
        RECT 53.360 202.765 53.575 202.815 ;
        RECT 51.780 202.355 52.675 202.730 ;
        RECT 53.185 202.685 53.575 202.765 ;
        RECT 50.725 201.925 51.610 202.095 ;
        RECT 51.790 201.625 52.105 202.125 ;
        RECT 52.335 201.795 52.675 202.355 ;
        RECT 52.845 201.625 53.015 202.635 ;
        RECT 53.185 201.840 53.515 202.685 ;
        RECT 53.750 202.635 54.100 203.285 ;
        RECT 54.270 202.465 54.500 203.455 ;
        RECT 53.835 202.295 54.500 202.465 ;
        RECT 53.835 201.795 54.005 202.295 ;
        RECT 54.175 201.625 54.505 202.125 ;
        RECT 54.675 201.795 54.860 203.915 ;
        RECT 55.115 203.715 55.365 204.175 ;
        RECT 55.535 203.725 55.870 203.895 ;
        RECT 56.065 203.725 56.740 203.895 ;
        RECT 55.535 203.585 55.705 203.725 ;
        RECT 55.030 202.595 55.310 203.545 ;
        RECT 55.480 203.455 55.705 203.585 ;
        RECT 55.480 202.350 55.650 203.455 ;
        RECT 55.875 203.305 56.400 203.525 ;
        RECT 55.820 202.540 56.060 203.135 ;
        RECT 56.230 202.605 56.400 203.305 ;
        RECT 56.570 202.945 56.740 203.725 ;
        RECT 57.060 203.675 57.430 204.175 ;
        RECT 57.610 203.725 58.015 203.895 ;
        RECT 58.185 203.725 58.970 203.895 ;
        RECT 57.610 203.495 57.780 203.725 ;
        RECT 56.950 203.195 57.780 203.495 ;
        RECT 58.165 203.225 58.630 203.555 ;
        RECT 56.950 203.165 57.150 203.195 ;
        RECT 57.270 202.945 57.440 203.015 ;
        RECT 56.570 202.775 57.440 202.945 ;
        RECT 56.930 202.685 57.440 202.775 ;
        RECT 55.480 202.220 55.785 202.350 ;
        RECT 56.230 202.240 56.760 202.605 ;
        RECT 55.100 201.625 55.365 202.085 ;
        RECT 55.535 201.795 55.785 202.220 ;
        RECT 56.930 202.070 57.100 202.685 ;
        RECT 55.995 201.900 57.100 202.070 ;
        RECT 57.270 201.625 57.440 202.425 ;
        RECT 57.610 202.125 57.780 203.195 ;
        RECT 57.950 202.295 58.140 203.015 ;
        RECT 58.310 202.265 58.630 203.225 ;
        RECT 58.800 203.265 58.970 203.725 ;
        RECT 59.245 203.645 59.455 204.175 ;
        RECT 59.715 203.435 60.045 203.960 ;
        RECT 60.215 203.565 60.385 204.175 ;
        RECT 60.555 203.520 60.885 203.955 ;
        RECT 60.555 203.435 60.935 203.520 ;
        RECT 59.845 203.265 60.045 203.435 ;
        RECT 60.710 203.395 60.935 203.435 ;
        RECT 58.800 202.935 59.675 203.265 ;
        RECT 59.845 202.935 60.595 203.265 ;
        RECT 57.610 201.795 57.860 202.125 ;
        RECT 58.800 202.095 58.970 202.935 ;
        RECT 59.845 202.730 60.035 202.935 ;
        RECT 60.765 202.815 60.935 203.395 ;
        RECT 60.720 202.765 60.935 202.815 ;
        RECT 59.140 202.355 60.035 202.730 ;
        RECT 60.545 202.685 60.935 202.765 ;
        RECT 61.105 203.435 61.490 204.005 ;
        RECT 61.660 203.715 61.985 204.175 ;
        RECT 62.505 203.545 62.785 204.005 ;
        RECT 61.105 202.765 61.385 203.435 ;
        RECT 61.660 203.375 62.785 203.545 ;
        RECT 61.660 203.265 62.110 203.375 ;
        RECT 61.555 202.935 62.110 203.265 ;
        RECT 62.975 203.205 63.375 204.005 ;
        RECT 63.775 203.715 64.045 204.175 ;
        RECT 64.215 203.545 64.500 204.005 ;
        RECT 58.085 201.925 58.970 202.095 ;
        RECT 59.150 201.625 59.465 202.125 ;
        RECT 59.695 201.795 60.035 202.355 ;
        RECT 60.205 201.625 60.375 202.635 ;
        RECT 60.545 201.840 60.875 202.685 ;
        RECT 61.105 201.795 61.490 202.765 ;
        RECT 61.660 202.475 62.110 202.935 ;
        RECT 62.280 202.645 63.375 203.205 ;
        RECT 61.660 202.255 62.785 202.475 ;
        RECT 61.660 201.625 61.985 202.085 ;
        RECT 62.505 201.795 62.785 202.255 ;
        RECT 62.975 201.795 63.375 202.645 ;
        RECT 63.545 203.375 64.500 203.545 ;
        RECT 65.360 203.545 65.645 204.005 ;
        RECT 65.815 203.715 66.085 204.175 ;
        RECT 65.360 203.375 66.315 203.545 ;
        RECT 63.545 202.475 63.755 203.375 ;
        RECT 63.925 202.645 64.615 203.205 ;
        RECT 65.245 202.645 65.935 203.205 ;
        RECT 66.105 202.475 66.315 203.375 ;
        RECT 63.545 202.255 64.500 202.475 ;
        RECT 63.775 201.625 64.045 202.085 ;
        RECT 64.215 201.795 64.500 202.255 ;
        RECT 65.360 202.255 66.315 202.475 ;
        RECT 66.485 203.205 66.885 204.005 ;
        RECT 67.075 203.545 67.355 204.005 ;
        RECT 67.875 203.715 68.200 204.175 ;
        RECT 67.075 203.375 68.200 203.545 ;
        RECT 68.370 203.435 68.755 204.005 ;
        RECT 68.925 203.450 69.215 204.175 ;
        RECT 69.540 203.525 69.870 203.990 ;
        RECT 70.040 203.705 70.210 204.175 ;
        RECT 70.380 203.525 70.710 204.005 ;
        RECT 67.750 203.265 68.200 203.375 ;
        RECT 66.485 202.645 67.580 203.205 ;
        RECT 67.750 202.935 68.305 203.265 ;
        RECT 65.360 201.795 65.645 202.255 ;
        RECT 65.815 201.625 66.085 202.085 ;
        RECT 66.485 201.795 66.885 202.645 ;
        RECT 67.750 202.475 68.200 202.935 ;
        RECT 68.475 202.765 68.755 203.435 ;
        RECT 69.540 203.355 70.710 203.525 ;
        RECT 69.385 202.975 70.030 203.185 ;
        RECT 70.200 202.975 70.770 203.185 ;
        RECT 70.940 202.805 71.110 204.005 ;
        RECT 71.650 203.605 71.820 203.810 ;
        RECT 67.075 202.255 68.200 202.475 ;
        RECT 67.075 201.795 67.355 202.255 ;
        RECT 67.875 201.625 68.200 202.085 ;
        RECT 68.370 201.795 68.755 202.765 ;
        RECT 68.925 201.625 69.215 202.790 ;
        RECT 69.600 201.625 69.930 202.725 ;
        RECT 70.405 202.395 71.110 202.805 ;
        RECT 71.280 203.435 71.820 203.605 ;
        RECT 72.100 203.435 72.270 204.175 ;
        RECT 72.535 203.435 72.895 203.810 ;
        RECT 73.155 203.625 73.325 203.915 ;
        RECT 73.495 203.795 73.825 204.175 ;
        RECT 73.155 203.455 73.820 203.625 ;
        RECT 71.280 202.735 71.450 203.435 ;
        RECT 71.620 202.935 71.950 203.265 ;
        RECT 72.120 202.935 72.470 203.265 ;
        RECT 71.280 202.565 71.905 202.735 ;
        RECT 72.120 202.395 72.385 202.935 ;
        RECT 72.640 202.780 72.895 203.435 ;
        RECT 70.405 202.225 72.385 202.395 ;
        RECT 70.405 201.795 70.730 202.225 ;
        RECT 70.900 201.625 71.230 202.045 ;
        RECT 71.975 201.625 72.385 202.055 ;
        RECT 72.555 201.795 72.895 202.780 ;
        RECT 73.070 202.635 73.420 203.285 ;
        RECT 73.590 202.465 73.820 203.455 ;
        RECT 73.155 202.295 73.820 202.465 ;
        RECT 73.155 201.795 73.325 202.295 ;
        RECT 73.495 201.625 73.825 202.125 ;
        RECT 73.995 201.795 74.180 203.915 ;
        RECT 74.435 203.715 74.685 204.175 ;
        RECT 74.855 203.725 75.190 203.895 ;
        RECT 75.385 203.725 76.060 203.895 ;
        RECT 74.855 203.585 75.025 203.725 ;
        RECT 74.350 202.595 74.630 203.545 ;
        RECT 74.800 203.455 75.025 203.585 ;
        RECT 74.800 202.350 74.970 203.455 ;
        RECT 75.195 203.305 75.720 203.525 ;
        RECT 75.140 202.540 75.380 203.135 ;
        RECT 75.550 202.605 75.720 203.305 ;
        RECT 75.890 202.945 76.060 203.725 ;
        RECT 76.380 203.675 76.750 204.175 ;
        RECT 76.930 203.725 77.335 203.895 ;
        RECT 77.505 203.725 78.290 203.895 ;
        RECT 76.930 203.495 77.100 203.725 ;
        RECT 76.270 203.195 77.100 203.495 ;
        RECT 77.485 203.225 77.950 203.555 ;
        RECT 76.270 203.165 76.470 203.195 ;
        RECT 76.590 202.945 76.760 203.015 ;
        RECT 75.890 202.775 76.760 202.945 ;
        RECT 76.250 202.685 76.760 202.775 ;
        RECT 74.800 202.220 75.105 202.350 ;
        RECT 75.550 202.240 76.080 202.605 ;
        RECT 74.420 201.625 74.685 202.085 ;
        RECT 74.855 201.795 75.105 202.220 ;
        RECT 76.250 202.070 76.420 202.685 ;
        RECT 75.315 201.900 76.420 202.070 ;
        RECT 76.590 201.625 76.760 202.425 ;
        RECT 76.930 202.125 77.100 203.195 ;
        RECT 77.270 202.295 77.460 203.015 ;
        RECT 77.630 202.265 77.950 203.225 ;
        RECT 78.120 203.265 78.290 203.725 ;
        RECT 78.565 203.645 78.775 204.175 ;
        RECT 79.035 203.435 79.365 203.960 ;
        RECT 79.535 203.565 79.705 204.175 ;
        RECT 79.875 203.520 80.205 203.955 ;
        RECT 80.515 203.625 80.685 203.915 ;
        RECT 80.855 203.795 81.185 204.175 ;
        RECT 79.875 203.435 80.255 203.520 ;
        RECT 80.515 203.455 81.180 203.625 ;
        RECT 79.165 203.265 79.365 203.435 ;
        RECT 80.030 203.395 80.255 203.435 ;
        RECT 78.120 202.935 78.995 203.265 ;
        RECT 79.165 202.935 79.915 203.265 ;
        RECT 76.930 201.795 77.180 202.125 ;
        RECT 78.120 202.095 78.290 202.935 ;
        RECT 79.165 202.730 79.355 202.935 ;
        RECT 80.085 202.815 80.255 203.395 ;
        RECT 80.040 202.765 80.255 202.815 ;
        RECT 78.460 202.355 79.355 202.730 ;
        RECT 79.865 202.685 80.255 202.765 ;
        RECT 77.405 201.925 78.290 202.095 ;
        RECT 78.470 201.625 78.785 202.125 ;
        RECT 79.015 201.795 79.355 202.355 ;
        RECT 79.525 201.625 79.695 202.635 ;
        RECT 79.865 201.840 80.195 202.685 ;
        RECT 80.430 202.635 80.780 203.285 ;
        RECT 80.950 202.465 81.180 203.455 ;
        RECT 80.515 202.295 81.180 202.465 ;
        RECT 80.515 201.795 80.685 202.295 ;
        RECT 80.855 201.625 81.185 202.125 ;
        RECT 81.355 201.795 81.540 203.915 ;
        RECT 81.795 203.715 82.045 204.175 ;
        RECT 82.215 203.725 82.550 203.895 ;
        RECT 82.745 203.725 83.420 203.895 ;
        RECT 82.215 203.585 82.385 203.725 ;
        RECT 81.710 202.595 81.990 203.545 ;
        RECT 82.160 203.455 82.385 203.585 ;
        RECT 82.160 202.350 82.330 203.455 ;
        RECT 82.555 203.305 83.080 203.525 ;
        RECT 82.500 202.540 82.740 203.135 ;
        RECT 82.910 202.605 83.080 203.305 ;
        RECT 83.250 202.945 83.420 203.725 ;
        RECT 83.740 203.675 84.110 204.175 ;
        RECT 84.290 203.725 84.695 203.895 ;
        RECT 84.865 203.725 85.650 203.895 ;
        RECT 84.290 203.495 84.460 203.725 ;
        RECT 83.630 203.195 84.460 203.495 ;
        RECT 84.845 203.225 85.310 203.555 ;
        RECT 83.630 203.165 83.830 203.195 ;
        RECT 83.950 202.945 84.120 203.015 ;
        RECT 83.250 202.775 84.120 202.945 ;
        RECT 83.610 202.685 84.120 202.775 ;
        RECT 82.160 202.220 82.465 202.350 ;
        RECT 82.910 202.240 83.440 202.605 ;
        RECT 81.780 201.625 82.045 202.085 ;
        RECT 82.215 201.795 82.465 202.220 ;
        RECT 83.610 202.070 83.780 202.685 ;
        RECT 82.675 201.900 83.780 202.070 ;
        RECT 83.950 201.625 84.120 202.425 ;
        RECT 84.290 202.125 84.460 203.195 ;
        RECT 84.630 202.295 84.820 203.015 ;
        RECT 84.990 202.265 85.310 203.225 ;
        RECT 85.480 203.265 85.650 203.725 ;
        RECT 85.925 203.645 86.135 204.175 ;
        RECT 86.395 203.435 86.725 203.960 ;
        RECT 86.895 203.565 87.065 204.175 ;
        RECT 87.235 203.520 87.565 203.955 ;
        RECT 88.795 203.525 88.965 204.005 ;
        RECT 89.135 203.695 89.465 204.175 ;
        RECT 89.690 203.755 91.225 204.005 ;
        RECT 89.690 203.525 89.860 203.755 ;
        RECT 87.235 203.435 87.615 203.520 ;
        RECT 86.525 203.265 86.725 203.435 ;
        RECT 87.390 203.395 87.615 203.435 ;
        RECT 85.480 202.935 86.355 203.265 ;
        RECT 86.525 202.935 87.275 203.265 ;
        RECT 84.290 201.795 84.540 202.125 ;
        RECT 85.480 202.095 85.650 202.935 ;
        RECT 86.525 202.730 86.715 202.935 ;
        RECT 87.445 202.815 87.615 203.395 ;
        RECT 88.795 203.355 89.860 203.525 ;
        RECT 90.040 203.185 90.320 203.585 ;
        RECT 88.710 202.975 89.060 203.185 ;
        RECT 89.230 202.985 89.675 203.185 ;
        RECT 89.845 202.985 90.320 203.185 ;
        RECT 90.590 203.185 90.875 203.585 ;
        RECT 91.055 203.525 91.225 203.755 ;
        RECT 91.395 203.695 91.725 204.175 ;
        RECT 91.940 203.675 92.195 204.005 ;
        RECT 91.985 203.665 92.195 203.675 ;
        RECT 92.010 203.595 92.195 203.665 ;
        RECT 91.055 203.355 91.855 203.525 ;
        RECT 90.590 202.985 90.920 203.185 ;
        RECT 91.090 202.985 91.455 203.185 ;
        RECT 87.400 202.765 87.615 202.815 ;
        RECT 91.685 202.805 91.855 203.355 ;
        RECT 85.820 202.355 86.715 202.730 ;
        RECT 87.225 202.685 87.615 202.765 ;
        RECT 84.765 201.925 85.650 202.095 ;
        RECT 85.830 201.625 86.145 202.125 ;
        RECT 86.375 201.795 86.715 202.355 ;
        RECT 86.885 201.625 87.055 202.635 ;
        RECT 87.225 201.840 87.555 202.685 ;
        RECT 88.795 202.635 91.855 202.805 ;
        RECT 88.795 201.795 88.965 202.635 ;
        RECT 92.025 202.465 92.195 203.595 ;
        RECT 92.445 203.355 92.655 204.175 ;
        RECT 92.825 203.375 93.155 204.005 ;
        RECT 92.825 202.775 93.075 203.375 ;
        RECT 93.325 203.355 93.555 204.175 ;
        RECT 94.685 203.450 94.975 204.175 ;
        RECT 95.160 203.605 95.415 203.955 ;
        RECT 95.585 203.775 95.915 204.175 ;
        RECT 96.085 203.605 96.255 203.955 ;
        RECT 96.425 203.775 96.805 204.175 ;
        RECT 95.160 203.435 96.825 203.605 ;
        RECT 96.995 203.500 97.270 203.845 ;
        RECT 96.655 203.265 96.825 203.435 ;
        RECT 93.245 202.935 93.575 203.185 ;
        RECT 95.145 202.935 95.490 203.265 ;
        RECT 95.660 202.935 96.485 203.265 ;
        RECT 96.655 202.935 96.930 203.265 ;
        RECT 89.135 201.965 89.465 202.465 ;
        RECT 89.635 202.225 91.270 202.465 ;
        RECT 89.635 202.135 89.865 202.225 ;
        RECT 89.975 201.965 90.305 202.005 ;
        RECT 89.135 201.795 90.305 201.965 ;
        RECT 90.495 201.625 90.850 202.045 ;
        RECT 91.020 201.795 91.270 202.225 ;
        RECT 91.440 201.625 91.770 202.385 ;
        RECT 91.940 201.795 92.195 202.465 ;
        RECT 92.445 201.625 92.655 202.765 ;
        RECT 92.825 201.795 93.155 202.775 ;
        RECT 93.325 201.625 93.555 202.765 ;
        RECT 94.685 201.625 94.975 202.790 ;
        RECT 95.165 202.475 95.490 202.765 ;
        RECT 95.660 202.645 95.855 202.935 ;
        RECT 96.655 202.765 96.825 202.935 ;
        RECT 97.100 202.765 97.270 203.500 ;
        RECT 96.165 202.595 96.825 202.765 ;
        RECT 96.165 202.475 96.335 202.595 ;
        RECT 95.165 202.305 96.335 202.475 ;
        RECT 95.145 201.845 96.335 202.135 ;
        RECT 96.505 201.625 96.785 202.425 ;
        RECT 96.995 201.795 97.270 202.765 ;
        RECT 97.445 203.450 97.705 204.005 ;
        RECT 97.875 203.730 98.305 204.175 ;
        RECT 98.540 203.605 98.710 204.005 ;
        RECT 98.880 203.775 99.600 204.175 ;
        RECT 97.445 202.735 97.620 203.450 ;
        RECT 98.540 203.435 99.420 203.605 ;
        RECT 99.770 203.560 99.940 204.005 ;
        RECT 100.515 203.665 100.915 204.175 ;
        RECT 97.790 202.935 98.045 203.265 ;
        RECT 97.445 201.795 97.705 202.735 ;
        RECT 97.875 202.455 98.045 202.935 ;
        RECT 98.270 202.645 98.600 203.265 ;
        RECT 98.770 202.885 99.060 203.265 ;
        RECT 99.250 202.715 99.420 203.435 ;
        RECT 98.900 202.545 99.420 202.715 ;
        RECT 99.590 203.390 99.940 203.560 ;
        RECT 101.175 203.520 101.505 203.955 ;
        RECT 101.675 203.565 101.845 204.175 ;
        RECT 97.875 202.285 98.635 202.455 ;
        RECT 98.900 202.355 99.070 202.545 ;
        RECT 99.590 202.365 99.760 203.390 ;
        RECT 100.180 202.905 100.440 203.495 ;
        RECT 99.960 202.605 100.440 202.905 ;
        RECT 100.640 202.605 100.900 203.495 ;
        RECT 101.125 203.435 101.505 203.520 ;
        RECT 102.015 203.435 102.345 203.960 ;
        RECT 102.605 203.645 102.815 204.175 ;
        RECT 103.090 203.725 103.875 203.895 ;
        RECT 104.045 203.725 104.450 203.895 ;
        RECT 101.125 203.395 101.350 203.435 ;
        RECT 101.125 202.815 101.295 203.395 ;
        RECT 102.015 203.265 102.215 203.435 ;
        RECT 103.090 203.265 103.260 203.725 ;
        RECT 101.465 202.935 102.215 203.265 ;
        RECT 102.385 202.935 103.260 203.265 ;
        RECT 101.125 202.765 101.340 202.815 ;
        RECT 101.125 202.685 101.515 202.765 ;
        RECT 98.465 202.060 98.635 202.285 ;
        RECT 99.350 202.195 99.760 202.365 ;
        RECT 99.935 202.255 100.875 202.425 ;
        RECT 99.350 202.060 99.605 202.195 ;
        RECT 97.875 201.625 98.205 202.025 ;
        RECT 98.465 201.890 99.605 202.060 ;
        RECT 99.935 202.005 100.105 202.255 ;
        RECT 99.350 201.795 99.605 201.890 ;
        RECT 99.775 201.835 100.105 202.005 ;
        RECT 100.275 201.625 100.525 202.085 ;
        RECT 100.695 201.795 100.875 202.255 ;
        RECT 101.185 201.840 101.515 202.685 ;
        RECT 102.025 202.730 102.215 202.935 ;
        RECT 101.685 201.625 101.855 202.635 ;
        RECT 102.025 202.355 102.920 202.730 ;
        RECT 102.025 201.795 102.365 202.355 ;
        RECT 102.595 201.625 102.910 202.125 ;
        RECT 103.090 202.095 103.260 202.935 ;
        RECT 103.430 203.225 103.895 203.555 ;
        RECT 104.280 203.495 104.450 203.725 ;
        RECT 104.630 203.675 105.000 204.175 ;
        RECT 105.320 203.725 105.995 203.895 ;
        RECT 106.190 203.725 106.525 203.895 ;
        RECT 103.430 202.265 103.750 203.225 ;
        RECT 104.280 203.195 105.110 203.495 ;
        RECT 103.920 202.295 104.110 203.015 ;
        RECT 104.280 202.125 104.450 203.195 ;
        RECT 104.910 203.165 105.110 203.195 ;
        RECT 104.620 202.945 104.790 203.015 ;
        RECT 105.320 202.945 105.490 203.725 ;
        RECT 106.355 203.585 106.525 203.725 ;
        RECT 106.695 203.715 106.945 204.175 ;
        RECT 104.620 202.775 105.490 202.945 ;
        RECT 105.660 203.305 106.185 203.525 ;
        RECT 106.355 203.455 106.580 203.585 ;
        RECT 104.620 202.685 105.130 202.775 ;
        RECT 103.090 201.925 103.975 202.095 ;
        RECT 104.200 201.795 104.450 202.125 ;
        RECT 104.620 201.625 104.790 202.425 ;
        RECT 104.960 202.070 105.130 202.685 ;
        RECT 105.660 202.605 105.830 203.305 ;
        RECT 105.300 202.240 105.830 202.605 ;
        RECT 106.000 202.540 106.240 203.135 ;
        RECT 106.410 202.350 106.580 203.455 ;
        RECT 106.750 202.595 107.030 203.545 ;
        RECT 106.275 202.220 106.580 202.350 ;
        RECT 104.960 201.900 106.065 202.070 ;
        RECT 106.275 201.795 106.525 202.220 ;
        RECT 106.695 201.625 106.960 202.085 ;
        RECT 107.200 201.795 107.385 203.915 ;
        RECT 107.555 203.795 107.885 204.175 ;
        RECT 108.055 203.625 108.225 203.915 ;
        RECT 108.485 203.630 113.830 204.175 ;
        RECT 114.005 203.630 119.350 204.175 ;
        RECT 107.560 203.455 108.225 203.625 ;
        RECT 107.560 202.465 107.790 203.455 ;
        RECT 107.960 202.635 108.310 203.285 ;
        RECT 110.070 202.800 110.410 203.630 ;
        RECT 107.560 202.295 108.225 202.465 ;
        RECT 107.555 201.625 107.885 202.125 ;
        RECT 108.055 201.795 108.225 202.295 ;
        RECT 111.890 202.060 112.240 203.310 ;
        RECT 115.590 202.800 115.930 203.630 ;
        RECT 120.445 203.450 120.735 204.175 ;
        RECT 120.905 203.630 126.250 204.175 ;
        RECT 126.425 203.630 131.770 204.175 ;
        RECT 131.945 203.630 137.290 204.175 ;
        RECT 137.465 203.630 142.810 204.175 ;
        RECT 117.410 202.060 117.760 203.310 ;
        RECT 122.490 202.800 122.830 203.630 ;
        RECT 108.485 201.625 113.830 202.060 ;
        RECT 114.005 201.625 119.350 202.060 ;
        RECT 120.445 201.625 120.735 202.790 ;
        RECT 124.310 202.060 124.660 203.310 ;
        RECT 128.010 202.800 128.350 203.630 ;
        RECT 129.830 202.060 130.180 203.310 ;
        RECT 133.530 202.800 133.870 203.630 ;
        RECT 135.350 202.060 135.700 203.310 ;
        RECT 139.050 202.800 139.390 203.630 ;
        RECT 142.985 203.405 145.575 204.175 ;
        RECT 145.745 203.425 146.955 204.175 ;
        RECT 140.870 202.060 141.220 203.310 ;
        RECT 142.985 202.885 144.195 203.405 ;
        RECT 144.365 202.715 145.575 203.235 ;
        RECT 120.905 201.625 126.250 202.060 ;
        RECT 126.425 201.625 131.770 202.060 ;
        RECT 131.945 201.625 137.290 202.060 ;
        RECT 137.465 201.625 142.810 202.060 ;
        RECT 142.985 201.625 145.575 202.715 ;
        RECT 145.745 202.715 146.265 203.255 ;
        RECT 146.435 202.885 146.955 203.425 ;
        RECT 145.745 201.625 146.955 202.715 ;
        RECT 17.320 201.455 147.040 201.625 ;
        RECT 17.405 200.365 18.615 201.455 ;
        RECT 18.785 201.020 24.130 201.455 ;
        RECT 24.305 201.020 29.650 201.455 ;
        RECT 17.405 199.655 17.925 200.195 ;
        RECT 18.095 199.825 18.615 200.365 ;
        RECT 17.405 198.905 18.615 199.655 ;
        RECT 20.370 199.450 20.710 200.280 ;
        RECT 22.190 199.770 22.540 201.020 ;
        RECT 25.890 199.450 26.230 200.280 ;
        RECT 27.710 199.770 28.060 201.020 ;
        RECT 30.285 200.290 30.575 201.455 ;
        RECT 30.745 201.020 36.090 201.455 ;
        RECT 36.265 201.020 41.610 201.455 ;
        RECT 18.785 198.905 24.130 199.450 ;
        RECT 24.305 198.905 29.650 199.450 ;
        RECT 30.285 198.905 30.575 199.630 ;
        RECT 32.330 199.450 32.670 200.280 ;
        RECT 34.150 199.770 34.500 201.020 ;
        RECT 37.850 199.450 38.190 200.280 ;
        RECT 39.670 199.770 40.020 201.020 ;
        RECT 41.785 200.365 45.295 201.455 ;
        RECT 46.015 200.785 46.185 201.285 ;
        RECT 46.355 200.955 46.685 201.455 ;
        RECT 46.015 200.615 46.680 200.785 ;
        RECT 41.785 199.675 43.435 200.195 ;
        RECT 43.605 199.845 45.295 200.365 ;
        RECT 45.930 199.795 46.280 200.445 ;
        RECT 30.745 198.905 36.090 199.450 ;
        RECT 36.265 198.905 41.610 199.450 ;
        RECT 41.785 198.905 45.295 199.675 ;
        RECT 46.450 199.625 46.680 200.615 ;
        RECT 46.015 199.455 46.680 199.625 ;
        RECT 46.015 199.165 46.185 199.455 ;
        RECT 46.355 198.905 46.685 199.285 ;
        RECT 46.855 199.165 47.040 201.285 ;
        RECT 47.280 200.995 47.545 201.455 ;
        RECT 47.715 200.860 47.965 201.285 ;
        RECT 48.175 201.010 49.280 201.180 ;
        RECT 47.660 200.730 47.965 200.860 ;
        RECT 47.210 199.535 47.490 200.485 ;
        RECT 47.660 199.625 47.830 200.730 ;
        RECT 48.000 199.945 48.240 200.540 ;
        RECT 48.410 200.475 48.940 200.840 ;
        RECT 48.410 199.775 48.580 200.475 ;
        RECT 49.110 200.395 49.280 201.010 ;
        RECT 49.450 200.655 49.620 201.455 ;
        RECT 49.790 200.955 50.040 201.285 ;
        RECT 50.265 200.985 51.150 201.155 ;
        RECT 49.110 200.305 49.620 200.395 ;
        RECT 47.660 199.495 47.885 199.625 ;
        RECT 48.055 199.555 48.580 199.775 ;
        RECT 48.750 200.135 49.620 200.305 ;
        RECT 47.295 198.905 47.545 199.365 ;
        RECT 47.715 199.355 47.885 199.495 ;
        RECT 48.750 199.355 48.920 200.135 ;
        RECT 49.450 200.065 49.620 200.135 ;
        RECT 49.130 199.885 49.330 199.915 ;
        RECT 49.790 199.885 49.960 200.955 ;
        RECT 50.130 200.065 50.320 200.785 ;
        RECT 49.130 199.585 49.960 199.885 ;
        RECT 50.490 199.855 50.810 200.815 ;
        RECT 47.715 199.185 48.050 199.355 ;
        RECT 48.245 199.185 48.920 199.355 ;
        RECT 49.240 198.905 49.610 199.405 ;
        RECT 49.790 199.355 49.960 199.585 ;
        RECT 50.345 199.525 50.810 199.855 ;
        RECT 50.980 200.145 51.150 200.985 ;
        RECT 51.330 200.955 51.645 201.455 ;
        RECT 51.875 200.725 52.215 201.285 ;
        RECT 51.320 200.350 52.215 200.725 ;
        RECT 52.385 200.445 52.555 201.455 ;
        RECT 52.025 200.145 52.215 200.350 ;
        RECT 52.725 200.395 53.055 201.240 ;
        RECT 54.215 200.845 54.545 201.275 ;
        RECT 54.725 201.015 54.920 201.455 ;
        RECT 55.090 200.845 55.420 201.275 ;
        RECT 54.215 200.675 55.420 200.845 ;
        RECT 52.725 200.315 53.115 200.395 ;
        RECT 54.215 200.345 55.110 200.675 ;
        RECT 55.590 200.505 55.865 201.275 ;
        RECT 52.900 200.265 53.115 200.315 ;
        RECT 50.980 199.815 51.855 200.145 ;
        RECT 52.025 199.815 52.775 200.145 ;
        RECT 50.980 199.355 51.150 199.815 ;
        RECT 52.025 199.645 52.225 199.815 ;
        RECT 52.945 199.685 53.115 200.265 ;
        RECT 55.280 200.315 55.865 200.505 ;
        RECT 54.220 199.815 54.515 200.145 ;
        RECT 54.695 199.815 55.110 200.145 ;
        RECT 52.890 199.645 53.115 199.685 ;
        RECT 49.790 199.185 50.195 199.355 ;
        RECT 50.365 199.185 51.150 199.355 ;
        RECT 51.425 198.905 51.635 199.435 ;
        RECT 51.895 199.120 52.225 199.645 ;
        RECT 52.735 199.560 53.115 199.645 ;
        RECT 52.395 198.905 52.565 199.515 ;
        RECT 52.735 199.125 53.065 199.560 ;
        RECT 54.215 198.905 54.515 199.635 ;
        RECT 54.695 199.195 54.925 199.815 ;
        RECT 55.280 199.645 55.455 200.315 ;
        RECT 56.045 200.290 56.335 201.455 ;
        RECT 56.510 201.075 56.845 201.455 ;
        RECT 55.125 199.465 55.455 199.645 ;
        RECT 55.625 199.495 55.865 200.145 ;
        RECT 55.125 199.085 55.350 199.465 ;
        RECT 55.520 198.905 55.850 199.295 ;
        RECT 56.045 198.905 56.335 199.630 ;
        RECT 56.505 199.585 56.745 200.895 ;
        RECT 57.015 200.485 57.265 201.285 ;
        RECT 57.485 200.735 57.815 201.455 ;
        RECT 58.000 200.485 58.250 201.285 ;
        RECT 58.715 200.655 59.045 201.455 ;
        RECT 59.215 201.025 59.555 201.285 ;
        RECT 56.915 200.315 59.105 200.485 ;
        RECT 56.915 199.405 57.085 200.315 ;
        RECT 58.790 200.145 59.105 200.315 ;
        RECT 56.590 199.075 57.085 199.405 ;
        RECT 57.305 199.180 57.655 200.145 ;
        RECT 57.835 199.175 58.135 200.145 ;
        RECT 58.315 199.175 58.595 200.145 ;
        RECT 58.790 199.895 59.120 200.145 ;
        RECT 58.775 198.905 59.045 199.705 ;
        RECT 59.295 199.625 59.555 201.025 ;
        RECT 59.215 199.115 59.555 199.625 ;
        RECT 60.185 200.585 60.460 201.285 ;
        RECT 60.630 200.910 60.885 201.455 ;
        RECT 61.055 200.945 61.535 201.285 ;
        RECT 61.710 200.900 62.315 201.455 ;
        RECT 62.485 200.945 62.785 201.455 ;
        RECT 61.700 200.800 62.315 200.900 ;
        RECT 61.700 200.775 61.885 200.800 ;
        RECT 62.955 200.775 63.285 201.285 ;
        RECT 63.455 200.945 64.085 201.455 ;
        RECT 64.665 200.945 65.045 201.115 ;
        RECT 65.215 200.945 65.515 201.455 ;
        RECT 64.875 200.775 65.045 200.945 ;
        RECT 65.795 200.785 65.965 201.285 ;
        RECT 66.135 200.955 66.465 201.455 ;
        RECT 60.185 199.555 60.355 200.585 ;
        RECT 60.630 200.455 61.385 200.705 ;
        RECT 61.555 200.530 61.885 200.775 ;
        RECT 60.630 200.420 61.400 200.455 ;
        RECT 60.630 200.410 61.415 200.420 ;
        RECT 60.525 200.395 61.420 200.410 ;
        RECT 60.525 200.380 61.440 200.395 ;
        RECT 60.525 200.370 61.460 200.380 ;
        RECT 60.525 200.360 61.485 200.370 ;
        RECT 60.525 200.330 61.555 200.360 ;
        RECT 60.525 200.300 61.575 200.330 ;
        RECT 60.525 200.270 61.595 200.300 ;
        RECT 60.525 200.245 61.625 200.270 ;
        RECT 60.525 200.210 61.660 200.245 ;
        RECT 60.525 200.205 61.690 200.210 ;
        RECT 60.525 199.810 60.755 200.205 ;
        RECT 61.300 200.200 61.690 200.205 ;
        RECT 61.325 200.190 61.690 200.200 ;
        RECT 61.340 200.185 61.690 200.190 ;
        RECT 61.355 200.180 61.690 200.185 ;
        RECT 62.055 200.180 62.315 200.630 ;
        RECT 61.355 200.175 62.315 200.180 ;
        RECT 61.365 200.165 62.315 200.175 ;
        RECT 61.375 200.160 62.315 200.165 ;
        RECT 61.385 200.150 62.315 200.160 ;
        RECT 61.390 200.140 62.315 200.150 ;
        RECT 61.395 200.135 62.315 200.140 ;
        RECT 61.405 200.120 62.315 200.135 ;
        RECT 61.410 200.105 62.315 200.120 ;
        RECT 61.420 200.080 62.315 200.105 ;
        RECT 60.925 199.610 61.255 200.035 ;
        RECT 60.185 199.075 60.445 199.555 ;
        RECT 60.615 198.905 60.865 199.445 ;
        RECT 61.035 199.125 61.255 199.610 ;
        RECT 61.425 200.010 62.315 200.080 ;
        RECT 62.485 200.605 64.705 200.775 ;
        RECT 61.425 199.285 61.595 200.010 ;
        RECT 61.765 199.455 62.315 199.840 ;
        RECT 62.485 199.645 62.655 200.605 ;
        RECT 62.825 200.265 64.365 200.435 ;
        RECT 62.825 199.815 63.070 200.265 ;
        RECT 63.330 199.895 64.025 200.095 ;
        RECT 64.195 200.065 64.365 200.265 ;
        RECT 64.535 200.405 64.705 200.605 ;
        RECT 64.875 200.575 65.535 200.775 ;
        RECT 65.795 200.615 66.460 200.785 ;
        RECT 64.535 200.235 65.195 200.405 ;
        RECT 64.195 199.895 64.795 200.065 ;
        RECT 65.025 199.815 65.195 200.235 ;
        RECT 61.425 199.115 62.315 199.285 ;
        RECT 62.485 199.100 62.950 199.645 ;
        RECT 63.455 198.905 63.625 199.725 ;
        RECT 63.795 199.645 64.705 199.725 ;
        RECT 65.365 199.645 65.535 200.575 ;
        RECT 65.710 199.795 66.060 200.445 ;
        RECT 63.795 199.555 65.045 199.645 ;
        RECT 63.795 199.075 64.125 199.555 ;
        RECT 64.535 199.475 65.045 199.555 ;
        RECT 64.295 198.905 64.645 199.295 ;
        RECT 64.815 199.075 65.045 199.475 ;
        RECT 65.215 199.165 65.535 199.645 ;
        RECT 66.230 199.625 66.460 200.615 ;
        RECT 65.795 199.455 66.460 199.625 ;
        RECT 65.795 199.165 65.965 199.455 ;
        RECT 66.135 198.905 66.465 199.285 ;
        RECT 66.635 199.165 66.820 201.285 ;
        RECT 67.060 200.995 67.325 201.455 ;
        RECT 67.495 200.860 67.745 201.285 ;
        RECT 67.955 201.010 69.060 201.180 ;
        RECT 67.440 200.730 67.745 200.860 ;
        RECT 66.990 199.535 67.270 200.485 ;
        RECT 67.440 199.625 67.610 200.730 ;
        RECT 67.780 199.945 68.020 200.540 ;
        RECT 68.190 200.475 68.720 200.840 ;
        RECT 68.190 199.775 68.360 200.475 ;
        RECT 68.890 200.395 69.060 201.010 ;
        RECT 69.230 200.655 69.400 201.455 ;
        RECT 69.570 200.955 69.820 201.285 ;
        RECT 70.045 200.985 70.930 201.155 ;
        RECT 68.890 200.305 69.400 200.395 ;
        RECT 67.440 199.495 67.665 199.625 ;
        RECT 67.835 199.555 68.360 199.775 ;
        RECT 68.530 200.135 69.400 200.305 ;
        RECT 67.075 198.905 67.325 199.365 ;
        RECT 67.495 199.355 67.665 199.495 ;
        RECT 68.530 199.355 68.700 200.135 ;
        RECT 69.230 200.065 69.400 200.135 ;
        RECT 68.910 199.885 69.110 199.915 ;
        RECT 69.570 199.885 69.740 200.955 ;
        RECT 69.910 200.065 70.100 200.785 ;
        RECT 68.910 199.585 69.740 199.885 ;
        RECT 70.270 199.855 70.590 200.815 ;
        RECT 67.495 199.185 67.830 199.355 ;
        RECT 68.025 199.185 68.700 199.355 ;
        RECT 69.020 198.905 69.390 199.405 ;
        RECT 69.570 199.355 69.740 199.585 ;
        RECT 70.125 199.525 70.590 199.855 ;
        RECT 70.760 200.145 70.930 200.985 ;
        RECT 71.110 200.955 71.425 201.455 ;
        RECT 71.655 200.725 71.995 201.285 ;
        RECT 71.100 200.350 71.995 200.725 ;
        RECT 72.165 200.445 72.335 201.455 ;
        RECT 71.805 200.145 71.995 200.350 ;
        RECT 72.505 200.395 72.835 201.240 ;
        RECT 73.065 200.945 74.255 201.235 ;
        RECT 73.085 200.605 74.255 200.775 ;
        RECT 74.425 200.655 74.705 201.455 ;
        RECT 72.505 200.315 72.895 200.395 ;
        RECT 73.085 200.315 73.410 200.605 ;
        RECT 74.085 200.485 74.255 200.605 ;
        RECT 72.680 200.265 72.895 200.315 ;
        RECT 70.760 199.815 71.635 200.145 ;
        RECT 71.805 199.815 72.555 200.145 ;
        RECT 70.760 199.355 70.930 199.815 ;
        RECT 71.805 199.645 72.005 199.815 ;
        RECT 72.725 199.685 72.895 200.265 ;
        RECT 73.580 200.145 73.775 200.435 ;
        RECT 74.085 200.315 74.745 200.485 ;
        RECT 74.915 200.315 75.190 201.285 ;
        RECT 75.365 201.020 80.710 201.455 ;
        RECT 74.575 200.145 74.745 200.315 ;
        RECT 73.065 199.815 73.410 200.145 ;
        RECT 73.580 199.815 74.405 200.145 ;
        RECT 74.575 199.815 74.850 200.145 ;
        RECT 72.670 199.645 72.895 199.685 ;
        RECT 74.575 199.645 74.745 199.815 ;
        RECT 69.570 199.185 69.975 199.355 ;
        RECT 70.145 199.185 70.930 199.355 ;
        RECT 71.205 198.905 71.415 199.435 ;
        RECT 71.675 199.120 72.005 199.645 ;
        RECT 72.515 199.560 72.895 199.645 ;
        RECT 72.175 198.905 72.345 199.515 ;
        RECT 72.515 199.125 72.845 199.560 ;
        RECT 73.080 199.475 74.745 199.645 ;
        RECT 75.020 199.580 75.190 200.315 ;
        RECT 73.080 199.125 73.335 199.475 ;
        RECT 73.505 198.905 73.835 199.305 ;
        RECT 74.005 199.125 74.175 199.475 ;
        RECT 74.345 198.905 74.725 199.305 ;
        RECT 74.915 199.235 75.190 199.580 ;
        RECT 76.950 199.450 77.290 200.280 ;
        RECT 78.770 199.770 79.120 201.020 ;
        RECT 81.805 200.290 82.095 201.455 ;
        RECT 75.365 198.905 80.710 199.450 ;
        RECT 81.805 198.905 82.095 199.630 ;
        RECT 82.740 199.085 83.020 201.275 ;
        RECT 83.210 200.315 83.495 201.455 ;
        RECT 83.760 200.805 83.930 201.275 ;
        RECT 84.105 200.975 84.435 201.455 ;
        RECT 84.605 200.805 84.785 201.275 ;
        RECT 83.760 200.605 84.785 200.805 ;
        RECT 83.220 199.635 83.480 200.145 ;
        RECT 83.690 199.815 83.950 200.435 ;
        RECT 84.145 199.815 84.570 200.435 ;
        RECT 84.955 200.165 85.285 201.275 ;
        RECT 85.455 201.045 85.805 201.455 ;
        RECT 85.975 200.865 86.215 201.255 ;
        RECT 84.740 199.865 85.285 200.165 ;
        RECT 85.465 200.665 86.215 200.865 ;
        RECT 85.465 199.985 85.805 200.665 ;
        RECT 84.740 199.635 84.960 199.865 ;
        RECT 83.220 199.445 84.960 199.635 ;
        RECT 83.220 198.905 83.950 199.275 ;
        RECT 84.530 199.085 84.960 199.445 ;
        RECT 85.130 198.905 85.375 199.685 ;
        RECT 85.575 199.085 85.805 199.985 ;
        RECT 85.985 199.145 86.215 200.485 ;
        RECT 86.405 200.315 86.790 201.285 ;
        RECT 86.960 200.995 87.285 201.455 ;
        RECT 87.805 200.825 88.085 201.285 ;
        RECT 86.960 200.605 88.085 200.825 ;
        RECT 86.405 199.645 86.685 200.315 ;
        RECT 86.960 200.145 87.410 200.605 ;
        RECT 88.275 200.435 88.675 201.285 ;
        RECT 89.075 200.995 89.345 201.455 ;
        RECT 89.515 200.825 89.800 201.285 ;
        RECT 86.855 199.815 87.410 200.145 ;
        RECT 87.580 199.875 88.675 200.435 ;
        RECT 86.960 199.705 87.410 199.815 ;
        RECT 86.405 199.075 86.790 199.645 ;
        RECT 86.960 199.535 88.085 199.705 ;
        RECT 86.960 198.905 87.285 199.365 ;
        RECT 87.805 199.075 88.085 199.535 ;
        RECT 88.275 199.075 88.675 199.875 ;
        RECT 88.845 200.605 89.800 200.825 ;
        RECT 88.845 199.705 89.055 200.605 ;
        RECT 89.225 199.875 89.915 200.435 ;
        RECT 90.085 200.315 90.360 201.285 ;
        RECT 90.570 200.655 90.850 201.455 ;
        RECT 91.020 200.945 92.635 201.275 ;
        RECT 91.020 200.605 92.195 200.775 ;
        RECT 91.020 200.485 91.190 200.605 ;
        RECT 90.530 200.315 91.190 200.485 ;
        RECT 88.845 199.535 89.800 199.705 ;
        RECT 89.075 198.905 89.345 199.365 ;
        RECT 89.515 199.075 89.800 199.535 ;
        RECT 90.085 199.580 90.255 200.315 ;
        RECT 90.530 200.145 90.700 200.315 ;
        RECT 91.450 200.145 91.695 200.435 ;
        RECT 91.865 200.315 92.195 200.605 ;
        RECT 92.455 200.145 92.625 200.705 ;
        RECT 92.875 200.315 93.135 201.455 ;
        RECT 93.490 200.485 93.880 200.660 ;
        RECT 94.365 200.655 94.695 201.455 ;
        RECT 94.865 200.665 95.400 201.285 ;
        RECT 93.490 200.315 94.915 200.485 ;
        RECT 90.425 199.815 90.700 200.145 ;
        RECT 90.870 199.815 91.695 200.145 ;
        RECT 91.910 199.815 92.625 200.145 ;
        RECT 92.795 199.895 93.130 200.145 ;
        RECT 90.530 199.645 90.700 199.815 ;
        RECT 92.375 199.725 92.625 199.815 ;
        RECT 90.085 199.235 90.360 199.580 ;
        RECT 90.530 199.475 92.195 199.645 ;
        RECT 90.550 198.905 90.925 199.305 ;
        RECT 91.095 199.125 91.265 199.475 ;
        RECT 91.435 198.905 91.765 199.305 ;
        RECT 91.935 199.075 92.195 199.475 ;
        RECT 92.375 199.305 92.705 199.725 ;
        RECT 92.875 198.905 93.135 199.725 ;
        RECT 93.365 199.585 93.720 200.145 ;
        RECT 93.890 199.415 94.060 200.315 ;
        RECT 94.230 199.585 94.495 200.145 ;
        RECT 94.745 199.815 94.915 200.315 ;
        RECT 95.085 199.645 95.400 200.665 ;
        RECT 95.605 200.365 97.275 201.455 ;
        RECT 93.470 198.905 93.710 199.415 ;
        RECT 93.890 199.085 94.170 199.415 ;
        RECT 94.400 198.905 94.615 199.415 ;
        RECT 94.785 199.075 95.400 199.645 ;
        RECT 95.605 199.675 96.355 200.195 ;
        RECT 96.525 199.845 97.275 200.365 ;
        RECT 97.445 200.485 97.735 201.285 ;
        RECT 97.905 200.655 98.140 201.455 ;
        RECT 98.325 201.115 99.860 201.285 ;
        RECT 98.325 200.485 98.655 201.115 ;
        RECT 97.445 200.315 98.655 200.485 ;
        RECT 97.445 199.815 97.690 200.145 ;
        RECT 95.605 198.905 97.275 199.675 ;
        RECT 97.860 199.645 98.030 200.315 ;
        RECT 98.825 200.145 99.060 200.890 ;
        RECT 98.200 199.815 98.600 200.145 ;
        RECT 98.770 199.815 99.060 200.145 ;
        RECT 99.250 200.145 99.520 200.890 ;
        RECT 99.690 200.485 99.860 201.115 ;
        RECT 100.030 200.655 100.435 201.455 ;
        RECT 99.690 200.315 100.435 200.485 ;
        RECT 99.250 199.815 99.590 200.145 ;
        RECT 99.760 199.815 100.095 200.145 ;
        RECT 100.265 199.815 100.435 200.315 ;
        RECT 100.605 199.890 100.955 201.285 ;
        RECT 101.125 201.020 106.470 201.455 ;
        RECT 97.445 199.075 98.030 199.645 ;
        RECT 98.280 199.475 99.675 199.645 ;
        RECT 98.280 199.130 98.610 199.475 ;
        RECT 98.825 198.905 99.200 199.305 ;
        RECT 99.380 199.130 99.675 199.475 ;
        RECT 99.845 198.905 100.515 199.645 ;
        RECT 100.685 199.075 100.955 199.890 ;
        RECT 102.710 199.450 103.050 200.280 ;
        RECT 104.530 199.770 104.880 201.020 ;
        RECT 107.565 200.290 107.855 201.455 ;
        RECT 108.025 201.020 113.370 201.455 ;
        RECT 113.545 201.020 118.890 201.455 ;
        RECT 119.065 201.020 124.410 201.455 ;
        RECT 124.585 201.020 129.930 201.455 ;
        RECT 101.125 198.905 106.470 199.450 ;
        RECT 107.565 198.905 107.855 199.630 ;
        RECT 109.610 199.450 109.950 200.280 ;
        RECT 111.430 199.770 111.780 201.020 ;
        RECT 115.130 199.450 115.470 200.280 ;
        RECT 116.950 199.770 117.300 201.020 ;
        RECT 120.650 199.450 120.990 200.280 ;
        RECT 122.470 199.770 122.820 201.020 ;
        RECT 126.170 199.450 126.510 200.280 ;
        RECT 127.990 199.770 128.340 201.020 ;
        RECT 130.105 200.365 132.695 201.455 ;
        RECT 130.105 199.675 131.315 200.195 ;
        RECT 131.485 199.845 132.695 200.365 ;
        RECT 133.325 200.290 133.615 201.455 ;
        RECT 133.785 201.020 139.130 201.455 ;
        RECT 139.305 201.020 144.650 201.455 ;
        RECT 108.025 198.905 113.370 199.450 ;
        RECT 113.545 198.905 118.890 199.450 ;
        RECT 119.065 198.905 124.410 199.450 ;
        RECT 124.585 198.905 129.930 199.450 ;
        RECT 130.105 198.905 132.695 199.675 ;
        RECT 133.325 198.905 133.615 199.630 ;
        RECT 135.370 199.450 135.710 200.280 ;
        RECT 137.190 199.770 137.540 201.020 ;
        RECT 140.890 199.450 141.230 200.280 ;
        RECT 142.710 199.770 143.060 201.020 ;
        RECT 145.745 200.365 146.955 201.455 ;
        RECT 145.745 199.825 146.265 200.365 ;
        RECT 146.435 199.655 146.955 200.195 ;
        RECT 133.785 198.905 139.130 199.450 ;
        RECT 139.305 198.905 144.650 199.450 ;
        RECT 145.745 198.905 146.955 199.655 ;
        RECT 17.320 198.735 147.040 198.905 ;
        RECT 17.405 197.985 18.615 198.735 ;
        RECT 18.785 198.190 24.130 198.735 ;
        RECT 24.305 198.190 29.650 198.735 ;
        RECT 29.825 198.190 35.170 198.735 ;
        RECT 35.345 198.190 40.690 198.735 ;
        RECT 17.405 197.445 17.925 197.985 ;
        RECT 18.095 197.275 18.615 197.815 ;
        RECT 20.370 197.360 20.710 198.190 ;
        RECT 17.405 196.185 18.615 197.275 ;
        RECT 22.190 196.620 22.540 197.870 ;
        RECT 25.890 197.360 26.230 198.190 ;
        RECT 27.710 196.620 28.060 197.870 ;
        RECT 31.410 197.360 31.750 198.190 ;
        RECT 33.230 196.620 33.580 197.870 ;
        RECT 36.930 197.360 37.270 198.190 ;
        RECT 40.865 197.965 42.535 198.735 ;
        RECT 43.165 198.010 43.455 198.735 ;
        RECT 43.625 198.190 48.970 198.735 ;
        RECT 38.750 196.620 39.100 197.870 ;
        RECT 40.865 197.445 41.615 197.965 ;
        RECT 41.785 197.275 42.535 197.795 ;
        RECT 45.210 197.360 45.550 198.190 ;
        RECT 49.145 197.985 50.355 198.735 ;
        RECT 18.785 196.185 24.130 196.620 ;
        RECT 24.305 196.185 29.650 196.620 ;
        RECT 29.825 196.185 35.170 196.620 ;
        RECT 35.345 196.185 40.690 196.620 ;
        RECT 40.865 196.185 42.535 197.275 ;
        RECT 43.165 196.185 43.455 197.350 ;
        RECT 47.030 196.620 47.380 197.870 ;
        RECT 49.145 197.445 49.665 197.985 ;
        RECT 50.545 197.925 50.785 198.735 ;
        RECT 50.955 197.925 51.285 198.565 ;
        RECT 51.455 197.925 51.725 198.735 ;
        RECT 51.905 197.965 54.495 198.735 ;
        RECT 49.835 197.275 50.355 197.815 ;
        RECT 50.525 197.495 50.875 197.745 ;
        RECT 51.045 197.325 51.215 197.925 ;
        RECT 51.385 197.495 51.735 197.745 ;
        RECT 51.905 197.445 53.115 197.965 ;
        RECT 55.185 197.915 55.395 198.735 ;
        RECT 55.565 197.935 55.895 198.565 ;
        RECT 43.625 196.185 48.970 196.620 ;
        RECT 49.145 196.185 50.355 197.275 ;
        RECT 50.535 197.155 51.215 197.325 ;
        RECT 50.535 196.370 50.865 197.155 ;
        RECT 51.395 196.185 51.725 197.325 ;
        RECT 53.285 197.275 54.495 197.795 ;
        RECT 55.565 197.335 55.815 197.935 ;
        RECT 56.065 197.915 56.295 198.735 ;
        RECT 56.505 198.190 61.850 198.735 ;
        RECT 55.985 197.495 56.315 197.745 ;
        RECT 58.090 197.360 58.430 198.190 ;
        RECT 62.025 197.965 63.695 198.735 ;
        RECT 63.935 198.335 64.265 198.735 ;
        RECT 64.435 198.165 64.605 198.435 ;
        RECT 64.775 198.335 65.105 198.735 ;
        RECT 65.275 198.165 65.530 198.435 ;
        RECT 51.905 196.185 54.495 197.275 ;
        RECT 55.185 196.185 55.395 197.325 ;
        RECT 55.565 196.355 55.895 197.335 ;
        RECT 56.065 196.185 56.295 197.325 ;
        RECT 59.910 196.620 60.260 197.870 ;
        RECT 62.025 197.445 62.775 197.965 ;
        RECT 62.945 197.275 63.695 197.795 ;
        RECT 56.505 196.185 61.850 196.620 ;
        RECT 62.025 196.185 63.695 197.275 ;
        RECT 63.865 197.155 64.135 198.165 ;
        RECT 64.305 197.995 65.530 198.165 ;
        RECT 66.625 198.085 66.885 198.565 ;
        RECT 67.055 198.195 67.305 198.735 ;
        RECT 64.305 197.325 64.475 197.995 ;
        RECT 64.645 197.495 65.025 197.825 ;
        RECT 65.195 197.495 65.530 197.825 ;
        RECT 64.305 197.155 64.620 197.325 ;
        RECT 63.870 196.185 64.185 196.985 ;
        RECT 64.450 196.540 64.620 197.155 ;
        RECT 64.790 196.815 65.025 197.495 ;
        RECT 65.195 196.540 65.530 197.325 ;
        RECT 64.450 196.370 65.530 196.540 ;
        RECT 66.625 197.055 66.795 198.085 ;
        RECT 67.475 198.030 67.695 198.515 ;
        RECT 66.965 197.435 67.195 197.830 ;
        RECT 67.365 197.605 67.695 198.030 ;
        RECT 67.865 198.355 68.755 198.525 ;
        RECT 67.865 197.630 68.035 198.355 ;
        RECT 68.205 197.800 68.755 198.185 ;
        RECT 68.925 198.010 69.215 198.735 ;
        RECT 69.390 197.895 69.650 198.735 ;
        RECT 69.825 197.990 70.080 198.565 ;
        RECT 70.250 198.355 70.580 198.735 ;
        RECT 70.795 198.185 70.965 198.565 ;
        RECT 71.225 198.190 76.570 198.735 ;
        RECT 76.745 198.190 82.090 198.735 ;
        RECT 70.250 198.015 70.965 198.185 ;
        RECT 67.865 197.560 68.755 197.630 ;
        RECT 67.860 197.535 68.755 197.560 ;
        RECT 67.850 197.520 68.755 197.535 ;
        RECT 67.845 197.505 68.755 197.520 ;
        RECT 67.835 197.500 68.755 197.505 ;
        RECT 67.830 197.490 68.755 197.500 ;
        RECT 67.825 197.480 68.755 197.490 ;
        RECT 67.815 197.475 68.755 197.480 ;
        RECT 67.805 197.465 68.755 197.475 ;
        RECT 67.795 197.460 68.755 197.465 ;
        RECT 67.795 197.455 68.130 197.460 ;
        RECT 67.780 197.450 68.130 197.455 ;
        RECT 67.765 197.440 68.130 197.450 ;
        RECT 67.740 197.435 68.130 197.440 ;
        RECT 66.965 197.430 68.130 197.435 ;
        RECT 66.965 197.395 68.100 197.430 ;
        RECT 66.965 197.370 68.065 197.395 ;
        RECT 66.965 197.340 68.035 197.370 ;
        RECT 66.965 197.310 68.015 197.340 ;
        RECT 66.965 197.280 67.995 197.310 ;
        RECT 66.965 197.270 67.925 197.280 ;
        RECT 66.965 197.260 67.900 197.270 ;
        RECT 66.965 197.245 67.880 197.260 ;
        RECT 66.965 197.230 67.860 197.245 ;
        RECT 67.070 197.220 67.855 197.230 ;
        RECT 67.070 197.185 67.840 197.220 ;
        RECT 66.625 196.355 66.900 197.055 ;
        RECT 67.070 196.935 67.825 197.185 ;
        RECT 67.995 196.865 68.325 197.110 ;
        RECT 68.495 197.010 68.755 197.460 ;
        RECT 68.140 196.840 68.325 196.865 ;
        RECT 68.140 196.740 68.755 196.840 ;
        RECT 67.070 196.185 67.325 196.730 ;
        RECT 67.495 196.355 67.975 196.695 ;
        RECT 68.150 196.185 68.755 196.740 ;
        RECT 68.925 196.185 69.215 197.350 ;
        RECT 69.390 196.185 69.650 197.335 ;
        RECT 69.825 197.260 69.995 197.990 ;
        RECT 70.250 197.825 70.420 198.015 ;
        RECT 70.165 197.495 70.420 197.825 ;
        RECT 70.250 197.285 70.420 197.495 ;
        RECT 70.700 197.465 71.055 197.835 ;
        RECT 72.810 197.360 73.150 198.190 ;
        RECT 69.825 196.355 70.080 197.260 ;
        RECT 70.250 197.115 70.965 197.285 ;
        RECT 70.250 196.185 70.580 196.945 ;
        RECT 70.795 196.355 70.965 197.115 ;
        RECT 74.630 196.620 74.980 197.870 ;
        RECT 78.330 197.360 78.670 198.190 ;
        RECT 82.265 197.965 84.855 198.735 ;
        RECT 80.150 196.620 80.500 197.870 ;
        RECT 82.265 197.445 83.475 197.965 ;
        RECT 83.645 197.275 84.855 197.795 ;
        RECT 71.225 196.185 76.570 196.620 ;
        RECT 76.745 196.185 82.090 196.620 ;
        RECT 82.265 196.185 84.855 197.275 ;
        RECT 85.485 197.790 85.825 198.565 ;
        RECT 85.995 198.275 86.165 198.735 ;
        RECT 86.405 198.300 86.765 198.565 ;
        RECT 86.405 198.295 86.760 198.300 ;
        RECT 86.405 198.285 86.755 198.295 ;
        RECT 86.405 198.280 86.750 198.285 ;
        RECT 86.405 198.270 86.745 198.280 ;
        RECT 87.395 198.275 87.565 198.735 ;
        RECT 86.405 198.265 86.740 198.270 ;
        RECT 86.405 198.255 86.730 198.265 ;
        RECT 86.405 198.245 86.720 198.255 ;
        RECT 86.405 198.105 86.705 198.245 ;
        RECT 85.995 197.915 86.705 198.105 ;
        RECT 86.895 198.105 87.225 198.185 ;
        RECT 87.735 198.105 88.075 198.565 ;
        RECT 88.245 198.190 93.590 198.735 ;
        RECT 86.895 197.915 88.075 198.105 ;
        RECT 85.485 196.355 85.765 197.790 ;
        RECT 85.995 197.345 86.280 197.915 ;
        RECT 86.465 197.515 86.935 197.745 ;
        RECT 87.105 197.725 87.435 197.745 ;
        RECT 87.105 197.545 87.555 197.725 ;
        RECT 87.745 197.545 88.075 197.745 ;
        RECT 85.995 197.130 87.145 197.345 ;
        RECT 85.935 196.185 86.645 196.960 ;
        RECT 86.815 196.355 87.145 197.130 ;
        RECT 87.340 196.430 87.555 197.545 ;
        RECT 87.845 197.205 88.075 197.545 ;
        RECT 89.830 197.360 90.170 198.190 ;
        RECT 94.685 198.010 94.975 198.735 ;
        RECT 95.165 197.925 95.405 198.735 ;
        RECT 95.575 197.925 95.905 198.565 ;
        RECT 96.075 197.925 96.345 198.735 ;
        RECT 96.525 198.190 101.870 198.735 ;
        RECT 102.045 198.190 107.390 198.735 ;
        RECT 87.735 196.185 88.065 196.905 ;
        RECT 91.650 196.620 92.000 197.870 ;
        RECT 95.145 197.495 95.495 197.745 ;
        RECT 88.245 196.185 93.590 196.620 ;
        RECT 94.685 196.185 94.975 197.350 ;
        RECT 95.665 197.325 95.835 197.925 ;
        RECT 96.005 197.495 96.355 197.745 ;
        RECT 98.110 197.360 98.450 198.190 ;
        RECT 95.155 197.155 95.835 197.325 ;
        RECT 95.155 196.370 95.485 197.155 ;
        RECT 96.015 196.185 96.345 197.325 ;
        RECT 99.930 196.620 100.280 197.870 ;
        RECT 103.630 197.360 103.970 198.190 ;
        RECT 107.565 197.965 110.155 198.735 ;
        RECT 110.900 198.105 111.185 198.565 ;
        RECT 111.355 198.275 111.625 198.735 ;
        RECT 105.450 196.620 105.800 197.870 ;
        RECT 107.565 197.445 108.775 197.965 ;
        RECT 110.900 197.935 111.855 198.105 ;
        RECT 108.945 197.275 110.155 197.795 ;
        RECT 96.525 196.185 101.870 196.620 ;
        RECT 102.045 196.185 107.390 196.620 ;
        RECT 107.565 196.185 110.155 197.275 ;
        RECT 110.785 197.205 111.475 197.765 ;
        RECT 111.645 197.035 111.855 197.935 ;
        RECT 110.900 196.815 111.855 197.035 ;
        RECT 112.025 197.765 112.425 198.565 ;
        RECT 112.615 198.105 112.895 198.565 ;
        RECT 113.415 198.275 113.740 198.735 ;
        RECT 112.615 197.935 113.740 198.105 ;
        RECT 113.910 197.995 114.295 198.565 ;
        RECT 114.465 198.190 119.810 198.735 ;
        RECT 113.290 197.825 113.740 197.935 ;
        RECT 112.025 197.205 113.120 197.765 ;
        RECT 113.290 197.495 113.845 197.825 ;
        RECT 110.900 196.355 111.185 196.815 ;
        RECT 111.355 196.185 111.625 196.645 ;
        RECT 112.025 196.355 112.425 197.205 ;
        RECT 113.290 197.035 113.740 197.495 ;
        RECT 114.015 197.325 114.295 197.995 ;
        RECT 116.050 197.360 116.390 198.190 ;
        RECT 120.445 198.010 120.735 198.735 ;
        RECT 120.905 198.190 126.250 198.735 ;
        RECT 126.425 198.190 131.770 198.735 ;
        RECT 131.945 198.190 137.290 198.735 ;
        RECT 137.465 198.190 142.810 198.735 ;
        RECT 112.615 196.815 113.740 197.035 ;
        RECT 112.615 196.355 112.895 196.815 ;
        RECT 113.415 196.185 113.740 196.645 ;
        RECT 113.910 196.355 114.295 197.325 ;
        RECT 117.870 196.620 118.220 197.870 ;
        RECT 122.490 197.360 122.830 198.190 ;
        RECT 114.465 196.185 119.810 196.620 ;
        RECT 120.445 196.185 120.735 197.350 ;
        RECT 124.310 196.620 124.660 197.870 ;
        RECT 128.010 197.360 128.350 198.190 ;
        RECT 129.830 196.620 130.180 197.870 ;
        RECT 133.530 197.360 133.870 198.190 ;
        RECT 135.350 196.620 135.700 197.870 ;
        RECT 139.050 197.360 139.390 198.190 ;
        RECT 142.985 197.965 145.575 198.735 ;
        RECT 145.745 197.985 146.955 198.735 ;
        RECT 140.870 196.620 141.220 197.870 ;
        RECT 142.985 197.445 144.195 197.965 ;
        RECT 144.365 197.275 145.575 197.795 ;
        RECT 120.905 196.185 126.250 196.620 ;
        RECT 126.425 196.185 131.770 196.620 ;
        RECT 131.945 196.185 137.290 196.620 ;
        RECT 137.465 196.185 142.810 196.620 ;
        RECT 142.985 196.185 145.575 197.275 ;
        RECT 145.745 197.275 146.265 197.815 ;
        RECT 146.435 197.445 146.955 197.985 ;
        RECT 145.745 196.185 146.955 197.275 ;
        RECT 17.320 196.015 147.040 196.185 ;
        RECT 17.405 194.925 18.615 196.015 ;
        RECT 18.785 195.580 24.130 196.015 ;
        RECT 17.405 194.215 17.925 194.755 ;
        RECT 18.095 194.385 18.615 194.925 ;
        RECT 17.405 193.465 18.615 194.215 ;
        RECT 20.370 194.010 20.710 194.840 ;
        RECT 22.190 194.330 22.540 195.580 ;
        RECT 24.305 194.925 25.975 196.015 ;
        RECT 24.305 194.235 25.055 194.755 ;
        RECT 25.225 194.405 25.975 194.925 ;
        RECT 26.155 195.045 26.485 195.845 ;
        RECT 26.655 195.215 26.885 196.015 ;
        RECT 27.055 195.045 27.385 195.845 ;
        RECT 26.155 194.875 27.385 195.045 ;
        RECT 27.555 194.875 27.810 196.015 ;
        RECT 27.985 194.925 29.655 196.015 ;
        RECT 26.145 194.375 26.455 194.705 ;
        RECT 18.785 193.465 24.130 194.010 ;
        RECT 24.305 193.465 25.975 194.235 ;
        RECT 26.155 193.975 26.485 194.205 ;
        RECT 26.660 194.145 27.035 194.705 ;
        RECT 27.205 193.975 27.385 194.875 ;
        RECT 27.570 194.125 27.790 194.705 ;
        RECT 27.985 194.235 28.735 194.755 ;
        RECT 28.905 194.405 29.655 194.925 ;
        RECT 30.285 194.850 30.575 196.015 ;
        RECT 30.745 195.580 36.090 196.015 ;
        RECT 26.155 193.635 27.385 193.975 ;
        RECT 27.555 193.465 27.810 193.955 ;
        RECT 27.985 193.465 29.655 194.235 ;
        RECT 30.285 193.465 30.575 194.190 ;
        RECT 32.330 194.010 32.670 194.840 ;
        RECT 34.150 194.330 34.500 195.580 ;
        RECT 36.265 194.925 38.855 196.015 ;
        RECT 36.265 194.235 37.475 194.755 ;
        RECT 37.645 194.405 38.855 194.925 ;
        RECT 39.025 195.045 39.295 195.815 ;
        RECT 39.465 195.235 39.795 196.015 ;
        RECT 40.000 195.410 40.185 195.815 ;
        RECT 40.355 195.590 40.690 196.015 ;
        RECT 40.865 195.580 46.210 196.015 ;
        RECT 46.385 195.580 51.730 196.015 ;
        RECT 40.000 195.235 40.665 195.410 ;
        RECT 39.025 194.875 40.155 195.045 ;
        RECT 30.745 193.465 36.090 194.010 ;
        RECT 36.265 193.465 38.855 194.235 ;
        RECT 39.025 193.965 39.195 194.875 ;
        RECT 39.365 194.125 39.725 194.705 ;
        RECT 39.905 194.375 40.155 194.875 ;
        RECT 40.325 194.205 40.665 195.235 ;
        RECT 39.980 194.035 40.665 194.205 ;
        RECT 39.025 193.635 39.285 193.965 ;
        RECT 39.495 193.465 39.770 193.945 ;
        RECT 39.980 193.635 40.185 194.035 ;
        RECT 42.450 194.010 42.790 194.840 ;
        RECT 44.270 194.330 44.620 195.580 ;
        RECT 47.970 194.010 48.310 194.840 ;
        RECT 49.790 194.330 50.140 195.580 ;
        RECT 51.905 194.925 53.575 196.015 ;
        RECT 51.905 194.235 52.655 194.755 ;
        RECT 52.825 194.405 53.575 194.925 ;
        RECT 53.930 195.045 54.320 195.220 ;
        RECT 54.805 195.215 55.135 196.015 ;
        RECT 55.305 195.225 55.840 195.845 ;
        RECT 53.930 194.875 55.355 195.045 ;
        RECT 40.355 193.465 40.690 193.865 ;
        RECT 40.865 193.465 46.210 194.010 ;
        RECT 46.385 193.465 51.730 194.010 ;
        RECT 51.905 193.465 53.575 194.235 ;
        RECT 53.805 194.145 54.160 194.705 ;
        RECT 54.330 193.975 54.500 194.875 ;
        RECT 54.670 194.145 54.935 194.705 ;
        RECT 55.185 194.375 55.355 194.875 ;
        RECT 55.525 194.205 55.840 195.225 ;
        RECT 56.045 194.850 56.335 196.015 ;
        RECT 56.515 195.295 56.845 196.015 ;
        RECT 56.505 194.655 56.735 194.995 ;
        RECT 57.025 194.655 57.240 195.770 ;
        RECT 57.435 195.070 57.765 195.845 ;
        RECT 57.935 195.240 58.645 196.015 ;
        RECT 57.435 194.855 58.585 195.070 ;
        RECT 56.505 194.455 56.835 194.655 ;
        RECT 57.025 194.475 57.475 194.655 ;
        RECT 57.145 194.455 57.475 194.475 ;
        RECT 57.645 194.455 58.115 194.685 ;
        RECT 58.300 194.285 58.585 194.855 ;
        RECT 58.815 194.410 59.095 195.845 ;
        RECT 59.275 195.065 59.550 195.835 ;
        RECT 59.720 195.405 60.050 195.835 ;
        RECT 60.220 195.575 60.415 196.015 ;
        RECT 60.595 195.405 60.925 195.835 ;
        RECT 61.105 195.580 66.450 196.015 ;
        RECT 66.625 195.580 71.970 196.015 ;
        RECT 72.145 195.580 77.490 196.015 ;
        RECT 59.720 195.235 60.925 195.405 ;
        RECT 59.275 194.875 59.860 195.065 ;
        RECT 60.030 194.905 60.925 195.235 ;
        RECT 53.910 193.465 54.150 193.975 ;
        RECT 54.330 193.645 54.610 193.975 ;
        RECT 54.840 193.465 55.055 193.975 ;
        RECT 55.225 193.635 55.840 194.205 ;
        RECT 56.045 193.465 56.335 194.190 ;
        RECT 56.505 194.095 57.685 194.285 ;
        RECT 56.505 193.635 56.845 194.095 ;
        RECT 57.355 194.015 57.685 194.095 ;
        RECT 57.875 194.095 58.585 194.285 ;
        RECT 57.875 193.955 58.175 194.095 ;
        RECT 57.860 193.945 58.175 193.955 ;
        RECT 57.850 193.935 58.175 193.945 ;
        RECT 57.840 193.930 58.175 193.935 ;
        RECT 57.015 193.465 57.185 193.925 ;
        RECT 57.835 193.920 58.175 193.930 ;
        RECT 57.830 193.915 58.175 193.920 ;
        RECT 57.825 193.905 58.175 193.915 ;
        RECT 57.820 193.900 58.175 193.905 ;
        RECT 57.815 193.635 58.175 193.900 ;
        RECT 58.415 193.465 58.585 193.925 ;
        RECT 58.755 193.635 59.095 194.410 ;
        RECT 59.275 194.055 59.515 194.705 ;
        RECT 59.685 194.205 59.860 194.875 ;
        RECT 60.030 194.375 60.445 194.705 ;
        RECT 60.625 194.375 60.920 194.705 ;
        RECT 59.685 194.025 60.015 194.205 ;
        RECT 59.290 193.465 59.620 193.855 ;
        RECT 59.790 193.645 60.015 194.025 ;
        RECT 60.215 193.755 60.445 194.375 ;
        RECT 60.625 193.465 60.925 194.195 ;
        RECT 62.690 194.010 63.030 194.840 ;
        RECT 64.510 194.330 64.860 195.580 ;
        RECT 68.210 194.010 68.550 194.840 ;
        RECT 70.030 194.330 70.380 195.580 ;
        RECT 73.730 194.010 74.070 194.840 ;
        RECT 75.550 194.330 75.900 195.580 ;
        RECT 77.665 194.925 79.335 196.015 ;
        RECT 77.665 194.235 78.415 194.755 ;
        RECT 78.585 194.405 79.335 194.925 ;
        RECT 79.970 194.875 80.290 196.015 ;
        RECT 80.470 194.705 80.665 195.755 ;
        RECT 80.845 195.165 81.175 195.845 ;
        RECT 81.375 195.215 81.630 196.015 ;
        RECT 80.845 194.885 81.195 195.165 ;
        RECT 80.030 194.655 80.290 194.705 ;
        RECT 80.025 194.485 80.290 194.655 ;
        RECT 80.030 194.375 80.290 194.485 ;
        RECT 80.470 194.375 80.855 194.705 ;
        RECT 81.025 194.505 81.195 194.885 ;
        RECT 81.385 194.675 81.630 195.035 ;
        RECT 81.805 194.850 82.095 196.015 ;
        RECT 82.355 195.345 82.525 195.845 ;
        RECT 82.695 195.515 83.025 196.015 ;
        RECT 82.355 195.175 83.020 195.345 ;
        RECT 81.025 194.335 81.545 194.505 ;
        RECT 82.270 194.355 82.620 195.005 ;
        RECT 61.105 193.465 66.450 194.010 ;
        RECT 66.625 193.465 71.970 194.010 ;
        RECT 72.145 193.465 77.490 194.010 ;
        RECT 77.665 193.465 79.335 194.235 ;
        RECT 79.970 193.995 81.185 194.165 ;
        RECT 79.970 193.645 80.260 193.995 ;
        RECT 80.455 193.465 80.785 193.825 ;
        RECT 80.955 193.690 81.185 193.995 ;
        RECT 81.375 193.975 81.545 194.335 ;
        RECT 81.375 193.805 81.575 193.975 ;
        RECT 81.375 193.770 81.545 193.805 ;
        RECT 81.805 193.465 82.095 194.190 ;
        RECT 82.790 194.185 83.020 195.175 ;
        RECT 82.355 194.015 83.020 194.185 ;
        RECT 82.355 193.725 82.525 194.015 ;
        RECT 82.695 193.465 83.025 193.845 ;
        RECT 83.195 193.725 83.380 195.845 ;
        RECT 83.620 195.555 83.885 196.015 ;
        RECT 84.055 195.420 84.305 195.845 ;
        RECT 84.515 195.570 85.620 195.740 ;
        RECT 84.000 195.290 84.305 195.420 ;
        RECT 83.550 194.095 83.830 195.045 ;
        RECT 84.000 194.185 84.170 195.290 ;
        RECT 84.340 194.505 84.580 195.100 ;
        RECT 84.750 195.035 85.280 195.400 ;
        RECT 84.750 194.335 84.920 195.035 ;
        RECT 85.450 194.955 85.620 195.570 ;
        RECT 85.790 195.215 85.960 196.015 ;
        RECT 86.130 195.515 86.380 195.845 ;
        RECT 86.605 195.545 87.490 195.715 ;
        RECT 85.450 194.865 85.960 194.955 ;
        RECT 84.000 194.055 84.225 194.185 ;
        RECT 84.395 194.115 84.920 194.335 ;
        RECT 85.090 194.695 85.960 194.865 ;
        RECT 83.635 193.465 83.885 193.925 ;
        RECT 84.055 193.915 84.225 194.055 ;
        RECT 85.090 193.915 85.260 194.695 ;
        RECT 85.790 194.625 85.960 194.695 ;
        RECT 85.470 194.445 85.670 194.475 ;
        RECT 86.130 194.445 86.300 195.515 ;
        RECT 86.470 194.625 86.660 195.345 ;
        RECT 85.470 194.145 86.300 194.445 ;
        RECT 86.830 194.415 87.150 195.375 ;
        RECT 84.055 193.745 84.390 193.915 ;
        RECT 84.585 193.745 85.260 193.915 ;
        RECT 85.580 193.465 85.950 193.965 ;
        RECT 86.130 193.915 86.300 194.145 ;
        RECT 86.685 194.085 87.150 194.415 ;
        RECT 87.320 194.705 87.490 195.545 ;
        RECT 87.670 195.515 87.985 196.015 ;
        RECT 88.215 195.285 88.555 195.845 ;
        RECT 87.660 194.910 88.555 195.285 ;
        RECT 88.725 195.005 88.895 196.015 ;
        RECT 88.365 194.705 88.555 194.910 ;
        RECT 89.065 194.955 89.395 195.800 ;
        RECT 89.065 194.875 89.455 194.955 ;
        RECT 89.240 194.825 89.455 194.875 ;
        RECT 87.320 194.375 88.195 194.705 ;
        RECT 88.365 194.375 89.115 194.705 ;
        RECT 87.320 193.915 87.490 194.375 ;
        RECT 88.365 194.205 88.565 194.375 ;
        RECT 89.285 194.245 89.455 194.825 ;
        RECT 89.230 194.205 89.455 194.245 ;
        RECT 86.130 193.745 86.535 193.915 ;
        RECT 86.705 193.745 87.490 193.915 ;
        RECT 87.765 193.465 87.975 193.995 ;
        RECT 88.235 193.680 88.565 194.205 ;
        RECT 89.075 194.120 89.455 194.205 ;
        RECT 89.625 194.875 90.010 195.845 ;
        RECT 90.180 195.555 90.505 196.015 ;
        RECT 91.025 195.385 91.305 195.845 ;
        RECT 90.180 195.165 91.305 195.385 ;
        RECT 89.625 194.205 89.905 194.875 ;
        RECT 90.180 194.705 90.630 195.165 ;
        RECT 91.495 194.995 91.895 195.845 ;
        RECT 92.295 195.555 92.565 196.015 ;
        RECT 92.735 195.385 93.020 195.845 ;
        RECT 90.075 194.375 90.630 194.705 ;
        RECT 90.800 194.435 91.895 194.995 ;
        RECT 90.180 194.265 90.630 194.375 ;
        RECT 88.735 193.465 88.905 194.075 ;
        RECT 89.075 193.685 89.405 194.120 ;
        RECT 89.625 193.635 90.010 194.205 ;
        RECT 90.180 194.095 91.305 194.265 ;
        RECT 90.180 193.465 90.505 193.925 ;
        RECT 91.025 193.635 91.305 194.095 ;
        RECT 91.495 193.635 91.895 194.435 ;
        RECT 92.065 195.165 93.020 195.385 ;
        RECT 92.065 194.265 92.275 195.165 ;
        RECT 92.445 194.435 93.135 194.995 ;
        RECT 93.305 194.875 93.580 195.845 ;
        RECT 93.790 195.215 94.070 196.015 ;
        RECT 94.240 195.505 95.855 195.835 ;
        RECT 94.240 195.165 95.415 195.335 ;
        RECT 94.240 195.045 94.410 195.165 ;
        RECT 93.750 194.875 94.410 195.045 ;
        RECT 92.065 194.095 93.020 194.265 ;
        RECT 92.295 193.465 92.565 193.925 ;
        RECT 92.735 193.635 93.020 194.095 ;
        RECT 93.305 194.140 93.475 194.875 ;
        RECT 93.750 194.705 93.920 194.875 ;
        RECT 94.670 194.705 94.915 194.995 ;
        RECT 95.085 194.875 95.415 195.165 ;
        RECT 95.675 194.705 95.845 195.265 ;
        RECT 96.095 194.875 96.355 196.015 ;
        RECT 96.615 195.345 96.785 195.845 ;
        RECT 96.955 195.515 97.285 196.015 ;
        RECT 96.615 195.175 97.280 195.345 ;
        RECT 93.645 194.375 93.920 194.705 ;
        RECT 94.090 194.375 94.915 194.705 ;
        RECT 95.130 194.375 95.845 194.705 ;
        RECT 96.015 194.455 96.350 194.705 ;
        RECT 93.750 194.205 93.920 194.375 ;
        RECT 95.595 194.285 95.845 194.375 ;
        RECT 96.530 194.355 96.880 195.005 ;
        RECT 93.305 193.795 93.580 194.140 ;
        RECT 93.750 194.035 95.415 194.205 ;
        RECT 93.770 193.465 94.145 193.865 ;
        RECT 94.315 193.685 94.485 194.035 ;
        RECT 94.655 193.465 94.985 193.865 ;
        RECT 95.155 193.635 95.415 194.035 ;
        RECT 95.595 193.865 95.925 194.285 ;
        RECT 96.095 193.465 96.355 194.285 ;
        RECT 97.050 194.185 97.280 195.175 ;
        RECT 96.615 194.015 97.280 194.185 ;
        RECT 96.615 193.725 96.785 194.015 ;
        RECT 96.955 193.465 97.285 193.845 ;
        RECT 97.455 193.725 97.640 195.845 ;
        RECT 97.880 195.555 98.145 196.015 ;
        RECT 98.315 195.420 98.565 195.845 ;
        RECT 98.775 195.570 99.880 195.740 ;
        RECT 98.260 195.290 98.565 195.420 ;
        RECT 97.810 194.095 98.090 195.045 ;
        RECT 98.260 194.185 98.430 195.290 ;
        RECT 98.600 194.505 98.840 195.100 ;
        RECT 99.010 195.035 99.540 195.400 ;
        RECT 99.010 194.335 99.180 195.035 ;
        RECT 99.710 194.955 99.880 195.570 ;
        RECT 100.050 195.215 100.220 196.015 ;
        RECT 100.390 195.515 100.640 195.845 ;
        RECT 100.865 195.545 101.750 195.715 ;
        RECT 99.710 194.865 100.220 194.955 ;
        RECT 98.260 194.055 98.485 194.185 ;
        RECT 98.655 194.115 99.180 194.335 ;
        RECT 99.350 194.695 100.220 194.865 ;
        RECT 97.895 193.465 98.145 193.925 ;
        RECT 98.315 193.915 98.485 194.055 ;
        RECT 99.350 193.915 99.520 194.695 ;
        RECT 100.050 194.625 100.220 194.695 ;
        RECT 99.730 194.445 99.930 194.475 ;
        RECT 100.390 194.445 100.560 195.515 ;
        RECT 100.730 194.625 100.920 195.345 ;
        RECT 99.730 194.145 100.560 194.445 ;
        RECT 101.090 194.415 101.410 195.375 ;
        RECT 98.315 193.745 98.650 193.915 ;
        RECT 98.845 193.745 99.520 193.915 ;
        RECT 99.840 193.465 100.210 193.965 ;
        RECT 100.390 193.915 100.560 194.145 ;
        RECT 100.945 194.085 101.410 194.415 ;
        RECT 101.580 194.705 101.750 195.545 ;
        RECT 101.930 195.515 102.245 196.015 ;
        RECT 102.475 195.285 102.815 195.845 ;
        RECT 101.920 194.910 102.815 195.285 ;
        RECT 102.985 195.005 103.155 196.015 ;
        RECT 102.625 194.705 102.815 194.910 ;
        RECT 103.325 194.955 103.655 195.800 ;
        RECT 103.325 194.875 103.715 194.955 ;
        RECT 103.500 194.825 103.715 194.875 ;
        RECT 101.580 194.375 102.455 194.705 ;
        RECT 102.625 194.375 103.375 194.705 ;
        RECT 101.580 193.915 101.750 194.375 ;
        RECT 102.625 194.205 102.825 194.375 ;
        RECT 103.545 194.245 103.715 194.825 ;
        RECT 103.490 194.205 103.715 194.245 ;
        RECT 100.390 193.745 100.795 193.915 ;
        RECT 100.965 193.745 101.750 193.915 ;
        RECT 102.025 193.465 102.235 193.995 ;
        RECT 102.495 193.680 102.825 194.205 ;
        RECT 103.335 194.120 103.715 194.205 ;
        RECT 103.885 194.875 104.270 195.845 ;
        RECT 104.440 195.555 104.765 196.015 ;
        RECT 105.285 195.385 105.565 195.845 ;
        RECT 104.440 195.165 105.565 195.385 ;
        RECT 103.885 194.205 104.165 194.875 ;
        RECT 104.440 194.705 104.890 195.165 ;
        RECT 105.755 194.995 106.155 195.845 ;
        RECT 106.555 195.555 106.825 196.015 ;
        RECT 106.995 195.385 107.280 195.845 ;
        RECT 104.335 194.375 104.890 194.705 ;
        RECT 105.060 194.435 106.155 194.995 ;
        RECT 104.440 194.265 104.890 194.375 ;
        RECT 102.995 193.465 103.165 194.075 ;
        RECT 103.335 193.685 103.665 194.120 ;
        RECT 103.885 193.635 104.270 194.205 ;
        RECT 104.440 194.095 105.565 194.265 ;
        RECT 104.440 193.465 104.765 193.925 ;
        RECT 105.285 193.635 105.565 194.095 ;
        RECT 105.755 193.635 106.155 194.435 ;
        RECT 106.325 195.165 107.280 195.385 ;
        RECT 106.325 194.265 106.535 195.165 ;
        RECT 106.705 194.435 107.395 194.995 ;
        RECT 107.565 194.850 107.855 196.015 ;
        RECT 108.545 194.955 108.875 195.800 ;
        RECT 109.045 195.005 109.215 196.015 ;
        RECT 109.385 195.285 109.725 195.845 ;
        RECT 109.955 195.515 110.270 196.015 ;
        RECT 110.450 195.545 111.335 195.715 ;
        RECT 108.485 194.875 108.875 194.955 ;
        RECT 109.385 194.910 110.280 195.285 ;
        RECT 108.485 194.825 108.700 194.875 ;
        RECT 106.325 194.095 107.280 194.265 ;
        RECT 108.485 194.245 108.655 194.825 ;
        RECT 109.385 194.705 109.575 194.910 ;
        RECT 110.450 194.705 110.620 195.545 ;
        RECT 111.560 195.515 111.810 195.845 ;
        RECT 108.825 194.375 109.575 194.705 ;
        RECT 109.745 194.375 110.620 194.705 ;
        RECT 108.485 194.205 108.710 194.245 ;
        RECT 109.375 194.205 109.575 194.375 ;
        RECT 106.555 193.465 106.825 193.925 ;
        RECT 106.995 193.635 107.280 194.095 ;
        RECT 107.565 193.465 107.855 194.190 ;
        RECT 108.485 194.120 108.865 194.205 ;
        RECT 108.535 193.685 108.865 194.120 ;
        RECT 109.035 193.465 109.205 194.075 ;
        RECT 109.375 193.680 109.705 194.205 ;
        RECT 109.965 193.465 110.175 193.995 ;
        RECT 110.450 193.915 110.620 194.375 ;
        RECT 110.790 194.415 111.110 195.375 ;
        RECT 111.280 194.625 111.470 195.345 ;
        RECT 111.640 194.445 111.810 195.515 ;
        RECT 111.980 195.215 112.150 196.015 ;
        RECT 112.320 195.570 113.425 195.740 ;
        RECT 112.320 194.955 112.490 195.570 ;
        RECT 113.635 195.420 113.885 195.845 ;
        RECT 114.055 195.555 114.320 196.015 ;
        RECT 112.660 195.035 113.190 195.400 ;
        RECT 113.635 195.290 113.940 195.420 ;
        RECT 111.980 194.865 112.490 194.955 ;
        RECT 111.980 194.695 112.850 194.865 ;
        RECT 111.980 194.625 112.150 194.695 ;
        RECT 112.270 194.445 112.470 194.475 ;
        RECT 110.790 194.085 111.255 194.415 ;
        RECT 111.640 194.145 112.470 194.445 ;
        RECT 111.640 193.915 111.810 194.145 ;
        RECT 110.450 193.745 111.235 193.915 ;
        RECT 111.405 193.745 111.810 193.915 ;
        RECT 111.990 193.465 112.360 193.965 ;
        RECT 112.680 193.915 112.850 194.695 ;
        RECT 113.020 194.335 113.190 195.035 ;
        RECT 113.360 194.505 113.600 195.100 ;
        RECT 113.020 194.115 113.545 194.335 ;
        RECT 113.770 194.185 113.940 195.290 ;
        RECT 113.715 194.055 113.940 194.185 ;
        RECT 114.110 194.095 114.390 195.045 ;
        RECT 113.715 193.915 113.885 194.055 ;
        RECT 112.680 193.745 113.355 193.915 ;
        RECT 113.550 193.745 113.885 193.915 ;
        RECT 114.055 193.465 114.305 193.925 ;
        RECT 114.560 193.725 114.745 195.845 ;
        RECT 114.915 195.515 115.245 196.015 ;
        RECT 115.415 195.345 115.585 195.845 ;
        RECT 115.845 195.580 121.190 196.015 ;
        RECT 121.365 195.580 126.710 196.015 ;
        RECT 126.885 195.580 132.230 196.015 ;
        RECT 114.920 195.175 115.585 195.345 ;
        RECT 114.920 194.185 115.150 195.175 ;
        RECT 115.320 194.355 115.670 195.005 ;
        RECT 114.920 194.015 115.585 194.185 ;
        RECT 114.915 193.465 115.245 193.845 ;
        RECT 115.415 193.725 115.585 194.015 ;
        RECT 117.430 194.010 117.770 194.840 ;
        RECT 119.250 194.330 119.600 195.580 ;
        RECT 122.950 194.010 123.290 194.840 ;
        RECT 124.770 194.330 125.120 195.580 ;
        RECT 128.470 194.010 128.810 194.840 ;
        RECT 130.290 194.330 130.640 195.580 ;
        RECT 133.325 194.850 133.615 196.015 ;
        RECT 133.785 195.580 139.130 196.015 ;
        RECT 139.305 195.580 144.650 196.015 ;
        RECT 115.845 193.465 121.190 194.010 ;
        RECT 121.365 193.465 126.710 194.010 ;
        RECT 126.885 193.465 132.230 194.010 ;
        RECT 133.325 193.465 133.615 194.190 ;
        RECT 135.370 194.010 135.710 194.840 ;
        RECT 137.190 194.330 137.540 195.580 ;
        RECT 140.890 194.010 141.230 194.840 ;
        RECT 142.710 194.330 143.060 195.580 ;
        RECT 145.745 194.925 146.955 196.015 ;
        RECT 145.745 194.385 146.265 194.925 ;
        RECT 146.435 194.215 146.955 194.755 ;
        RECT 133.785 193.465 139.130 194.010 ;
        RECT 139.305 193.465 144.650 194.010 ;
        RECT 145.745 193.465 146.955 194.215 ;
        RECT 17.320 193.295 147.040 193.465 ;
        RECT 17.405 192.545 18.615 193.295 ;
        RECT 18.875 192.745 19.045 193.125 ;
        RECT 19.225 192.915 19.555 193.295 ;
        RECT 18.875 192.575 19.540 192.745 ;
        RECT 19.735 192.620 19.995 193.125 ;
        RECT 17.405 192.005 17.925 192.545 ;
        RECT 18.095 191.835 18.615 192.375 ;
        RECT 18.805 192.025 19.135 192.395 ;
        RECT 19.370 192.320 19.540 192.575 ;
        RECT 19.370 191.990 19.655 192.320 ;
        RECT 19.370 191.845 19.540 191.990 ;
        RECT 17.405 190.745 18.615 191.835 ;
        RECT 18.875 191.675 19.540 191.845 ;
        RECT 19.825 191.820 19.995 192.620 ;
        RECT 20.165 192.545 21.375 193.295 ;
        RECT 21.550 192.790 21.885 193.295 ;
        RECT 22.055 192.725 22.295 193.100 ;
        RECT 22.575 192.965 22.745 193.110 ;
        RECT 22.575 192.770 22.950 192.965 ;
        RECT 23.310 192.800 23.705 193.295 ;
        RECT 20.165 192.005 20.685 192.545 ;
        RECT 20.855 191.835 21.375 192.375 ;
        RECT 18.875 190.915 19.045 191.675 ;
        RECT 19.225 190.745 19.555 191.505 ;
        RECT 19.725 190.915 19.995 191.820 ;
        RECT 20.165 190.745 21.375 191.835 ;
        RECT 21.605 191.765 21.905 192.615 ;
        RECT 22.075 192.575 22.295 192.725 ;
        RECT 22.075 192.245 22.610 192.575 ;
        RECT 22.780 192.435 22.950 192.770 ;
        RECT 23.875 192.605 24.115 193.125 ;
        RECT 22.075 191.595 22.310 192.245 ;
        RECT 22.780 192.075 23.765 192.435 ;
        RECT 21.635 191.365 22.310 191.595 ;
        RECT 22.480 192.055 23.765 192.075 ;
        RECT 22.480 191.905 23.340 192.055 ;
        RECT 21.635 190.935 21.805 191.365 ;
        RECT 21.975 190.745 22.305 191.195 ;
        RECT 22.480 190.960 22.765 191.905 ;
        RECT 23.940 191.800 24.115 192.605 ;
        RECT 25.315 192.745 25.485 193.035 ;
        RECT 25.655 192.915 25.985 193.295 ;
        RECT 25.315 192.575 25.980 192.745 ;
        RECT 22.940 191.425 23.635 191.735 ;
        RECT 22.945 190.745 23.630 191.215 ;
        RECT 23.810 191.015 24.115 191.800 ;
        RECT 25.230 191.755 25.580 192.405 ;
        RECT 25.750 191.585 25.980 192.575 ;
        RECT 25.315 191.415 25.980 191.585 ;
        RECT 25.315 190.915 25.485 191.415 ;
        RECT 25.655 190.745 25.985 191.245 ;
        RECT 26.155 190.915 26.340 193.035 ;
        RECT 26.595 192.835 26.845 193.295 ;
        RECT 27.015 192.845 27.350 193.015 ;
        RECT 27.545 192.845 28.220 193.015 ;
        RECT 27.015 192.705 27.185 192.845 ;
        RECT 26.510 191.715 26.790 192.665 ;
        RECT 26.960 192.575 27.185 192.705 ;
        RECT 26.960 191.470 27.130 192.575 ;
        RECT 27.355 192.425 27.880 192.645 ;
        RECT 27.300 191.660 27.540 192.255 ;
        RECT 27.710 191.725 27.880 192.425 ;
        RECT 28.050 192.065 28.220 192.845 ;
        RECT 28.540 192.795 28.910 193.295 ;
        RECT 29.090 192.845 29.495 193.015 ;
        RECT 29.665 192.845 30.450 193.015 ;
        RECT 29.090 192.615 29.260 192.845 ;
        RECT 28.430 192.315 29.260 192.615 ;
        RECT 29.645 192.345 30.110 192.675 ;
        RECT 28.430 192.285 28.630 192.315 ;
        RECT 28.750 192.065 28.920 192.135 ;
        RECT 28.050 191.895 28.920 192.065 ;
        RECT 28.410 191.805 28.920 191.895 ;
        RECT 26.960 191.340 27.265 191.470 ;
        RECT 27.710 191.360 28.240 191.725 ;
        RECT 26.580 190.745 26.845 191.205 ;
        RECT 27.015 190.915 27.265 191.340 ;
        RECT 28.410 191.190 28.580 191.805 ;
        RECT 27.475 191.020 28.580 191.190 ;
        RECT 28.750 190.745 28.920 191.545 ;
        RECT 29.090 191.245 29.260 192.315 ;
        RECT 29.430 191.415 29.620 192.135 ;
        RECT 29.790 191.385 30.110 192.345 ;
        RECT 30.280 192.385 30.450 192.845 ;
        RECT 30.725 192.765 30.935 193.295 ;
        RECT 31.195 192.555 31.525 193.080 ;
        RECT 31.695 192.685 31.865 193.295 ;
        RECT 32.035 192.640 32.365 193.075 ;
        RECT 32.675 192.745 32.845 193.035 ;
        RECT 33.015 192.915 33.345 193.295 ;
        RECT 32.035 192.555 32.415 192.640 ;
        RECT 32.675 192.575 33.340 192.745 ;
        RECT 31.325 192.385 31.525 192.555 ;
        RECT 32.190 192.515 32.415 192.555 ;
        RECT 30.280 192.055 31.155 192.385 ;
        RECT 31.325 192.055 32.075 192.385 ;
        RECT 29.090 190.915 29.340 191.245 ;
        RECT 30.280 191.215 30.450 192.055 ;
        RECT 31.325 191.850 31.515 192.055 ;
        RECT 32.245 191.935 32.415 192.515 ;
        RECT 32.200 191.885 32.415 191.935 ;
        RECT 30.620 191.475 31.515 191.850 ;
        RECT 32.025 191.805 32.415 191.885 ;
        RECT 29.565 191.045 30.450 191.215 ;
        RECT 30.630 190.745 30.945 191.245 ;
        RECT 31.175 190.915 31.515 191.475 ;
        RECT 31.685 190.745 31.855 191.755 ;
        RECT 32.025 190.960 32.355 191.805 ;
        RECT 32.590 191.755 32.940 192.405 ;
        RECT 33.110 191.585 33.340 192.575 ;
        RECT 32.675 191.415 33.340 191.585 ;
        RECT 32.675 190.915 32.845 191.415 ;
        RECT 33.015 190.745 33.345 191.245 ;
        RECT 33.515 190.915 33.700 193.035 ;
        RECT 33.955 192.835 34.205 193.295 ;
        RECT 34.375 192.845 34.710 193.015 ;
        RECT 34.905 192.845 35.580 193.015 ;
        RECT 34.375 192.705 34.545 192.845 ;
        RECT 33.870 191.715 34.150 192.665 ;
        RECT 34.320 192.575 34.545 192.705 ;
        RECT 34.320 191.470 34.490 192.575 ;
        RECT 34.715 192.425 35.240 192.645 ;
        RECT 34.660 191.660 34.900 192.255 ;
        RECT 35.070 191.725 35.240 192.425 ;
        RECT 35.410 192.065 35.580 192.845 ;
        RECT 35.900 192.795 36.270 193.295 ;
        RECT 36.450 192.845 36.855 193.015 ;
        RECT 37.025 192.845 37.810 193.015 ;
        RECT 36.450 192.615 36.620 192.845 ;
        RECT 35.790 192.315 36.620 192.615 ;
        RECT 37.005 192.345 37.470 192.675 ;
        RECT 35.790 192.285 35.990 192.315 ;
        RECT 36.110 192.065 36.280 192.135 ;
        RECT 35.410 191.895 36.280 192.065 ;
        RECT 35.770 191.805 36.280 191.895 ;
        RECT 34.320 191.340 34.625 191.470 ;
        RECT 35.070 191.360 35.600 191.725 ;
        RECT 33.940 190.745 34.205 191.205 ;
        RECT 34.375 190.915 34.625 191.340 ;
        RECT 35.770 191.190 35.940 191.805 ;
        RECT 34.835 191.020 35.940 191.190 ;
        RECT 36.110 190.745 36.280 191.545 ;
        RECT 36.450 191.245 36.620 192.315 ;
        RECT 36.790 191.415 36.980 192.135 ;
        RECT 37.150 191.385 37.470 192.345 ;
        RECT 37.640 192.385 37.810 192.845 ;
        RECT 38.085 192.765 38.295 193.295 ;
        RECT 38.555 192.555 38.885 193.080 ;
        RECT 39.055 192.685 39.225 193.295 ;
        RECT 39.395 192.640 39.725 193.075 ;
        RECT 39.395 192.555 39.775 192.640 ;
        RECT 38.685 192.385 38.885 192.555 ;
        RECT 39.550 192.515 39.775 192.555 ;
        RECT 37.640 192.055 38.515 192.385 ;
        RECT 38.685 192.055 39.435 192.385 ;
        RECT 36.450 190.915 36.700 191.245 ;
        RECT 37.640 191.215 37.810 192.055 ;
        RECT 38.685 191.850 38.875 192.055 ;
        RECT 39.605 191.935 39.775 192.515 ;
        RECT 39.965 192.485 40.205 193.295 ;
        RECT 40.375 192.485 40.705 193.125 ;
        RECT 40.875 192.485 41.145 193.295 ;
        RECT 39.945 192.055 40.295 192.305 ;
        RECT 39.560 191.885 39.775 191.935 ;
        RECT 40.465 191.885 40.635 192.485 ;
        RECT 41.330 192.455 41.590 193.295 ;
        RECT 41.765 192.550 42.020 193.125 ;
        RECT 42.190 192.915 42.520 193.295 ;
        RECT 42.735 192.745 42.905 193.125 ;
        RECT 42.190 192.575 42.905 192.745 ;
        RECT 40.805 192.055 41.155 192.305 ;
        RECT 37.980 191.475 38.875 191.850 ;
        RECT 39.385 191.805 39.775 191.885 ;
        RECT 36.925 191.045 37.810 191.215 ;
        RECT 37.990 190.745 38.305 191.245 ;
        RECT 38.535 190.915 38.875 191.475 ;
        RECT 39.045 190.745 39.215 191.755 ;
        RECT 39.385 190.960 39.715 191.805 ;
        RECT 39.955 191.715 40.635 191.885 ;
        RECT 39.955 190.930 40.285 191.715 ;
        RECT 40.815 190.745 41.145 191.885 ;
        RECT 41.330 190.745 41.590 191.895 ;
        RECT 41.765 191.820 41.935 192.550 ;
        RECT 42.190 192.385 42.360 192.575 ;
        RECT 43.165 192.570 43.455 193.295 ;
        RECT 43.865 192.825 44.035 193.295 ;
        RECT 44.705 192.825 44.875 193.295 ;
        RECT 45.140 192.905 46.370 193.125 ;
        RECT 44.205 192.655 44.535 192.735 ;
        RECT 45.565 192.655 45.895 192.735 ;
        RECT 43.625 192.475 45.895 192.655 ;
        RECT 46.120 192.655 46.370 192.905 ;
        RECT 46.540 192.825 46.710 193.295 ;
        RECT 46.880 192.655 47.210 193.125 ;
        RECT 47.480 192.825 47.650 193.295 ;
        RECT 46.120 192.475 47.210 192.655 ;
        RECT 47.820 192.655 48.150 193.125 ;
        RECT 48.320 192.825 48.490 193.295 ;
        RECT 48.660 192.655 48.990 193.125 ;
        RECT 49.160 192.825 49.330 193.295 ;
        RECT 47.820 192.475 49.400 192.655 ;
        RECT 42.105 192.055 42.360 192.385 ;
        RECT 42.190 191.845 42.360 192.055 ;
        RECT 42.640 192.025 42.995 192.395 ;
        RECT 43.625 191.965 44.035 192.475 ;
        RECT 44.245 192.135 44.905 192.305 ;
        RECT 41.765 190.915 42.020 191.820 ;
        RECT 42.190 191.675 42.905 191.845 ;
        RECT 42.190 190.745 42.520 191.505 ;
        RECT 42.735 190.915 42.905 191.675 ;
        RECT 43.165 190.745 43.455 191.910 ;
        RECT 43.625 191.755 44.495 191.965 ;
        RECT 44.735 191.935 44.905 192.135 ;
        RECT 45.430 192.105 46.100 192.305 ;
        RECT 46.290 192.105 47.810 192.305 ;
        RECT 47.980 192.105 48.475 192.305 ;
        RECT 48.645 192.105 48.975 192.305 ;
        RECT 47.640 191.935 47.810 192.105 ;
        RECT 48.645 191.935 48.815 192.105 ;
        RECT 44.735 191.765 47.470 191.935 ;
        RECT 47.640 191.765 48.815 191.935 ;
        RECT 43.825 191.085 44.075 191.585 ;
        RECT 44.245 191.255 44.495 191.755 ;
        RECT 47.300 191.595 47.470 191.765 ;
        RECT 49.230 191.595 49.400 192.475 ;
        RECT 49.605 192.545 50.815 193.295 ;
        RECT 50.985 192.785 51.325 193.295 ;
        RECT 49.605 192.005 50.125 192.545 ;
        RECT 50.295 191.835 50.815 192.375 ;
        RECT 50.995 192.055 51.335 192.615 ;
        RECT 51.505 192.385 51.755 193.115 ;
        RECT 52.080 192.755 52.265 193.115 ;
        RECT 52.445 192.925 52.775 193.295 ;
        RECT 52.955 192.755 53.180 193.115 ;
        RECT 53.830 192.795 54.325 193.125 ;
        RECT 52.080 192.565 53.560 192.755 ;
        RECT 51.505 192.055 52.145 192.385 ;
        RECT 52.325 192.055 52.655 192.385 ;
        RECT 44.665 191.425 47.130 191.595 ;
        RECT 47.300 191.425 49.400 191.595 ;
        RECT 44.665 191.085 45.435 191.425 ;
        RECT 43.825 190.915 45.435 191.085 ;
        RECT 45.605 190.745 45.910 191.245 ;
        RECT 46.080 190.915 46.330 191.425 ;
        RECT 46.920 191.255 47.130 191.425 ;
        RECT 47.860 191.255 48.110 191.425 ;
        RECT 46.500 190.745 46.750 191.245 ;
        RECT 46.920 190.915 47.235 191.255 ;
        RECT 48.285 191.245 48.455 191.255 ;
        RECT 49.205 191.245 49.375 191.255 ;
        RECT 47.440 191.085 47.690 191.245 ;
        RECT 48.280 191.085 48.530 191.245 ;
        RECT 47.440 190.915 48.530 191.085 ;
        RECT 48.700 190.745 48.950 191.245 ;
        RECT 49.120 190.915 49.400 191.245 ;
        RECT 49.605 190.745 50.815 191.835 ;
        RECT 51.150 191.655 52.255 191.855 ;
        RECT 51.150 190.925 51.400 191.655 ;
        RECT 51.570 190.745 51.900 191.475 ;
        RECT 52.070 190.925 52.255 191.655 ;
        RECT 52.425 190.925 52.655 192.055 ;
        RECT 52.835 191.765 53.135 192.385 ;
        RECT 53.345 191.595 53.560 192.565 ;
        RECT 52.835 190.925 53.560 191.595 ;
        RECT 53.745 191.305 53.985 192.615 ;
        RECT 54.155 191.885 54.325 192.795 ;
        RECT 54.545 192.055 54.895 193.020 ;
        RECT 55.075 192.055 55.375 193.025 ;
        RECT 55.555 192.055 55.835 193.025 ;
        RECT 56.015 192.495 56.285 193.295 ;
        RECT 56.455 192.575 56.795 193.085 ;
        RECT 56.965 192.795 57.305 193.295 ;
        RECT 56.030 192.055 56.360 192.305 ;
        RECT 56.030 191.885 56.345 192.055 ;
        RECT 54.155 191.715 56.345 191.885 ;
        RECT 53.750 190.745 54.085 191.125 ;
        RECT 54.255 190.915 54.505 191.715 ;
        RECT 54.725 190.745 55.055 191.465 ;
        RECT 55.240 190.915 55.490 191.715 ;
        RECT 55.955 190.745 56.285 191.545 ;
        RECT 56.535 191.175 56.795 192.575 ;
        RECT 56.965 192.055 57.305 192.625 ;
        RECT 57.475 192.385 57.720 193.075 ;
        RECT 57.915 192.795 58.245 193.295 ;
        RECT 58.445 192.725 58.615 193.075 ;
        RECT 58.790 192.895 59.120 193.295 ;
        RECT 59.290 192.725 59.460 193.075 ;
        RECT 59.630 192.895 60.010 193.295 ;
        RECT 58.445 192.555 60.030 192.725 ;
        RECT 60.200 192.620 60.475 192.965 ;
        RECT 59.860 192.385 60.030 192.555 ;
        RECT 57.475 192.055 58.130 192.385 ;
        RECT 56.455 190.915 56.795 191.175 ;
        RECT 56.965 190.745 57.305 191.820 ;
        RECT 57.475 191.460 57.715 192.055 ;
        RECT 57.910 191.595 58.230 191.885 ;
        RECT 58.400 191.765 59.140 192.385 ;
        RECT 59.310 192.055 59.690 192.385 ;
        RECT 59.860 192.055 60.135 192.385 ;
        RECT 59.860 191.885 60.030 192.055 ;
        RECT 60.305 191.885 60.475 192.620 ;
        RECT 59.370 191.715 60.030 191.885 ;
        RECT 59.370 191.595 59.540 191.715 ;
        RECT 57.910 191.425 59.540 191.595 ;
        RECT 57.485 191.085 59.540 191.255 ;
        RECT 57.490 190.965 59.540 191.085 ;
        RECT 59.710 190.745 59.990 191.545 ;
        RECT 60.200 190.915 60.475 191.885 ;
        RECT 60.645 192.350 60.985 193.125 ;
        RECT 61.155 192.835 61.325 193.295 ;
        RECT 61.565 192.860 61.925 193.125 ;
        RECT 61.565 192.855 61.920 192.860 ;
        RECT 61.565 192.845 61.915 192.855 ;
        RECT 61.565 192.840 61.910 192.845 ;
        RECT 61.565 192.830 61.905 192.840 ;
        RECT 62.555 192.835 62.725 193.295 ;
        RECT 61.565 192.825 61.900 192.830 ;
        RECT 61.565 192.815 61.890 192.825 ;
        RECT 61.565 192.805 61.880 192.815 ;
        RECT 61.565 192.665 61.865 192.805 ;
        RECT 61.155 192.475 61.865 192.665 ;
        RECT 62.055 192.665 62.385 192.745 ;
        RECT 62.895 192.665 63.235 193.125 ;
        RECT 62.055 192.475 63.235 192.665 ;
        RECT 63.465 192.475 63.675 193.295 ;
        RECT 63.845 192.495 64.175 193.125 ;
        RECT 60.645 190.915 60.925 192.350 ;
        RECT 61.155 191.905 61.440 192.475 ;
        RECT 61.625 192.075 62.095 192.305 ;
        RECT 62.265 192.285 62.595 192.305 ;
        RECT 62.265 192.105 62.715 192.285 ;
        RECT 62.905 192.105 63.235 192.305 ;
        RECT 61.155 191.690 62.305 191.905 ;
        RECT 61.095 190.745 61.805 191.520 ;
        RECT 61.975 190.915 62.305 191.690 ;
        RECT 62.500 190.990 62.715 192.105 ;
        RECT 63.005 191.765 63.235 192.105 ;
        RECT 63.845 191.895 64.095 192.495 ;
        RECT 64.345 192.475 64.575 193.295 ;
        RECT 64.785 192.525 68.295 193.295 ;
        RECT 68.925 192.570 69.215 193.295 ;
        RECT 69.845 192.555 70.230 193.125 ;
        RECT 70.400 192.835 70.725 193.295 ;
        RECT 71.245 192.665 71.525 193.125 ;
        RECT 64.265 192.055 64.595 192.305 ;
        RECT 64.785 192.005 66.435 192.525 ;
        RECT 62.895 190.745 63.225 191.465 ;
        RECT 63.465 190.745 63.675 191.885 ;
        RECT 63.845 190.915 64.175 191.895 ;
        RECT 64.345 190.745 64.575 191.885 ;
        RECT 66.605 191.835 68.295 192.355 ;
        RECT 64.785 190.745 68.295 191.835 ;
        RECT 68.925 190.745 69.215 191.910 ;
        RECT 69.845 191.885 70.125 192.555 ;
        RECT 70.400 192.495 71.525 192.665 ;
        RECT 70.400 192.385 70.850 192.495 ;
        RECT 70.295 192.055 70.850 192.385 ;
        RECT 71.715 192.325 72.115 193.125 ;
        RECT 72.515 192.835 72.785 193.295 ;
        RECT 72.955 192.665 73.240 193.125 ;
        RECT 69.845 190.915 70.230 191.885 ;
        RECT 70.400 191.595 70.850 192.055 ;
        RECT 71.020 191.765 72.115 192.325 ;
        RECT 70.400 191.375 71.525 191.595 ;
        RECT 70.400 190.745 70.725 191.205 ;
        RECT 71.245 190.915 71.525 191.375 ;
        RECT 71.715 190.915 72.115 191.765 ;
        RECT 72.285 192.495 73.240 192.665 ;
        RECT 73.525 192.835 74.085 193.125 ;
        RECT 74.255 192.835 74.505 193.295 ;
        RECT 72.285 191.595 72.495 192.495 ;
        RECT 72.665 191.765 73.355 192.325 ;
        RECT 72.285 191.375 73.240 191.595 ;
        RECT 72.515 190.745 72.785 191.205 ;
        RECT 72.955 190.915 73.240 191.375 ;
        RECT 73.525 191.465 73.775 192.835 ;
        RECT 75.125 192.665 75.455 193.025 ;
        RECT 76.530 192.815 76.830 193.295 ;
        RECT 74.065 192.475 75.455 192.665 ;
        RECT 77.000 192.645 77.260 193.100 ;
        RECT 77.430 192.815 77.690 193.295 ;
        RECT 77.860 192.645 78.120 193.100 ;
        RECT 78.290 192.815 78.550 193.295 ;
        RECT 78.720 192.645 78.980 193.100 ;
        RECT 79.150 192.815 79.410 193.295 ;
        RECT 79.580 192.645 79.840 193.100 ;
        RECT 80.010 192.770 80.270 193.295 ;
        RECT 76.530 192.475 79.840 192.645 ;
        RECT 74.065 192.385 74.235 192.475 ;
        RECT 73.945 192.055 74.235 192.385 ;
        RECT 74.405 192.055 74.745 192.305 ;
        RECT 74.965 192.055 75.640 192.305 ;
        RECT 74.065 191.805 74.235 192.055 ;
        RECT 74.065 191.635 75.005 191.805 ;
        RECT 75.375 191.695 75.640 192.055 ;
        RECT 76.530 191.885 77.500 192.475 ;
        RECT 80.440 192.305 80.690 193.115 ;
        RECT 80.870 192.835 81.115 193.295 ;
        RECT 77.670 192.055 80.690 192.305 ;
        RECT 80.860 192.055 81.175 192.665 ;
        RECT 81.405 192.475 81.615 193.295 ;
        RECT 81.785 192.495 82.115 193.125 ;
        RECT 76.530 191.645 79.840 191.885 ;
        RECT 73.525 190.915 73.985 191.465 ;
        RECT 74.175 190.745 74.505 191.465 ;
        RECT 74.705 191.085 75.005 191.635 ;
        RECT 75.175 190.745 75.455 191.415 ;
        RECT 76.535 190.745 76.830 191.475 ;
        RECT 77.000 190.920 77.260 191.645 ;
        RECT 77.430 190.745 77.690 191.475 ;
        RECT 77.860 190.920 78.120 191.645 ;
        RECT 78.290 190.745 78.550 191.475 ;
        RECT 78.720 190.920 78.980 191.645 ;
        RECT 79.150 190.745 79.410 191.475 ;
        RECT 79.580 190.920 79.840 191.645 ;
        RECT 80.010 190.745 80.270 191.855 ;
        RECT 80.440 190.920 80.690 192.055 ;
        RECT 81.785 191.895 82.035 192.495 ;
        RECT 82.285 192.475 82.515 193.295 ;
        RECT 82.840 192.665 83.125 193.125 ;
        RECT 83.295 192.835 83.565 193.295 ;
        RECT 82.840 192.495 83.795 192.665 ;
        RECT 82.205 192.055 82.535 192.305 ;
        RECT 80.870 190.745 81.165 191.855 ;
        RECT 81.405 190.745 81.615 191.885 ;
        RECT 81.785 190.915 82.115 191.895 ;
        RECT 82.285 190.745 82.515 191.885 ;
        RECT 82.725 191.765 83.415 192.325 ;
        RECT 83.585 191.595 83.795 192.495 ;
        RECT 82.840 191.375 83.795 191.595 ;
        RECT 83.965 192.325 84.365 193.125 ;
        RECT 84.555 192.665 84.835 193.125 ;
        RECT 85.355 192.835 85.680 193.295 ;
        RECT 84.555 192.495 85.680 192.665 ;
        RECT 85.850 192.555 86.235 193.125 ;
        RECT 87.415 192.745 87.585 193.035 ;
        RECT 87.755 192.915 88.085 193.295 ;
        RECT 87.415 192.575 88.080 192.745 ;
        RECT 85.230 192.385 85.680 192.495 ;
        RECT 83.965 191.765 85.060 192.325 ;
        RECT 85.230 192.055 85.785 192.385 ;
        RECT 82.840 190.915 83.125 191.375 ;
        RECT 83.295 190.745 83.565 191.205 ;
        RECT 83.965 190.915 84.365 191.765 ;
        RECT 85.230 191.595 85.680 192.055 ;
        RECT 85.955 191.885 86.235 192.555 ;
        RECT 84.555 191.375 85.680 191.595 ;
        RECT 84.555 190.915 84.835 191.375 ;
        RECT 85.355 190.745 85.680 191.205 ;
        RECT 85.850 190.915 86.235 191.885 ;
        RECT 87.330 191.755 87.680 192.405 ;
        RECT 87.850 191.585 88.080 192.575 ;
        RECT 87.415 191.415 88.080 191.585 ;
        RECT 87.415 190.915 87.585 191.415 ;
        RECT 87.755 190.745 88.085 191.245 ;
        RECT 88.255 190.915 88.440 193.035 ;
        RECT 88.695 192.835 88.945 193.295 ;
        RECT 89.115 192.845 89.450 193.015 ;
        RECT 89.645 192.845 90.320 193.015 ;
        RECT 89.115 192.705 89.285 192.845 ;
        RECT 88.610 191.715 88.890 192.665 ;
        RECT 89.060 192.575 89.285 192.705 ;
        RECT 89.060 191.470 89.230 192.575 ;
        RECT 89.455 192.425 89.980 192.645 ;
        RECT 89.400 191.660 89.640 192.255 ;
        RECT 89.810 191.725 89.980 192.425 ;
        RECT 90.150 192.065 90.320 192.845 ;
        RECT 90.640 192.795 91.010 193.295 ;
        RECT 91.190 192.845 91.595 193.015 ;
        RECT 91.765 192.845 92.550 193.015 ;
        RECT 91.190 192.615 91.360 192.845 ;
        RECT 90.530 192.315 91.360 192.615 ;
        RECT 91.745 192.345 92.210 192.675 ;
        RECT 90.530 192.285 90.730 192.315 ;
        RECT 90.850 192.065 91.020 192.135 ;
        RECT 90.150 191.895 91.020 192.065 ;
        RECT 90.510 191.805 91.020 191.895 ;
        RECT 89.060 191.340 89.365 191.470 ;
        RECT 89.810 191.360 90.340 191.725 ;
        RECT 88.680 190.745 88.945 191.205 ;
        RECT 89.115 190.915 89.365 191.340 ;
        RECT 90.510 191.190 90.680 191.805 ;
        RECT 89.575 191.020 90.680 191.190 ;
        RECT 90.850 190.745 91.020 191.545 ;
        RECT 91.190 191.245 91.360 192.315 ;
        RECT 91.530 191.415 91.720 192.135 ;
        RECT 91.890 191.385 92.210 192.345 ;
        RECT 92.380 192.385 92.550 192.845 ;
        RECT 92.825 192.765 93.035 193.295 ;
        RECT 93.295 192.555 93.625 193.080 ;
        RECT 93.795 192.685 93.965 193.295 ;
        RECT 94.135 192.640 94.465 193.075 ;
        RECT 94.135 192.555 94.515 192.640 ;
        RECT 94.685 192.570 94.975 193.295 ;
        RECT 93.425 192.385 93.625 192.555 ;
        RECT 94.290 192.515 94.515 192.555 ;
        RECT 92.380 192.055 93.255 192.385 ;
        RECT 93.425 192.055 94.175 192.385 ;
        RECT 91.190 190.915 91.440 191.245 ;
        RECT 92.380 191.215 92.550 192.055 ;
        RECT 93.425 191.850 93.615 192.055 ;
        RECT 94.345 191.935 94.515 192.515 ;
        RECT 94.300 191.885 94.515 191.935 ;
        RECT 95.150 192.555 95.405 193.125 ;
        RECT 95.575 192.895 95.905 193.295 ;
        RECT 96.330 192.760 96.860 193.125 ;
        RECT 96.330 192.725 96.505 192.760 ;
        RECT 95.575 192.555 96.505 192.725 ;
        RECT 97.050 192.615 97.325 193.125 ;
        RECT 92.720 191.475 93.615 191.850 ;
        RECT 94.125 191.805 94.515 191.885 ;
        RECT 91.665 191.045 92.550 191.215 ;
        RECT 92.730 190.745 93.045 191.245 ;
        RECT 93.275 190.915 93.615 191.475 ;
        RECT 93.785 190.745 93.955 191.755 ;
        RECT 94.125 190.960 94.455 191.805 ;
        RECT 94.685 190.745 94.975 191.910 ;
        RECT 95.150 191.885 95.320 192.555 ;
        RECT 95.575 192.385 95.745 192.555 ;
        RECT 95.490 192.055 95.745 192.385 ;
        RECT 95.970 192.055 96.165 192.385 ;
        RECT 95.150 190.915 95.485 191.885 ;
        RECT 95.655 190.745 95.825 191.885 ;
        RECT 95.995 191.085 96.165 192.055 ;
        RECT 96.335 191.425 96.505 192.555 ;
        RECT 96.675 191.765 96.845 192.565 ;
        RECT 97.045 192.445 97.325 192.615 ;
        RECT 97.050 191.965 97.325 192.445 ;
        RECT 97.495 191.765 97.685 193.125 ;
        RECT 97.865 192.760 98.375 193.295 ;
        RECT 98.595 192.485 98.840 193.090 ;
        RECT 99.285 192.555 99.795 193.125 ;
        RECT 99.965 192.735 100.135 193.295 ;
        RECT 100.340 192.725 100.670 193.125 ;
        RECT 100.845 192.895 101.175 193.295 ;
        RECT 101.410 192.915 102.795 193.125 ;
        RECT 101.410 192.725 101.740 192.915 ;
        RECT 100.340 192.555 101.740 192.725 ;
        RECT 101.910 192.555 102.335 192.745 ;
        RECT 102.505 192.645 102.795 192.915 ;
        RECT 97.885 192.315 99.115 192.485 ;
        RECT 96.675 191.595 97.685 191.765 ;
        RECT 97.855 191.750 98.605 191.940 ;
        RECT 96.335 191.255 97.460 191.425 ;
        RECT 97.855 191.085 98.025 191.750 ;
        RECT 98.775 191.505 99.115 192.315 ;
        RECT 95.995 190.915 98.025 191.085 ;
        RECT 98.195 190.745 98.365 191.505 ;
        RECT 98.600 191.095 99.115 191.505 ;
        RECT 99.285 191.885 99.460 192.555 ;
        RECT 99.645 192.305 99.835 192.385 ;
        RECT 100.205 192.305 100.375 192.385 ;
        RECT 99.645 192.055 100.010 192.305 ;
        RECT 100.205 192.055 100.455 192.305 ;
        RECT 100.665 192.055 101.010 192.385 ;
        RECT 99.840 191.885 100.010 192.055 ;
        RECT 99.285 190.925 99.670 191.885 ;
        RECT 99.840 191.715 100.515 191.885 ;
        RECT 99.885 190.745 100.175 191.545 ;
        RECT 100.345 191.085 100.515 191.715 ;
        RECT 100.685 191.255 101.010 192.055 ;
        RECT 101.180 191.720 101.455 192.385 ;
        RECT 101.640 191.720 101.995 192.385 ;
        RECT 102.165 191.545 102.335 192.555 ;
        RECT 102.975 192.570 103.305 193.080 ;
        RECT 103.475 192.895 103.805 193.295 ;
        RECT 104.855 192.725 105.185 193.065 ;
        RECT 105.355 192.895 105.685 193.295 ;
        RECT 102.520 192.055 102.795 192.385 ;
        RECT 101.380 191.295 102.335 191.545 ;
        RECT 101.380 191.085 101.710 191.295 ;
        RECT 100.345 190.915 101.710 191.085 ;
        RECT 102.505 190.745 102.795 191.885 ;
        RECT 102.975 191.805 103.165 192.570 ;
        RECT 103.475 192.555 105.840 192.725 ;
        RECT 103.475 192.385 103.645 192.555 ;
        RECT 103.335 192.055 103.645 192.385 ;
        RECT 103.815 192.055 104.120 192.385 ;
        RECT 102.975 190.955 103.305 191.805 ;
        RECT 103.475 190.745 103.725 191.885 ;
        RECT 103.905 191.725 104.120 192.055 ;
        RECT 104.295 191.725 104.580 192.385 ;
        RECT 104.775 191.725 105.040 192.385 ;
        RECT 105.255 191.725 105.500 192.385 ;
        RECT 105.670 191.555 105.840 192.555 ;
        RECT 106.225 192.475 106.455 193.295 ;
        RECT 106.625 192.495 106.955 193.125 ;
        RECT 106.205 192.055 106.535 192.305 ;
        RECT 106.705 191.895 106.955 192.495 ;
        RECT 107.125 192.475 107.335 193.295 ;
        RECT 107.565 192.525 111.075 193.295 ;
        RECT 107.565 192.005 109.215 192.525 ;
        RECT 111.520 192.485 111.765 193.090 ;
        RECT 111.985 192.760 112.495 193.295 ;
        RECT 103.915 191.385 105.205 191.555 ;
        RECT 103.915 190.965 104.165 191.385 ;
        RECT 104.395 190.745 104.725 191.215 ;
        RECT 104.955 190.965 105.205 191.385 ;
        RECT 105.385 191.385 105.840 191.555 ;
        RECT 105.385 190.955 105.715 191.385 ;
        RECT 106.225 190.745 106.455 191.885 ;
        RECT 106.625 190.915 106.955 191.895 ;
        RECT 107.125 190.745 107.335 191.885 ;
        RECT 109.385 191.835 111.075 192.355 ;
        RECT 107.565 190.745 111.075 191.835 ;
        RECT 111.245 192.315 112.475 192.485 ;
        RECT 111.245 191.505 111.585 192.315 ;
        RECT 111.755 191.750 112.505 191.940 ;
        RECT 111.245 191.095 111.760 191.505 ;
        RECT 111.995 190.745 112.165 191.505 ;
        RECT 112.335 191.085 112.505 191.750 ;
        RECT 112.675 191.765 112.865 193.125 ;
        RECT 113.035 192.275 113.310 193.125 ;
        RECT 113.500 192.760 114.030 193.125 ;
        RECT 114.455 192.895 114.785 193.295 ;
        RECT 113.855 192.725 114.030 192.760 ;
        RECT 113.035 192.105 113.315 192.275 ;
        RECT 113.035 191.965 113.310 192.105 ;
        RECT 113.515 191.765 113.685 192.565 ;
        RECT 112.675 191.595 113.685 191.765 ;
        RECT 113.855 192.555 114.785 192.725 ;
        RECT 114.955 192.555 115.210 193.125 ;
        RECT 113.855 191.425 114.025 192.555 ;
        RECT 114.615 192.385 114.785 192.555 ;
        RECT 112.900 191.255 114.025 191.425 ;
        RECT 114.195 192.055 114.390 192.385 ;
        RECT 114.615 192.055 114.870 192.385 ;
        RECT 114.195 191.085 114.365 192.055 ;
        RECT 115.040 191.885 115.210 192.555 ;
        RECT 115.385 192.525 118.895 193.295 ;
        RECT 119.065 192.545 120.275 193.295 ;
        RECT 120.445 192.570 120.735 193.295 ;
        RECT 120.905 192.750 126.250 193.295 ;
        RECT 126.425 192.750 131.770 193.295 ;
        RECT 131.945 192.750 137.290 193.295 ;
        RECT 137.465 192.750 142.810 193.295 ;
        RECT 115.385 192.005 117.035 192.525 ;
        RECT 112.335 190.915 114.365 191.085 ;
        RECT 114.535 190.745 114.705 191.885 ;
        RECT 114.875 190.915 115.210 191.885 ;
        RECT 117.205 191.835 118.895 192.355 ;
        RECT 119.065 192.005 119.585 192.545 ;
        RECT 119.755 191.835 120.275 192.375 ;
        RECT 122.490 191.920 122.830 192.750 ;
        RECT 115.385 190.745 118.895 191.835 ;
        RECT 119.065 190.745 120.275 191.835 ;
        RECT 120.445 190.745 120.735 191.910 ;
        RECT 124.310 191.180 124.660 192.430 ;
        RECT 128.010 191.920 128.350 192.750 ;
        RECT 129.830 191.180 130.180 192.430 ;
        RECT 133.530 191.920 133.870 192.750 ;
        RECT 135.350 191.180 135.700 192.430 ;
        RECT 139.050 191.920 139.390 192.750 ;
        RECT 142.985 192.525 145.575 193.295 ;
        RECT 145.745 192.545 146.955 193.295 ;
        RECT 140.870 191.180 141.220 192.430 ;
        RECT 142.985 192.005 144.195 192.525 ;
        RECT 144.365 191.835 145.575 192.355 ;
        RECT 120.905 190.745 126.250 191.180 ;
        RECT 126.425 190.745 131.770 191.180 ;
        RECT 131.945 190.745 137.290 191.180 ;
        RECT 137.465 190.745 142.810 191.180 ;
        RECT 142.985 190.745 145.575 191.835 ;
        RECT 145.745 191.835 146.265 192.375 ;
        RECT 146.435 192.005 146.955 192.545 ;
        RECT 145.745 190.745 146.955 191.835 ;
        RECT 17.320 190.575 147.040 190.745 ;
        RECT 17.405 189.485 18.615 190.575 ;
        RECT 18.785 189.485 21.375 190.575 ;
        RECT 21.635 189.905 21.805 190.405 ;
        RECT 21.975 190.075 22.305 190.575 ;
        RECT 21.635 189.735 22.300 189.905 ;
        RECT 17.405 188.775 17.925 189.315 ;
        RECT 18.095 188.945 18.615 189.485 ;
        RECT 18.785 188.795 19.995 189.315 ;
        RECT 20.165 188.965 21.375 189.485 ;
        RECT 21.550 188.915 21.900 189.565 ;
        RECT 17.405 188.025 18.615 188.775 ;
        RECT 18.785 188.025 21.375 188.795 ;
        RECT 22.070 188.745 22.300 189.735 ;
        RECT 21.635 188.575 22.300 188.745 ;
        RECT 21.635 188.285 21.805 188.575 ;
        RECT 21.975 188.025 22.305 188.405 ;
        RECT 22.475 188.285 22.660 190.405 ;
        RECT 22.900 190.115 23.165 190.575 ;
        RECT 23.335 189.980 23.585 190.405 ;
        RECT 23.795 190.130 24.900 190.300 ;
        RECT 23.280 189.850 23.585 189.980 ;
        RECT 22.830 188.655 23.110 189.605 ;
        RECT 23.280 188.745 23.450 189.850 ;
        RECT 23.620 189.065 23.860 189.660 ;
        RECT 24.030 189.595 24.560 189.960 ;
        RECT 24.030 188.895 24.200 189.595 ;
        RECT 24.730 189.515 24.900 190.130 ;
        RECT 25.070 189.775 25.240 190.575 ;
        RECT 25.410 190.075 25.660 190.405 ;
        RECT 25.885 190.105 26.770 190.275 ;
        RECT 24.730 189.425 25.240 189.515 ;
        RECT 23.280 188.615 23.505 188.745 ;
        RECT 23.675 188.675 24.200 188.895 ;
        RECT 24.370 189.255 25.240 189.425 ;
        RECT 22.915 188.025 23.165 188.485 ;
        RECT 23.335 188.475 23.505 188.615 ;
        RECT 24.370 188.475 24.540 189.255 ;
        RECT 25.070 189.185 25.240 189.255 ;
        RECT 24.750 189.005 24.950 189.035 ;
        RECT 25.410 189.005 25.580 190.075 ;
        RECT 25.750 189.185 25.940 189.905 ;
        RECT 24.750 188.705 25.580 189.005 ;
        RECT 26.110 188.975 26.430 189.935 ;
        RECT 23.335 188.305 23.670 188.475 ;
        RECT 23.865 188.305 24.540 188.475 ;
        RECT 24.860 188.025 25.230 188.525 ;
        RECT 25.410 188.475 25.580 188.705 ;
        RECT 25.965 188.645 26.430 188.975 ;
        RECT 26.600 189.265 26.770 190.105 ;
        RECT 26.950 190.075 27.265 190.575 ;
        RECT 27.495 189.845 27.835 190.405 ;
        RECT 26.940 189.470 27.835 189.845 ;
        RECT 28.005 189.565 28.175 190.575 ;
        RECT 27.645 189.265 27.835 189.470 ;
        RECT 28.345 189.515 28.675 190.360 ;
        RECT 28.345 189.435 28.735 189.515 ;
        RECT 28.905 189.435 29.185 190.575 ;
        RECT 28.520 189.385 28.735 189.435 ;
        RECT 29.355 189.425 29.685 190.405 ;
        RECT 29.855 189.435 30.115 190.575 ;
        RECT 26.600 188.935 27.475 189.265 ;
        RECT 27.645 188.935 28.395 189.265 ;
        RECT 26.600 188.475 26.770 188.935 ;
        RECT 27.645 188.765 27.845 188.935 ;
        RECT 28.565 188.805 28.735 189.385 ;
        RECT 28.915 188.995 29.250 189.265 ;
        RECT 29.420 188.825 29.590 189.425 ;
        RECT 30.285 189.410 30.575 190.575 ;
        RECT 29.760 189.015 30.095 189.265 ;
        RECT 28.510 188.765 28.735 188.805 ;
        RECT 25.410 188.305 25.815 188.475 ;
        RECT 25.985 188.305 26.770 188.475 ;
        RECT 27.045 188.025 27.255 188.555 ;
        RECT 27.515 188.240 27.845 188.765 ;
        RECT 28.355 188.680 28.735 188.765 ;
        RECT 28.015 188.025 28.185 188.635 ;
        RECT 28.355 188.245 28.685 188.680 ;
        RECT 28.905 188.025 29.215 188.825 ;
        RECT 29.420 188.195 30.115 188.825 ;
        RECT 30.285 188.025 30.575 188.750 ;
        RECT 30.755 188.205 31.015 190.395 ;
        RECT 31.185 189.845 31.525 190.575 ;
        RECT 31.705 189.665 31.975 190.395 ;
        RECT 31.205 189.445 31.975 189.665 ;
        RECT 32.155 189.685 32.385 190.395 ;
        RECT 32.555 189.865 32.885 190.575 ;
        RECT 33.055 189.685 33.315 190.395 ;
        RECT 32.155 189.445 33.315 189.685 ;
        RECT 33.690 189.605 34.080 189.780 ;
        RECT 34.565 189.775 34.895 190.575 ;
        RECT 35.065 189.785 35.600 190.405 ;
        RECT 31.205 188.775 31.495 189.445 ;
        RECT 33.690 189.435 35.115 189.605 ;
        RECT 31.675 188.955 32.140 189.265 ;
        RECT 32.320 188.955 32.845 189.265 ;
        RECT 31.205 188.575 32.435 188.775 ;
        RECT 31.275 188.025 31.945 188.395 ;
        RECT 32.125 188.205 32.435 188.575 ;
        RECT 32.615 188.315 32.845 188.955 ;
        RECT 33.025 188.935 33.325 189.265 ;
        RECT 33.025 188.025 33.315 188.755 ;
        RECT 33.565 188.705 33.920 189.265 ;
        RECT 34.090 188.535 34.260 189.435 ;
        RECT 34.430 188.705 34.695 189.265 ;
        RECT 34.945 188.935 35.115 189.435 ;
        RECT 35.285 188.765 35.600 189.785 ;
        RECT 33.670 188.025 33.910 188.535 ;
        RECT 34.090 188.205 34.370 188.535 ;
        RECT 34.600 188.025 34.815 188.535 ;
        RECT 34.985 188.195 35.600 188.765 ;
        RECT 35.805 189.705 36.080 190.405 ;
        RECT 36.250 190.030 36.505 190.575 ;
        RECT 36.675 190.065 37.155 190.405 ;
        RECT 37.330 190.020 37.935 190.575 ;
        RECT 37.320 189.920 37.935 190.020 ;
        RECT 37.320 189.895 37.505 189.920 ;
        RECT 35.805 188.675 35.975 189.705 ;
        RECT 36.250 189.575 37.005 189.825 ;
        RECT 37.175 189.650 37.505 189.895 ;
        RECT 36.250 189.540 37.020 189.575 ;
        RECT 36.250 189.530 37.035 189.540 ;
        RECT 36.145 189.515 37.040 189.530 ;
        RECT 36.145 189.500 37.060 189.515 ;
        RECT 36.145 189.490 37.080 189.500 ;
        RECT 36.145 189.480 37.105 189.490 ;
        RECT 36.145 189.450 37.175 189.480 ;
        RECT 36.145 189.420 37.195 189.450 ;
        RECT 36.145 189.390 37.215 189.420 ;
        RECT 36.145 189.365 37.245 189.390 ;
        RECT 36.145 189.330 37.280 189.365 ;
        RECT 36.145 189.325 37.310 189.330 ;
        RECT 36.145 188.930 36.375 189.325 ;
        RECT 36.920 189.320 37.310 189.325 ;
        RECT 36.945 189.310 37.310 189.320 ;
        RECT 36.960 189.305 37.310 189.310 ;
        RECT 36.975 189.300 37.310 189.305 ;
        RECT 37.675 189.300 37.935 189.750 ;
        RECT 39.035 189.595 39.365 190.405 ;
        RECT 39.535 189.775 39.775 190.575 ;
        RECT 39.035 189.425 39.750 189.595 ;
        RECT 36.975 189.295 37.935 189.300 ;
        RECT 36.985 189.285 37.935 189.295 ;
        RECT 36.995 189.280 37.935 189.285 ;
        RECT 37.005 189.270 37.935 189.280 ;
        RECT 37.010 189.260 37.935 189.270 ;
        RECT 37.015 189.255 37.935 189.260 ;
        RECT 37.025 189.240 37.935 189.255 ;
        RECT 37.030 189.225 37.935 189.240 ;
        RECT 37.040 189.200 37.935 189.225 ;
        RECT 36.545 188.730 36.875 189.155 ;
        RECT 36.625 188.705 36.875 188.730 ;
        RECT 35.805 188.195 36.065 188.675 ;
        RECT 36.235 188.025 36.485 188.565 ;
        RECT 36.655 188.245 36.875 188.705 ;
        RECT 37.045 189.130 37.935 189.200 ;
        RECT 37.045 188.405 37.215 189.130 ;
        RECT 39.030 189.015 39.410 189.255 ;
        RECT 39.580 189.185 39.750 189.425 ;
        RECT 39.955 189.555 40.125 190.405 ;
        RECT 40.295 189.775 40.625 190.575 ;
        RECT 40.795 189.555 40.965 190.405 ;
        RECT 39.955 189.385 40.965 189.555 ;
        RECT 41.135 189.425 41.465 190.575 ;
        RECT 42.270 189.605 42.570 189.800 ;
        RECT 42.740 189.775 42.995 190.575 ;
        RECT 43.195 189.945 43.525 190.405 ;
        RECT 43.695 190.115 44.270 190.575 ;
        RECT 44.440 189.945 44.795 190.405 ;
        RECT 43.195 189.775 44.795 189.945 ;
        RECT 42.270 189.435 43.520 189.605 ;
        RECT 40.470 189.215 40.965 189.385 ;
        RECT 39.580 189.015 40.080 189.185 ;
        RECT 40.465 189.045 40.965 189.215 ;
        RECT 37.385 188.575 37.935 188.960 ;
        RECT 39.580 188.845 39.750 189.015 ;
        RECT 40.470 188.845 40.965 189.045 ;
        RECT 39.115 188.675 39.750 188.845 ;
        RECT 39.955 188.675 40.965 188.845 ;
        RECT 37.045 188.235 37.935 188.405 ;
        RECT 39.115 188.195 39.285 188.675 ;
        RECT 39.465 188.025 39.705 188.505 ;
        RECT 39.955 188.195 40.125 188.675 ;
        RECT 40.295 188.025 40.625 188.505 ;
        RECT 40.795 188.195 40.965 188.675 ;
        RECT 41.135 188.025 41.465 188.825 ;
        RECT 42.270 188.780 42.440 189.435 ;
        RECT 42.615 188.935 42.960 189.265 ;
        RECT 43.190 189.015 43.520 189.435 ;
        RECT 43.690 188.845 43.970 189.775 ;
        RECT 44.150 189.555 44.340 189.595 ;
        RECT 44.145 189.385 44.340 189.555 ;
        RECT 44.520 189.435 44.795 189.775 ;
        RECT 44.965 189.435 45.295 190.575 ;
        RECT 45.650 189.605 46.040 189.780 ;
        RECT 46.525 189.775 46.855 190.575 ;
        RECT 47.025 189.785 47.560 190.405 ;
        RECT 45.650 189.435 47.075 189.605 ;
        RECT 44.605 189.385 44.775 189.435 ;
        RECT 44.150 189.215 44.340 189.385 ;
        RECT 44.150 189.015 45.295 189.215 ;
        RECT 42.270 188.450 42.505 188.780 ;
        RECT 42.675 188.025 43.005 188.765 ;
        RECT 43.240 188.405 43.515 188.845 ;
        RECT 43.690 188.745 44.015 188.845 ;
        RECT 43.685 188.575 44.015 188.745 ;
        RECT 44.185 188.635 45.295 188.845 ;
        RECT 45.525 188.705 45.880 189.265 ;
        RECT 44.185 188.405 44.435 188.635 ;
        RECT 43.240 188.195 44.435 188.405 ;
        RECT 44.605 188.025 44.775 188.465 ;
        RECT 44.945 188.195 45.295 188.635 ;
        RECT 46.050 188.535 46.220 189.435 ;
        RECT 46.390 188.705 46.655 189.265 ;
        RECT 46.905 188.935 47.075 189.435 ;
        RECT 47.245 188.765 47.560 189.785 ;
        RECT 48.695 189.625 48.970 190.395 ;
        RECT 49.140 189.965 49.470 190.395 ;
        RECT 49.640 190.135 49.835 190.575 ;
        RECT 50.015 189.965 50.345 190.395 ;
        RECT 49.140 189.795 50.345 189.965 ;
        RECT 50.725 189.905 51.005 190.575 ;
        RECT 48.695 189.435 49.280 189.625 ;
        RECT 49.450 189.465 50.345 189.795 ;
        RECT 51.175 189.685 51.475 190.235 ;
        RECT 51.675 189.855 52.005 190.575 ;
        RECT 52.195 189.855 52.655 190.405 ;
        RECT 53.125 189.935 53.455 190.365 ;
        RECT 45.630 188.025 45.870 188.535 ;
        RECT 46.050 188.205 46.330 188.535 ;
        RECT 46.560 188.025 46.775 188.535 ;
        RECT 46.945 188.195 47.560 188.765 ;
        RECT 48.695 188.615 48.935 189.265 ;
        RECT 49.105 188.765 49.280 189.435 ;
        RECT 50.540 189.265 50.805 189.625 ;
        RECT 51.175 189.515 52.115 189.685 ;
        RECT 51.945 189.265 52.115 189.515 ;
        RECT 49.450 188.935 49.865 189.265 ;
        RECT 50.045 188.935 50.340 189.265 ;
        RECT 50.540 189.015 51.215 189.265 ;
        RECT 51.435 189.015 51.775 189.265 ;
        RECT 51.945 188.935 52.235 189.265 ;
        RECT 49.105 188.585 49.435 188.765 ;
        RECT 48.710 188.025 49.040 188.415 ;
        RECT 49.210 188.205 49.435 188.585 ;
        RECT 49.635 188.315 49.865 188.935 ;
        RECT 51.945 188.845 52.115 188.935 ;
        RECT 50.045 188.025 50.345 188.755 ;
        RECT 50.725 188.655 52.115 188.845 ;
        RECT 50.725 188.295 51.055 188.655 ;
        RECT 52.405 188.485 52.655 189.855 ;
        RECT 53.000 189.765 53.455 189.935 ;
        RECT 53.635 189.935 53.885 190.355 ;
        RECT 54.115 190.105 54.445 190.575 ;
        RECT 54.675 189.935 54.925 190.355 ;
        RECT 53.635 189.765 54.925 189.935 ;
        RECT 53.000 188.765 53.170 189.765 ;
        RECT 53.340 188.935 53.585 189.595 ;
        RECT 53.800 188.935 54.065 189.595 ;
        RECT 54.260 188.935 54.545 189.595 ;
        RECT 54.720 189.265 54.935 189.595 ;
        RECT 55.115 189.435 55.365 190.575 ;
        RECT 55.535 189.515 55.865 190.365 ;
        RECT 54.720 188.935 55.025 189.265 ;
        RECT 55.195 188.935 55.505 189.265 ;
        RECT 55.195 188.765 55.365 188.935 ;
        RECT 53.000 188.595 55.365 188.765 ;
        RECT 55.675 188.750 55.865 189.515 ;
        RECT 56.045 189.410 56.335 190.575 ;
        RECT 56.565 189.435 56.775 190.575 ;
        RECT 56.945 189.425 57.275 190.405 ;
        RECT 57.445 189.435 57.675 190.575 ;
        RECT 57.885 190.075 58.145 190.405 ;
        RECT 58.455 190.195 58.785 190.575 ;
        RECT 51.675 188.025 51.925 188.485 ;
        RECT 52.095 188.195 52.655 188.485 ;
        RECT 53.155 188.025 53.485 188.425 ;
        RECT 53.655 188.255 53.985 188.595 ;
        RECT 55.035 188.025 55.365 188.425 ;
        RECT 55.535 188.240 55.865 188.750 ;
        RECT 56.045 188.025 56.335 188.750 ;
        RECT 56.565 188.025 56.775 188.845 ;
        RECT 56.945 188.825 57.195 189.425 ;
        RECT 57.885 189.395 58.055 190.075 ;
        RECT 59.025 190.025 59.215 190.405 ;
        RECT 59.465 190.195 59.795 190.575 ;
        RECT 60.005 190.025 60.175 190.405 ;
        RECT 60.370 190.195 60.700 190.575 ;
        RECT 60.960 190.025 61.130 190.405 ;
        RECT 61.555 190.195 61.885 190.575 ;
        RECT 58.225 189.565 58.575 189.895 ;
        RECT 59.025 189.855 59.765 190.025 ;
        RECT 58.845 189.515 59.425 189.685 ;
        RECT 58.845 189.395 59.015 189.515 ;
        RECT 57.365 189.015 57.695 189.265 ;
        RECT 57.885 189.225 59.015 189.395 ;
        RECT 59.595 189.345 59.765 189.855 ;
        RECT 56.945 188.195 57.275 188.825 ;
        RECT 57.445 188.025 57.675 188.845 ;
        RECT 57.885 188.525 58.055 189.225 ;
        RECT 59.195 189.175 59.765 189.345 ;
        RECT 59.935 189.855 61.885 190.025 ;
        RECT 58.405 188.885 59.025 189.055 ;
        RECT 58.405 188.705 58.615 188.885 ;
        RECT 59.195 188.695 59.365 189.175 ;
        RECT 59.935 188.865 60.105 189.855 ;
        RECT 60.695 189.265 60.880 189.575 ;
        RECT 61.150 189.265 61.345 189.575 ;
        RECT 57.885 188.195 58.145 188.525 ;
        RECT 58.455 188.025 58.785 188.405 ;
        RECT 58.965 188.365 59.365 188.695 ;
        RECT 59.555 188.535 60.105 188.865 ;
        RECT 60.275 188.365 60.445 189.265 ;
        RECT 58.965 188.195 60.445 188.365 ;
        RECT 60.695 188.935 60.925 189.265 ;
        RECT 61.150 188.935 61.405 189.265 ;
        RECT 61.715 188.935 61.885 189.855 ;
        RECT 60.695 188.355 60.880 188.935 ;
        RECT 61.150 188.360 61.345 188.935 ;
        RECT 61.555 188.025 61.885 188.405 ;
        RECT 62.055 188.195 62.315 190.405 ;
        RECT 62.485 189.435 62.760 190.405 ;
        RECT 62.970 189.775 63.250 190.575 ;
        RECT 63.420 190.065 65.035 190.395 ;
        RECT 63.420 189.725 64.595 189.895 ;
        RECT 63.420 189.605 63.590 189.725 ;
        RECT 62.930 189.435 63.590 189.605 ;
        RECT 62.485 188.700 62.655 189.435 ;
        RECT 62.930 189.265 63.100 189.435 ;
        RECT 63.850 189.265 64.095 189.555 ;
        RECT 64.265 189.435 64.595 189.725 ;
        RECT 64.855 189.265 65.025 189.825 ;
        RECT 65.275 189.435 65.535 190.575 ;
        RECT 65.710 189.435 66.030 190.575 ;
        RECT 66.210 189.265 66.405 190.315 ;
        RECT 66.585 189.725 66.915 190.405 ;
        RECT 67.115 189.775 67.370 190.575 ;
        RECT 66.585 189.445 66.935 189.725 ;
        RECT 62.825 188.935 63.100 189.265 ;
        RECT 63.270 188.935 64.095 189.265 ;
        RECT 64.310 188.935 65.025 189.265 ;
        RECT 65.195 189.015 65.530 189.265 ;
        RECT 65.770 189.215 66.030 189.265 ;
        RECT 65.765 189.045 66.030 189.215 ;
        RECT 65.770 188.935 66.030 189.045 ;
        RECT 66.210 188.935 66.595 189.265 ;
        RECT 66.765 189.065 66.935 189.445 ;
        RECT 67.125 189.235 67.370 189.595 ;
        RECT 67.545 189.485 68.755 190.575 ;
        RECT 62.930 188.765 63.100 188.935 ;
        RECT 64.775 188.845 65.025 188.935 ;
        RECT 66.765 188.895 67.285 189.065 ;
        RECT 62.485 188.355 62.760 188.700 ;
        RECT 62.930 188.595 64.595 188.765 ;
        RECT 62.950 188.025 63.325 188.425 ;
        RECT 63.495 188.245 63.665 188.595 ;
        RECT 63.835 188.025 64.165 188.425 ;
        RECT 64.335 188.195 64.595 188.595 ;
        RECT 64.775 188.425 65.105 188.845 ;
        RECT 65.275 188.025 65.535 188.845 ;
        RECT 65.710 188.555 66.925 188.725 ;
        RECT 65.710 188.205 66.000 188.555 ;
        RECT 66.195 188.025 66.525 188.385 ;
        RECT 66.695 188.250 66.925 188.555 ;
        RECT 67.115 188.330 67.285 188.895 ;
        RECT 67.545 188.775 68.065 189.315 ;
        RECT 68.235 188.945 68.755 189.485 ;
        RECT 68.935 189.605 69.265 190.390 ;
        RECT 68.935 189.435 69.615 189.605 ;
        RECT 69.795 189.435 70.125 190.575 ;
        RECT 70.395 189.905 70.565 190.405 ;
        RECT 70.735 190.075 71.065 190.575 ;
        RECT 70.395 189.735 71.060 189.905 ;
        RECT 68.925 189.015 69.275 189.265 ;
        RECT 69.445 188.835 69.615 189.435 ;
        RECT 69.785 189.015 70.135 189.265 ;
        RECT 70.310 188.915 70.660 189.565 ;
        RECT 67.545 188.025 68.755 188.775 ;
        RECT 68.945 188.025 69.185 188.835 ;
        RECT 69.355 188.195 69.685 188.835 ;
        RECT 69.855 188.025 70.125 188.835 ;
        RECT 70.830 188.745 71.060 189.735 ;
        RECT 70.395 188.575 71.060 188.745 ;
        RECT 70.395 188.285 70.565 188.575 ;
        RECT 70.735 188.025 71.065 188.405 ;
        RECT 71.235 188.285 71.420 190.405 ;
        RECT 71.660 190.115 71.925 190.575 ;
        RECT 72.095 189.980 72.345 190.405 ;
        RECT 72.555 190.130 73.660 190.300 ;
        RECT 72.040 189.850 72.345 189.980 ;
        RECT 71.590 188.655 71.870 189.605 ;
        RECT 72.040 188.745 72.210 189.850 ;
        RECT 72.380 189.065 72.620 189.660 ;
        RECT 72.790 189.595 73.320 189.960 ;
        RECT 72.790 188.895 72.960 189.595 ;
        RECT 73.490 189.515 73.660 190.130 ;
        RECT 73.830 189.775 74.000 190.575 ;
        RECT 74.170 190.075 74.420 190.405 ;
        RECT 74.645 190.105 75.530 190.275 ;
        RECT 73.490 189.425 74.000 189.515 ;
        RECT 72.040 188.615 72.265 188.745 ;
        RECT 72.435 188.675 72.960 188.895 ;
        RECT 73.130 189.255 74.000 189.425 ;
        RECT 71.675 188.025 71.925 188.485 ;
        RECT 72.095 188.475 72.265 188.615 ;
        RECT 73.130 188.475 73.300 189.255 ;
        RECT 73.830 189.185 74.000 189.255 ;
        RECT 73.510 189.005 73.710 189.035 ;
        RECT 74.170 189.005 74.340 190.075 ;
        RECT 74.510 189.185 74.700 189.905 ;
        RECT 73.510 188.705 74.340 189.005 ;
        RECT 74.870 188.975 75.190 189.935 ;
        RECT 72.095 188.305 72.430 188.475 ;
        RECT 72.625 188.305 73.300 188.475 ;
        RECT 73.620 188.025 73.990 188.525 ;
        RECT 74.170 188.475 74.340 188.705 ;
        RECT 74.725 188.645 75.190 188.975 ;
        RECT 75.360 189.265 75.530 190.105 ;
        RECT 75.710 190.075 76.025 190.575 ;
        RECT 76.255 189.845 76.595 190.405 ;
        RECT 75.700 189.470 76.595 189.845 ;
        RECT 76.765 189.565 76.935 190.575 ;
        RECT 76.405 189.265 76.595 189.470 ;
        RECT 77.105 189.515 77.435 190.360 ;
        RECT 77.735 189.570 77.990 190.375 ;
        RECT 78.160 189.740 78.420 190.575 ;
        RECT 78.590 189.570 78.850 190.375 ;
        RECT 79.020 189.740 79.275 190.575 ;
        RECT 77.105 189.435 77.495 189.515 ;
        RECT 77.280 189.385 77.495 189.435 ;
        RECT 77.735 189.400 79.335 189.570 ;
        RECT 79.505 189.485 81.175 190.575 ;
        RECT 75.360 188.935 76.235 189.265 ;
        RECT 76.405 188.935 77.155 189.265 ;
        RECT 75.360 188.475 75.530 188.935 ;
        RECT 76.405 188.765 76.605 188.935 ;
        RECT 77.325 188.805 77.495 189.385 ;
        RECT 77.665 189.005 78.885 189.230 ;
        RECT 79.055 188.835 79.335 189.400 ;
        RECT 77.270 188.765 77.495 188.805 ;
        RECT 74.170 188.305 74.575 188.475 ;
        RECT 74.745 188.305 75.530 188.475 ;
        RECT 75.805 188.025 76.015 188.555 ;
        RECT 76.275 188.240 76.605 188.765 ;
        RECT 77.115 188.680 77.495 188.765 ;
        RECT 76.775 188.025 76.945 188.635 ;
        RECT 77.115 188.245 77.445 188.680 ;
        RECT 78.605 188.665 79.335 188.835 ;
        RECT 79.505 188.795 80.255 189.315 ;
        RECT 80.425 188.965 81.175 189.485 ;
        RECT 81.805 189.410 82.095 190.575 ;
        RECT 82.265 189.485 83.935 190.575 ;
        RECT 82.265 188.795 83.015 189.315 ;
        RECT 83.185 188.965 83.935 189.485 ;
        RECT 78.140 188.025 78.435 188.550 ;
        RECT 78.605 188.220 78.830 188.665 ;
        RECT 79.000 188.025 79.330 188.495 ;
        RECT 79.505 188.025 81.175 188.795 ;
        RECT 81.805 188.025 82.095 188.750 ;
        RECT 82.265 188.025 83.935 188.795 ;
        RECT 84.115 188.205 84.375 190.395 ;
        RECT 84.545 189.845 84.885 190.575 ;
        RECT 85.065 189.665 85.335 190.395 ;
        RECT 84.565 189.445 85.335 189.665 ;
        RECT 85.515 189.685 85.745 190.395 ;
        RECT 85.915 189.865 86.245 190.575 ;
        RECT 86.415 189.685 86.675 190.395 ;
        RECT 85.515 189.445 86.675 189.685 ;
        RECT 86.865 189.485 88.535 190.575 ;
        RECT 84.565 188.775 84.855 189.445 ;
        RECT 85.035 188.955 85.500 189.265 ;
        RECT 85.680 188.955 86.205 189.265 ;
        RECT 84.565 188.575 85.795 188.775 ;
        RECT 84.635 188.025 85.305 188.395 ;
        RECT 85.485 188.205 85.795 188.575 ;
        RECT 85.975 188.315 86.205 188.955 ;
        RECT 86.385 188.935 86.685 189.265 ;
        RECT 86.865 188.795 87.615 189.315 ;
        RECT 87.785 188.965 88.535 189.485 ;
        RECT 89.165 189.435 89.425 190.575 ;
        RECT 89.595 189.425 89.925 190.405 ;
        RECT 90.095 189.435 90.375 190.575 ;
        RECT 90.555 189.435 90.885 190.575 ;
        RECT 91.415 189.605 91.745 190.390 ;
        RECT 91.065 189.435 91.745 189.605 ;
        RECT 91.985 189.435 92.195 190.575 ;
        RECT 89.185 189.015 89.520 189.265 ;
        RECT 89.690 188.875 89.860 189.425 ;
        RECT 90.030 188.995 90.365 189.265 ;
        RECT 90.545 189.015 90.895 189.265 ;
        RECT 89.685 188.825 89.860 188.875 ;
        RECT 91.065 188.835 91.235 189.435 ;
        RECT 92.365 189.425 92.695 190.405 ;
        RECT 92.865 189.435 93.095 190.575 ;
        RECT 93.325 189.685 93.585 190.395 ;
        RECT 93.755 189.865 94.085 190.575 ;
        RECT 94.255 189.685 94.485 190.395 ;
        RECT 93.325 189.445 94.485 189.685 ;
        RECT 94.665 189.665 94.935 190.395 ;
        RECT 95.115 189.845 95.455 190.575 ;
        RECT 94.665 189.445 95.435 189.665 ;
        RECT 91.405 189.015 91.755 189.265 ;
        RECT 86.385 188.025 86.675 188.755 ;
        RECT 86.865 188.025 88.535 188.795 ;
        RECT 89.165 188.195 89.860 188.825 ;
        RECT 90.065 188.025 90.375 188.825 ;
        RECT 90.555 188.025 90.825 188.835 ;
        RECT 90.995 188.195 91.325 188.835 ;
        RECT 91.495 188.025 91.735 188.835 ;
        RECT 91.985 188.025 92.195 188.845 ;
        RECT 92.365 188.825 92.615 189.425 ;
        RECT 92.785 189.015 93.115 189.265 ;
        RECT 93.315 188.935 93.615 189.265 ;
        RECT 93.795 188.955 94.320 189.265 ;
        RECT 94.500 188.955 94.965 189.265 ;
        RECT 92.365 188.195 92.695 188.825 ;
        RECT 92.865 188.025 93.095 188.845 ;
        RECT 93.325 188.025 93.615 188.755 ;
        RECT 93.795 188.315 94.025 188.955 ;
        RECT 95.145 188.775 95.435 189.445 ;
        RECT 94.205 188.575 95.435 188.775 ;
        RECT 94.205 188.205 94.515 188.575 ;
        RECT 94.695 188.025 95.365 188.395 ;
        RECT 95.625 188.205 95.885 190.395 ;
        RECT 96.065 189.725 96.405 190.365 ;
        RECT 96.575 190.115 96.820 190.575 ;
        RECT 96.995 189.945 97.245 190.405 ;
        RECT 97.435 190.195 98.105 190.575 ;
        RECT 98.305 189.945 98.555 190.405 ;
        RECT 96.995 189.775 98.555 189.945 ;
        RECT 96.065 188.610 96.235 189.725 ;
        RECT 99.315 189.605 99.485 190.405 ;
        RECT 96.545 189.435 99.485 189.605 ;
        RECT 99.780 189.785 100.315 190.405 ;
        RECT 96.545 189.265 96.715 189.435 ;
        RECT 96.405 188.935 96.715 189.265 ;
        RECT 96.885 188.935 97.220 189.265 ;
        RECT 96.545 188.765 96.715 188.935 ;
        RECT 96.065 188.195 96.375 188.610 ;
        RECT 96.545 188.595 97.240 188.765 ;
        RECT 97.490 188.690 97.685 189.265 ;
        RECT 97.945 188.935 98.290 189.265 ;
        RECT 98.600 188.935 99.075 189.265 ;
        RECT 99.330 188.935 99.515 189.265 ;
        RECT 97.945 188.705 98.135 188.935 ;
        RECT 99.780 188.765 100.095 189.785 ;
        RECT 100.485 189.775 100.815 190.575 ;
        RECT 101.300 189.605 101.690 189.780 ;
        RECT 100.265 189.435 101.690 189.605 ;
        RECT 102.065 189.735 102.320 190.405 ;
        RECT 102.490 189.815 102.820 190.575 ;
        RECT 102.990 189.975 103.240 190.405 ;
        RECT 103.410 190.155 103.765 190.575 ;
        RECT 103.955 190.235 105.125 190.405 ;
        RECT 103.955 190.195 104.285 190.235 ;
        RECT 104.395 189.975 104.625 190.065 ;
        RECT 102.990 189.735 104.625 189.975 ;
        RECT 104.795 189.735 105.125 190.235 ;
        RECT 100.265 188.935 100.435 189.435 ;
        RECT 96.570 188.025 96.900 188.405 ;
        RECT 97.070 188.365 97.240 188.595 ;
        RECT 98.305 188.595 99.485 188.765 ;
        RECT 98.305 188.365 98.475 188.595 ;
        RECT 97.070 188.195 98.475 188.365 ;
        RECT 98.745 188.025 99.075 188.425 ;
        RECT 99.315 188.195 99.485 188.595 ;
        RECT 99.780 188.195 100.395 188.765 ;
        RECT 100.685 188.705 100.950 189.265 ;
        RECT 101.120 188.535 101.290 189.435 ;
        RECT 101.460 188.705 101.815 189.265 ;
        RECT 102.065 188.605 102.235 189.735 ;
        RECT 105.295 189.565 105.465 190.405 ;
        RECT 102.405 189.395 105.465 189.565 ;
        RECT 105.765 189.435 105.995 190.575 ;
        RECT 106.165 189.425 106.495 190.405 ;
        RECT 106.665 189.435 106.875 190.575 ;
        RECT 102.405 188.845 102.575 189.395 ;
        RECT 102.805 189.015 103.170 189.215 ;
        RECT 103.340 189.015 103.670 189.215 ;
        RECT 102.405 188.675 103.205 188.845 ;
        RECT 102.065 188.535 102.250 188.605 ;
        RECT 100.565 188.025 100.780 188.535 ;
        RECT 101.010 188.205 101.290 188.535 ;
        RECT 101.470 188.025 101.710 188.535 ;
        RECT 102.065 188.525 102.275 188.535 ;
        RECT 102.065 188.195 102.320 188.525 ;
        RECT 102.535 188.025 102.865 188.505 ;
        RECT 103.035 188.445 103.205 188.675 ;
        RECT 103.385 188.615 103.670 189.015 ;
        RECT 103.940 189.015 104.415 189.215 ;
        RECT 104.585 189.015 105.030 189.215 ;
        RECT 105.200 189.015 105.550 189.225 ;
        RECT 105.745 189.015 106.075 189.265 ;
        RECT 103.940 188.615 104.220 189.015 ;
        RECT 104.400 188.675 105.465 188.845 ;
        RECT 104.400 188.445 104.570 188.675 ;
        RECT 103.035 188.195 104.570 188.445 ;
        RECT 104.795 188.025 105.125 188.505 ;
        RECT 105.295 188.195 105.465 188.675 ;
        RECT 105.765 188.025 105.995 188.845 ;
        RECT 106.245 188.825 106.495 189.425 ;
        RECT 107.565 189.410 107.855 190.575 ;
        RECT 108.035 189.605 108.365 190.390 ;
        RECT 108.035 189.435 108.715 189.605 ;
        RECT 108.895 189.435 109.225 190.575 ;
        RECT 110.330 189.435 110.665 190.405 ;
        RECT 110.835 189.435 111.005 190.575 ;
        RECT 111.175 190.235 113.205 190.405 ;
        RECT 108.025 189.015 108.375 189.265 ;
        RECT 106.165 188.195 106.495 188.825 ;
        RECT 106.665 188.025 106.875 188.845 ;
        RECT 108.545 188.835 108.715 189.435 ;
        RECT 108.885 189.015 109.235 189.265 ;
        RECT 107.565 188.025 107.855 188.750 ;
        RECT 108.045 188.025 108.285 188.835 ;
        RECT 108.455 188.195 108.785 188.835 ;
        RECT 108.955 188.025 109.225 188.835 ;
        RECT 110.330 188.765 110.500 189.435 ;
        RECT 111.175 189.265 111.345 190.235 ;
        RECT 110.670 188.935 110.925 189.265 ;
        RECT 111.150 188.935 111.345 189.265 ;
        RECT 111.515 189.895 112.640 190.065 ;
        RECT 110.755 188.765 110.925 188.935 ;
        RECT 111.515 188.765 111.685 189.895 ;
        RECT 110.330 188.195 110.585 188.765 ;
        RECT 110.755 188.595 111.685 188.765 ;
        RECT 111.855 189.555 112.865 189.725 ;
        RECT 111.855 188.755 112.025 189.555 ;
        RECT 112.230 188.875 112.505 189.355 ;
        RECT 112.225 188.705 112.505 188.875 ;
        RECT 111.510 188.560 111.685 188.595 ;
        RECT 110.755 188.025 111.085 188.425 ;
        RECT 111.510 188.195 112.040 188.560 ;
        RECT 112.230 188.195 112.505 188.705 ;
        RECT 112.675 188.195 112.865 189.555 ;
        RECT 113.035 189.570 113.205 190.235 ;
        RECT 113.375 189.815 113.545 190.575 ;
        RECT 113.780 189.815 114.295 190.225 ;
        RECT 113.035 189.380 113.785 189.570 ;
        RECT 113.955 189.005 114.295 189.815 ;
        RECT 113.065 188.835 114.295 189.005 ;
        RECT 114.465 189.435 114.850 190.405 ;
        RECT 115.020 190.115 115.345 190.575 ;
        RECT 115.865 189.945 116.145 190.405 ;
        RECT 115.020 189.725 116.145 189.945 ;
        RECT 113.045 188.025 113.555 188.560 ;
        RECT 113.775 188.230 114.020 188.835 ;
        RECT 114.465 188.765 114.745 189.435 ;
        RECT 115.020 189.265 115.470 189.725 ;
        RECT 116.335 189.555 116.735 190.405 ;
        RECT 117.135 190.115 117.405 190.575 ;
        RECT 117.575 189.945 117.860 190.405 ;
        RECT 114.915 188.935 115.470 189.265 ;
        RECT 115.640 188.995 116.735 189.555 ;
        RECT 115.020 188.825 115.470 188.935 ;
        RECT 114.465 188.195 114.850 188.765 ;
        RECT 115.020 188.655 116.145 188.825 ;
        RECT 115.020 188.025 115.345 188.485 ;
        RECT 115.865 188.195 116.145 188.655 ;
        RECT 116.335 188.195 116.735 188.995 ;
        RECT 116.905 189.725 117.860 189.945 ;
        RECT 116.905 188.825 117.115 189.725 ;
        RECT 117.285 188.995 117.975 189.555 ;
        RECT 118.145 189.485 121.655 190.575 ;
        RECT 116.905 188.655 117.860 188.825 ;
        RECT 117.135 188.025 117.405 188.485 ;
        RECT 117.575 188.195 117.860 188.655 ;
        RECT 118.145 188.795 119.795 189.315 ;
        RECT 119.965 188.965 121.655 189.485 ;
        RECT 122.285 189.725 122.545 190.405 ;
        RECT 122.715 189.795 122.965 190.575 ;
        RECT 123.215 190.025 123.465 190.405 ;
        RECT 123.635 190.195 123.990 190.575 ;
        RECT 124.995 190.185 125.330 190.405 ;
        RECT 124.595 190.025 124.825 190.065 ;
        RECT 123.215 189.825 124.825 190.025 ;
        RECT 123.215 189.815 124.050 189.825 ;
        RECT 124.640 189.735 124.825 189.825 ;
        RECT 118.145 188.025 121.655 188.795 ;
        RECT 122.285 188.535 122.455 189.725 ;
        RECT 124.155 189.625 124.485 189.655 ;
        RECT 122.685 189.565 124.485 189.625 ;
        RECT 125.075 189.565 125.330 190.185 ;
        RECT 125.505 190.140 130.850 190.575 ;
        RECT 122.625 189.455 125.330 189.565 ;
        RECT 122.625 189.420 122.825 189.455 ;
        RECT 122.625 188.845 122.795 189.420 ;
        RECT 124.155 189.395 125.330 189.455 ;
        RECT 123.025 188.980 123.435 189.285 ;
        RECT 123.605 189.015 123.935 189.225 ;
        RECT 122.625 188.725 122.895 188.845 ;
        RECT 122.625 188.680 123.470 188.725 ;
        RECT 122.715 188.555 123.470 188.680 ;
        RECT 123.725 188.615 123.935 189.015 ;
        RECT 124.180 189.015 124.655 189.225 ;
        RECT 124.845 189.015 125.335 189.215 ;
        RECT 124.180 188.615 124.400 189.015 ;
        RECT 122.285 188.525 122.515 188.535 ;
        RECT 122.285 188.195 122.545 188.525 ;
        RECT 123.300 188.405 123.470 188.555 ;
        RECT 122.715 188.025 123.045 188.385 ;
        RECT 123.300 188.195 124.600 188.405 ;
        RECT 124.875 188.025 125.330 188.790 ;
        RECT 127.090 188.570 127.430 189.400 ;
        RECT 128.910 188.890 129.260 190.140 ;
        RECT 131.025 189.485 132.695 190.575 ;
        RECT 131.025 188.795 131.775 189.315 ;
        RECT 131.945 188.965 132.695 189.485 ;
        RECT 133.325 189.410 133.615 190.575 ;
        RECT 133.785 190.140 139.130 190.575 ;
        RECT 139.305 190.140 144.650 190.575 ;
        RECT 125.505 188.025 130.850 188.570 ;
        RECT 131.025 188.025 132.695 188.795 ;
        RECT 133.325 188.025 133.615 188.750 ;
        RECT 135.370 188.570 135.710 189.400 ;
        RECT 137.190 188.890 137.540 190.140 ;
        RECT 140.890 188.570 141.230 189.400 ;
        RECT 142.710 188.890 143.060 190.140 ;
        RECT 145.745 189.485 146.955 190.575 ;
        RECT 145.745 188.945 146.265 189.485 ;
        RECT 146.435 188.775 146.955 189.315 ;
        RECT 133.785 188.025 139.130 188.570 ;
        RECT 139.305 188.025 144.650 188.570 ;
        RECT 145.745 188.025 146.955 188.775 ;
        RECT 17.320 187.855 147.040 188.025 ;
        RECT 17.405 187.105 18.615 187.855 ;
        RECT 19.295 187.200 19.625 187.635 ;
        RECT 19.795 187.245 19.965 187.855 ;
        RECT 19.245 187.115 19.625 187.200 ;
        RECT 20.135 187.115 20.465 187.640 ;
        RECT 20.725 187.325 20.935 187.855 ;
        RECT 21.210 187.405 21.995 187.575 ;
        RECT 22.165 187.405 22.570 187.575 ;
        RECT 17.405 186.565 17.925 187.105 ;
        RECT 19.245 187.075 19.470 187.115 ;
        RECT 18.095 186.395 18.615 186.935 ;
        RECT 17.405 185.305 18.615 186.395 ;
        RECT 19.245 186.495 19.415 187.075 ;
        RECT 20.135 186.945 20.335 187.115 ;
        RECT 21.210 186.945 21.380 187.405 ;
        RECT 19.585 186.615 20.335 186.945 ;
        RECT 20.505 186.615 21.380 186.945 ;
        RECT 19.245 186.445 19.460 186.495 ;
        RECT 19.245 186.365 19.635 186.445 ;
        RECT 19.305 185.520 19.635 186.365 ;
        RECT 20.145 186.410 20.335 186.615 ;
        RECT 19.805 185.305 19.975 186.315 ;
        RECT 20.145 186.035 21.040 186.410 ;
        RECT 20.145 185.475 20.485 186.035 ;
        RECT 20.715 185.305 21.030 185.805 ;
        RECT 21.210 185.775 21.380 186.615 ;
        RECT 21.550 186.905 22.015 187.235 ;
        RECT 22.400 187.175 22.570 187.405 ;
        RECT 22.750 187.355 23.120 187.855 ;
        RECT 23.440 187.405 24.115 187.575 ;
        RECT 24.310 187.405 24.645 187.575 ;
        RECT 21.550 185.945 21.870 186.905 ;
        RECT 22.400 186.875 23.230 187.175 ;
        RECT 22.040 185.975 22.230 186.695 ;
        RECT 22.400 185.805 22.570 186.875 ;
        RECT 23.030 186.845 23.230 186.875 ;
        RECT 22.740 186.625 22.910 186.695 ;
        RECT 23.440 186.625 23.610 187.405 ;
        RECT 24.475 187.265 24.645 187.405 ;
        RECT 24.815 187.395 25.065 187.855 ;
        RECT 22.740 186.455 23.610 186.625 ;
        RECT 23.780 186.985 24.305 187.205 ;
        RECT 24.475 187.135 24.700 187.265 ;
        RECT 22.740 186.365 23.250 186.455 ;
        RECT 21.210 185.605 22.095 185.775 ;
        RECT 22.320 185.475 22.570 185.805 ;
        RECT 22.740 185.305 22.910 186.105 ;
        RECT 23.080 185.750 23.250 186.365 ;
        RECT 23.780 186.285 23.950 186.985 ;
        RECT 23.420 185.920 23.950 186.285 ;
        RECT 24.120 186.220 24.360 186.815 ;
        RECT 24.530 186.030 24.700 187.135 ;
        RECT 24.870 186.275 25.150 187.225 ;
        RECT 24.395 185.900 24.700 186.030 ;
        RECT 23.080 185.580 24.185 185.750 ;
        RECT 24.395 185.475 24.645 185.900 ;
        RECT 24.815 185.305 25.080 185.765 ;
        RECT 25.320 185.475 25.505 187.595 ;
        RECT 25.675 187.475 26.005 187.855 ;
        RECT 26.175 187.305 26.345 187.595 ;
        RECT 25.680 187.135 26.345 187.305 ;
        RECT 26.605 187.135 26.945 187.645 ;
        RECT 25.680 186.145 25.910 187.135 ;
        RECT 26.080 186.315 26.430 186.965 ;
        RECT 25.680 185.975 26.345 186.145 ;
        RECT 25.675 185.305 26.005 185.805 ;
        RECT 26.175 185.475 26.345 185.975 ;
        RECT 26.605 185.735 26.865 187.135 ;
        RECT 27.115 187.055 27.385 187.855 ;
        RECT 27.040 186.615 27.370 186.865 ;
        RECT 27.565 186.615 27.845 187.585 ;
        RECT 28.025 186.615 28.325 187.585 ;
        RECT 28.505 186.615 28.855 187.580 ;
        RECT 29.075 187.355 29.570 187.685 ;
        RECT 27.055 186.445 27.370 186.615 ;
        RECT 29.075 186.445 29.245 187.355 ;
        RECT 27.055 186.275 29.245 186.445 ;
        RECT 26.605 185.475 26.945 185.735 ;
        RECT 27.115 185.305 27.445 186.105 ;
        RECT 27.910 185.475 28.160 186.275 ;
        RECT 28.345 185.305 28.675 186.025 ;
        RECT 28.895 185.475 29.145 186.275 ;
        RECT 29.415 185.865 29.655 187.175 ;
        RECT 29.835 187.130 30.165 187.640 ;
        RECT 30.335 187.455 30.665 187.855 ;
        RECT 31.715 187.285 32.045 187.625 ;
        RECT 32.215 187.455 32.545 187.855 ;
        RECT 33.520 187.285 33.775 187.635 ;
        RECT 33.945 187.455 34.275 187.855 ;
        RECT 34.445 187.285 34.615 187.635 ;
        RECT 34.785 187.455 35.165 187.855 ;
        RECT 29.835 186.365 30.025 187.130 ;
        RECT 30.335 187.115 32.700 187.285 ;
        RECT 33.520 187.115 35.185 187.285 ;
        RECT 35.355 187.180 35.630 187.525 ;
        RECT 30.335 186.945 30.505 187.115 ;
        RECT 30.195 186.615 30.505 186.945 ;
        RECT 30.675 186.615 30.980 186.945 ;
        RECT 29.315 185.305 29.650 185.685 ;
        RECT 29.835 185.515 30.165 186.365 ;
        RECT 30.335 185.305 30.585 186.445 ;
        RECT 30.765 186.285 30.980 186.615 ;
        RECT 31.155 186.285 31.440 186.945 ;
        RECT 31.635 186.285 31.900 186.945 ;
        RECT 32.115 186.285 32.360 186.945 ;
        RECT 32.530 186.115 32.700 187.115 ;
        RECT 35.015 186.945 35.185 187.115 ;
        RECT 33.505 186.615 33.850 186.945 ;
        RECT 34.020 186.615 34.845 186.945 ;
        RECT 35.015 186.615 35.290 186.945 ;
        RECT 30.775 185.945 32.065 186.115 ;
        RECT 30.775 185.525 31.025 185.945 ;
        RECT 31.255 185.305 31.585 185.775 ;
        RECT 31.815 185.525 32.065 185.945 ;
        RECT 32.245 185.945 32.700 186.115 ;
        RECT 33.525 186.155 33.850 186.445 ;
        RECT 34.020 186.325 34.215 186.615 ;
        RECT 35.015 186.445 35.185 186.615 ;
        RECT 35.460 186.445 35.630 187.180 ;
        RECT 35.805 187.245 36.145 187.660 ;
        RECT 36.315 187.415 36.485 187.855 ;
        RECT 36.655 187.465 37.905 187.645 ;
        RECT 36.655 187.245 36.985 187.465 ;
        RECT 38.175 187.395 38.345 187.855 ;
        RECT 35.805 187.075 36.985 187.245 ;
        RECT 37.155 187.225 37.520 187.295 ;
        RECT 37.155 187.045 38.405 187.225 ;
        RECT 35.805 186.665 36.270 186.865 ;
        RECT 36.445 186.615 36.775 186.865 ;
        RECT 36.945 186.835 37.410 186.865 ;
        RECT 36.945 186.665 37.415 186.835 ;
        RECT 36.945 186.615 37.410 186.665 ;
        RECT 37.605 186.615 37.960 186.865 ;
        RECT 36.445 186.495 36.625 186.615 ;
        RECT 34.525 186.275 35.185 186.445 ;
        RECT 34.525 186.155 34.695 186.275 ;
        RECT 33.525 185.985 34.695 186.155 ;
        RECT 32.245 185.515 32.575 185.945 ;
        RECT 33.505 185.525 34.695 185.815 ;
        RECT 34.865 185.305 35.145 186.105 ;
        RECT 35.355 185.475 35.630 186.445 ;
        RECT 35.805 185.305 36.125 186.485 ;
        RECT 36.295 186.325 36.625 186.495 ;
        RECT 38.130 186.445 38.405 187.045 ;
        RECT 36.295 185.535 36.495 186.325 ;
        RECT 36.795 186.235 38.405 186.445 ;
        RECT 36.795 186.135 37.205 186.235 ;
        RECT 36.820 185.475 37.205 186.135 ;
        RECT 37.600 185.305 38.385 186.065 ;
        RECT 38.575 185.475 38.855 187.575 ;
        RECT 39.030 187.090 39.485 187.855 ;
        RECT 39.760 187.475 41.060 187.685 ;
        RECT 41.315 187.495 41.645 187.855 ;
        RECT 40.890 187.325 41.060 187.475 ;
        RECT 41.815 187.355 42.075 187.685 ;
        RECT 39.960 186.865 40.180 187.265 ;
        RECT 39.025 186.665 39.515 186.865 ;
        RECT 39.705 186.655 40.180 186.865 ;
        RECT 40.425 186.865 40.635 187.265 ;
        RECT 40.890 187.200 41.645 187.325 ;
        RECT 40.890 187.155 41.735 187.200 ;
        RECT 41.465 187.035 41.735 187.155 ;
        RECT 40.425 186.655 40.755 186.865 ;
        RECT 40.925 186.595 41.335 186.900 ;
        RECT 39.030 186.425 40.205 186.485 ;
        RECT 41.565 186.460 41.735 187.035 ;
        RECT 41.535 186.425 41.735 186.460 ;
        RECT 39.030 186.315 41.735 186.425 ;
        RECT 39.030 185.695 39.285 186.315 ;
        RECT 39.875 186.255 41.675 186.315 ;
        RECT 39.875 186.225 40.205 186.255 ;
        RECT 41.905 186.155 42.075 187.355 ;
        RECT 43.165 187.130 43.455 187.855 ;
        RECT 43.630 187.205 43.900 187.415 ;
        RECT 44.120 187.395 44.450 187.855 ;
        RECT 44.960 187.395 45.710 187.685 ;
        RECT 45.930 187.455 46.265 187.855 ;
        RECT 43.630 187.035 44.965 187.205 ;
        RECT 44.795 186.865 44.965 187.035 ;
        RECT 43.630 186.625 43.980 186.865 ;
        RECT 44.150 186.625 44.625 186.865 ;
        RECT 44.795 186.615 45.170 186.865 ;
        RECT 39.535 186.055 39.720 186.145 ;
        RECT 40.310 186.055 41.145 186.065 ;
        RECT 39.535 185.855 41.145 186.055 ;
        RECT 39.535 185.815 39.765 185.855 ;
        RECT 39.030 185.475 39.365 185.695 ;
        RECT 40.370 185.305 40.725 185.685 ;
        RECT 40.895 185.475 41.145 185.855 ;
        RECT 41.395 185.305 41.645 186.085 ;
        RECT 41.815 185.475 42.075 186.155 ;
        RECT 43.165 185.305 43.455 186.470 ;
        RECT 44.795 186.445 44.965 186.615 ;
        RECT 43.630 186.275 44.965 186.445 ;
        RECT 43.630 186.115 43.910 186.275 ;
        RECT 45.340 186.105 45.710 187.395 ;
        RECT 46.435 187.285 46.640 187.685 ;
        RECT 46.850 187.375 47.125 187.855 ;
        RECT 47.335 187.355 47.595 187.685 ;
        RECT 44.120 185.305 44.370 186.105 ;
        RECT 44.540 185.935 45.710 186.105 ;
        RECT 45.955 187.115 46.640 187.285 ;
        RECT 45.955 186.085 46.295 187.115 ;
        RECT 46.465 186.445 46.715 186.945 ;
        RECT 46.895 186.615 47.255 187.195 ;
        RECT 47.425 186.445 47.595 187.355 ;
        RECT 47.765 187.085 50.355 187.855 ;
        RECT 47.765 186.565 48.975 187.085 ;
        RECT 50.985 187.055 51.295 187.855 ;
        RECT 51.500 187.055 52.195 187.685 ;
        RECT 52.380 187.285 52.635 187.635 ;
        RECT 52.805 187.455 53.135 187.855 ;
        RECT 53.305 187.285 53.475 187.635 ;
        RECT 53.645 187.455 54.025 187.855 ;
        RECT 52.380 187.115 54.045 187.285 ;
        RECT 54.215 187.180 54.490 187.525 ;
        RECT 46.465 186.275 47.595 186.445 ;
        RECT 49.145 186.395 50.355 186.915 ;
        RECT 50.995 186.615 51.330 186.885 ;
        RECT 51.500 186.455 51.670 187.055 ;
        RECT 53.875 186.945 54.045 187.115 ;
        RECT 51.840 186.615 52.175 186.865 ;
        RECT 52.365 186.615 52.710 186.945 ;
        RECT 52.880 186.615 53.705 186.945 ;
        RECT 53.875 186.615 54.150 186.945 ;
        RECT 44.540 185.475 44.870 185.935 ;
        RECT 45.955 185.910 46.620 186.085 ;
        RECT 45.040 185.305 45.255 185.765 ;
        RECT 45.930 185.305 46.265 185.730 ;
        RECT 46.435 185.505 46.620 185.910 ;
        RECT 46.825 185.305 47.155 186.085 ;
        RECT 47.325 185.505 47.595 186.275 ;
        RECT 47.765 185.305 50.355 186.395 ;
        RECT 50.985 185.305 51.265 186.445 ;
        RECT 51.435 185.475 51.765 186.455 ;
        RECT 51.935 185.305 52.195 186.445 ;
        RECT 52.385 186.155 52.710 186.445 ;
        RECT 52.880 186.325 53.075 186.615 ;
        RECT 53.875 186.445 54.045 186.615 ;
        RECT 54.320 186.445 54.490 187.180 ;
        RECT 53.385 186.275 54.045 186.445 ;
        RECT 53.385 186.155 53.555 186.275 ;
        RECT 52.385 185.985 53.555 186.155 ;
        RECT 52.365 185.525 53.555 185.815 ;
        RECT 53.725 185.305 54.005 186.105 ;
        RECT 54.215 185.475 54.490 186.445 ;
        RECT 54.665 185.475 54.945 187.575 ;
        RECT 55.175 187.395 55.345 187.855 ;
        RECT 55.615 187.465 56.865 187.645 ;
        RECT 56.000 187.225 56.365 187.295 ;
        RECT 55.115 187.045 56.365 187.225 ;
        RECT 56.535 187.245 56.865 187.465 ;
        RECT 57.035 187.415 57.205 187.855 ;
        RECT 57.375 187.245 57.715 187.660 ;
        RECT 56.535 187.075 57.715 187.245 ;
        RECT 58.090 187.075 58.590 187.685 ;
        RECT 55.115 186.445 55.390 187.045 ;
        RECT 55.560 186.615 55.915 186.865 ;
        RECT 56.110 186.835 56.575 186.865 ;
        RECT 56.105 186.665 56.575 186.835 ;
        RECT 56.110 186.615 56.575 186.665 ;
        RECT 56.745 186.615 57.075 186.865 ;
        RECT 57.250 186.665 57.715 186.865 ;
        RECT 57.885 186.615 58.235 186.865 ;
        RECT 56.895 186.495 57.075 186.615 ;
        RECT 55.115 186.235 56.725 186.445 ;
        RECT 56.895 186.325 57.225 186.495 ;
        RECT 56.315 186.135 56.725 186.235 ;
        RECT 55.135 185.305 55.920 186.065 ;
        RECT 56.315 185.475 56.700 186.135 ;
        RECT 57.025 185.535 57.225 186.325 ;
        RECT 57.395 185.305 57.715 186.485 ;
        RECT 58.420 186.445 58.590 187.075 ;
        RECT 59.220 187.205 59.550 187.685 ;
        RECT 59.720 187.395 59.945 187.855 ;
        RECT 60.115 187.205 60.445 187.685 ;
        RECT 59.220 187.035 60.445 187.205 ;
        RECT 60.635 187.055 60.885 187.855 ;
        RECT 61.055 187.055 61.395 187.685 ;
        RECT 61.585 187.125 61.875 187.855 ;
        RECT 58.760 186.665 59.090 186.865 ;
        RECT 59.260 186.665 59.590 186.865 ;
        RECT 59.760 186.665 60.180 186.865 ;
        RECT 60.355 186.695 61.050 186.865 ;
        RECT 60.355 186.445 60.525 186.695 ;
        RECT 61.220 186.445 61.395 187.055 ;
        RECT 61.575 186.615 61.875 186.945 ;
        RECT 62.055 186.925 62.285 187.565 ;
        RECT 62.465 187.305 62.775 187.675 ;
        RECT 62.955 187.485 63.625 187.855 ;
        RECT 62.465 187.105 63.695 187.305 ;
        RECT 62.055 186.615 62.580 186.925 ;
        RECT 62.760 186.615 63.225 186.925 ;
        RECT 58.090 186.275 60.525 186.445 ;
        RECT 58.090 185.475 58.420 186.275 ;
        RECT 58.590 185.305 58.920 186.105 ;
        RECT 59.220 185.475 59.550 186.275 ;
        RECT 60.195 185.305 60.445 186.105 ;
        RECT 60.715 185.305 60.885 186.445 ;
        RECT 61.055 185.475 61.395 186.445 ;
        RECT 63.405 186.435 63.695 187.105 ;
        RECT 61.585 186.195 62.745 186.435 ;
        RECT 61.585 185.485 61.845 186.195 ;
        RECT 62.015 185.305 62.345 186.015 ;
        RECT 62.515 185.485 62.745 186.195 ;
        RECT 62.925 186.215 63.695 186.435 ;
        RECT 62.925 185.485 63.195 186.215 ;
        RECT 63.375 185.305 63.715 186.035 ;
        RECT 63.885 185.485 64.145 187.675 ;
        RECT 64.325 187.085 67.835 187.855 ;
        RECT 68.925 187.130 69.215 187.855 ;
        RECT 69.385 187.085 71.055 187.855 ;
        RECT 71.230 187.285 71.485 187.555 ;
        RECT 71.655 187.455 71.985 187.855 ;
        RECT 72.155 187.285 72.325 187.555 ;
        RECT 72.495 187.455 72.825 187.855 ;
        RECT 71.230 187.115 72.455 187.285 ;
        RECT 64.325 186.565 65.975 187.085 ;
        RECT 66.145 186.395 67.835 186.915 ;
        RECT 69.385 186.565 70.135 187.085 ;
        RECT 64.325 185.305 67.835 186.395 ;
        RECT 68.925 185.305 69.215 186.470 ;
        RECT 70.305 186.395 71.055 186.915 ;
        RECT 71.230 186.615 71.565 186.945 ;
        RECT 71.735 186.615 72.115 186.945 ;
        RECT 69.385 185.305 71.055 186.395 ;
        RECT 71.230 185.660 71.565 186.445 ;
        RECT 71.735 185.935 71.970 186.615 ;
        RECT 72.285 186.445 72.455 187.115 ;
        RECT 72.140 186.275 72.455 186.445 ;
        RECT 72.625 186.275 72.895 187.285 ;
        RECT 73.115 187.200 73.445 187.635 ;
        RECT 73.615 187.245 73.785 187.855 ;
        RECT 73.065 187.115 73.445 187.200 ;
        RECT 73.955 187.115 74.285 187.640 ;
        RECT 74.545 187.325 74.755 187.855 ;
        RECT 75.030 187.405 75.815 187.575 ;
        RECT 75.985 187.405 76.390 187.575 ;
        RECT 73.065 187.075 73.290 187.115 ;
        RECT 73.065 186.495 73.235 187.075 ;
        RECT 73.955 186.945 74.155 187.115 ;
        RECT 75.030 186.945 75.200 187.405 ;
        RECT 73.405 186.615 74.155 186.945 ;
        RECT 74.325 186.615 75.200 186.945 ;
        RECT 73.065 186.445 73.280 186.495 ;
        RECT 73.065 186.365 73.455 186.445 ;
        RECT 72.140 185.660 72.310 186.275 ;
        RECT 71.230 185.490 72.310 185.660 ;
        RECT 72.575 185.305 72.890 186.105 ;
        RECT 73.125 185.520 73.455 186.365 ;
        RECT 73.965 186.410 74.155 186.615 ;
        RECT 73.625 185.305 73.795 186.315 ;
        RECT 73.965 186.035 74.860 186.410 ;
        RECT 73.965 185.475 74.305 186.035 ;
        RECT 74.535 185.305 74.850 185.805 ;
        RECT 75.030 185.775 75.200 186.615 ;
        RECT 75.370 186.905 75.835 187.235 ;
        RECT 76.220 187.175 76.390 187.405 ;
        RECT 76.570 187.355 76.940 187.855 ;
        RECT 77.260 187.405 77.935 187.575 ;
        RECT 78.130 187.405 78.465 187.575 ;
        RECT 75.370 185.945 75.690 186.905 ;
        RECT 76.220 186.875 77.050 187.175 ;
        RECT 75.860 185.975 76.050 186.695 ;
        RECT 76.220 185.805 76.390 186.875 ;
        RECT 76.850 186.845 77.050 186.875 ;
        RECT 76.560 186.625 76.730 186.695 ;
        RECT 77.260 186.625 77.430 187.405 ;
        RECT 78.295 187.265 78.465 187.405 ;
        RECT 78.635 187.395 78.885 187.855 ;
        RECT 76.560 186.455 77.430 186.625 ;
        RECT 77.600 186.985 78.125 187.205 ;
        RECT 78.295 187.135 78.520 187.265 ;
        RECT 76.560 186.365 77.070 186.455 ;
        RECT 75.030 185.605 75.915 185.775 ;
        RECT 76.140 185.475 76.390 185.805 ;
        RECT 76.560 185.305 76.730 186.105 ;
        RECT 76.900 185.750 77.070 186.365 ;
        RECT 77.600 186.285 77.770 186.985 ;
        RECT 77.240 185.920 77.770 186.285 ;
        RECT 77.940 186.220 78.180 186.815 ;
        RECT 78.350 186.030 78.520 187.135 ;
        RECT 78.690 186.275 78.970 187.225 ;
        RECT 78.215 185.900 78.520 186.030 ;
        RECT 76.900 185.580 78.005 185.750 ;
        RECT 78.215 185.475 78.465 185.900 ;
        RECT 78.635 185.305 78.900 185.765 ;
        RECT 79.140 185.475 79.325 187.595 ;
        RECT 79.495 187.475 79.825 187.855 ;
        RECT 79.995 187.305 80.165 187.595 ;
        RECT 79.500 187.135 80.165 187.305 ;
        RECT 80.975 187.305 81.145 187.595 ;
        RECT 81.315 187.475 81.645 187.855 ;
        RECT 80.975 187.135 81.640 187.305 ;
        RECT 79.500 186.145 79.730 187.135 ;
        RECT 79.900 186.315 80.250 186.965 ;
        RECT 80.890 186.315 81.240 186.965 ;
        RECT 81.410 186.145 81.640 187.135 ;
        RECT 79.500 185.975 80.165 186.145 ;
        RECT 79.495 185.305 79.825 185.805 ;
        RECT 79.995 185.475 80.165 185.975 ;
        RECT 80.975 185.975 81.640 186.145 ;
        RECT 80.975 185.475 81.145 185.975 ;
        RECT 81.315 185.305 81.645 185.805 ;
        RECT 81.815 185.475 82.000 187.595 ;
        RECT 82.255 187.395 82.505 187.855 ;
        RECT 82.675 187.405 83.010 187.575 ;
        RECT 83.205 187.405 83.880 187.575 ;
        RECT 82.675 187.265 82.845 187.405 ;
        RECT 82.170 186.275 82.450 187.225 ;
        RECT 82.620 187.135 82.845 187.265 ;
        RECT 82.620 186.030 82.790 187.135 ;
        RECT 83.015 186.985 83.540 187.205 ;
        RECT 82.960 186.220 83.200 186.815 ;
        RECT 83.370 186.285 83.540 186.985 ;
        RECT 83.710 186.625 83.880 187.405 ;
        RECT 84.200 187.355 84.570 187.855 ;
        RECT 84.750 187.405 85.155 187.575 ;
        RECT 85.325 187.405 86.110 187.575 ;
        RECT 84.750 187.175 84.920 187.405 ;
        RECT 84.090 186.875 84.920 187.175 ;
        RECT 85.305 186.905 85.770 187.235 ;
        RECT 84.090 186.845 84.290 186.875 ;
        RECT 84.410 186.625 84.580 186.695 ;
        RECT 83.710 186.455 84.580 186.625 ;
        RECT 84.070 186.365 84.580 186.455 ;
        RECT 82.620 185.900 82.925 186.030 ;
        RECT 83.370 185.920 83.900 186.285 ;
        RECT 82.240 185.305 82.505 185.765 ;
        RECT 82.675 185.475 82.925 185.900 ;
        RECT 84.070 185.750 84.240 186.365 ;
        RECT 83.135 185.580 84.240 185.750 ;
        RECT 84.410 185.305 84.580 186.105 ;
        RECT 84.750 185.805 84.920 186.875 ;
        RECT 85.090 185.975 85.280 186.695 ;
        RECT 85.450 185.945 85.770 186.905 ;
        RECT 85.940 186.945 86.110 187.405 ;
        RECT 86.385 187.325 86.595 187.855 ;
        RECT 86.855 187.115 87.185 187.640 ;
        RECT 87.355 187.245 87.525 187.855 ;
        RECT 87.695 187.200 88.025 187.635 ;
        RECT 88.245 187.310 93.590 187.855 ;
        RECT 87.695 187.115 88.075 187.200 ;
        RECT 86.985 186.945 87.185 187.115 ;
        RECT 87.850 187.075 88.075 187.115 ;
        RECT 85.940 186.615 86.815 186.945 ;
        RECT 86.985 186.615 87.735 186.945 ;
        RECT 84.750 185.475 85.000 185.805 ;
        RECT 85.940 185.775 86.110 186.615 ;
        RECT 86.985 186.410 87.175 186.615 ;
        RECT 87.905 186.495 88.075 187.075 ;
        RECT 87.860 186.445 88.075 186.495 ;
        RECT 89.830 186.480 90.170 187.310 ;
        RECT 94.685 187.130 94.975 187.855 ;
        RECT 95.145 187.085 97.735 187.855 ;
        RECT 97.910 187.090 98.365 187.855 ;
        RECT 98.640 187.475 99.940 187.685 ;
        RECT 100.195 187.495 100.525 187.855 ;
        RECT 99.770 187.325 99.940 187.475 ;
        RECT 100.695 187.355 100.955 187.685 ;
        RECT 101.915 187.455 102.245 187.855 ;
        RECT 100.725 187.345 100.955 187.355 ;
        RECT 86.280 186.035 87.175 186.410 ;
        RECT 87.685 186.365 88.075 186.445 ;
        RECT 85.225 185.605 86.110 185.775 ;
        RECT 86.290 185.305 86.605 185.805 ;
        RECT 86.835 185.475 87.175 186.035 ;
        RECT 87.345 185.305 87.515 186.315 ;
        RECT 87.685 185.520 88.015 186.365 ;
        RECT 91.650 185.740 92.000 186.990 ;
        RECT 95.145 186.565 96.355 187.085 ;
        RECT 88.245 185.305 93.590 185.740 ;
        RECT 94.685 185.305 94.975 186.470 ;
        RECT 96.525 186.395 97.735 186.915 ;
        RECT 98.840 186.865 99.060 187.265 ;
        RECT 97.905 186.665 98.395 186.865 ;
        RECT 98.585 186.655 99.060 186.865 ;
        RECT 99.305 186.865 99.515 187.265 ;
        RECT 99.770 187.200 100.525 187.325 ;
        RECT 99.770 187.155 100.615 187.200 ;
        RECT 100.345 187.035 100.615 187.155 ;
        RECT 99.305 186.655 99.635 186.865 ;
        RECT 99.805 186.595 100.215 186.900 ;
        RECT 95.145 185.305 97.735 186.395 ;
        RECT 97.910 186.425 99.085 186.485 ;
        RECT 100.445 186.460 100.615 187.035 ;
        RECT 100.415 186.425 100.615 186.460 ;
        RECT 97.910 186.315 100.615 186.425 ;
        RECT 97.910 185.695 98.165 186.315 ;
        RECT 98.755 186.255 100.555 186.315 ;
        RECT 98.755 186.225 99.085 186.255 ;
        RECT 100.785 186.155 100.955 187.345 ;
        RECT 102.415 187.285 102.745 187.625 ;
        RECT 103.795 187.455 104.125 187.855 ;
        RECT 98.415 186.055 98.600 186.145 ;
        RECT 99.190 186.055 100.025 186.065 ;
        RECT 98.415 185.855 100.025 186.055 ;
        RECT 98.415 185.815 98.645 185.855 ;
        RECT 97.910 185.475 98.245 185.695 ;
        RECT 99.250 185.305 99.605 185.685 ;
        RECT 99.775 185.475 100.025 185.855 ;
        RECT 100.275 185.305 100.525 186.085 ;
        RECT 100.695 185.475 100.955 186.155 ;
        RECT 101.760 187.115 104.125 187.285 ;
        RECT 104.295 187.130 104.625 187.640 ;
        RECT 101.760 186.115 101.930 187.115 ;
        RECT 103.955 186.945 104.125 187.115 ;
        RECT 102.100 186.285 102.345 186.945 ;
        RECT 102.560 186.285 102.825 186.945 ;
        RECT 103.020 186.285 103.305 186.945 ;
        RECT 103.480 186.615 103.785 186.945 ;
        RECT 103.955 186.615 104.265 186.945 ;
        RECT 103.480 186.285 103.695 186.615 ;
        RECT 101.760 185.945 102.215 186.115 ;
        RECT 101.885 185.515 102.215 185.945 ;
        RECT 102.395 185.945 103.685 186.115 ;
        RECT 102.395 185.525 102.645 185.945 ;
        RECT 102.875 185.305 103.205 185.775 ;
        RECT 103.435 185.525 103.685 185.945 ;
        RECT 103.875 185.305 104.125 186.445 ;
        RECT 104.435 186.365 104.625 187.130 ;
        RECT 104.845 187.035 105.075 187.855 ;
        RECT 105.245 187.055 105.575 187.685 ;
        RECT 104.825 186.615 105.155 186.865 ;
        RECT 105.325 186.455 105.575 187.055 ;
        RECT 105.745 187.035 105.955 187.855 ;
        RECT 106.185 187.105 107.395 187.855 ;
        RECT 107.655 187.305 107.825 187.595 ;
        RECT 107.995 187.475 108.325 187.855 ;
        RECT 107.655 187.135 108.320 187.305 ;
        RECT 106.185 186.565 106.705 187.105 ;
        RECT 104.295 185.515 104.625 186.365 ;
        RECT 104.845 185.305 105.075 186.445 ;
        RECT 105.245 185.475 105.575 186.455 ;
        RECT 105.745 185.305 105.955 186.445 ;
        RECT 106.875 186.395 107.395 186.935 ;
        RECT 106.185 185.305 107.395 186.395 ;
        RECT 107.570 186.315 107.920 186.965 ;
        RECT 108.090 186.145 108.320 187.135 ;
        RECT 107.655 185.975 108.320 186.145 ;
        RECT 107.655 185.475 107.825 185.975 ;
        RECT 107.995 185.305 108.325 185.805 ;
        RECT 108.495 185.475 108.680 187.595 ;
        RECT 108.935 187.395 109.185 187.855 ;
        RECT 109.355 187.405 109.690 187.575 ;
        RECT 109.885 187.405 110.560 187.575 ;
        RECT 109.355 187.265 109.525 187.405 ;
        RECT 108.850 186.275 109.130 187.225 ;
        RECT 109.300 187.135 109.525 187.265 ;
        RECT 109.300 186.030 109.470 187.135 ;
        RECT 109.695 186.985 110.220 187.205 ;
        RECT 109.640 186.220 109.880 186.815 ;
        RECT 110.050 186.285 110.220 186.985 ;
        RECT 110.390 186.625 110.560 187.405 ;
        RECT 110.880 187.355 111.250 187.855 ;
        RECT 111.430 187.405 111.835 187.575 ;
        RECT 112.005 187.405 112.790 187.575 ;
        RECT 111.430 187.175 111.600 187.405 ;
        RECT 110.770 186.875 111.600 187.175 ;
        RECT 111.985 186.905 112.450 187.235 ;
        RECT 110.770 186.845 110.970 186.875 ;
        RECT 111.090 186.625 111.260 186.695 ;
        RECT 110.390 186.455 111.260 186.625 ;
        RECT 110.750 186.365 111.260 186.455 ;
        RECT 109.300 185.900 109.605 186.030 ;
        RECT 110.050 185.920 110.580 186.285 ;
        RECT 108.920 185.305 109.185 185.765 ;
        RECT 109.355 185.475 109.605 185.900 ;
        RECT 110.750 185.750 110.920 186.365 ;
        RECT 109.815 185.580 110.920 185.750 ;
        RECT 111.090 185.305 111.260 186.105 ;
        RECT 111.430 185.805 111.600 186.875 ;
        RECT 111.770 185.975 111.960 186.695 ;
        RECT 112.130 185.945 112.450 186.905 ;
        RECT 112.620 186.945 112.790 187.405 ;
        RECT 113.065 187.325 113.275 187.855 ;
        RECT 113.535 187.115 113.865 187.640 ;
        RECT 114.035 187.245 114.205 187.855 ;
        RECT 114.375 187.200 114.705 187.635 ;
        RECT 114.925 187.310 120.270 187.855 ;
        RECT 114.375 187.115 114.755 187.200 ;
        RECT 113.665 186.945 113.865 187.115 ;
        RECT 114.530 187.075 114.755 187.115 ;
        RECT 112.620 186.615 113.495 186.945 ;
        RECT 113.665 186.615 114.415 186.945 ;
        RECT 111.430 185.475 111.680 185.805 ;
        RECT 112.620 185.775 112.790 186.615 ;
        RECT 113.665 186.410 113.855 186.615 ;
        RECT 114.585 186.495 114.755 187.075 ;
        RECT 114.540 186.445 114.755 186.495 ;
        RECT 116.510 186.480 116.850 187.310 ;
        RECT 120.445 187.130 120.735 187.855 ;
        RECT 120.910 187.115 121.165 187.685 ;
        RECT 121.335 187.455 121.665 187.855 ;
        RECT 122.090 187.320 122.620 187.685 ;
        RECT 122.090 187.285 122.265 187.320 ;
        RECT 121.335 187.115 122.265 187.285 ;
        RECT 112.960 186.035 113.855 186.410 ;
        RECT 114.365 186.365 114.755 186.445 ;
        RECT 111.905 185.605 112.790 185.775 ;
        RECT 112.970 185.305 113.285 185.805 ;
        RECT 113.515 185.475 113.855 186.035 ;
        RECT 114.025 185.305 114.195 186.315 ;
        RECT 114.365 185.520 114.695 186.365 ;
        RECT 118.330 185.740 118.680 186.990 ;
        RECT 114.925 185.305 120.270 185.740 ;
        RECT 120.445 185.305 120.735 186.470 ;
        RECT 120.910 186.445 121.080 187.115 ;
        RECT 121.335 186.945 121.505 187.115 ;
        RECT 121.250 186.615 121.505 186.945 ;
        RECT 121.730 186.615 121.925 186.945 ;
        RECT 120.910 185.475 121.245 186.445 ;
        RECT 121.415 185.305 121.585 186.445 ;
        RECT 121.755 185.645 121.925 186.615 ;
        RECT 122.095 185.985 122.265 187.115 ;
        RECT 122.435 186.325 122.605 187.125 ;
        RECT 122.810 186.835 123.085 187.685 ;
        RECT 122.805 186.665 123.085 186.835 ;
        RECT 122.810 186.525 123.085 186.665 ;
        RECT 123.255 186.325 123.445 187.685 ;
        RECT 123.625 187.320 124.135 187.855 ;
        RECT 124.355 187.045 124.600 187.650 ;
        RECT 126.015 187.200 126.345 187.635 ;
        RECT 126.515 187.245 126.685 187.855 ;
        RECT 125.965 187.115 126.345 187.200 ;
        RECT 126.855 187.115 127.185 187.640 ;
        RECT 127.445 187.325 127.655 187.855 ;
        RECT 127.930 187.405 128.715 187.575 ;
        RECT 128.885 187.405 129.290 187.575 ;
        RECT 125.965 187.075 126.190 187.115 ;
        RECT 123.645 186.875 124.875 187.045 ;
        RECT 122.435 186.155 123.445 186.325 ;
        RECT 123.615 186.310 124.365 186.500 ;
        RECT 122.095 185.815 123.220 185.985 ;
        RECT 123.615 185.645 123.785 186.310 ;
        RECT 124.535 186.065 124.875 186.875 ;
        RECT 125.965 186.495 126.135 187.075 ;
        RECT 126.855 186.945 127.055 187.115 ;
        RECT 127.930 186.945 128.100 187.405 ;
        RECT 126.305 186.615 127.055 186.945 ;
        RECT 127.225 186.615 128.100 186.945 ;
        RECT 125.965 186.445 126.180 186.495 ;
        RECT 125.965 186.365 126.355 186.445 ;
        RECT 121.755 185.475 123.785 185.645 ;
        RECT 123.955 185.305 124.125 186.065 ;
        RECT 124.360 185.655 124.875 186.065 ;
        RECT 126.025 185.520 126.355 186.365 ;
        RECT 126.865 186.410 127.055 186.615 ;
        RECT 126.525 185.305 126.695 186.315 ;
        RECT 126.865 186.035 127.760 186.410 ;
        RECT 126.865 185.475 127.205 186.035 ;
        RECT 127.435 185.305 127.750 185.805 ;
        RECT 127.930 185.775 128.100 186.615 ;
        RECT 128.270 186.905 128.735 187.235 ;
        RECT 129.120 187.175 129.290 187.405 ;
        RECT 129.470 187.355 129.840 187.855 ;
        RECT 130.160 187.405 130.835 187.575 ;
        RECT 131.030 187.405 131.365 187.575 ;
        RECT 128.270 185.945 128.590 186.905 ;
        RECT 129.120 186.875 129.950 187.175 ;
        RECT 128.760 185.975 128.950 186.695 ;
        RECT 129.120 185.805 129.290 186.875 ;
        RECT 129.750 186.845 129.950 186.875 ;
        RECT 129.460 186.625 129.630 186.695 ;
        RECT 130.160 186.625 130.330 187.405 ;
        RECT 131.195 187.265 131.365 187.405 ;
        RECT 131.535 187.395 131.785 187.855 ;
        RECT 129.460 186.455 130.330 186.625 ;
        RECT 130.500 186.985 131.025 187.205 ;
        RECT 131.195 187.135 131.420 187.265 ;
        RECT 129.460 186.365 129.970 186.455 ;
        RECT 127.930 185.605 128.815 185.775 ;
        RECT 129.040 185.475 129.290 185.805 ;
        RECT 129.460 185.305 129.630 186.105 ;
        RECT 129.800 185.750 129.970 186.365 ;
        RECT 130.500 186.285 130.670 186.985 ;
        RECT 130.140 185.920 130.670 186.285 ;
        RECT 130.840 186.220 131.080 186.815 ;
        RECT 131.250 186.030 131.420 187.135 ;
        RECT 131.590 186.275 131.870 187.225 ;
        RECT 131.115 185.900 131.420 186.030 ;
        RECT 129.800 185.580 130.905 185.750 ;
        RECT 131.115 185.475 131.365 185.900 ;
        RECT 131.535 185.305 131.800 185.765 ;
        RECT 132.040 185.475 132.225 187.595 ;
        RECT 132.395 187.475 132.725 187.855 ;
        RECT 132.895 187.305 133.065 187.595 ;
        RECT 133.330 187.455 133.665 187.855 ;
        RECT 132.400 187.135 133.065 187.305 ;
        RECT 133.835 187.285 134.040 187.685 ;
        RECT 134.250 187.375 134.525 187.855 ;
        RECT 134.735 187.355 134.995 187.685 ;
        RECT 132.400 186.145 132.630 187.135 ;
        RECT 133.355 187.115 134.040 187.285 ;
        RECT 132.800 186.315 133.150 186.965 ;
        RECT 132.400 185.975 133.065 186.145 ;
        RECT 132.395 185.305 132.725 185.805 ;
        RECT 132.895 185.475 133.065 185.975 ;
        RECT 133.355 186.085 133.695 187.115 ;
        RECT 133.865 186.445 134.115 186.945 ;
        RECT 134.295 186.615 134.655 187.195 ;
        RECT 134.825 186.445 134.995 187.355 ;
        RECT 135.165 187.310 140.510 187.855 ;
        RECT 136.750 186.480 137.090 187.310 ;
        RECT 140.685 187.085 144.195 187.855 ;
        RECT 144.365 187.105 145.575 187.855 ;
        RECT 145.745 187.105 146.955 187.855 ;
        RECT 133.865 186.275 134.995 186.445 ;
        RECT 133.355 185.910 134.020 186.085 ;
        RECT 133.330 185.305 133.665 185.730 ;
        RECT 133.835 185.505 134.020 185.910 ;
        RECT 134.225 185.305 134.555 186.085 ;
        RECT 134.725 185.505 134.995 186.275 ;
        RECT 138.570 185.740 138.920 186.990 ;
        RECT 140.685 186.565 142.335 187.085 ;
        RECT 142.505 186.395 144.195 186.915 ;
        RECT 144.365 186.565 144.885 187.105 ;
        RECT 145.055 186.395 145.575 186.935 ;
        RECT 135.165 185.305 140.510 185.740 ;
        RECT 140.685 185.305 144.195 186.395 ;
        RECT 144.365 185.305 145.575 186.395 ;
        RECT 145.745 186.395 146.265 186.935 ;
        RECT 146.435 186.565 146.955 187.105 ;
        RECT 145.745 185.305 146.955 186.395 ;
        RECT 17.320 185.135 147.040 185.305 ;
        RECT 17.405 184.045 18.615 185.135 ;
        RECT 18.785 184.045 22.295 185.135 ;
        RECT 17.405 183.335 17.925 183.875 ;
        RECT 18.095 183.505 18.615 184.045 ;
        RECT 18.785 183.355 20.435 183.875 ;
        RECT 20.605 183.525 22.295 184.045 ;
        RECT 22.925 184.265 23.200 184.965 ;
        RECT 23.370 184.590 23.625 185.135 ;
        RECT 23.795 184.625 24.275 184.965 ;
        RECT 24.450 184.580 25.055 185.135 ;
        RECT 24.440 184.480 25.055 184.580 ;
        RECT 24.440 184.455 24.625 184.480 ;
        RECT 17.405 182.585 18.615 183.335 ;
        RECT 18.785 182.585 22.295 183.355 ;
        RECT 22.925 183.235 23.095 184.265 ;
        RECT 23.370 184.135 24.125 184.385 ;
        RECT 24.295 184.210 24.625 184.455 ;
        RECT 23.370 184.100 24.140 184.135 ;
        RECT 23.370 184.090 24.155 184.100 ;
        RECT 23.265 184.075 24.160 184.090 ;
        RECT 23.265 184.060 24.180 184.075 ;
        RECT 23.265 184.050 24.200 184.060 ;
        RECT 23.265 184.040 24.225 184.050 ;
        RECT 23.265 184.010 24.295 184.040 ;
        RECT 23.265 183.980 24.315 184.010 ;
        RECT 23.265 183.950 24.335 183.980 ;
        RECT 23.265 183.925 24.365 183.950 ;
        RECT 23.265 183.890 24.400 183.925 ;
        RECT 23.265 183.885 24.430 183.890 ;
        RECT 23.265 183.490 23.495 183.885 ;
        RECT 24.040 183.880 24.430 183.885 ;
        RECT 24.065 183.870 24.430 183.880 ;
        RECT 24.080 183.865 24.430 183.870 ;
        RECT 24.095 183.860 24.430 183.865 ;
        RECT 24.795 183.860 25.055 184.310 ;
        RECT 24.095 183.855 25.055 183.860 ;
        RECT 24.105 183.845 25.055 183.855 ;
        RECT 24.115 183.840 25.055 183.845 ;
        RECT 24.125 183.830 25.055 183.840 ;
        RECT 24.130 183.820 25.055 183.830 ;
        RECT 24.135 183.815 25.055 183.820 ;
        RECT 24.145 183.800 25.055 183.815 ;
        RECT 24.150 183.785 25.055 183.800 ;
        RECT 24.160 183.760 25.055 183.785 ;
        RECT 23.665 183.290 23.995 183.715 ;
        RECT 22.925 182.755 23.185 183.235 ;
        RECT 23.355 182.585 23.605 183.125 ;
        RECT 23.775 182.805 23.995 183.290 ;
        RECT 24.165 183.690 25.055 183.760 ;
        RECT 26.145 184.265 26.420 184.965 ;
        RECT 26.590 184.590 26.845 185.135 ;
        RECT 27.015 184.625 27.495 184.965 ;
        RECT 27.670 184.580 28.275 185.135 ;
        RECT 27.660 184.480 28.275 184.580 ;
        RECT 27.660 184.455 27.845 184.480 ;
        RECT 24.165 182.965 24.335 183.690 ;
        RECT 24.505 183.135 25.055 183.520 ;
        RECT 26.145 183.235 26.315 184.265 ;
        RECT 26.590 184.135 27.345 184.385 ;
        RECT 27.515 184.210 27.845 184.455 ;
        RECT 26.590 184.100 27.360 184.135 ;
        RECT 26.590 184.090 27.375 184.100 ;
        RECT 26.485 184.075 27.380 184.090 ;
        RECT 26.485 184.060 27.400 184.075 ;
        RECT 26.485 184.050 27.420 184.060 ;
        RECT 26.485 184.040 27.445 184.050 ;
        RECT 26.485 184.010 27.515 184.040 ;
        RECT 26.485 183.980 27.535 184.010 ;
        RECT 26.485 183.950 27.555 183.980 ;
        RECT 26.485 183.925 27.585 183.950 ;
        RECT 26.485 183.890 27.620 183.925 ;
        RECT 26.485 183.885 27.650 183.890 ;
        RECT 26.485 183.490 26.715 183.885 ;
        RECT 27.260 183.880 27.650 183.885 ;
        RECT 27.285 183.870 27.650 183.880 ;
        RECT 27.300 183.865 27.650 183.870 ;
        RECT 27.315 183.860 27.650 183.865 ;
        RECT 28.015 183.860 28.275 184.310 ;
        RECT 28.485 183.995 28.715 185.135 ;
        RECT 28.885 183.985 29.215 184.965 ;
        RECT 29.385 183.995 29.595 185.135 ;
        RECT 27.315 183.855 28.275 183.860 ;
        RECT 27.325 183.845 28.275 183.855 ;
        RECT 27.335 183.840 28.275 183.845 ;
        RECT 27.345 183.830 28.275 183.840 ;
        RECT 27.350 183.820 28.275 183.830 ;
        RECT 27.355 183.815 28.275 183.820 ;
        RECT 27.365 183.800 28.275 183.815 ;
        RECT 27.370 183.785 28.275 183.800 ;
        RECT 27.380 183.760 28.275 183.785 ;
        RECT 26.885 183.290 27.215 183.715 ;
        RECT 24.165 182.795 25.055 182.965 ;
        RECT 26.145 182.755 26.405 183.235 ;
        RECT 26.575 182.585 26.825 183.125 ;
        RECT 26.995 182.805 27.215 183.290 ;
        RECT 27.385 183.690 28.275 183.760 ;
        RECT 27.385 182.965 27.555 183.690 ;
        RECT 28.465 183.575 28.795 183.825 ;
        RECT 27.725 183.135 28.275 183.520 ;
        RECT 27.385 182.795 28.275 182.965 ;
        RECT 28.485 182.585 28.715 183.405 ;
        RECT 28.965 183.385 29.215 183.985 ;
        RECT 30.285 183.970 30.575 185.135 ;
        RECT 30.745 184.700 36.090 185.135 ;
        RECT 28.885 182.755 29.215 183.385 ;
        RECT 29.385 182.585 29.595 183.405 ;
        RECT 30.285 182.585 30.575 183.310 ;
        RECT 32.330 183.130 32.670 183.960 ;
        RECT 34.150 183.450 34.500 184.700 ;
        RECT 36.265 184.045 37.475 185.135 ;
        RECT 36.265 183.335 36.785 183.875 ;
        RECT 36.955 183.505 37.475 184.045 ;
        RECT 37.655 184.795 38.825 184.965 ;
        RECT 37.655 184.125 37.985 184.795 ;
        RECT 38.495 184.755 38.825 184.795 ;
        RECT 38.995 184.755 39.370 185.135 ;
        RECT 38.155 184.585 38.385 184.625 ;
        RECT 38.155 184.535 38.770 184.585 ;
        RECT 39.515 184.535 39.685 184.665 ;
        RECT 38.155 184.335 39.685 184.535 ;
        RECT 39.920 184.355 40.185 185.135 ;
        RECT 38.155 184.295 39.035 184.335 ;
        RECT 39.175 184.125 40.235 184.165 ;
        RECT 37.655 183.995 40.235 184.125 ;
        RECT 40.405 183.995 40.685 185.135 ;
        RECT 37.655 183.945 39.400 183.995 ;
        RECT 30.745 182.585 36.090 183.130 ;
        RECT 36.265 182.585 37.475 183.335 ;
        RECT 37.685 183.265 38.135 183.775 ;
        RECT 38.325 183.575 38.800 183.775 ;
        RECT 38.550 183.175 38.800 183.575 ;
        RECT 39.050 183.575 39.400 183.775 ;
        RECT 39.050 183.175 39.260 183.575 ;
        RECT 39.570 183.495 39.895 183.825 ;
        RECT 40.065 183.325 40.235 183.995 ;
        RECT 40.855 183.985 41.185 184.965 ;
        RECT 41.355 183.995 41.615 185.135 ;
        RECT 41.785 184.415 42.245 184.965 ;
        RECT 42.435 184.415 42.765 185.135 ;
        RECT 40.415 183.555 40.750 183.825 ;
        RECT 40.920 183.385 41.090 183.985 ;
        RECT 41.260 183.575 41.595 183.825 ;
        RECT 39.505 183.155 40.235 183.325 ;
        RECT 37.655 182.585 38.105 183.095 ;
        RECT 39.505 183.005 39.685 183.155 ;
        RECT 38.380 182.755 39.685 183.005 ;
        RECT 39.865 182.585 40.195 182.985 ;
        RECT 40.405 182.585 40.715 183.385 ;
        RECT 40.920 182.755 41.615 183.385 ;
        RECT 41.785 183.045 42.035 184.415 ;
        RECT 42.965 184.245 43.265 184.795 ;
        RECT 43.435 184.465 43.715 185.135 ;
        RECT 42.325 184.075 43.265 184.245 ;
        RECT 42.325 183.825 42.495 184.075 ;
        RECT 43.635 183.825 43.900 184.185 ;
        RECT 42.205 183.495 42.495 183.825 ;
        RECT 42.665 183.575 43.005 183.825 ;
        RECT 43.225 183.575 43.900 183.825 ;
        RECT 44.085 184.115 44.460 184.965 ;
        RECT 44.630 184.335 44.880 185.135 ;
        RECT 45.050 184.505 45.300 184.965 ;
        RECT 45.470 184.675 45.720 185.135 ;
        RECT 45.890 184.505 46.140 184.965 ;
        RECT 46.310 184.675 46.560 185.135 ;
        RECT 46.730 184.505 46.980 184.965 ;
        RECT 47.150 184.675 47.400 185.135 ;
        RECT 47.570 184.505 47.820 184.965 ;
        RECT 45.050 184.285 47.820 184.505 ;
        RECT 48.035 184.505 48.350 184.965 ;
        RECT 48.520 184.675 48.770 185.135 ;
        RECT 48.940 184.505 49.190 184.965 ;
        RECT 49.360 184.675 49.610 185.135 ;
        RECT 49.780 184.715 51.750 184.965 ;
        RECT 49.780 184.505 49.990 184.715 ;
        RECT 51.960 184.545 52.250 184.965 ;
        RECT 48.035 184.285 49.990 184.505 ;
        RECT 50.160 184.285 52.250 184.545 ;
        RECT 52.420 184.335 52.670 185.135 ;
        RECT 45.050 184.115 45.300 184.285 ;
        RECT 51.960 184.165 52.250 184.285 ;
        RECT 52.840 184.165 53.090 184.965 ;
        RECT 53.260 184.335 53.510 185.135 ;
        RECT 53.680 184.165 54.035 184.965 ;
        RECT 44.085 183.945 45.300 184.115 ;
        RECT 45.685 183.945 49.730 184.115 ;
        RECT 49.900 183.945 51.770 184.115 ;
        RECT 51.960 183.945 54.035 184.165 ;
        RECT 54.205 184.045 55.875 185.135 ;
        RECT 42.325 183.405 42.495 183.495 ;
        RECT 44.085 183.405 44.320 183.945 ;
        RECT 45.685 183.775 45.855 183.945 ;
        RECT 49.560 183.775 49.730 183.945 ;
        RECT 51.600 183.775 51.770 183.945 ;
        RECT 44.490 183.575 45.855 183.775 ;
        RECT 46.175 183.575 49.390 183.775 ;
        RECT 49.560 183.575 51.430 183.775 ;
        RECT 51.600 183.575 53.645 183.775 ;
        RECT 53.815 183.405 54.035 183.945 ;
        RECT 42.325 183.215 43.715 183.405 ;
        RECT 41.785 182.755 42.345 183.045 ;
        RECT 42.515 182.585 42.765 183.045 ;
        RECT 43.385 182.855 43.715 183.215 ;
        RECT 44.085 183.145 45.760 183.405 ;
        RECT 45.930 183.225 47.860 183.405 ;
        RECT 45.930 182.975 46.180 183.225 ;
        RECT 44.170 182.755 46.180 182.975 ;
        RECT 46.350 182.585 46.520 183.055 ;
        RECT 46.690 182.755 47.020 183.225 ;
        RECT 47.190 182.585 47.360 183.055 ;
        RECT 47.530 182.755 47.860 183.225 ;
        RECT 48.035 182.585 48.310 183.405 ;
        RECT 48.480 183.235 52.210 183.405 ;
        RECT 48.480 183.225 51.430 183.235 ;
        RECT 48.480 182.755 48.810 183.225 ;
        RECT 48.980 182.585 49.150 183.055 ;
        RECT 49.320 182.755 49.650 183.225 ;
        RECT 49.820 182.585 49.990 183.055 ;
        RECT 50.160 182.755 50.490 183.225 ;
        RECT 50.660 182.585 50.830 183.055 ;
        RECT 51.000 182.755 51.330 183.225 ;
        RECT 51.500 182.585 51.770 183.055 ;
        RECT 51.960 182.975 52.210 183.235 ;
        RECT 52.380 183.145 54.035 183.405 ;
        RECT 54.205 183.355 54.955 183.875 ;
        RECT 55.125 183.525 55.875 184.045 ;
        RECT 56.045 183.970 56.335 185.135 ;
        RECT 56.510 184.745 56.845 184.965 ;
        RECT 57.850 184.755 58.205 185.135 ;
        RECT 56.510 184.125 56.765 184.745 ;
        RECT 57.015 184.585 57.245 184.625 ;
        RECT 58.375 184.585 58.625 184.965 ;
        RECT 57.015 184.385 58.625 184.585 ;
        RECT 57.015 184.295 57.200 184.385 ;
        RECT 57.790 184.375 58.625 184.385 ;
        RECT 58.875 184.355 59.125 185.135 ;
        RECT 59.295 184.285 59.555 184.965 ;
        RECT 57.355 184.185 57.685 184.215 ;
        RECT 57.355 184.125 59.155 184.185 ;
        RECT 56.510 184.015 59.215 184.125 ;
        RECT 56.510 183.955 57.685 184.015 ;
        RECT 59.015 183.980 59.215 184.015 ;
        RECT 56.505 183.575 56.995 183.775 ;
        RECT 57.185 183.575 57.660 183.785 ;
        RECT 51.960 182.805 53.970 182.975 ;
        RECT 54.205 182.585 55.875 183.355 ;
        RECT 56.045 182.585 56.335 183.310 ;
        RECT 56.510 182.585 56.965 183.350 ;
        RECT 57.440 183.175 57.660 183.575 ;
        RECT 57.905 183.575 58.235 183.785 ;
        RECT 57.905 183.175 58.115 183.575 ;
        RECT 58.405 183.540 58.815 183.845 ;
        RECT 59.045 183.405 59.215 183.980 ;
        RECT 58.945 183.285 59.215 183.405 ;
        RECT 58.370 183.240 59.215 183.285 ;
        RECT 58.370 183.115 59.125 183.240 ;
        RECT 58.370 182.965 58.540 183.115 ;
        RECT 59.385 183.085 59.555 184.285 ;
        RECT 57.240 182.755 58.540 182.965 ;
        RECT 58.795 182.585 59.125 182.945 ;
        RECT 59.295 182.755 59.555 183.085 ;
        RECT 59.725 184.415 60.185 184.965 ;
        RECT 60.375 184.415 60.705 185.135 ;
        RECT 59.725 183.045 59.975 184.415 ;
        RECT 60.905 184.245 61.205 184.795 ;
        RECT 61.375 184.465 61.655 185.135 ;
        RECT 62.025 184.700 67.370 185.135 ;
        RECT 60.265 184.075 61.205 184.245 ;
        RECT 60.265 183.825 60.435 184.075 ;
        RECT 61.575 183.825 61.840 184.185 ;
        RECT 60.145 183.495 60.435 183.825 ;
        RECT 60.605 183.575 60.945 183.825 ;
        RECT 61.165 183.575 61.840 183.825 ;
        RECT 60.265 183.405 60.435 183.495 ;
        RECT 60.265 183.215 61.655 183.405 ;
        RECT 59.725 182.755 60.285 183.045 ;
        RECT 60.455 182.585 60.705 183.045 ;
        RECT 61.325 182.855 61.655 183.215 ;
        RECT 63.610 183.130 63.950 183.960 ;
        RECT 65.430 183.450 65.780 184.700 ;
        RECT 67.545 184.045 71.055 185.135 ;
        RECT 71.225 184.045 72.435 185.135 ;
        RECT 72.605 184.625 72.905 185.135 ;
        RECT 73.075 184.455 73.405 184.965 ;
        RECT 73.575 184.625 74.205 185.135 ;
        RECT 74.785 184.625 75.165 184.795 ;
        RECT 75.335 184.625 75.635 185.135 ;
        RECT 74.995 184.455 75.165 184.625 ;
        RECT 67.545 183.355 69.195 183.875 ;
        RECT 69.365 183.525 71.055 184.045 ;
        RECT 62.025 182.585 67.370 183.130 ;
        RECT 67.545 182.585 71.055 183.355 ;
        RECT 71.225 183.335 71.745 183.875 ;
        RECT 71.915 183.505 72.435 184.045 ;
        RECT 72.605 184.285 74.825 184.455 ;
        RECT 71.225 182.585 72.435 183.335 ;
        RECT 72.605 183.325 72.775 184.285 ;
        RECT 72.945 183.945 74.485 184.115 ;
        RECT 72.945 183.495 73.190 183.945 ;
        RECT 73.450 183.575 74.145 183.775 ;
        RECT 74.315 183.745 74.485 183.945 ;
        RECT 74.655 184.085 74.825 184.285 ;
        RECT 74.995 184.255 75.655 184.455 ;
        RECT 76.995 184.405 77.290 185.135 ;
        RECT 74.655 183.915 75.315 184.085 ;
        RECT 74.315 183.575 74.915 183.745 ;
        RECT 75.145 183.495 75.315 183.915 ;
        RECT 72.605 182.780 73.070 183.325 ;
        RECT 73.575 182.585 73.745 183.405 ;
        RECT 73.915 183.325 74.825 183.405 ;
        RECT 75.485 183.325 75.655 184.255 ;
        RECT 77.460 184.235 77.720 184.960 ;
        RECT 77.890 184.405 78.150 185.135 ;
        RECT 78.320 184.235 78.580 184.960 ;
        RECT 78.750 184.405 79.010 185.135 ;
        RECT 79.180 184.235 79.440 184.960 ;
        RECT 79.610 184.405 79.870 185.135 ;
        RECT 80.040 184.235 80.300 184.960 ;
        RECT 73.915 183.235 75.165 183.325 ;
        RECT 73.915 182.755 74.245 183.235 ;
        RECT 74.655 183.155 75.165 183.235 ;
        RECT 74.415 182.585 74.765 182.975 ;
        RECT 74.935 182.755 75.165 183.155 ;
        RECT 75.335 182.845 75.655 183.325 ;
        RECT 76.990 183.995 80.300 184.235 ;
        RECT 80.470 184.025 80.730 185.135 ;
        RECT 76.990 183.405 77.960 183.995 ;
        RECT 80.900 183.825 81.150 184.960 ;
        RECT 81.330 184.025 81.625 185.135 ;
        RECT 81.805 183.970 82.095 185.135 ;
        RECT 82.265 184.700 87.610 185.135 ;
        RECT 78.130 183.575 81.150 183.825 ;
        RECT 76.990 183.235 80.300 183.405 ;
        RECT 76.990 182.585 77.290 183.065 ;
        RECT 77.460 182.780 77.720 183.235 ;
        RECT 77.890 182.585 78.150 183.065 ;
        RECT 78.320 182.780 78.580 183.235 ;
        RECT 78.750 182.585 79.010 183.065 ;
        RECT 79.180 182.780 79.440 183.235 ;
        RECT 79.610 182.585 79.870 183.065 ;
        RECT 80.040 182.780 80.300 183.235 ;
        RECT 80.470 182.585 80.730 183.110 ;
        RECT 80.900 182.765 81.150 183.575 ;
        RECT 81.320 183.215 81.635 183.825 ;
        RECT 81.330 182.585 81.575 183.045 ;
        RECT 81.805 182.585 82.095 183.310 ;
        RECT 83.850 183.130 84.190 183.960 ;
        RECT 85.670 183.450 86.020 184.700 ;
        RECT 87.785 184.045 91.295 185.135 ;
        RECT 87.785 183.355 89.435 183.875 ;
        RECT 89.605 183.525 91.295 184.045 ;
        RECT 91.465 183.995 91.850 184.965 ;
        RECT 92.020 184.675 92.345 185.135 ;
        RECT 92.865 184.505 93.145 184.965 ;
        RECT 92.020 184.285 93.145 184.505 ;
        RECT 82.265 182.585 87.610 183.130 ;
        RECT 87.785 182.585 91.295 183.355 ;
        RECT 91.465 183.325 91.745 183.995 ;
        RECT 92.020 183.825 92.470 184.285 ;
        RECT 93.335 184.115 93.735 184.965 ;
        RECT 94.135 184.675 94.405 185.135 ;
        RECT 94.575 184.505 94.860 184.965 ;
        RECT 91.915 183.495 92.470 183.825 ;
        RECT 92.640 183.555 93.735 184.115 ;
        RECT 92.020 183.385 92.470 183.495 ;
        RECT 91.465 182.755 91.850 183.325 ;
        RECT 92.020 183.215 93.145 183.385 ;
        RECT 92.020 182.585 92.345 183.045 ;
        RECT 92.865 182.755 93.145 183.215 ;
        RECT 93.335 182.755 93.735 183.555 ;
        RECT 93.905 184.285 94.860 184.505 ;
        RECT 95.235 184.465 95.405 184.965 ;
        RECT 95.575 184.635 95.905 185.135 ;
        RECT 95.235 184.295 95.900 184.465 ;
        RECT 93.905 183.385 94.115 184.285 ;
        RECT 94.285 183.555 94.975 184.115 ;
        RECT 95.150 183.475 95.500 184.125 ;
        RECT 93.905 183.215 94.860 183.385 ;
        RECT 95.670 183.305 95.900 184.295 ;
        RECT 94.135 182.585 94.405 183.045 ;
        RECT 94.575 182.755 94.860 183.215 ;
        RECT 95.235 183.135 95.900 183.305 ;
        RECT 95.235 182.845 95.405 183.135 ;
        RECT 95.575 182.585 95.905 182.965 ;
        RECT 96.075 182.845 96.260 184.965 ;
        RECT 96.500 184.675 96.765 185.135 ;
        RECT 96.935 184.540 97.185 184.965 ;
        RECT 97.395 184.690 98.500 184.860 ;
        RECT 96.880 184.410 97.185 184.540 ;
        RECT 96.430 183.215 96.710 184.165 ;
        RECT 96.880 183.305 97.050 184.410 ;
        RECT 97.220 183.625 97.460 184.220 ;
        RECT 97.630 184.155 98.160 184.520 ;
        RECT 97.630 183.455 97.800 184.155 ;
        RECT 98.330 184.075 98.500 184.690 ;
        RECT 98.670 184.335 98.840 185.135 ;
        RECT 99.010 184.635 99.260 184.965 ;
        RECT 99.485 184.665 100.370 184.835 ;
        RECT 98.330 183.985 98.840 184.075 ;
        RECT 96.880 183.175 97.105 183.305 ;
        RECT 97.275 183.235 97.800 183.455 ;
        RECT 97.970 183.815 98.840 183.985 ;
        RECT 96.515 182.585 96.765 183.045 ;
        RECT 96.935 183.035 97.105 183.175 ;
        RECT 97.970 183.035 98.140 183.815 ;
        RECT 98.670 183.745 98.840 183.815 ;
        RECT 98.350 183.565 98.550 183.595 ;
        RECT 99.010 183.565 99.180 184.635 ;
        RECT 99.350 183.745 99.540 184.465 ;
        RECT 98.350 183.265 99.180 183.565 ;
        RECT 99.710 183.535 100.030 184.495 ;
        RECT 96.935 182.865 97.270 183.035 ;
        RECT 97.465 182.865 98.140 183.035 ;
        RECT 98.460 182.585 98.830 183.085 ;
        RECT 99.010 183.035 99.180 183.265 ;
        RECT 99.565 183.205 100.030 183.535 ;
        RECT 100.200 183.825 100.370 184.665 ;
        RECT 100.550 184.635 100.865 185.135 ;
        RECT 101.095 184.405 101.435 184.965 ;
        RECT 100.540 184.030 101.435 184.405 ;
        RECT 101.605 184.125 101.775 185.135 ;
        RECT 101.245 183.825 101.435 184.030 ;
        RECT 101.945 184.075 102.275 184.920 ;
        RECT 101.945 183.995 102.335 184.075 ;
        RECT 102.120 183.945 102.335 183.995 ;
        RECT 100.200 183.495 101.075 183.825 ;
        RECT 101.245 183.495 101.995 183.825 ;
        RECT 100.200 183.035 100.370 183.495 ;
        RECT 101.245 183.325 101.445 183.495 ;
        RECT 102.165 183.365 102.335 183.945 ;
        RECT 102.110 183.325 102.335 183.365 ;
        RECT 99.010 182.865 99.415 183.035 ;
        RECT 99.585 182.865 100.370 183.035 ;
        RECT 100.645 182.585 100.855 183.115 ;
        RECT 101.115 182.800 101.445 183.325 ;
        RECT 101.955 183.240 102.335 183.325 ;
        RECT 102.510 183.995 102.845 184.965 ;
        RECT 103.015 183.995 103.185 185.135 ;
        RECT 103.355 184.795 105.385 184.965 ;
        RECT 102.510 183.325 102.680 183.995 ;
        RECT 103.355 183.825 103.525 184.795 ;
        RECT 102.850 183.495 103.105 183.825 ;
        RECT 103.330 183.495 103.525 183.825 ;
        RECT 103.695 184.455 104.820 184.625 ;
        RECT 102.935 183.325 103.105 183.495 ;
        RECT 103.695 183.325 103.865 184.455 ;
        RECT 101.615 182.585 101.785 183.195 ;
        RECT 101.955 182.805 102.285 183.240 ;
        RECT 102.510 182.755 102.765 183.325 ;
        RECT 102.935 183.155 103.865 183.325 ;
        RECT 104.035 184.115 105.045 184.285 ;
        RECT 104.035 183.315 104.205 184.115 ;
        RECT 104.410 183.435 104.685 183.915 ;
        RECT 104.405 183.265 104.685 183.435 ;
        RECT 103.690 183.120 103.865 183.155 ;
        RECT 102.935 182.585 103.265 182.985 ;
        RECT 103.690 182.755 104.220 183.120 ;
        RECT 104.410 182.755 104.685 183.265 ;
        RECT 104.855 182.755 105.045 184.115 ;
        RECT 105.215 184.130 105.385 184.795 ;
        RECT 105.555 184.375 105.725 185.135 ;
        RECT 105.960 184.375 106.475 184.785 ;
        RECT 105.215 183.940 105.965 184.130 ;
        RECT 106.135 183.565 106.475 184.375 ;
        RECT 107.565 183.970 107.855 185.135 ;
        RECT 108.115 184.465 108.285 184.965 ;
        RECT 108.455 184.635 108.785 185.135 ;
        RECT 108.115 184.295 108.780 184.465 ;
        RECT 105.245 183.395 106.475 183.565 ;
        RECT 108.030 183.475 108.380 184.125 ;
        RECT 105.225 182.585 105.735 183.120 ;
        RECT 105.955 182.790 106.200 183.395 ;
        RECT 107.565 182.585 107.855 183.310 ;
        RECT 108.550 183.305 108.780 184.295 ;
        RECT 108.115 183.135 108.780 183.305 ;
        RECT 108.115 182.845 108.285 183.135 ;
        RECT 108.455 182.585 108.785 182.965 ;
        RECT 108.955 182.845 109.140 184.965 ;
        RECT 109.380 184.675 109.645 185.135 ;
        RECT 109.815 184.540 110.065 184.965 ;
        RECT 110.275 184.690 111.380 184.860 ;
        RECT 109.760 184.410 110.065 184.540 ;
        RECT 109.310 183.215 109.590 184.165 ;
        RECT 109.760 183.305 109.930 184.410 ;
        RECT 110.100 183.625 110.340 184.220 ;
        RECT 110.510 184.155 111.040 184.520 ;
        RECT 110.510 183.455 110.680 184.155 ;
        RECT 111.210 184.075 111.380 184.690 ;
        RECT 111.550 184.335 111.720 185.135 ;
        RECT 111.890 184.635 112.140 184.965 ;
        RECT 112.365 184.665 113.250 184.835 ;
        RECT 111.210 183.985 111.720 184.075 ;
        RECT 109.760 183.175 109.985 183.305 ;
        RECT 110.155 183.235 110.680 183.455 ;
        RECT 110.850 183.815 111.720 183.985 ;
        RECT 109.395 182.585 109.645 183.045 ;
        RECT 109.815 183.035 109.985 183.175 ;
        RECT 110.850 183.035 111.020 183.815 ;
        RECT 111.550 183.745 111.720 183.815 ;
        RECT 111.230 183.565 111.430 183.595 ;
        RECT 111.890 183.565 112.060 184.635 ;
        RECT 112.230 183.745 112.420 184.465 ;
        RECT 111.230 183.265 112.060 183.565 ;
        RECT 112.590 183.535 112.910 184.495 ;
        RECT 109.815 182.865 110.150 183.035 ;
        RECT 110.345 182.865 111.020 183.035 ;
        RECT 111.340 182.585 111.710 183.085 ;
        RECT 111.890 183.035 112.060 183.265 ;
        RECT 112.445 183.205 112.910 183.535 ;
        RECT 113.080 183.825 113.250 184.665 ;
        RECT 113.430 184.635 113.745 185.135 ;
        RECT 113.975 184.405 114.315 184.965 ;
        RECT 113.420 184.030 114.315 184.405 ;
        RECT 114.485 184.125 114.655 185.135 ;
        RECT 114.125 183.825 114.315 184.030 ;
        RECT 114.825 184.075 115.155 184.920 ;
        RECT 114.825 183.995 115.215 184.075 ;
        RECT 115.385 184.045 117.975 185.135 ;
        RECT 115.000 183.945 115.215 183.995 ;
        RECT 113.080 183.495 113.955 183.825 ;
        RECT 114.125 183.495 114.875 183.825 ;
        RECT 113.080 183.035 113.250 183.495 ;
        RECT 114.125 183.325 114.325 183.495 ;
        RECT 115.045 183.365 115.215 183.945 ;
        RECT 114.990 183.325 115.215 183.365 ;
        RECT 111.890 182.865 112.295 183.035 ;
        RECT 112.465 182.865 113.250 183.035 ;
        RECT 113.525 182.585 113.735 183.115 ;
        RECT 113.995 182.800 114.325 183.325 ;
        RECT 114.835 183.240 115.215 183.325 ;
        RECT 115.385 183.355 116.595 183.875 ;
        RECT 116.765 183.525 117.975 184.045 ;
        RECT 118.150 183.995 118.485 184.965 ;
        RECT 118.655 183.995 118.825 185.135 ;
        RECT 118.995 184.795 121.025 184.965 ;
        RECT 114.495 182.585 114.665 183.195 ;
        RECT 114.835 182.805 115.165 183.240 ;
        RECT 115.385 182.585 117.975 183.355 ;
        RECT 118.150 183.325 118.320 183.995 ;
        RECT 118.995 183.825 119.165 184.795 ;
        RECT 118.490 183.495 118.745 183.825 ;
        RECT 118.970 183.495 119.165 183.825 ;
        RECT 119.335 184.455 120.460 184.625 ;
        RECT 118.575 183.325 118.745 183.495 ;
        RECT 119.335 183.325 119.505 184.455 ;
        RECT 118.150 182.755 118.405 183.325 ;
        RECT 118.575 183.155 119.505 183.325 ;
        RECT 119.675 184.115 120.685 184.285 ;
        RECT 119.675 183.315 119.845 184.115 ;
        RECT 119.330 183.120 119.505 183.155 ;
        RECT 118.575 182.585 118.905 182.985 ;
        RECT 119.330 182.755 119.860 183.120 ;
        RECT 120.050 183.095 120.325 183.915 ;
        RECT 120.045 182.925 120.325 183.095 ;
        RECT 120.050 182.755 120.325 182.925 ;
        RECT 120.495 182.755 120.685 184.115 ;
        RECT 120.855 184.130 121.025 184.795 ;
        RECT 121.195 184.375 121.365 185.135 ;
        RECT 121.600 184.375 122.115 184.785 ;
        RECT 120.855 183.940 121.605 184.130 ;
        RECT 121.775 183.565 122.115 184.375 ;
        RECT 122.400 184.505 122.685 184.965 ;
        RECT 122.855 184.675 123.125 185.135 ;
        RECT 122.400 184.285 123.355 184.505 ;
        RECT 120.885 183.395 122.115 183.565 ;
        RECT 122.285 183.555 122.975 184.115 ;
        RECT 120.865 182.585 121.375 183.120 ;
        RECT 121.595 182.790 121.840 183.395 ;
        RECT 123.145 183.385 123.355 184.285 ;
        RECT 122.400 183.215 123.355 183.385 ;
        RECT 123.525 184.115 123.925 184.965 ;
        RECT 124.115 184.505 124.395 184.965 ;
        RECT 124.915 184.675 125.240 185.135 ;
        RECT 124.115 184.285 125.240 184.505 ;
        RECT 123.525 183.555 124.620 184.115 ;
        RECT 124.790 183.825 125.240 184.285 ;
        RECT 125.410 183.995 125.795 184.965 ;
        RECT 125.965 184.045 127.175 185.135 ;
        RECT 127.460 184.505 127.745 184.965 ;
        RECT 127.915 184.675 128.185 185.135 ;
        RECT 127.460 184.285 128.415 184.505 ;
        RECT 122.400 182.755 122.685 183.215 ;
        RECT 122.855 182.585 123.125 183.045 ;
        RECT 123.525 182.755 123.925 183.555 ;
        RECT 124.790 183.495 125.345 183.825 ;
        RECT 124.790 183.385 125.240 183.495 ;
        RECT 124.115 183.215 125.240 183.385 ;
        RECT 125.515 183.325 125.795 183.995 ;
        RECT 124.115 182.755 124.395 183.215 ;
        RECT 124.915 182.585 125.240 183.045 ;
        RECT 125.410 182.755 125.795 183.325 ;
        RECT 125.965 183.335 126.485 183.875 ;
        RECT 126.655 183.505 127.175 184.045 ;
        RECT 127.345 183.555 128.035 184.115 ;
        RECT 128.205 183.385 128.415 184.285 ;
        RECT 125.965 182.585 127.175 183.335 ;
        RECT 127.460 183.215 128.415 183.385 ;
        RECT 128.585 184.115 128.985 184.965 ;
        RECT 129.175 184.505 129.455 184.965 ;
        RECT 129.975 184.675 130.300 185.135 ;
        RECT 129.175 184.285 130.300 184.505 ;
        RECT 128.585 183.555 129.680 184.115 ;
        RECT 129.850 183.825 130.300 184.285 ;
        RECT 130.470 183.995 130.855 184.965 ;
        RECT 131.115 184.205 131.285 184.965 ;
        RECT 131.500 184.375 131.830 185.135 ;
        RECT 131.115 184.035 131.830 184.205 ;
        RECT 132.000 184.060 132.255 184.965 ;
        RECT 127.460 182.755 127.745 183.215 ;
        RECT 127.915 182.585 128.185 183.045 ;
        RECT 128.585 182.755 128.985 183.555 ;
        RECT 129.850 183.495 130.405 183.825 ;
        RECT 129.850 183.385 130.300 183.495 ;
        RECT 129.175 183.215 130.300 183.385 ;
        RECT 130.575 183.325 130.855 183.995 ;
        RECT 131.025 183.485 131.380 183.855 ;
        RECT 131.660 183.825 131.830 184.035 ;
        RECT 131.660 183.495 131.915 183.825 ;
        RECT 129.175 182.755 129.455 183.215 ;
        RECT 129.975 182.585 130.300 183.045 ;
        RECT 130.470 182.755 130.855 183.325 ;
        RECT 131.660 183.305 131.830 183.495 ;
        RECT 132.085 183.330 132.255 184.060 ;
        RECT 132.430 183.985 132.690 185.135 ;
        RECT 133.325 183.970 133.615 185.135 ;
        RECT 133.785 184.285 134.045 184.965 ;
        RECT 134.215 184.355 134.465 185.135 ;
        RECT 134.715 184.585 134.965 184.965 ;
        RECT 135.135 184.755 135.490 185.135 ;
        RECT 136.495 184.745 136.830 184.965 ;
        RECT 136.095 184.585 136.325 184.625 ;
        RECT 134.715 184.385 136.325 184.585 ;
        RECT 134.715 184.375 135.550 184.385 ;
        RECT 136.140 184.295 136.325 184.385 ;
        RECT 131.115 183.135 131.830 183.305 ;
        RECT 131.115 182.755 131.285 183.135 ;
        RECT 131.500 182.585 131.830 182.965 ;
        RECT 132.000 182.755 132.255 183.330 ;
        RECT 132.430 182.585 132.690 183.425 ;
        RECT 133.325 182.585 133.615 183.310 ;
        RECT 133.785 183.085 133.955 184.285 ;
        RECT 135.655 184.185 135.985 184.215 ;
        RECT 134.185 184.125 135.985 184.185 ;
        RECT 136.575 184.125 136.830 184.745 ;
        RECT 137.005 184.700 142.350 185.135 ;
        RECT 134.125 184.015 136.830 184.125 ;
        RECT 134.125 183.980 134.325 184.015 ;
        RECT 134.125 183.405 134.295 183.980 ;
        RECT 135.655 183.955 136.830 184.015 ;
        RECT 134.525 183.540 134.935 183.845 ;
        RECT 135.105 183.575 135.435 183.785 ;
        RECT 134.125 183.285 134.395 183.405 ;
        RECT 134.125 183.240 134.970 183.285 ;
        RECT 134.215 183.115 134.970 183.240 ;
        RECT 135.225 183.175 135.435 183.575 ;
        RECT 135.680 183.575 136.155 183.785 ;
        RECT 136.345 183.575 136.835 183.775 ;
        RECT 135.680 183.175 135.900 183.575 ;
        RECT 133.785 182.755 134.045 183.085 ;
        RECT 134.800 182.965 134.970 183.115 ;
        RECT 134.215 182.585 134.545 182.945 ;
        RECT 134.800 182.755 136.100 182.965 ;
        RECT 136.375 182.585 136.830 183.350 ;
        RECT 138.590 183.130 138.930 183.960 ;
        RECT 140.410 183.450 140.760 184.700 ;
        RECT 142.525 184.045 145.115 185.135 ;
        RECT 142.525 183.355 143.735 183.875 ;
        RECT 143.905 183.525 145.115 184.045 ;
        RECT 145.745 184.045 146.955 185.135 ;
        RECT 145.745 183.505 146.265 184.045 ;
        RECT 137.005 182.585 142.350 183.130 ;
        RECT 142.525 182.585 145.115 183.355 ;
        RECT 146.435 183.335 146.955 183.875 ;
        RECT 145.745 182.585 146.955 183.335 ;
        RECT 17.320 182.415 147.040 182.585 ;
        RECT 17.405 181.665 18.615 182.415 ;
        RECT 18.785 181.870 24.130 182.415 ;
        RECT 17.405 181.125 17.925 181.665 ;
        RECT 18.095 180.955 18.615 181.495 ;
        RECT 20.370 181.040 20.710 181.870 ;
        RECT 24.765 181.615 25.075 182.415 ;
        RECT 25.280 181.615 25.975 182.245 ;
        RECT 26.145 181.870 31.490 182.415 ;
        RECT 17.405 179.865 18.615 180.955 ;
        RECT 22.190 180.300 22.540 181.550 ;
        RECT 24.775 181.175 25.110 181.445 ;
        RECT 25.280 181.015 25.450 181.615 ;
        RECT 25.620 181.175 25.955 181.425 ;
        RECT 27.730 181.040 28.070 181.870 ;
        RECT 31.665 181.645 35.175 182.415 ;
        RECT 18.785 179.865 24.130 180.300 ;
        RECT 24.765 179.865 25.045 181.005 ;
        RECT 25.215 180.035 25.545 181.015 ;
        RECT 25.715 179.865 25.975 181.005 ;
        RECT 29.550 180.300 29.900 181.550 ;
        RECT 31.665 181.125 33.315 181.645 ;
        RECT 35.550 181.635 36.050 182.245 ;
        RECT 33.485 180.955 35.175 181.475 ;
        RECT 35.345 181.175 35.695 181.425 ;
        RECT 35.880 181.005 36.050 181.635 ;
        RECT 36.680 181.765 37.010 182.245 ;
        RECT 37.180 181.955 37.405 182.415 ;
        RECT 37.575 181.765 37.905 182.245 ;
        RECT 36.680 181.595 37.905 181.765 ;
        RECT 38.095 181.615 38.345 182.415 ;
        RECT 38.515 181.615 38.855 182.245 ;
        RECT 39.230 181.635 39.730 182.245 ;
        RECT 38.625 181.565 38.855 181.615 ;
        RECT 36.220 181.225 36.550 181.425 ;
        RECT 36.720 181.225 37.050 181.425 ;
        RECT 37.220 181.225 37.640 181.425 ;
        RECT 37.815 181.255 38.510 181.425 ;
        RECT 37.815 181.005 37.985 181.255 ;
        RECT 38.680 181.005 38.855 181.565 ;
        RECT 39.025 181.175 39.375 181.425 ;
        RECT 39.560 181.005 39.730 181.635 ;
        RECT 40.360 181.765 40.690 182.245 ;
        RECT 40.860 181.955 41.085 182.415 ;
        RECT 41.255 181.765 41.585 182.245 ;
        RECT 40.360 181.595 41.585 181.765 ;
        RECT 41.775 181.615 42.025 182.415 ;
        RECT 42.195 181.615 42.535 182.245 ;
        RECT 43.165 181.690 43.455 182.415 ;
        RECT 43.685 181.955 43.930 182.415 ;
        RECT 39.900 181.225 40.230 181.425 ;
        RECT 40.400 181.225 40.730 181.425 ;
        RECT 40.900 181.225 41.320 181.425 ;
        RECT 41.495 181.255 42.190 181.425 ;
        RECT 41.495 181.005 41.665 181.255 ;
        RECT 42.360 181.005 42.535 181.615 ;
        RECT 43.625 181.175 43.940 181.785 ;
        RECT 44.110 181.425 44.360 182.235 ;
        RECT 44.530 181.890 44.790 182.415 ;
        RECT 44.960 181.765 45.220 182.220 ;
        RECT 45.390 181.935 45.650 182.415 ;
        RECT 45.820 181.765 46.080 182.220 ;
        RECT 46.250 181.935 46.510 182.415 ;
        RECT 46.680 181.765 46.940 182.220 ;
        RECT 47.110 181.935 47.370 182.415 ;
        RECT 47.540 181.765 47.800 182.220 ;
        RECT 47.970 181.935 48.270 182.415 ;
        RECT 48.730 181.955 48.995 182.415 ;
        RECT 49.365 181.775 49.535 182.245 ;
        RECT 49.785 181.955 49.955 182.415 ;
        RECT 50.205 181.775 50.375 182.245 ;
        RECT 50.625 181.955 50.795 182.415 ;
        RECT 51.045 181.775 51.215 182.245 ;
        RECT 51.385 181.950 51.635 182.415 ;
        RECT 44.960 181.595 48.270 181.765 ;
        RECT 49.365 181.595 51.735 181.775 ;
        RECT 52.575 181.725 52.905 182.415 ;
        RECT 53.365 181.820 53.985 182.245 ;
        RECT 54.155 181.925 54.485 182.415 ;
        RECT 44.110 181.175 47.130 181.425 ;
        RECT 26.145 179.865 31.490 180.300 ;
        RECT 31.665 179.865 35.175 180.955 ;
        RECT 35.550 180.835 37.985 181.005 ;
        RECT 35.550 180.035 35.880 180.835 ;
        RECT 36.050 179.865 36.380 180.665 ;
        RECT 36.680 180.035 37.010 180.835 ;
        RECT 37.655 179.865 37.905 180.665 ;
        RECT 38.175 179.865 38.345 181.005 ;
        RECT 38.515 180.035 38.855 181.005 ;
        RECT 39.230 180.835 41.665 181.005 ;
        RECT 39.230 180.035 39.560 180.835 ;
        RECT 39.730 179.865 40.060 180.665 ;
        RECT 40.360 180.035 40.690 180.835 ;
        RECT 41.335 179.865 41.585 180.665 ;
        RECT 41.855 179.865 42.025 181.005 ;
        RECT 42.195 180.035 42.535 181.005 ;
        RECT 43.165 179.865 43.455 181.030 ;
        RECT 43.635 179.865 43.930 180.975 ;
        RECT 44.110 180.040 44.360 181.175 ;
        RECT 47.300 181.005 48.270 181.595 ;
        RECT 48.705 181.175 51.215 181.425 ;
        RECT 51.385 181.005 51.735 181.595 ;
        RECT 53.625 181.485 53.985 181.820 ;
        RECT 52.565 181.205 53.985 181.485 ;
        RECT 44.530 179.865 44.790 180.975 ;
        RECT 44.960 180.765 48.270 181.005 ;
        RECT 44.960 180.040 45.220 180.765 ;
        RECT 45.390 179.865 45.650 180.595 ;
        RECT 45.820 180.040 46.080 180.765 ;
        RECT 46.250 179.865 46.510 180.595 ;
        RECT 46.680 180.040 46.940 180.765 ;
        RECT 47.110 179.865 47.370 180.595 ;
        RECT 47.540 180.040 47.800 180.765 ;
        RECT 47.970 179.865 48.265 180.595 ;
        RECT 48.730 179.865 49.025 181.005 ;
        RECT 49.285 180.835 51.735 181.005 ;
        RECT 49.285 180.035 49.615 180.835 ;
        RECT 49.785 179.865 49.955 180.665 ;
        RECT 50.125 180.035 50.455 180.835 ;
        RECT 50.965 180.815 51.735 180.835 ;
        RECT 50.625 179.865 50.795 180.665 ;
        RECT 50.965 180.035 51.295 180.815 ;
        RECT 51.465 179.865 51.635 180.325 ;
        RECT 52.035 179.865 52.365 181.035 ;
        RECT 52.565 180.035 52.895 181.205 ;
        RECT 53.095 179.865 53.425 181.035 ;
        RECT 53.625 180.035 53.985 181.205 ;
        RECT 54.155 181.175 54.495 181.755 ;
        RECT 54.665 181.645 56.335 182.415 ;
        RECT 54.665 181.125 55.415 181.645 ;
        RECT 56.545 181.595 56.775 182.415 ;
        RECT 56.945 181.615 57.275 182.245 ;
        RECT 54.155 179.865 54.485 181.005 ;
        RECT 55.585 180.955 56.335 181.475 ;
        RECT 56.525 181.175 56.855 181.425 ;
        RECT 57.025 181.015 57.275 181.615 ;
        RECT 57.445 181.595 57.655 182.415 ;
        RECT 57.910 182.015 58.240 182.415 ;
        RECT 58.410 181.845 58.580 182.115 ;
        RECT 58.750 181.905 59.065 182.415 ;
        RECT 59.295 181.905 59.585 182.245 ;
        RECT 59.755 181.905 59.995 182.415 ;
        RECT 60.655 181.915 60.985 182.415 ;
        RECT 57.885 181.675 58.580 181.845 ;
        RECT 54.665 179.865 56.335 180.955 ;
        RECT 56.545 179.865 56.775 181.005 ;
        RECT 56.945 180.035 57.275 181.015 ;
        RECT 57.445 179.865 57.655 181.005 ;
        RECT 57.885 180.665 58.315 181.675 ;
        RECT 58.485 181.005 58.655 181.505 ;
        RECT 58.825 181.175 59.235 181.735 ;
        RECT 59.405 181.005 59.585 181.905 ;
        RECT 61.185 181.845 61.355 182.195 ;
        RECT 61.555 182.015 61.885 182.415 ;
        RECT 62.055 181.845 62.225 182.195 ;
        RECT 62.395 182.015 62.775 182.415 ;
        RECT 59.755 181.565 59.955 181.735 ;
        RECT 59.755 181.175 59.950 181.565 ;
        RECT 60.650 181.175 61.000 181.745 ;
        RECT 61.185 181.675 62.795 181.845 ;
        RECT 62.965 181.740 63.235 182.085 ;
        RECT 62.625 181.505 62.795 181.675 ;
        RECT 61.170 181.055 61.880 181.505 ;
        RECT 62.050 181.175 62.455 181.505 ;
        RECT 62.625 181.175 62.895 181.505 ;
        RECT 58.485 180.835 59.945 181.005 ;
        RECT 57.885 180.495 58.660 180.665 ;
        RECT 57.990 179.865 58.160 180.325 ;
        RECT 58.330 180.035 58.660 180.495 ;
        RECT 58.830 179.865 59.000 180.665 ;
        RECT 59.585 180.660 59.945 180.835 ;
        RECT 60.650 180.715 60.970 181.005 ;
        RECT 61.165 180.885 61.880 181.055 ;
        RECT 62.625 181.005 62.795 181.175 ;
        RECT 63.065 181.005 63.235 181.740 ;
        RECT 63.410 181.650 63.865 182.415 ;
        RECT 64.140 182.035 65.440 182.245 ;
        RECT 65.695 182.055 66.025 182.415 ;
        RECT 65.270 181.885 65.440 182.035 ;
        RECT 66.195 181.915 66.455 182.245 ;
        RECT 66.225 181.905 66.455 181.915 ;
        RECT 66.790 181.905 67.030 182.415 ;
        RECT 67.210 181.905 67.490 182.235 ;
        RECT 67.720 181.905 67.935 182.415 ;
        RECT 64.340 181.425 64.560 181.825 ;
        RECT 63.405 181.225 63.895 181.425 ;
        RECT 64.085 181.215 64.560 181.425 ;
        RECT 64.805 181.425 65.015 181.825 ;
        RECT 65.270 181.760 66.025 181.885 ;
        RECT 65.270 181.715 66.115 181.760 ;
        RECT 65.845 181.595 66.115 181.715 ;
        RECT 64.805 181.215 65.135 181.425 ;
        RECT 65.305 181.155 65.715 181.460 ;
        RECT 62.070 180.835 62.795 181.005 ;
        RECT 62.070 180.715 62.240 180.835 ;
        RECT 60.650 180.545 62.240 180.715 ;
        RECT 60.650 180.085 62.305 180.375 ;
        RECT 62.475 179.865 62.755 180.665 ;
        RECT 62.965 180.035 63.235 181.005 ;
        RECT 63.410 180.985 64.585 181.045 ;
        RECT 65.945 181.020 66.115 181.595 ;
        RECT 65.915 180.985 66.115 181.020 ;
        RECT 63.410 180.875 66.115 180.985 ;
        RECT 63.410 180.255 63.665 180.875 ;
        RECT 64.255 180.815 66.055 180.875 ;
        RECT 64.255 180.785 64.585 180.815 ;
        RECT 66.285 180.715 66.455 181.905 ;
        RECT 66.685 181.175 67.040 181.735 ;
        RECT 67.210 181.005 67.380 181.905 ;
        RECT 67.550 181.175 67.815 181.735 ;
        RECT 68.105 181.675 68.720 182.245 ;
        RECT 68.925 181.690 69.215 182.415 ;
        RECT 69.395 181.685 69.695 182.415 ;
        RECT 68.065 181.005 68.235 181.505 ;
        RECT 63.915 180.615 64.100 180.705 ;
        RECT 64.690 180.615 65.525 180.625 ;
        RECT 63.915 180.415 65.525 180.615 ;
        RECT 63.915 180.375 64.145 180.415 ;
        RECT 63.410 180.035 63.745 180.255 ;
        RECT 64.750 179.865 65.105 180.245 ;
        RECT 65.275 180.035 65.525 180.415 ;
        RECT 65.775 179.865 66.025 180.645 ;
        RECT 66.195 180.035 66.455 180.715 ;
        RECT 66.810 180.835 68.235 181.005 ;
        RECT 66.810 180.660 67.200 180.835 ;
        RECT 67.685 179.865 68.015 180.665 ;
        RECT 68.405 180.655 68.720 181.675 ;
        RECT 69.875 181.505 70.105 182.125 ;
        RECT 70.305 181.855 70.530 182.235 ;
        RECT 70.700 182.025 71.030 182.415 ;
        RECT 71.225 182.035 72.115 182.205 ;
        RECT 70.305 181.675 70.635 181.855 ;
        RECT 69.400 181.175 69.695 181.505 ;
        RECT 69.875 181.175 70.290 181.505 ;
        RECT 68.185 180.035 68.720 180.655 ;
        RECT 68.925 179.865 69.215 181.030 ;
        RECT 70.460 181.005 70.635 181.675 ;
        RECT 70.805 181.175 71.045 181.825 ;
        RECT 71.225 181.480 71.775 181.865 ;
        RECT 71.945 181.310 72.115 182.035 ;
        RECT 71.225 181.240 72.115 181.310 ;
        RECT 72.285 181.710 72.505 182.195 ;
        RECT 72.675 181.875 72.925 182.415 ;
        RECT 73.095 181.765 73.355 182.245 ;
        RECT 72.285 181.285 72.615 181.710 ;
        RECT 71.225 181.215 72.120 181.240 ;
        RECT 71.225 181.200 72.130 181.215 ;
        RECT 71.225 181.185 72.135 181.200 ;
        RECT 71.225 181.180 72.145 181.185 ;
        RECT 71.225 181.170 72.150 181.180 ;
        RECT 71.225 181.160 72.155 181.170 ;
        RECT 71.225 181.155 72.165 181.160 ;
        RECT 71.225 181.145 72.175 181.155 ;
        RECT 71.225 181.140 72.185 181.145 ;
        RECT 69.395 180.645 70.290 180.975 ;
        RECT 70.460 180.815 71.045 181.005 ;
        RECT 69.395 180.475 70.600 180.645 ;
        RECT 69.395 180.045 69.725 180.475 ;
        RECT 69.905 179.865 70.100 180.305 ;
        RECT 70.270 180.045 70.600 180.475 ;
        RECT 70.770 180.045 71.045 180.815 ;
        RECT 71.225 180.690 71.485 181.140 ;
        RECT 71.850 181.135 72.185 181.140 ;
        RECT 71.850 181.130 72.200 181.135 ;
        RECT 71.850 181.120 72.215 181.130 ;
        RECT 71.850 181.115 72.240 181.120 ;
        RECT 72.785 181.115 73.015 181.510 ;
        RECT 71.850 181.110 73.015 181.115 ;
        RECT 71.880 181.075 73.015 181.110 ;
        RECT 71.915 181.050 73.015 181.075 ;
        RECT 71.945 181.020 73.015 181.050 ;
        RECT 71.965 180.990 73.015 181.020 ;
        RECT 71.985 180.960 73.015 180.990 ;
        RECT 72.055 180.950 73.015 180.960 ;
        RECT 72.080 180.940 73.015 180.950 ;
        RECT 72.100 180.925 73.015 180.940 ;
        RECT 72.120 180.910 73.015 180.925 ;
        RECT 72.125 180.900 72.910 180.910 ;
        RECT 72.140 180.865 72.910 180.900 ;
        RECT 71.655 180.545 71.985 180.790 ;
        RECT 72.155 180.615 72.910 180.865 ;
        RECT 73.185 180.735 73.355 181.765 ;
        RECT 71.655 180.520 71.840 180.545 ;
        RECT 71.225 180.420 71.840 180.520 ;
        RECT 71.225 179.865 71.830 180.420 ;
        RECT 72.005 180.035 72.485 180.375 ;
        RECT 72.655 179.865 72.910 180.410 ;
        RECT 73.080 180.035 73.355 180.735 ;
        RECT 73.525 181.675 73.910 182.245 ;
        RECT 74.080 181.955 74.405 182.415 ;
        RECT 74.925 181.785 75.205 182.245 ;
        RECT 73.525 181.005 73.805 181.675 ;
        RECT 74.080 181.615 75.205 181.785 ;
        RECT 74.080 181.505 74.530 181.615 ;
        RECT 73.975 181.175 74.530 181.505 ;
        RECT 75.395 181.445 75.795 182.245 ;
        RECT 76.195 181.955 76.465 182.415 ;
        RECT 76.635 181.785 76.920 182.245 ;
        RECT 78.145 181.945 78.440 182.415 ;
        RECT 73.525 180.035 73.910 181.005 ;
        RECT 74.080 180.715 74.530 181.175 ;
        RECT 74.700 180.885 75.795 181.445 ;
        RECT 74.080 180.495 75.205 180.715 ;
        RECT 74.080 179.865 74.405 180.325 ;
        RECT 74.925 180.035 75.205 180.495 ;
        RECT 75.395 180.035 75.795 180.885 ;
        RECT 75.965 181.615 76.920 181.785 ;
        RECT 78.610 181.775 78.870 182.220 ;
        RECT 79.040 181.945 79.300 182.415 ;
        RECT 79.470 181.775 79.725 182.220 ;
        RECT 79.895 181.945 80.195 182.415 ;
        RECT 75.965 180.715 76.175 181.615 ;
        RECT 77.685 181.605 80.715 181.775 ;
        RECT 80.905 181.605 81.145 182.415 ;
        RECT 81.315 181.605 81.645 182.245 ;
        RECT 81.815 181.605 82.085 182.415 ;
        RECT 82.265 181.870 87.610 182.415 ;
        RECT 76.345 180.885 77.035 181.445 ;
        RECT 77.685 181.040 77.855 181.605 ;
        RECT 78.025 181.210 80.240 181.435 ;
        RECT 80.415 181.040 80.715 181.605 ;
        RECT 80.885 181.175 81.235 181.425 ;
        RECT 77.685 180.870 80.715 181.040 ;
        RECT 81.405 181.005 81.575 181.605 ;
        RECT 81.745 181.175 82.095 181.425 ;
        RECT 83.850 181.040 84.190 181.870 ;
        RECT 88.710 181.675 88.965 182.245 ;
        RECT 89.135 182.015 89.465 182.415 ;
        RECT 89.890 181.880 90.420 182.245 ;
        RECT 89.890 181.845 90.065 181.880 ;
        RECT 89.135 181.675 90.065 181.845 ;
        RECT 75.965 180.495 76.920 180.715 ;
        RECT 76.195 179.865 76.465 180.325 ;
        RECT 76.635 180.035 76.920 180.495 ;
        RECT 77.665 179.865 78.010 180.700 ;
        RECT 78.185 180.065 78.440 180.870 ;
        RECT 78.610 179.865 78.870 180.700 ;
        RECT 79.045 180.065 79.300 180.870 ;
        RECT 79.470 179.865 79.730 180.700 ;
        RECT 79.900 180.065 80.160 180.870 ;
        RECT 80.895 180.835 81.575 181.005 ;
        RECT 80.330 179.865 80.715 180.700 ;
        RECT 80.895 180.050 81.225 180.835 ;
        RECT 81.755 179.865 82.085 181.005 ;
        RECT 85.670 180.300 86.020 181.550 ;
        RECT 88.710 181.005 88.880 181.675 ;
        RECT 89.135 181.505 89.305 181.675 ;
        RECT 89.050 181.175 89.305 181.505 ;
        RECT 89.530 181.175 89.725 181.505 ;
        RECT 82.265 179.865 87.610 180.300 ;
        RECT 88.710 180.035 89.045 181.005 ;
        RECT 89.215 179.865 89.385 181.005 ;
        RECT 89.555 180.205 89.725 181.175 ;
        RECT 89.895 180.545 90.065 181.675 ;
        RECT 90.235 180.885 90.405 181.685 ;
        RECT 90.610 181.395 90.885 182.245 ;
        RECT 90.605 181.225 90.885 181.395 ;
        RECT 90.610 181.085 90.885 181.225 ;
        RECT 91.055 180.885 91.245 182.245 ;
        RECT 91.425 181.880 91.935 182.415 ;
        RECT 92.155 181.605 92.400 182.210 ;
        RECT 92.845 181.645 94.515 182.415 ;
        RECT 94.685 181.690 94.975 182.415 ;
        RECT 95.610 181.675 95.865 182.245 ;
        RECT 96.035 182.015 96.365 182.415 ;
        RECT 96.790 181.880 97.320 182.245 ;
        RECT 96.790 181.845 96.965 181.880 ;
        RECT 96.035 181.675 96.965 181.845 ;
        RECT 91.445 181.435 92.675 181.605 ;
        RECT 90.235 180.715 91.245 180.885 ;
        RECT 91.415 180.870 92.165 181.060 ;
        RECT 89.895 180.375 91.020 180.545 ;
        RECT 91.415 180.205 91.585 180.870 ;
        RECT 92.335 180.625 92.675 181.435 ;
        RECT 92.845 181.125 93.595 181.645 ;
        RECT 93.765 180.955 94.515 181.475 ;
        RECT 89.555 180.035 91.585 180.205 ;
        RECT 91.755 179.865 91.925 180.625 ;
        RECT 92.160 180.215 92.675 180.625 ;
        RECT 92.845 179.865 94.515 180.955 ;
        RECT 94.685 179.865 94.975 181.030 ;
        RECT 95.610 181.005 95.780 181.675 ;
        RECT 96.035 181.505 96.205 181.675 ;
        RECT 95.950 181.175 96.205 181.505 ;
        RECT 96.430 181.175 96.625 181.505 ;
        RECT 95.610 180.035 95.945 181.005 ;
        RECT 96.115 179.865 96.285 181.005 ;
        RECT 96.455 180.205 96.625 181.175 ;
        RECT 96.795 180.545 96.965 181.675 ;
        RECT 97.135 180.885 97.305 181.685 ;
        RECT 97.510 181.395 97.785 182.245 ;
        RECT 97.505 181.225 97.785 181.395 ;
        RECT 97.510 181.085 97.785 181.225 ;
        RECT 97.955 180.885 98.145 182.245 ;
        RECT 98.325 181.880 98.835 182.415 ;
        RECT 99.055 181.605 99.300 182.210 ;
        RECT 99.860 181.785 100.145 182.245 ;
        RECT 100.315 181.955 100.585 182.415 ;
        RECT 99.860 181.615 100.815 181.785 ;
        RECT 98.345 181.435 99.575 181.605 ;
        RECT 97.135 180.715 98.145 180.885 ;
        RECT 98.315 180.870 99.065 181.060 ;
        RECT 96.795 180.375 97.920 180.545 ;
        RECT 98.315 180.205 98.485 180.870 ;
        RECT 99.235 180.625 99.575 181.435 ;
        RECT 99.745 180.885 100.435 181.445 ;
        RECT 100.605 180.715 100.815 181.615 ;
        RECT 96.455 180.035 98.485 180.205 ;
        RECT 98.655 179.865 98.825 180.625 ;
        RECT 99.060 180.215 99.575 180.625 ;
        RECT 99.860 180.495 100.815 180.715 ;
        RECT 100.985 181.445 101.385 182.245 ;
        RECT 101.575 181.785 101.855 182.245 ;
        RECT 102.375 181.955 102.700 182.415 ;
        RECT 101.575 181.615 102.700 181.785 ;
        RECT 102.870 181.675 103.255 182.245 ;
        RECT 102.250 181.505 102.700 181.615 ;
        RECT 100.985 180.885 102.080 181.445 ;
        RECT 102.250 181.175 102.805 181.505 ;
        RECT 99.860 180.035 100.145 180.495 ;
        RECT 100.315 179.865 100.585 180.325 ;
        RECT 100.985 180.035 101.385 180.885 ;
        RECT 102.250 180.715 102.700 181.175 ;
        RECT 102.975 181.005 103.255 181.675 ;
        RECT 103.540 181.785 103.825 182.245 ;
        RECT 103.995 181.955 104.265 182.415 ;
        RECT 103.540 181.615 104.495 181.785 ;
        RECT 101.575 180.495 102.700 180.715 ;
        RECT 101.575 180.035 101.855 180.495 ;
        RECT 102.375 179.865 102.700 180.325 ;
        RECT 102.870 180.035 103.255 181.005 ;
        RECT 103.425 180.885 104.115 181.445 ;
        RECT 104.285 180.715 104.495 181.615 ;
        RECT 103.540 180.495 104.495 180.715 ;
        RECT 104.665 181.445 105.065 182.245 ;
        RECT 105.255 181.785 105.535 182.245 ;
        RECT 106.055 181.955 106.380 182.415 ;
        RECT 105.255 181.615 106.380 181.785 ;
        RECT 106.550 181.675 106.935 182.245 ;
        RECT 105.930 181.505 106.380 181.615 ;
        RECT 104.665 180.885 105.760 181.445 ;
        RECT 105.930 181.175 106.485 181.505 ;
        RECT 103.540 180.035 103.825 180.495 ;
        RECT 103.995 179.865 104.265 180.325 ;
        RECT 104.665 180.035 105.065 180.885 ;
        RECT 105.930 180.715 106.380 181.175 ;
        RECT 106.655 181.005 106.935 181.675 ;
        RECT 107.105 181.665 108.315 182.415 ;
        RECT 108.490 181.675 108.745 182.245 ;
        RECT 108.915 182.015 109.245 182.415 ;
        RECT 109.670 181.880 110.200 182.245 ;
        RECT 110.390 182.075 110.665 182.245 ;
        RECT 110.385 181.905 110.665 182.075 ;
        RECT 109.670 181.845 109.845 181.880 ;
        RECT 108.915 181.675 109.845 181.845 ;
        RECT 107.105 181.125 107.625 181.665 ;
        RECT 105.255 180.495 106.380 180.715 ;
        RECT 105.255 180.035 105.535 180.495 ;
        RECT 106.055 179.865 106.380 180.325 ;
        RECT 106.550 180.035 106.935 181.005 ;
        RECT 107.795 180.955 108.315 181.495 ;
        RECT 107.105 179.865 108.315 180.955 ;
        RECT 108.490 181.005 108.660 181.675 ;
        RECT 108.915 181.505 109.085 181.675 ;
        RECT 108.830 181.175 109.085 181.505 ;
        RECT 109.310 181.175 109.505 181.505 ;
        RECT 108.490 180.035 108.825 181.005 ;
        RECT 108.995 179.865 109.165 181.005 ;
        RECT 109.335 180.205 109.505 181.175 ;
        RECT 109.675 180.545 109.845 181.675 ;
        RECT 110.015 180.885 110.185 181.685 ;
        RECT 110.390 181.085 110.665 181.905 ;
        RECT 110.835 180.885 111.025 182.245 ;
        RECT 111.205 181.880 111.715 182.415 ;
        RECT 111.935 181.605 112.180 182.210 ;
        RECT 112.625 181.675 113.010 182.245 ;
        RECT 113.180 181.955 113.505 182.415 ;
        RECT 114.025 181.785 114.305 182.245 ;
        RECT 111.225 181.435 112.455 181.605 ;
        RECT 110.015 180.715 111.025 180.885 ;
        RECT 111.195 180.870 111.945 181.060 ;
        RECT 109.675 180.375 110.800 180.545 ;
        RECT 111.195 180.205 111.365 180.870 ;
        RECT 112.115 180.625 112.455 181.435 ;
        RECT 109.335 180.035 111.365 180.205 ;
        RECT 111.535 179.865 111.705 180.625 ;
        RECT 111.940 180.215 112.455 180.625 ;
        RECT 112.625 181.005 112.905 181.675 ;
        RECT 113.180 181.615 114.305 181.785 ;
        RECT 113.180 181.505 113.630 181.615 ;
        RECT 113.075 181.175 113.630 181.505 ;
        RECT 114.495 181.445 114.895 182.245 ;
        RECT 115.295 181.955 115.565 182.415 ;
        RECT 115.735 181.785 116.020 182.245 ;
        RECT 112.625 180.035 113.010 181.005 ;
        RECT 113.180 180.715 113.630 181.175 ;
        RECT 113.800 180.885 114.895 181.445 ;
        RECT 113.180 180.495 114.305 180.715 ;
        RECT 113.180 179.865 113.505 180.325 ;
        RECT 114.025 180.035 114.305 180.495 ;
        RECT 114.495 180.035 114.895 180.885 ;
        RECT 115.065 181.615 116.020 181.785 ;
        RECT 116.310 181.675 116.565 182.245 ;
        RECT 116.735 182.015 117.065 182.415 ;
        RECT 117.490 181.880 118.020 182.245 ;
        RECT 117.490 181.845 117.665 181.880 ;
        RECT 116.735 181.675 117.665 181.845 ;
        RECT 115.065 180.715 115.275 181.615 ;
        RECT 115.445 180.885 116.135 181.445 ;
        RECT 116.310 181.005 116.480 181.675 ;
        RECT 116.735 181.505 116.905 181.675 ;
        RECT 116.650 181.175 116.905 181.505 ;
        RECT 117.130 181.175 117.325 181.505 ;
        RECT 115.065 180.495 116.020 180.715 ;
        RECT 115.295 179.865 115.565 180.325 ;
        RECT 115.735 180.035 116.020 180.495 ;
        RECT 116.310 180.035 116.645 181.005 ;
        RECT 116.815 179.865 116.985 181.005 ;
        RECT 117.155 180.205 117.325 181.175 ;
        RECT 117.495 180.545 117.665 181.675 ;
        RECT 117.835 180.885 118.005 181.685 ;
        RECT 118.210 181.395 118.485 182.245 ;
        RECT 118.205 181.225 118.485 181.395 ;
        RECT 118.210 181.085 118.485 181.225 ;
        RECT 118.655 180.885 118.845 182.245 ;
        RECT 119.025 181.880 119.535 182.415 ;
        RECT 119.755 181.605 120.000 182.210 ;
        RECT 120.445 181.690 120.735 182.415 ;
        RECT 120.995 181.865 121.165 182.155 ;
        RECT 121.335 182.035 121.665 182.415 ;
        RECT 120.995 181.695 121.660 181.865 ;
        RECT 119.045 181.435 120.275 181.605 ;
        RECT 117.835 180.715 118.845 180.885 ;
        RECT 119.015 180.870 119.765 181.060 ;
        RECT 117.495 180.375 118.620 180.545 ;
        RECT 119.015 180.205 119.185 180.870 ;
        RECT 119.935 180.625 120.275 181.435 ;
        RECT 117.155 180.035 119.185 180.205 ;
        RECT 119.355 179.865 119.525 180.625 ;
        RECT 119.760 180.215 120.275 180.625 ;
        RECT 120.445 179.865 120.735 181.030 ;
        RECT 120.910 180.875 121.260 181.525 ;
        RECT 121.430 180.705 121.660 181.695 ;
        RECT 120.995 180.535 121.660 180.705 ;
        RECT 120.995 180.035 121.165 180.535 ;
        RECT 121.335 179.865 121.665 180.365 ;
        RECT 121.835 180.035 122.020 182.155 ;
        RECT 122.275 181.955 122.525 182.415 ;
        RECT 122.695 181.965 123.030 182.135 ;
        RECT 123.225 181.965 123.900 182.135 ;
        RECT 122.695 181.825 122.865 181.965 ;
        RECT 122.190 180.835 122.470 181.785 ;
        RECT 122.640 181.695 122.865 181.825 ;
        RECT 122.640 180.590 122.810 181.695 ;
        RECT 123.035 181.545 123.560 181.765 ;
        RECT 122.980 180.780 123.220 181.375 ;
        RECT 123.390 180.845 123.560 181.545 ;
        RECT 123.730 181.185 123.900 181.965 ;
        RECT 124.220 181.915 124.590 182.415 ;
        RECT 124.770 181.965 125.175 182.135 ;
        RECT 125.345 181.965 126.130 182.135 ;
        RECT 124.770 181.735 124.940 181.965 ;
        RECT 124.110 181.435 124.940 181.735 ;
        RECT 125.325 181.465 125.790 181.795 ;
        RECT 124.110 181.405 124.310 181.435 ;
        RECT 124.430 181.185 124.600 181.255 ;
        RECT 123.730 181.015 124.600 181.185 ;
        RECT 124.090 180.925 124.600 181.015 ;
        RECT 122.640 180.460 122.945 180.590 ;
        RECT 123.390 180.480 123.920 180.845 ;
        RECT 122.260 179.865 122.525 180.325 ;
        RECT 122.695 180.035 122.945 180.460 ;
        RECT 124.090 180.310 124.260 180.925 ;
        RECT 123.155 180.140 124.260 180.310 ;
        RECT 124.430 179.865 124.600 180.665 ;
        RECT 124.770 180.365 124.940 181.435 ;
        RECT 125.110 180.535 125.300 181.255 ;
        RECT 125.470 180.505 125.790 181.465 ;
        RECT 125.960 181.505 126.130 181.965 ;
        RECT 126.405 181.885 126.615 182.415 ;
        RECT 126.875 181.675 127.205 182.200 ;
        RECT 127.375 181.805 127.545 182.415 ;
        RECT 127.715 181.760 128.045 182.195 ;
        RECT 127.715 181.675 128.095 181.760 ;
        RECT 127.005 181.505 127.205 181.675 ;
        RECT 127.870 181.635 128.095 181.675 ;
        RECT 125.960 181.175 126.835 181.505 ;
        RECT 127.005 181.175 127.755 181.505 ;
        RECT 124.770 180.035 125.020 180.365 ;
        RECT 125.960 180.335 126.130 181.175 ;
        RECT 127.005 180.970 127.195 181.175 ;
        RECT 127.925 181.055 128.095 181.635 ;
        RECT 127.880 181.005 128.095 181.055 ;
        RECT 126.300 180.595 127.195 180.970 ;
        RECT 127.705 180.925 128.095 181.005 ;
        RECT 128.265 181.675 128.650 182.245 ;
        RECT 128.820 181.955 129.145 182.415 ;
        RECT 129.665 181.785 129.945 182.245 ;
        RECT 128.265 181.005 128.545 181.675 ;
        RECT 128.820 181.615 129.945 181.785 ;
        RECT 128.820 181.505 129.270 181.615 ;
        RECT 128.715 181.175 129.270 181.505 ;
        RECT 130.135 181.445 130.535 182.245 ;
        RECT 130.935 181.955 131.205 182.415 ;
        RECT 131.375 181.785 131.660 182.245 ;
        RECT 132.110 181.905 132.350 182.415 ;
        RECT 132.530 181.905 132.810 182.235 ;
        RECT 133.040 181.905 133.255 182.415 ;
        RECT 125.245 180.165 126.130 180.335 ;
        RECT 126.310 179.865 126.625 180.365 ;
        RECT 126.855 180.035 127.195 180.595 ;
        RECT 127.365 179.865 127.535 180.875 ;
        RECT 127.705 180.080 128.035 180.925 ;
        RECT 128.265 180.035 128.650 181.005 ;
        RECT 128.820 180.715 129.270 181.175 ;
        RECT 129.440 180.885 130.535 181.445 ;
        RECT 128.820 180.495 129.945 180.715 ;
        RECT 128.820 179.865 129.145 180.325 ;
        RECT 129.665 180.035 129.945 180.495 ;
        RECT 130.135 180.035 130.535 180.885 ;
        RECT 130.705 181.615 131.660 181.785 ;
        RECT 130.705 180.715 130.915 181.615 ;
        RECT 131.085 180.885 131.775 181.445 ;
        RECT 132.005 181.175 132.360 181.735 ;
        RECT 132.530 181.005 132.700 181.905 ;
        RECT 132.870 181.175 133.135 181.735 ;
        RECT 133.425 181.675 134.040 182.245 ;
        RECT 134.295 181.760 134.625 182.195 ;
        RECT 134.795 181.805 134.965 182.415 ;
        RECT 133.385 181.005 133.555 181.505 ;
        RECT 132.130 180.835 133.555 181.005 ;
        RECT 130.705 180.495 131.660 180.715 ;
        RECT 132.130 180.660 132.520 180.835 ;
        RECT 130.935 179.865 131.205 180.325 ;
        RECT 131.375 180.035 131.660 180.495 ;
        RECT 133.005 179.865 133.335 180.665 ;
        RECT 133.725 180.655 134.040 181.675 ;
        RECT 134.245 181.675 134.625 181.760 ;
        RECT 135.135 181.675 135.465 182.200 ;
        RECT 135.725 181.885 135.935 182.415 ;
        RECT 136.210 181.965 136.995 182.135 ;
        RECT 137.165 181.965 137.570 182.135 ;
        RECT 134.245 181.635 134.470 181.675 ;
        RECT 134.245 181.055 134.415 181.635 ;
        RECT 135.135 181.505 135.335 181.675 ;
        RECT 136.210 181.505 136.380 181.965 ;
        RECT 134.585 181.175 135.335 181.505 ;
        RECT 135.505 181.175 136.380 181.505 ;
        RECT 134.245 181.005 134.460 181.055 ;
        RECT 134.245 180.925 134.635 181.005 ;
        RECT 133.505 180.035 134.040 180.655 ;
        RECT 134.305 180.080 134.635 180.925 ;
        RECT 135.145 180.970 135.335 181.175 ;
        RECT 134.805 179.865 134.975 180.875 ;
        RECT 135.145 180.595 136.040 180.970 ;
        RECT 135.145 180.035 135.485 180.595 ;
        RECT 135.715 179.865 136.030 180.365 ;
        RECT 136.210 180.335 136.380 181.175 ;
        RECT 136.550 181.465 137.015 181.795 ;
        RECT 137.400 181.735 137.570 181.965 ;
        RECT 137.750 181.915 138.120 182.415 ;
        RECT 138.440 181.965 139.115 182.135 ;
        RECT 139.310 181.965 139.645 182.135 ;
        RECT 136.550 180.505 136.870 181.465 ;
        RECT 137.400 181.435 138.230 181.735 ;
        RECT 137.040 180.535 137.230 181.255 ;
        RECT 137.400 180.365 137.570 181.435 ;
        RECT 138.030 181.405 138.230 181.435 ;
        RECT 137.740 181.185 137.910 181.255 ;
        RECT 138.440 181.185 138.610 181.965 ;
        RECT 139.475 181.825 139.645 181.965 ;
        RECT 139.815 181.955 140.065 182.415 ;
        RECT 137.740 181.015 138.610 181.185 ;
        RECT 138.780 181.545 139.305 181.765 ;
        RECT 139.475 181.695 139.700 181.825 ;
        RECT 137.740 180.925 138.250 181.015 ;
        RECT 136.210 180.165 137.095 180.335 ;
        RECT 137.320 180.035 137.570 180.365 ;
        RECT 137.740 179.865 137.910 180.665 ;
        RECT 138.080 180.310 138.250 180.925 ;
        RECT 138.780 180.845 138.950 181.545 ;
        RECT 138.420 180.480 138.950 180.845 ;
        RECT 139.120 180.780 139.360 181.375 ;
        RECT 139.530 180.590 139.700 181.695 ;
        RECT 139.870 180.835 140.150 181.785 ;
        RECT 139.395 180.460 139.700 180.590 ;
        RECT 138.080 180.140 139.185 180.310 ;
        RECT 139.395 180.035 139.645 180.460 ;
        RECT 139.815 179.865 140.080 180.325 ;
        RECT 140.320 180.035 140.505 182.155 ;
        RECT 140.675 182.035 141.005 182.415 ;
        RECT 141.175 181.865 141.345 182.155 ;
        RECT 140.680 181.695 141.345 181.865 ;
        RECT 140.680 180.705 140.910 181.695 ;
        RECT 141.605 181.645 145.115 182.415 ;
        RECT 145.745 181.665 146.955 182.415 ;
        RECT 141.080 180.875 141.430 181.525 ;
        RECT 141.605 181.125 143.255 181.645 ;
        RECT 143.425 180.955 145.115 181.475 ;
        RECT 140.680 180.535 141.345 180.705 ;
        RECT 140.675 179.865 141.005 180.365 ;
        RECT 141.175 180.035 141.345 180.535 ;
        RECT 141.605 179.865 145.115 180.955 ;
        RECT 145.745 180.955 146.265 181.495 ;
        RECT 146.435 181.125 146.955 181.665 ;
        RECT 145.745 179.865 146.955 180.955 ;
        RECT 17.320 179.695 147.040 179.865 ;
        RECT 17.405 178.605 18.615 179.695 ;
        RECT 18.785 178.605 22.295 179.695 ;
        RECT 17.405 177.895 17.925 178.435 ;
        RECT 18.095 178.065 18.615 178.605 ;
        RECT 18.785 177.915 20.435 178.435 ;
        RECT 20.605 178.085 22.295 178.605 ;
        RECT 22.465 178.825 22.740 179.525 ;
        RECT 22.910 179.150 23.165 179.695 ;
        RECT 23.335 179.185 23.815 179.525 ;
        RECT 23.990 179.140 24.595 179.695 ;
        RECT 23.980 179.040 24.595 179.140 ;
        RECT 23.980 179.015 24.165 179.040 ;
        RECT 17.405 177.145 18.615 177.895 ;
        RECT 18.785 177.145 22.295 177.915 ;
        RECT 22.465 177.795 22.635 178.825 ;
        RECT 22.910 178.695 23.665 178.945 ;
        RECT 23.835 178.770 24.165 179.015 ;
        RECT 22.910 178.660 23.680 178.695 ;
        RECT 22.910 178.650 23.695 178.660 ;
        RECT 22.805 178.635 23.700 178.650 ;
        RECT 22.805 178.620 23.720 178.635 ;
        RECT 22.805 178.610 23.740 178.620 ;
        RECT 22.805 178.600 23.765 178.610 ;
        RECT 22.805 178.570 23.835 178.600 ;
        RECT 22.805 178.540 23.855 178.570 ;
        RECT 22.805 178.510 23.875 178.540 ;
        RECT 22.805 178.485 23.905 178.510 ;
        RECT 22.805 178.450 23.940 178.485 ;
        RECT 22.805 178.445 23.970 178.450 ;
        RECT 22.805 178.050 23.035 178.445 ;
        RECT 23.580 178.440 23.970 178.445 ;
        RECT 23.605 178.430 23.970 178.440 ;
        RECT 23.620 178.425 23.970 178.430 ;
        RECT 23.635 178.420 23.970 178.425 ;
        RECT 24.335 178.420 24.595 178.870 ;
        RECT 24.950 178.725 25.340 178.900 ;
        RECT 25.825 178.895 26.155 179.695 ;
        RECT 26.325 178.905 26.860 179.525 ;
        RECT 24.950 178.555 26.375 178.725 ;
        RECT 23.635 178.415 24.595 178.420 ;
        RECT 23.645 178.405 24.595 178.415 ;
        RECT 23.655 178.400 24.595 178.405 ;
        RECT 23.665 178.390 24.595 178.400 ;
        RECT 23.670 178.380 24.595 178.390 ;
        RECT 23.675 178.375 24.595 178.380 ;
        RECT 23.685 178.360 24.595 178.375 ;
        RECT 23.690 178.345 24.595 178.360 ;
        RECT 23.700 178.320 24.595 178.345 ;
        RECT 23.205 177.850 23.535 178.275 ;
        RECT 22.465 177.315 22.725 177.795 ;
        RECT 22.895 177.145 23.145 177.685 ;
        RECT 23.315 177.365 23.535 177.850 ;
        RECT 23.705 178.250 24.595 178.320 ;
        RECT 23.705 177.525 23.875 178.250 ;
        RECT 24.045 177.695 24.595 178.080 ;
        RECT 24.825 177.825 25.180 178.385 ;
        RECT 25.350 177.655 25.520 178.555 ;
        RECT 25.690 177.825 25.955 178.385 ;
        RECT 26.205 178.055 26.375 178.555 ;
        RECT 26.545 177.885 26.860 178.905 ;
        RECT 27.105 178.555 27.335 179.695 ;
        RECT 27.505 178.545 27.835 179.525 ;
        RECT 28.005 178.555 28.215 179.695 ;
        RECT 28.445 178.555 28.705 179.695 ;
        RECT 28.875 178.545 29.205 179.525 ;
        RECT 29.375 178.555 29.655 179.695 ;
        RECT 27.085 178.135 27.415 178.385 ;
        RECT 23.705 177.355 24.595 177.525 ;
        RECT 24.930 177.145 25.170 177.655 ;
        RECT 25.350 177.325 25.630 177.655 ;
        RECT 25.860 177.145 26.075 177.655 ;
        RECT 26.245 177.315 26.860 177.885 ;
        RECT 27.105 177.145 27.335 177.965 ;
        RECT 27.585 177.945 27.835 178.545 ;
        RECT 28.465 178.135 28.800 178.385 ;
        RECT 27.505 177.315 27.835 177.945 ;
        RECT 28.005 177.145 28.215 177.965 ;
        RECT 28.970 177.945 29.140 178.545 ;
        RECT 30.285 178.530 30.575 179.695 ;
        RECT 30.745 178.605 34.255 179.695 ;
        RECT 29.310 178.115 29.645 178.385 ;
        RECT 28.445 177.315 29.140 177.945 ;
        RECT 29.345 177.145 29.655 177.945 ;
        RECT 30.745 177.915 32.395 178.435 ;
        RECT 32.565 178.085 34.255 178.605 ;
        RECT 35.090 178.725 35.420 179.525 ;
        RECT 35.590 178.895 35.920 179.695 ;
        RECT 36.220 178.725 36.550 179.525 ;
        RECT 37.195 178.895 37.445 179.695 ;
        RECT 35.090 178.555 37.525 178.725 ;
        RECT 37.715 178.555 37.885 179.695 ;
        RECT 38.055 178.555 38.395 179.525 ;
        RECT 38.565 178.555 38.845 179.695 ;
        RECT 34.885 178.135 35.235 178.385 ;
        RECT 35.420 177.925 35.590 178.555 ;
        RECT 35.760 178.135 36.090 178.335 ;
        RECT 36.260 178.135 36.590 178.335 ;
        RECT 36.760 178.135 37.180 178.335 ;
        RECT 37.355 178.305 37.525 178.555 ;
        RECT 37.355 178.135 38.050 178.305 ;
        RECT 30.285 177.145 30.575 177.870 ;
        RECT 30.745 177.145 34.255 177.915 ;
        RECT 35.090 177.315 35.590 177.925 ;
        RECT 36.220 177.795 37.445 177.965 ;
        RECT 38.220 177.945 38.395 178.555 ;
        RECT 39.015 178.545 39.345 179.525 ;
        RECT 39.515 178.555 39.775 179.695 ;
        RECT 39.945 178.555 40.205 179.695 ;
        RECT 40.445 179.185 42.060 179.515 ;
        RECT 38.575 178.115 38.910 178.385 ;
        RECT 39.080 177.995 39.250 178.545 ;
        RECT 40.455 178.385 40.625 178.945 ;
        RECT 40.885 178.845 42.060 179.015 ;
        RECT 42.230 178.895 42.510 179.695 ;
        RECT 40.885 178.555 41.215 178.845 ;
        RECT 41.890 178.725 42.060 178.845 ;
        RECT 41.385 178.385 41.630 178.675 ;
        RECT 41.890 178.555 42.550 178.725 ;
        RECT 42.720 178.555 42.995 179.525 ;
        RECT 43.415 178.965 43.710 179.695 ;
        RECT 43.880 178.795 44.140 179.520 ;
        RECT 44.310 178.965 44.570 179.695 ;
        RECT 44.740 178.795 45.000 179.520 ;
        RECT 45.170 178.965 45.430 179.695 ;
        RECT 45.600 178.795 45.860 179.520 ;
        RECT 46.030 178.965 46.290 179.695 ;
        RECT 46.460 178.795 46.720 179.520 ;
        RECT 42.380 178.385 42.550 178.555 ;
        RECT 39.420 178.135 39.755 178.385 ;
        RECT 39.950 178.135 40.285 178.385 ;
        RECT 40.455 178.055 41.170 178.385 ;
        RECT 41.385 178.055 42.210 178.385 ;
        RECT 42.380 178.055 42.655 178.385 ;
        RECT 39.080 177.945 39.255 177.995 ;
        RECT 40.455 177.965 40.705 178.055 ;
        RECT 36.220 177.315 36.550 177.795 ;
        RECT 36.720 177.145 36.945 177.605 ;
        RECT 37.115 177.315 37.445 177.795 ;
        RECT 37.635 177.145 37.885 177.945 ;
        RECT 38.055 177.315 38.395 177.945 ;
        RECT 38.565 177.145 38.875 177.945 ;
        RECT 39.080 177.315 39.775 177.945 ;
        RECT 39.945 177.145 40.205 177.965 ;
        RECT 40.375 177.545 40.705 177.965 ;
        RECT 42.380 177.885 42.550 178.055 ;
        RECT 40.885 177.715 42.550 177.885 ;
        RECT 42.825 177.820 42.995 178.555 ;
        RECT 40.885 177.315 41.145 177.715 ;
        RECT 41.315 177.145 41.645 177.545 ;
        RECT 41.815 177.365 41.985 177.715 ;
        RECT 42.155 177.145 42.530 177.545 ;
        RECT 42.720 177.475 42.995 177.820 ;
        RECT 43.410 178.555 46.720 178.795 ;
        RECT 46.890 178.585 47.150 179.695 ;
        RECT 43.410 177.965 44.380 178.555 ;
        RECT 47.320 178.385 47.570 179.520 ;
        RECT 47.750 178.585 48.045 179.695 ;
        RECT 48.225 179.260 53.570 179.695 ;
        RECT 44.550 178.135 47.570 178.385 ;
        RECT 43.410 177.795 46.720 177.965 ;
        RECT 43.410 177.145 43.710 177.625 ;
        RECT 43.880 177.340 44.140 177.795 ;
        RECT 44.310 177.145 44.570 177.625 ;
        RECT 44.740 177.340 45.000 177.795 ;
        RECT 45.170 177.145 45.430 177.625 ;
        RECT 45.600 177.340 45.860 177.795 ;
        RECT 46.030 177.145 46.290 177.625 ;
        RECT 46.460 177.340 46.720 177.795 ;
        RECT 46.890 177.145 47.150 177.670 ;
        RECT 47.320 177.325 47.570 178.135 ;
        RECT 47.740 177.775 48.055 178.385 ;
        RECT 49.810 177.690 50.150 178.520 ;
        RECT 51.630 178.010 51.980 179.260 ;
        RECT 53.745 178.605 55.415 179.695 ;
        RECT 53.745 177.915 54.495 178.435 ;
        RECT 54.665 178.085 55.415 178.605 ;
        RECT 56.045 178.530 56.335 179.695 ;
        RECT 56.970 178.555 57.290 179.695 ;
        RECT 57.470 178.385 57.665 179.435 ;
        RECT 57.845 178.845 58.175 179.525 ;
        RECT 58.375 178.895 58.630 179.695 ;
        RECT 57.845 178.565 58.195 178.845 ;
        RECT 58.970 178.785 59.220 179.515 ;
        RECT 59.390 178.965 59.720 179.695 ;
        RECT 59.890 178.785 60.075 179.515 ;
        RECT 57.030 178.335 57.290 178.385 ;
        RECT 57.025 178.165 57.290 178.335 ;
        RECT 57.030 178.055 57.290 178.165 ;
        RECT 57.470 178.055 57.855 178.385 ;
        RECT 58.025 178.185 58.195 178.565 ;
        RECT 58.385 178.355 58.630 178.715 ;
        RECT 58.970 178.585 60.075 178.785 ;
        RECT 60.245 178.385 60.475 179.515 ;
        RECT 60.655 178.845 61.380 179.515 ;
        RECT 58.025 178.015 58.545 178.185 ;
        RECT 47.750 177.145 47.995 177.605 ;
        RECT 48.225 177.145 53.570 177.690 ;
        RECT 53.745 177.145 55.415 177.915 ;
        RECT 56.045 177.145 56.335 177.870 ;
        RECT 56.970 177.675 58.185 177.845 ;
        RECT 56.970 177.325 57.260 177.675 ;
        RECT 57.455 177.145 57.785 177.505 ;
        RECT 57.955 177.370 58.185 177.675 ;
        RECT 58.375 177.450 58.545 178.015 ;
        RECT 58.815 177.825 59.155 178.385 ;
        RECT 59.325 178.055 59.965 178.385 ;
        RECT 60.145 178.055 60.475 178.385 ;
        RECT 60.655 178.055 60.955 178.675 ;
        RECT 58.805 177.145 59.145 177.655 ;
        RECT 59.325 177.325 59.575 178.055 ;
        RECT 61.165 177.875 61.380 178.845 ;
        RECT 61.565 178.725 61.855 179.525 ;
        RECT 62.025 178.895 62.260 179.695 ;
        RECT 62.445 179.355 63.980 179.525 ;
        RECT 62.445 178.725 62.775 179.355 ;
        RECT 61.565 178.555 62.775 178.725 ;
        RECT 61.565 178.055 61.810 178.385 ;
        RECT 61.980 177.885 62.150 178.555 ;
        RECT 62.945 178.385 63.180 179.130 ;
        RECT 62.320 178.055 62.720 178.385 ;
        RECT 62.890 178.055 63.180 178.385 ;
        RECT 63.370 178.385 63.640 179.130 ;
        RECT 63.810 178.725 63.980 179.355 ;
        RECT 64.150 178.895 64.555 179.695 ;
        RECT 63.810 178.555 64.555 178.725 ;
        RECT 63.370 178.055 63.710 178.385 ;
        RECT 63.880 178.055 64.215 178.385 ;
        RECT 64.385 178.055 64.555 178.555 ;
        RECT 64.725 178.130 65.075 179.525 ;
        RECT 65.245 179.260 70.590 179.695 ;
        RECT 59.900 177.685 61.380 177.875 ;
        RECT 59.900 177.325 60.085 177.685 ;
        RECT 60.265 177.145 60.595 177.515 ;
        RECT 60.775 177.325 61.000 177.685 ;
        RECT 61.565 177.315 62.150 177.885 ;
        RECT 62.400 177.715 63.795 177.885 ;
        RECT 62.400 177.370 62.730 177.715 ;
        RECT 62.945 177.145 63.320 177.545 ;
        RECT 63.500 177.370 63.795 177.715 ;
        RECT 63.965 177.145 64.635 177.885 ;
        RECT 64.805 177.315 65.075 178.130 ;
        RECT 66.830 177.690 67.170 178.520 ;
        RECT 68.650 178.010 69.000 179.260 ;
        RECT 70.765 178.605 71.975 179.695 ;
        RECT 70.765 177.895 71.285 178.435 ;
        RECT 71.455 178.065 71.975 178.605 ;
        RECT 72.150 179.340 73.230 179.510 ;
        RECT 72.150 178.555 72.485 179.340 ;
        RECT 72.655 178.385 72.890 179.065 ;
        RECT 73.060 178.725 73.230 179.340 ;
        RECT 73.495 178.895 73.810 179.695 ;
        RECT 73.060 178.555 73.375 178.725 ;
        RECT 72.150 178.055 72.485 178.385 ;
        RECT 72.655 178.055 73.035 178.385 ;
        RECT 65.245 177.145 70.590 177.690 ;
        RECT 70.765 177.145 71.975 177.895 ;
        RECT 73.205 177.885 73.375 178.555 ;
        RECT 72.150 177.715 73.375 177.885 ;
        RECT 73.545 177.715 73.815 178.725 ;
        RECT 74.045 178.635 74.375 179.480 ;
        RECT 74.545 178.685 74.715 179.695 ;
        RECT 74.885 178.965 75.225 179.525 ;
        RECT 75.455 179.195 75.770 179.695 ;
        RECT 75.950 179.225 76.835 179.395 ;
        RECT 73.985 178.555 74.375 178.635 ;
        RECT 74.885 178.590 75.780 178.965 ;
        RECT 73.985 178.505 74.200 178.555 ;
        RECT 73.985 177.925 74.155 178.505 ;
        RECT 74.885 178.385 75.075 178.590 ;
        RECT 75.950 178.385 76.120 179.225 ;
        RECT 77.060 179.195 77.310 179.525 ;
        RECT 74.325 178.055 75.075 178.385 ;
        RECT 75.245 178.055 76.120 178.385 ;
        RECT 73.985 177.885 74.210 177.925 ;
        RECT 74.875 177.885 75.075 178.055 ;
        RECT 73.985 177.800 74.365 177.885 ;
        RECT 72.150 177.445 72.405 177.715 ;
        RECT 72.575 177.145 72.905 177.545 ;
        RECT 73.075 177.445 73.245 177.715 ;
        RECT 73.415 177.145 73.745 177.545 ;
        RECT 74.035 177.365 74.365 177.800 ;
        RECT 74.535 177.145 74.705 177.755 ;
        RECT 74.875 177.360 75.205 177.885 ;
        RECT 75.465 177.145 75.675 177.675 ;
        RECT 75.950 177.595 76.120 178.055 ;
        RECT 76.290 178.095 76.610 179.055 ;
        RECT 76.780 178.305 76.970 179.025 ;
        RECT 77.140 178.125 77.310 179.195 ;
        RECT 77.480 178.895 77.650 179.695 ;
        RECT 77.820 179.250 78.925 179.420 ;
        RECT 77.820 178.635 77.990 179.250 ;
        RECT 79.135 179.100 79.385 179.525 ;
        RECT 79.555 179.235 79.820 179.695 ;
        RECT 78.160 178.715 78.690 179.080 ;
        RECT 79.135 178.970 79.440 179.100 ;
        RECT 77.480 178.545 77.990 178.635 ;
        RECT 77.480 178.375 78.350 178.545 ;
        RECT 77.480 178.305 77.650 178.375 ;
        RECT 77.770 178.125 77.970 178.155 ;
        RECT 76.290 177.765 76.755 178.095 ;
        RECT 77.140 177.825 77.970 178.125 ;
        RECT 77.140 177.595 77.310 177.825 ;
        RECT 75.950 177.425 76.735 177.595 ;
        RECT 76.905 177.425 77.310 177.595 ;
        RECT 77.490 177.145 77.860 177.645 ;
        RECT 78.180 177.595 78.350 178.375 ;
        RECT 78.520 178.015 78.690 178.715 ;
        RECT 78.860 178.185 79.100 178.780 ;
        RECT 78.520 177.795 79.045 178.015 ;
        RECT 79.270 177.865 79.440 178.970 ;
        RECT 79.215 177.735 79.440 177.865 ;
        RECT 79.610 177.775 79.890 178.725 ;
        RECT 79.215 177.595 79.385 177.735 ;
        RECT 78.180 177.425 78.855 177.595 ;
        RECT 79.050 177.425 79.385 177.595 ;
        RECT 79.555 177.145 79.805 177.605 ;
        RECT 80.060 177.405 80.245 179.525 ;
        RECT 80.415 179.195 80.745 179.695 ;
        RECT 80.915 179.025 81.085 179.525 ;
        RECT 80.420 178.855 81.085 179.025 ;
        RECT 80.420 177.865 80.650 178.855 ;
        RECT 80.820 178.035 81.170 178.685 ;
        RECT 81.805 178.530 82.095 179.695 ;
        RECT 82.265 178.605 83.935 179.695 ;
        RECT 84.655 179.025 84.825 179.525 ;
        RECT 84.995 179.195 85.325 179.695 ;
        RECT 84.655 178.855 85.320 179.025 ;
        RECT 82.265 177.915 83.015 178.435 ;
        RECT 83.185 178.085 83.935 178.605 ;
        RECT 84.570 178.035 84.920 178.685 ;
        RECT 80.420 177.695 81.085 177.865 ;
        RECT 80.415 177.145 80.745 177.525 ;
        RECT 80.915 177.405 81.085 177.695 ;
        RECT 81.805 177.145 82.095 177.870 ;
        RECT 82.265 177.145 83.935 177.915 ;
        RECT 85.090 177.865 85.320 178.855 ;
        RECT 84.655 177.695 85.320 177.865 ;
        RECT 84.655 177.405 84.825 177.695 ;
        RECT 84.995 177.145 85.325 177.525 ;
        RECT 85.495 177.405 85.680 179.525 ;
        RECT 85.920 179.235 86.185 179.695 ;
        RECT 86.355 179.100 86.605 179.525 ;
        RECT 86.815 179.250 87.920 179.420 ;
        RECT 86.300 178.970 86.605 179.100 ;
        RECT 85.850 177.775 86.130 178.725 ;
        RECT 86.300 177.865 86.470 178.970 ;
        RECT 86.640 178.185 86.880 178.780 ;
        RECT 87.050 178.715 87.580 179.080 ;
        RECT 87.050 178.015 87.220 178.715 ;
        RECT 87.750 178.635 87.920 179.250 ;
        RECT 88.090 178.895 88.260 179.695 ;
        RECT 88.430 179.195 88.680 179.525 ;
        RECT 88.905 179.225 89.790 179.395 ;
        RECT 87.750 178.545 88.260 178.635 ;
        RECT 86.300 177.735 86.525 177.865 ;
        RECT 86.695 177.795 87.220 178.015 ;
        RECT 87.390 178.375 88.260 178.545 ;
        RECT 85.935 177.145 86.185 177.605 ;
        RECT 86.355 177.595 86.525 177.735 ;
        RECT 87.390 177.595 87.560 178.375 ;
        RECT 88.090 178.305 88.260 178.375 ;
        RECT 87.770 178.125 87.970 178.155 ;
        RECT 88.430 178.125 88.600 179.195 ;
        RECT 88.770 178.305 88.960 179.025 ;
        RECT 87.770 177.825 88.600 178.125 ;
        RECT 89.130 178.095 89.450 179.055 ;
        RECT 86.355 177.425 86.690 177.595 ;
        RECT 86.885 177.425 87.560 177.595 ;
        RECT 87.880 177.145 88.250 177.645 ;
        RECT 88.430 177.595 88.600 177.825 ;
        RECT 88.985 177.765 89.450 178.095 ;
        RECT 89.620 178.385 89.790 179.225 ;
        RECT 89.970 179.195 90.285 179.695 ;
        RECT 90.515 178.965 90.855 179.525 ;
        RECT 89.960 178.590 90.855 178.965 ;
        RECT 91.025 178.685 91.195 179.695 ;
        RECT 90.665 178.385 90.855 178.590 ;
        RECT 91.365 178.635 91.695 179.480 ;
        RECT 92.905 178.635 93.235 179.480 ;
        RECT 93.405 178.685 93.575 179.695 ;
        RECT 93.745 178.965 94.085 179.525 ;
        RECT 94.315 179.195 94.630 179.695 ;
        RECT 94.810 179.225 95.695 179.395 ;
        RECT 91.365 178.555 91.755 178.635 ;
        RECT 91.540 178.505 91.755 178.555 ;
        RECT 89.620 178.055 90.495 178.385 ;
        RECT 90.665 178.055 91.415 178.385 ;
        RECT 89.620 177.595 89.790 178.055 ;
        RECT 90.665 177.885 90.865 178.055 ;
        RECT 91.585 177.925 91.755 178.505 ;
        RECT 91.530 177.885 91.755 177.925 ;
        RECT 88.430 177.425 88.835 177.595 ;
        RECT 89.005 177.425 89.790 177.595 ;
        RECT 90.065 177.145 90.275 177.675 ;
        RECT 90.535 177.360 90.865 177.885 ;
        RECT 91.375 177.800 91.755 177.885 ;
        RECT 92.845 178.555 93.235 178.635 ;
        RECT 93.745 178.590 94.640 178.965 ;
        RECT 92.845 178.505 93.060 178.555 ;
        RECT 92.845 177.925 93.015 178.505 ;
        RECT 93.745 178.385 93.935 178.590 ;
        RECT 94.810 178.385 94.980 179.225 ;
        RECT 95.920 179.195 96.170 179.525 ;
        RECT 93.185 178.055 93.935 178.385 ;
        RECT 94.105 178.055 94.980 178.385 ;
        RECT 92.845 177.885 93.070 177.925 ;
        RECT 93.735 177.885 93.935 178.055 ;
        RECT 92.845 177.800 93.225 177.885 ;
        RECT 91.035 177.145 91.205 177.755 ;
        RECT 91.375 177.365 91.705 177.800 ;
        RECT 92.895 177.365 93.225 177.800 ;
        RECT 93.395 177.145 93.565 177.755 ;
        RECT 93.735 177.360 94.065 177.885 ;
        RECT 94.325 177.145 94.535 177.675 ;
        RECT 94.810 177.595 94.980 178.055 ;
        RECT 95.150 178.095 95.470 179.055 ;
        RECT 95.640 178.305 95.830 179.025 ;
        RECT 96.000 178.125 96.170 179.195 ;
        RECT 96.340 178.895 96.510 179.695 ;
        RECT 96.680 179.250 97.785 179.420 ;
        RECT 96.680 178.635 96.850 179.250 ;
        RECT 97.995 179.100 98.245 179.525 ;
        RECT 98.415 179.235 98.680 179.695 ;
        RECT 97.020 178.715 97.550 179.080 ;
        RECT 97.995 178.970 98.300 179.100 ;
        RECT 96.340 178.545 96.850 178.635 ;
        RECT 96.340 178.375 97.210 178.545 ;
        RECT 96.340 178.305 96.510 178.375 ;
        RECT 96.630 178.125 96.830 178.155 ;
        RECT 95.150 177.765 95.615 178.095 ;
        RECT 96.000 177.825 96.830 178.125 ;
        RECT 96.000 177.595 96.170 177.825 ;
        RECT 94.810 177.425 95.595 177.595 ;
        RECT 95.765 177.425 96.170 177.595 ;
        RECT 96.350 177.145 96.720 177.645 ;
        RECT 97.040 177.595 97.210 178.375 ;
        RECT 97.380 178.015 97.550 178.715 ;
        RECT 97.720 178.185 97.960 178.780 ;
        RECT 97.380 177.795 97.905 178.015 ;
        RECT 98.130 177.865 98.300 178.970 ;
        RECT 98.075 177.735 98.300 177.865 ;
        RECT 98.470 177.775 98.750 178.725 ;
        RECT 98.075 177.595 98.245 177.735 ;
        RECT 97.040 177.425 97.715 177.595 ;
        RECT 97.910 177.425 98.245 177.595 ;
        RECT 98.415 177.145 98.665 177.605 ;
        RECT 98.920 177.405 99.105 179.525 ;
        RECT 99.275 179.195 99.605 179.695 ;
        RECT 99.775 179.025 99.945 179.525 ;
        RECT 99.280 178.855 99.945 179.025 ;
        RECT 99.280 177.865 99.510 178.855 ;
        RECT 99.680 178.035 100.030 178.685 ;
        RECT 100.210 178.555 100.545 179.525 ;
        RECT 100.715 178.555 100.885 179.695 ;
        RECT 101.055 179.355 103.085 179.525 ;
        RECT 100.210 177.885 100.380 178.555 ;
        RECT 101.055 178.385 101.225 179.355 ;
        RECT 100.550 178.055 100.805 178.385 ;
        RECT 101.030 178.055 101.225 178.385 ;
        RECT 101.395 179.015 102.520 179.185 ;
        RECT 100.635 177.885 100.805 178.055 ;
        RECT 101.395 177.885 101.565 179.015 ;
        RECT 99.280 177.695 99.945 177.865 ;
        RECT 99.275 177.145 99.605 177.525 ;
        RECT 99.775 177.405 99.945 177.695 ;
        RECT 100.210 177.315 100.465 177.885 ;
        RECT 100.635 177.715 101.565 177.885 ;
        RECT 101.735 178.675 102.745 178.845 ;
        RECT 101.735 177.875 101.905 178.675 ;
        RECT 101.390 177.680 101.565 177.715 ;
        RECT 100.635 177.145 100.965 177.545 ;
        RECT 101.390 177.315 101.920 177.680 ;
        RECT 102.110 177.655 102.385 178.475 ;
        RECT 102.105 177.485 102.385 177.655 ;
        RECT 102.110 177.315 102.385 177.485 ;
        RECT 102.555 177.315 102.745 178.675 ;
        RECT 102.915 178.690 103.085 179.355 ;
        RECT 103.255 178.935 103.425 179.695 ;
        RECT 103.660 178.935 104.175 179.345 ;
        RECT 102.915 178.500 103.665 178.690 ;
        RECT 103.835 178.125 104.175 178.935 ;
        RECT 104.345 178.605 106.935 179.695 ;
        RECT 102.945 177.955 104.175 178.125 ;
        RECT 102.925 177.145 103.435 177.680 ;
        RECT 103.655 177.350 103.900 177.955 ;
        RECT 104.345 177.915 105.555 178.435 ;
        RECT 105.725 178.085 106.935 178.605 ;
        RECT 107.565 178.530 107.855 179.695 ;
        RECT 108.025 178.845 108.285 179.525 ;
        RECT 108.455 178.915 108.705 179.695 ;
        RECT 108.955 179.145 109.205 179.525 ;
        RECT 109.375 179.315 109.730 179.695 ;
        RECT 110.735 179.305 111.070 179.525 ;
        RECT 110.335 179.145 110.565 179.185 ;
        RECT 108.955 178.945 110.565 179.145 ;
        RECT 108.955 178.935 109.790 178.945 ;
        RECT 110.380 178.855 110.565 178.945 ;
        RECT 104.345 177.145 106.935 177.915 ;
        RECT 107.565 177.145 107.855 177.870 ;
        RECT 108.025 177.655 108.195 178.845 ;
        RECT 109.895 178.745 110.225 178.775 ;
        RECT 108.425 178.685 110.225 178.745 ;
        RECT 110.815 178.685 111.070 179.305 ;
        RECT 111.245 179.260 116.590 179.695 ;
        RECT 108.365 178.575 111.070 178.685 ;
        RECT 108.365 178.540 108.565 178.575 ;
        RECT 108.365 177.965 108.535 178.540 ;
        RECT 109.895 178.515 111.070 178.575 ;
        RECT 108.765 178.100 109.175 178.405 ;
        RECT 109.345 178.135 109.675 178.345 ;
        RECT 108.365 177.845 108.635 177.965 ;
        RECT 108.365 177.800 109.210 177.845 ;
        RECT 108.455 177.675 109.210 177.800 ;
        RECT 109.465 177.735 109.675 178.135 ;
        RECT 109.920 178.135 110.395 178.345 ;
        RECT 110.585 178.135 111.075 178.335 ;
        RECT 109.920 177.735 110.140 178.135 ;
        RECT 108.025 177.645 108.255 177.655 ;
        RECT 108.025 177.315 108.285 177.645 ;
        RECT 109.040 177.525 109.210 177.675 ;
        RECT 108.455 177.145 108.785 177.505 ;
        RECT 109.040 177.315 110.340 177.525 ;
        RECT 110.615 177.145 111.070 177.910 ;
        RECT 112.830 177.690 113.170 178.520 ;
        RECT 114.650 178.010 115.000 179.260 ;
        RECT 116.825 178.635 117.155 179.480 ;
        RECT 117.325 178.685 117.495 179.695 ;
        RECT 117.665 178.965 118.005 179.525 ;
        RECT 118.235 179.195 118.550 179.695 ;
        RECT 118.730 179.225 119.615 179.395 ;
        RECT 116.765 178.555 117.155 178.635 ;
        RECT 117.665 178.590 118.560 178.965 ;
        RECT 116.765 178.505 116.980 178.555 ;
        RECT 116.765 177.925 116.935 178.505 ;
        RECT 117.665 178.385 117.855 178.590 ;
        RECT 118.730 178.385 118.900 179.225 ;
        RECT 119.840 179.195 120.090 179.525 ;
        RECT 117.105 178.055 117.855 178.385 ;
        RECT 118.025 178.055 118.900 178.385 ;
        RECT 116.765 177.885 116.990 177.925 ;
        RECT 117.655 177.885 117.855 178.055 ;
        RECT 116.765 177.800 117.145 177.885 ;
        RECT 111.245 177.145 116.590 177.690 ;
        RECT 116.815 177.365 117.145 177.800 ;
        RECT 117.315 177.145 117.485 177.755 ;
        RECT 117.655 177.360 117.985 177.885 ;
        RECT 118.245 177.145 118.455 177.675 ;
        RECT 118.730 177.595 118.900 178.055 ;
        RECT 119.070 178.095 119.390 179.055 ;
        RECT 119.560 178.305 119.750 179.025 ;
        RECT 119.920 178.125 120.090 179.195 ;
        RECT 120.260 178.895 120.430 179.695 ;
        RECT 120.600 179.250 121.705 179.420 ;
        RECT 120.600 178.635 120.770 179.250 ;
        RECT 121.915 179.100 122.165 179.525 ;
        RECT 122.335 179.235 122.600 179.695 ;
        RECT 120.940 178.715 121.470 179.080 ;
        RECT 121.915 178.970 122.220 179.100 ;
        RECT 120.260 178.545 120.770 178.635 ;
        RECT 120.260 178.375 121.130 178.545 ;
        RECT 120.260 178.305 120.430 178.375 ;
        RECT 120.550 178.125 120.750 178.155 ;
        RECT 119.070 177.765 119.535 178.095 ;
        RECT 119.920 177.825 120.750 178.125 ;
        RECT 119.920 177.595 120.090 177.825 ;
        RECT 118.730 177.425 119.515 177.595 ;
        RECT 119.685 177.425 120.090 177.595 ;
        RECT 120.270 177.145 120.640 177.645 ;
        RECT 120.960 177.595 121.130 178.375 ;
        RECT 121.300 178.015 121.470 178.715 ;
        RECT 121.640 178.185 121.880 178.780 ;
        RECT 121.300 177.795 121.825 178.015 ;
        RECT 122.050 177.865 122.220 178.970 ;
        RECT 121.995 177.735 122.220 177.865 ;
        RECT 122.390 177.775 122.670 178.725 ;
        RECT 121.995 177.595 122.165 177.735 ;
        RECT 120.960 177.425 121.635 177.595 ;
        RECT 121.830 177.425 122.165 177.595 ;
        RECT 122.335 177.145 122.585 177.605 ;
        RECT 122.840 177.405 123.025 179.525 ;
        RECT 123.195 179.195 123.525 179.695 ;
        RECT 123.695 179.025 123.865 179.525 ;
        RECT 123.200 178.855 123.865 179.025 ;
        RECT 123.200 177.865 123.430 178.855 ;
        RECT 124.125 178.845 124.385 179.525 ;
        RECT 124.555 178.915 124.805 179.695 ;
        RECT 125.055 179.145 125.305 179.525 ;
        RECT 125.475 179.315 125.830 179.695 ;
        RECT 126.835 179.305 127.170 179.525 ;
        RECT 126.435 179.145 126.665 179.185 ;
        RECT 125.055 178.945 126.665 179.145 ;
        RECT 125.055 178.935 125.890 178.945 ;
        RECT 126.480 178.855 126.665 178.945 ;
        RECT 123.600 178.035 123.950 178.685 ;
        RECT 123.200 177.695 123.865 177.865 ;
        RECT 123.195 177.145 123.525 177.525 ;
        RECT 123.695 177.405 123.865 177.695 ;
        RECT 124.125 177.645 124.295 178.845 ;
        RECT 125.995 178.745 126.325 178.775 ;
        RECT 124.525 178.685 126.325 178.745 ;
        RECT 126.915 178.685 127.170 179.305 ;
        RECT 124.465 178.575 127.170 178.685 ;
        RECT 124.465 178.540 124.665 178.575 ;
        RECT 124.465 177.965 124.635 178.540 ;
        RECT 125.995 178.515 127.170 178.575 ;
        RECT 127.350 178.555 127.625 179.525 ;
        RECT 127.835 178.895 128.115 179.695 ;
        RECT 128.285 179.185 129.475 179.475 ;
        RECT 129.735 179.355 130.895 179.525 ;
        RECT 128.285 178.845 129.455 179.015 ;
        RECT 129.735 178.855 129.905 179.355 ;
        RECT 128.285 178.725 128.455 178.845 ;
        RECT 127.795 178.555 128.455 178.725 ;
        RECT 124.865 178.100 125.275 178.405 ;
        RECT 125.445 178.135 125.775 178.345 ;
        RECT 124.465 177.845 124.735 177.965 ;
        RECT 124.465 177.800 125.310 177.845 ;
        RECT 124.555 177.675 125.310 177.800 ;
        RECT 125.565 177.735 125.775 178.135 ;
        RECT 126.020 178.135 126.495 178.345 ;
        RECT 126.685 178.135 127.175 178.335 ;
        RECT 126.020 177.735 126.240 178.135 ;
        RECT 124.125 177.315 124.385 177.645 ;
        RECT 125.140 177.525 125.310 177.675 ;
        RECT 124.555 177.145 124.885 177.505 ;
        RECT 125.140 177.315 126.440 177.525 ;
        RECT 126.715 177.145 127.170 177.910 ;
        RECT 127.350 177.820 127.520 178.555 ;
        RECT 127.795 178.385 127.965 178.555 ;
        RECT 128.765 178.385 128.960 178.675 ;
        RECT 129.130 178.555 129.455 178.845 ;
        RECT 130.165 178.725 130.335 179.185 ;
        RECT 130.565 179.105 130.895 179.355 ;
        RECT 131.120 179.275 131.450 179.695 ;
        RECT 131.705 179.105 131.990 179.525 ;
        RECT 130.565 178.935 131.990 179.105 ;
        RECT 132.235 178.895 132.565 179.695 ;
        RECT 132.815 178.975 133.150 179.485 ;
        RECT 129.710 178.385 129.915 178.675 ;
        RECT 130.165 178.555 132.535 178.725 ;
        RECT 132.365 178.385 132.535 178.555 ;
        RECT 127.690 178.055 127.965 178.385 ;
        RECT 128.135 178.055 128.960 178.385 ;
        RECT 129.130 178.055 129.475 178.385 ;
        RECT 129.710 178.335 130.060 178.385 ;
        RECT 129.705 178.165 130.060 178.335 ;
        RECT 129.710 178.055 130.060 178.165 ;
        RECT 127.795 177.885 127.965 178.055 ;
        RECT 127.350 177.475 127.625 177.820 ;
        RECT 127.795 177.715 129.460 177.885 ;
        RECT 127.815 177.145 128.195 177.545 ;
        RECT 128.365 177.365 128.535 177.715 ;
        RECT 128.705 177.145 129.035 177.545 ;
        RECT 129.205 177.365 129.460 177.715 ;
        RECT 129.655 177.145 129.985 177.865 ;
        RECT 130.370 177.720 130.790 178.385 ;
        RECT 130.960 177.995 131.250 178.385 ;
        RECT 131.440 177.995 131.710 178.385 ;
        RECT 131.920 178.335 132.170 178.385 ;
        RECT 131.920 178.165 132.175 178.335 ;
        RECT 131.920 178.055 132.170 178.165 ;
        RECT 132.365 178.055 132.670 178.385 ;
        RECT 130.960 177.825 131.255 177.995 ;
        RECT 131.440 177.825 131.715 177.995 ;
        RECT 132.365 177.885 132.535 178.055 ;
        RECT 130.960 177.725 131.250 177.825 ;
        RECT 131.440 177.725 131.710 177.825 ;
        RECT 131.975 177.715 132.535 177.885 ;
        RECT 131.975 177.545 132.145 177.715 ;
        RECT 132.895 177.620 133.150 178.975 ;
        RECT 133.325 178.530 133.615 179.695 ;
        RECT 133.875 179.025 134.045 179.525 ;
        RECT 134.215 179.195 134.545 179.695 ;
        RECT 133.875 178.855 134.540 179.025 ;
        RECT 133.790 178.035 134.140 178.685 ;
        RECT 130.530 177.375 132.145 177.545 ;
        RECT 132.315 177.145 132.645 177.545 ;
        RECT 132.815 177.360 133.150 177.620 ;
        RECT 133.325 177.145 133.615 177.870 ;
        RECT 134.310 177.865 134.540 178.855 ;
        RECT 133.875 177.695 134.540 177.865 ;
        RECT 133.875 177.405 134.045 177.695 ;
        RECT 134.215 177.145 134.545 177.525 ;
        RECT 134.715 177.405 134.900 179.525 ;
        RECT 135.140 179.235 135.405 179.695 ;
        RECT 135.575 179.100 135.825 179.525 ;
        RECT 136.035 179.250 137.140 179.420 ;
        RECT 135.520 178.970 135.825 179.100 ;
        RECT 135.070 177.775 135.350 178.725 ;
        RECT 135.520 177.865 135.690 178.970 ;
        RECT 135.860 178.185 136.100 178.780 ;
        RECT 136.270 178.715 136.800 179.080 ;
        RECT 136.270 178.015 136.440 178.715 ;
        RECT 136.970 178.635 137.140 179.250 ;
        RECT 137.310 178.895 137.480 179.695 ;
        RECT 137.650 179.195 137.900 179.525 ;
        RECT 138.125 179.225 139.010 179.395 ;
        RECT 136.970 178.545 137.480 178.635 ;
        RECT 135.520 177.735 135.745 177.865 ;
        RECT 135.915 177.795 136.440 178.015 ;
        RECT 136.610 178.375 137.480 178.545 ;
        RECT 135.155 177.145 135.405 177.605 ;
        RECT 135.575 177.595 135.745 177.735 ;
        RECT 136.610 177.595 136.780 178.375 ;
        RECT 137.310 178.305 137.480 178.375 ;
        RECT 136.990 178.125 137.190 178.155 ;
        RECT 137.650 178.125 137.820 179.195 ;
        RECT 137.990 178.305 138.180 179.025 ;
        RECT 136.990 177.825 137.820 178.125 ;
        RECT 138.350 178.095 138.670 179.055 ;
        RECT 135.575 177.425 135.910 177.595 ;
        RECT 136.105 177.425 136.780 177.595 ;
        RECT 137.100 177.145 137.470 177.645 ;
        RECT 137.650 177.595 137.820 177.825 ;
        RECT 138.205 177.765 138.670 178.095 ;
        RECT 138.840 178.385 139.010 179.225 ;
        RECT 139.190 179.195 139.505 179.695 ;
        RECT 139.735 178.965 140.075 179.525 ;
        RECT 139.180 178.590 140.075 178.965 ;
        RECT 140.245 178.685 140.415 179.695 ;
        RECT 139.885 178.385 140.075 178.590 ;
        RECT 140.585 178.635 140.915 179.480 ;
        RECT 141.145 178.845 141.405 179.525 ;
        RECT 141.575 178.915 141.825 179.695 ;
        RECT 142.075 179.145 142.325 179.525 ;
        RECT 142.495 179.315 142.850 179.695 ;
        RECT 143.855 179.305 144.190 179.525 ;
        RECT 143.455 179.145 143.685 179.185 ;
        RECT 142.075 178.945 143.685 179.145 ;
        RECT 142.075 178.935 142.910 178.945 ;
        RECT 143.500 178.855 143.685 178.945 ;
        RECT 140.585 178.555 140.975 178.635 ;
        RECT 140.760 178.505 140.975 178.555 ;
        RECT 138.840 178.055 139.715 178.385 ;
        RECT 139.885 178.055 140.635 178.385 ;
        RECT 138.840 177.595 139.010 178.055 ;
        RECT 139.885 177.885 140.085 178.055 ;
        RECT 140.805 177.925 140.975 178.505 ;
        RECT 140.750 177.885 140.975 177.925 ;
        RECT 137.650 177.425 138.055 177.595 ;
        RECT 138.225 177.425 139.010 177.595 ;
        RECT 139.285 177.145 139.495 177.675 ;
        RECT 139.755 177.360 140.085 177.885 ;
        RECT 140.595 177.800 140.975 177.885 ;
        RECT 140.255 177.145 140.425 177.755 ;
        RECT 140.595 177.365 140.925 177.800 ;
        RECT 141.145 177.645 141.315 178.845 ;
        RECT 143.015 178.745 143.345 178.775 ;
        RECT 141.545 178.685 143.345 178.745 ;
        RECT 143.935 178.685 144.190 179.305 ;
        RECT 141.485 178.575 144.190 178.685 ;
        RECT 144.365 178.605 145.575 179.695 ;
        RECT 141.485 178.540 141.685 178.575 ;
        RECT 141.485 177.965 141.655 178.540 ;
        RECT 143.015 178.515 144.190 178.575 ;
        RECT 141.885 178.100 142.295 178.405 ;
        RECT 142.465 178.135 142.795 178.345 ;
        RECT 141.485 177.845 141.755 177.965 ;
        RECT 141.485 177.800 142.330 177.845 ;
        RECT 141.575 177.675 142.330 177.800 ;
        RECT 142.585 177.735 142.795 178.135 ;
        RECT 143.040 178.135 143.515 178.345 ;
        RECT 143.705 178.135 144.195 178.335 ;
        RECT 143.040 177.735 143.260 178.135 ;
        RECT 141.145 177.315 141.405 177.645 ;
        RECT 142.160 177.525 142.330 177.675 ;
        RECT 141.575 177.145 141.905 177.505 ;
        RECT 142.160 177.315 143.460 177.525 ;
        RECT 143.735 177.145 144.190 177.910 ;
        RECT 144.365 177.895 144.885 178.435 ;
        RECT 145.055 178.065 145.575 178.605 ;
        RECT 145.745 178.605 146.955 179.695 ;
        RECT 145.745 178.065 146.265 178.605 ;
        RECT 146.435 177.895 146.955 178.435 ;
        RECT 144.365 177.145 145.575 177.895 ;
        RECT 145.745 177.145 146.955 177.895 ;
        RECT 17.320 176.975 147.040 177.145 ;
        RECT 17.405 176.225 18.615 176.975 ;
        RECT 19.795 176.425 19.965 176.715 ;
        RECT 20.135 176.595 20.465 176.975 ;
        RECT 19.795 176.255 20.460 176.425 ;
        RECT 17.405 175.685 17.925 176.225 ;
        RECT 18.095 175.515 18.615 176.055 ;
        RECT 17.405 174.425 18.615 175.515 ;
        RECT 19.710 175.435 20.060 176.085 ;
        RECT 20.230 175.265 20.460 176.255 ;
        RECT 19.795 175.095 20.460 175.265 ;
        RECT 19.795 174.595 19.965 175.095 ;
        RECT 20.135 174.425 20.465 174.925 ;
        RECT 20.635 174.595 20.820 176.715 ;
        RECT 21.075 176.515 21.325 176.975 ;
        RECT 21.495 176.525 21.830 176.695 ;
        RECT 22.025 176.525 22.700 176.695 ;
        RECT 21.495 176.385 21.665 176.525 ;
        RECT 20.990 175.395 21.270 176.345 ;
        RECT 21.440 176.255 21.665 176.385 ;
        RECT 21.440 175.150 21.610 176.255 ;
        RECT 21.835 176.105 22.360 176.325 ;
        RECT 21.780 175.340 22.020 175.935 ;
        RECT 22.190 175.405 22.360 176.105 ;
        RECT 22.530 175.745 22.700 176.525 ;
        RECT 23.020 176.475 23.390 176.975 ;
        RECT 23.570 176.525 23.975 176.695 ;
        RECT 24.145 176.525 24.930 176.695 ;
        RECT 23.570 176.295 23.740 176.525 ;
        RECT 22.910 175.995 23.740 176.295 ;
        RECT 24.125 176.025 24.590 176.355 ;
        RECT 22.910 175.965 23.110 175.995 ;
        RECT 23.230 175.745 23.400 175.815 ;
        RECT 22.530 175.575 23.400 175.745 ;
        RECT 22.890 175.485 23.400 175.575 ;
        RECT 21.440 175.020 21.745 175.150 ;
        RECT 22.190 175.040 22.720 175.405 ;
        RECT 21.060 174.425 21.325 174.885 ;
        RECT 21.495 174.595 21.745 175.020 ;
        RECT 22.890 174.870 23.060 175.485 ;
        RECT 21.955 174.700 23.060 174.870 ;
        RECT 23.230 174.425 23.400 175.225 ;
        RECT 23.570 174.925 23.740 175.995 ;
        RECT 23.910 175.095 24.100 175.815 ;
        RECT 24.270 175.065 24.590 176.025 ;
        RECT 24.760 176.065 24.930 176.525 ;
        RECT 25.205 176.445 25.415 176.975 ;
        RECT 25.675 176.235 26.005 176.760 ;
        RECT 26.175 176.365 26.345 176.975 ;
        RECT 26.515 176.320 26.845 176.755 ;
        RECT 27.065 176.595 27.955 176.765 ;
        RECT 26.515 176.235 26.895 176.320 ;
        RECT 25.805 176.065 26.005 176.235 ;
        RECT 26.670 176.195 26.895 176.235 ;
        RECT 24.760 175.735 25.635 176.065 ;
        RECT 25.805 175.735 26.555 176.065 ;
        RECT 23.570 174.595 23.820 174.925 ;
        RECT 24.760 174.895 24.930 175.735 ;
        RECT 25.805 175.530 25.995 175.735 ;
        RECT 26.725 175.615 26.895 176.195 ;
        RECT 27.065 176.040 27.615 176.425 ;
        RECT 27.785 175.870 27.955 176.595 ;
        RECT 26.680 175.565 26.895 175.615 ;
        RECT 25.100 175.155 25.995 175.530 ;
        RECT 26.505 175.485 26.895 175.565 ;
        RECT 27.065 175.800 27.955 175.870 ;
        RECT 28.125 176.270 28.345 176.755 ;
        RECT 28.515 176.435 28.765 176.975 ;
        RECT 28.935 176.325 29.195 176.805 ;
        RECT 28.125 175.845 28.455 176.270 ;
        RECT 27.065 175.775 27.960 175.800 ;
        RECT 27.065 175.760 27.970 175.775 ;
        RECT 27.065 175.745 27.975 175.760 ;
        RECT 27.065 175.740 27.985 175.745 ;
        RECT 27.065 175.730 27.990 175.740 ;
        RECT 27.065 175.720 27.995 175.730 ;
        RECT 27.065 175.715 28.005 175.720 ;
        RECT 27.065 175.705 28.015 175.715 ;
        RECT 27.065 175.700 28.025 175.705 ;
        RECT 24.045 174.725 24.930 174.895 ;
        RECT 25.110 174.425 25.425 174.925 ;
        RECT 25.655 174.595 25.995 175.155 ;
        RECT 26.165 174.425 26.335 175.435 ;
        RECT 26.505 174.640 26.835 175.485 ;
        RECT 27.065 175.250 27.325 175.700 ;
        RECT 27.690 175.695 28.025 175.700 ;
        RECT 27.690 175.690 28.040 175.695 ;
        RECT 27.690 175.680 28.055 175.690 ;
        RECT 27.690 175.675 28.080 175.680 ;
        RECT 28.625 175.675 28.855 176.070 ;
        RECT 27.690 175.670 28.855 175.675 ;
        RECT 27.720 175.635 28.855 175.670 ;
        RECT 27.755 175.610 28.855 175.635 ;
        RECT 27.785 175.580 28.855 175.610 ;
        RECT 27.805 175.550 28.855 175.580 ;
        RECT 27.825 175.520 28.855 175.550 ;
        RECT 27.895 175.510 28.855 175.520 ;
        RECT 27.920 175.500 28.855 175.510 ;
        RECT 27.940 175.485 28.855 175.500 ;
        RECT 27.960 175.470 28.855 175.485 ;
        RECT 27.965 175.460 28.750 175.470 ;
        RECT 27.980 175.425 28.750 175.460 ;
        RECT 27.495 175.105 27.825 175.350 ;
        RECT 27.995 175.175 28.750 175.425 ;
        RECT 29.025 175.295 29.195 176.325 ;
        RECT 27.495 175.080 27.680 175.105 ;
        RECT 27.065 174.980 27.680 175.080 ;
        RECT 27.065 174.425 27.670 174.980 ;
        RECT 27.845 174.595 28.325 174.935 ;
        RECT 28.495 174.425 28.750 174.970 ;
        RECT 28.920 174.595 29.195 175.295 ;
        RECT 29.365 176.325 29.625 176.805 ;
        RECT 29.795 176.435 30.045 176.975 ;
        RECT 29.365 175.295 29.535 176.325 ;
        RECT 30.215 176.270 30.435 176.755 ;
        RECT 29.705 175.675 29.935 176.070 ;
        RECT 30.105 175.845 30.435 176.270 ;
        RECT 30.605 176.595 31.495 176.765 ;
        RECT 30.605 175.870 30.775 176.595 ;
        RECT 30.945 176.040 31.495 176.425 ;
        RECT 31.705 176.155 31.935 176.975 ;
        RECT 32.105 176.175 32.435 176.805 ;
        RECT 30.605 175.800 31.495 175.870 ;
        RECT 30.600 175.775 31.495 175.800 ;
        RECT 30.590 175.760 31.495 175.775 ;
        RECT 30.585 175.745 31.495 175.760 ;
        RECT 30.575 175.740 31.495 175.745 ;
        RECT 30.570 175.730 31.495 175.740 ;
        RECT 31.685 175.735 32.015 175.985 ;
        RECT 30.565 175.720 31.495 175.730 ;
        RECT 30.555 175.715 31.495 175.720 ;
        RECT 30.545 175.705 31.495 175.715 ;
        RECT 30.535 175.700 31.495 175.705 ;
        RECT 30.535 175.695 30.870 175.700 ;
        RECT 30.520 175.690 30.870 175.695 ;
        RECT 30.505 175.680 30.870 175.690 ;
        RECT 30.480 175.675 30.870 175.680 ;
        RECT 29.705 175.670 30.870 175.675 ;
        RECT 29.705 175.635 30.840 175.670 ;
        RECT 29.705 175.610 30.805 175.635 ;
        RECT 29.705 175.580 30.775 175.610 ;
        RECT 29.705 175.550 30.755 175.580 ;
        RECT 29.705 175.520 30.735 175.550 ;
        RECT 29.705 175.510 30.665 175.520 ;
        RECT 29.705 175.500 30.640 175.510 ;
        RECT 29.705 175.485 30.620 175.500 ;
        RECT 29.705 175.470 30.600 175.485 ;
        RECT 29.810 175.460 30.595 175.470 ;
        RECT 29.810 175.425 30.580 175.460 ;
        RECT 29.365 174.595 29.640 175.295 ;
        RECT 29.810 175.175 30.565 175.425 ;
        RECT 30.735 175.105 31.065 175.350 ;
        RECT 31.235 175.250 31.495 175.700 ;
        RECT 32.185 175.575 32.435 176.175 ;
        RECT 32.605 176.155 32.815 176.975 ;
        RECT 33.045 176.205 36.555 176.975 ;
        RECT 37.345 176.415 37.675 176.805 ;
        RECT 37.845 176.585 39.030 176.755 ;
        RECT 39.290 176.505 39.460 176.975 ;
        RECT 37.345 176.235 37.855 176.415 ;
        RECT 33.045 175.685 34.695 176.205 ;
        RECT 30.880 175.080 31.065 175.105 ;
        RECT 30.880 174.980 31.495 175.080 ;
        RECT 29.810 174.425 30.065 174.970 ;
        RECT 30.235 174.595 30.715 174.935 ;
        RECT 30.890 174.425 31.495 174.980 ;
        RECT 31.705 174.425 31.935 175.565 ;
        RECT 32.105 174.595 32.435 175.575 ;
        RECT 32.605 174.425 32.815 175.565 ;
        RECT 34.865 175.515 36.555 176.035 ;
        RECT 37.185 175.775 37.515 176.065 ;
        RECT 37.685 175.605 37.855 176.235 ;
        RECT 38.260 176.325 38.645 176.415 ;
        RECT 39.630 176.325 39.960 176.790 ;
        RECT 38.260 176.155 39.960 176.325 ;
        RECT 40.130 176.155 40.300 176.975 ;
        RECT 40.470 176.155 41.155 176.795 ;
        RECT 41.345 176.165 41.585 176.975 ;
        RECT 41.755 176.165 42.085 176.805 ;
        RECT 42.255 176.165 42.525 176.975 ;
        RECT 43.165 176.250 43.455 176.975 ;
        RECT 43.625 176.235 44.065 176.795 ;
        RECT 44.235 176.235 44.685 176.975 ;
        RECT 44.855 176.405 45.025 176.805 ;
        RECT 45.195 176.575 45.615 176.975 ;
        RECT 45.785 176.405 46.015 176.805 ;
        RECT 44.855 176.235 46.015 176.405 ;
        RECT 46.185 176.235 46.675 176.805 ;
        RECT 46.845 176.430 52.190 176.975 ;
        RECT 52.365 176.430 57.710 176.975 ;
        RECT 38.025 175.775 38.355 175.985 ;
        RECT 38.535 175.735 38.915 175.985 ;
        RECT 39.105 175.955 39.590 175.985 ;
        RECT 39.085 175.785 39.590 175.955 ;
        RECT 33.045 174.425 36.555 175.515 ;
        RECT 37.340 175.435 38.425 175.605 ;
        RECT 37.340 174.595 37.640 175.435 ;
        RECT 37.835 174.425 38.085 175.265 ;
        RECT 38.255 175.185 38.425 175.435 ;
        RECT 38.595 175.355 38.915 175.735 ;
        RECT 39.105 175.775 39.590 175.785 ;
        RECT 39.780 175.775 40.230 175.985 ;
        RECT 40.400 175.775 40.735 175.985 ;
        RECT 39.105 175.355 39.480 175.775 ;
        RECT 40.400 175.605 40.570 175.775 ;
        RECT 39.650 175.435 40.570 175.605 ;
        RECT 39.650 175.185 39.820 175.435 ;
        RECT 38.255 175.015 39.820 175.185 ;
        RECT 38.675 174.595 39.480 175.015 ;
        RECT 39.990 174.425 40.320 175.265 ;
        RECT 40.905 175.185 41.155 176.155 ;
        RECT 41.325 175.735 41.675 175.985 ;
        RECT 41.845 175.565 42.015 176.165 ;
        RECT 42.185 175.735 42.535 175.985 ;
        RECT 40.490 174.595 41.155 175.185 ;
        RECT 41.335 175.395 42.015 175.565 ;
        RECT 41.335 174.610 41.665 175.395 ;
        RECT 42.195 174.425 42.525 175.565 ;
        RECT 43.165 174.425 43.455 175.590 ;
        RECT 43.625 175.225 43.935 176.235 ;
        RECT 44.105 175.615 44.275 176.065 ;
        RECT 44.445 175.785 44.835 176.065 ;
        RECT 45.020 175.735 45.265 176.065 ;
        RECT 44.105 175.445 44.895 175.615 ;
        RECT 43.625 174.595 44.065 175.225 ;
        RECT 44.240 174.425 44.555 175.275 ;
        RECT 44.725 174.765 44.895 175.445 ;
        RECT 45.065 174.935 45.265 175.735 ;
        RECT 45.465 174.935 45.715 176.065 ;
        RECT 45.930 175.735 46.335 176.065 ;
        RECT 46.505 175.565 46.675 176.235 ;
        RECT 48.430 175.600 48.770 176.430 ;
        RECT 45.905 175.395 46.675 175.565 ;
        RECT 45.905 174.765 46.155 175.395 ;
        RECT 44.725 174.595 46.155 174.765 ;
        RECT 46.335 174.425 46.665 175.225 ;
        RECT 50.250 174.860 50.600 176.110 ;
        RECT 53.950 175.600 54.290 176.430 ;
        RECT 57.885 176.205 60.475 176.975 ;
        RECT 55.770 174.860 56.120 176.110 ;
        RECT 57.885 175.685 59.095 176.205 ;
        RECT 61.125 176.165 61.365 176.975 ;
        RECT 61.535 176.165 61.865 176.805 ;
        RECT 62.035 176.165 62.305 176.975 ;
        RECT 59.265 175.515 60.475 176.035 ;
        RECT 61.105 175.735 61.455 175.985 ;
        RECT 61.625 175.565 61.795 176.165 ;
        RECT 61.965 175.735 62.315 175.985 ;
        RECT 46.845 174.425 52.190 174.860 ;
        RECT 52.365 174.425 57.710 174.860 ;
        RECT 57.885 174.425 60.475 175.515 ;
        RECT 61.115 175.395 61.795 175.565 ;
        RECT 61.115 174.610 61.445 175.395 ;
        RECT 61.975 174.425 62.305 175.565 ;
        RECT 62.950 175.375 63.285 176.795 ;
        RECT 63.465 176.605 64.210 176.975 ;
        RECT 64.775 176.435 65.030 176.795 ;
        RECT 65.210 176.605 65.540 176.975 ;
        RECT 65.720 176.435 65.945 176.795 ;
        RECT 63.460 176.245 65.945 176.435 ;
        RECT 63.460 175.555 63.685 176.245 ;
        RECT 66.165 176.205 68.755 176.975 ;
        RECT 68.925 176.250 69.215 176.975 ;
        RECT 69.385 176.205 72.895 176.975 ;
        RECT 73.065 176.225 74.275 176.975 ;
        RECT 74.560 176.345 74.845 176.805 ;
        RECT 75.015 176.515 75.285 176.975 ;
        RECT 63.885 175.735 64.165 176.065 ;
        RECT 64.345 175.735 64.920 176.065 ;
        RECT 65.100 175.735 65.535 176.065 ;
        RECT 65.715 175.735 65.985 176.065 ;
        RECT 66.165 175.685 67.375 176.205 ;
        RECT 63.460 175.375 65.955 175.555 ;
        RECT 67.545 175.515 68.755 176.035 ;
        RECT 69.385 175.685 71.035 176.205 ;
        RECT 62.950 174.605 63.215 175.375 ;
        RECT 63.385 174.425 63.715 175.145 ;
        RECT 63.905 174.965 65.095 175.195 ;
        RECT 63.905 174.605 64.165 174.965 ;
        RECT 64.335 174.425 64.665 174.795 ;
        RECT 64.835 174.605 65.095 174.965 ;
        RECT 65.665 174.605 65.955 175.375 ;
        RECT 66.165 174.425 68.755 175.515 ;
        RECT 68.925 174.425 69.215 175.590 ;
        RECT 71.205 175.515 72.895 176.035 ;
        RECT 73.065 175.685 73.585 176.225 ;
        RECT 74.560 176.175 75.515 176.345 ;
        RECT 73.755 175.515 74.275 176.055 ;
        RECT 69.385 174.425 72.895 175.515 ;
        RECT 73.065 174.425 74.275 175.515 ;
        RECT 74.445 175.445 75.135 176.005 ;
        RECT 75.305 175.275 75.515 176.175 ;
        RECT 74.560 175.055 75.515 175.275 ;
        RECT 75.685 176.005 76.085 176.805 ;
        RECT 76.275 176.345 76.555 176.805 ;
        RECT 77.075 176.515 77.400 176.975 ;
        RECT 76.275 176.175 77.400 176.345 ;
        RECT 77.570 176.235 77.955 176.805 ;
        RECT 76.950 176.065 77.400 176.175 ;
        RECT 75.685 175.445 76.780 176.005 ;
        RECT 76.950 175.735 77.505 176.065 ;
        RECT 74.560 174.595 74.845 175.055 ;
        RECT 75.015 174.425 75.285 174.885 ;
        RECT 75.685 174.595 76.085 175.445 ;
        RECT 76.950 175.275 77.400 175.735 ;
        RECT 77.675 175.565 77.955 176.235 ;
        RECT 78.145 176.165 78.385 176.975 ;
        RECT 78.555 176.165 78.885 176.805 ;
        RECT 79.055 176.165 79.325 176.975 ;
        RECT 79.505 176.430 84.850 176.975 ;
        RECT 78.125 175.735 78.475 175.985 ;
        RECT 78.645 175.565 78.815 176.165 ;
        RECT 78.985 175.735 79.335 175.985 ;
        RECT 81.090 175.600 81.430 176.430 ;
        RECT 85.025 176.205 86.695 176.975 ;
        RECT 87.415 176.425 87.585 176.715 ;
        RECT 87.755 176.595 88.085 176.975 ;
        RECT 87.415 176.255 88.080 176.425 ;
        RECT 76.275 175.055 77.400 175.275 ;
        RECT 76.275 174.595 76.555 175.055 ;
        RECT 77.075 174.425 77.400 174.885 ;
        RECT 77.570 174.595 77.955 175.565 ;
        RECT 78.135 175.395 78.815 175.565 ;
        RECT 78.135 174.610 78.465 175.395 ;
        RECT 78.995 174.425 79.325 175.565 ;
        RECT 82.910 174.860 83.260 176.110 ;
        RECT 85.025 175.685 85.775 176.205 ;
        RECT 85.945 175.515 86.695 176.035 ;
        RECT 79.505 174.425 84.850 174.860 ;
        RECT 85.025 174.425 86.695 175.515 ;
        RECT 87.330 175.435 87.680 176.085 ;
        RECT 87.850 175.265 88.080 176.255 ;
        RECT 87.415 175.095 88.080 175.265 ;
        RECT 87.415 174.595 87.585 175.095 ;
        RECT 87.755 174.425 88.085 174.925 ;
        RECT 88.255 174.595 88.440 176.715 ;
        RECT 88.695 176.515 88.945 176.975 ;
        RECT 89.115 176.525 89.450 176.695 ;
        RECT 89.645 176.525 90.320 176.695 ;
        RECT 89.115 176.385 89.285 176.525 ;
        RECT 88.610 175.395 88.890 176.345 ;
        RECT 89.060 176.255 89.285 176.385 ;
        RECT 89.060 175.150 89.230 176.255 ;
        RECT 89.455 176.105 89.980 176.325 ;
        RECT 89.400 175.340 89.640 175.935 ;
        RECT 89.810 175.405 89.980 176.105 ;
        RECT 90.150 175.745 90.320 176.525 ;
        RECT 90.640 176.475 91.010 176.975 ;
        RECT 91.190 176.525 91.595 176.695 ;
        RECT 91.765 176.525 92.550 176.695 ;
        RECT 91.190 176.295 91.360 176.525 ;
        RECT 90.530 175.995 91.360 176.295 ;
        RECT 91.745 176.025 92.210 176.355 ;
        RECT 90.530 175.965 90.730 175.995 ;
        RECT 90.850 175.745 91.020 175.815 ;
        RECT 90.150 175.575 91.020 175.745 ;
        RECT 90.510 175.485 91.020 175.575 ;
        RECT 89.060 175.020 89.365 175.150 ;
        RECT 89.810 175.040 90.340 175.405 ;
        RECT 88.680 174.425 88.945 174.885 ;
        RECT 89.115 174.595 89.365 175.020 ;
        RECT 90.510 174.870 90.680 175.485 ;
        RECT 89.575 174.700 90.680 174.870 ;
        RECT 90.850 174.425 91.020 175.225 ;
        RECT 91.190 174.925 91.360 175.995 ;
        RECT 91.530 175.095 91.720 175.815 ;
        RECT 91.890 175.065 92.210 176.025 ;
        RECT 92.380 176.065 92.550 176.525 ;
        RECT 92.825 176.445 93.035 176.975 ;
        RECT 93.295 176.235 93.625 176.760 ;
        RECT 93.795 176.365 93.965 176.975 ;
        RECT 94.135 176.320 94.465 176.755 ;
        RECT 94.135 176.235 94.515 176.320 ;
        RECT 94.685 176.250 94.975 176.975 ;
        RECT 93.425 176.065 93.625 176.235 ;
        RECT 94.290 176.195 94.515 176.235 ;
        RECT 92.380 175.735 93.255 176.065 ;
        RECT 93.425 175.735 94.175 176.065 ;
        RECT 91.190 174.595 91.440 174.925 ;
        RECT 92.380 174.895 92.550 175.735 ;
        RECT 93.425 175.530 93.615 175.735 ;
        RECT 94.345 175.615 94.515 176.195 ;
        RECT 94.300 175.565 94.515 175.615 ;
        RECT 95.145 176.235 95.530 176.805 ;
        RECT 95.700 176.515 96.025 176.975 ;
        RECT 96.545 176.345 96.825 176.805 ;
        RECT 92.720 175.155 93.615 175.530 ;
        RECT 94.125 175.485 94.515 175.565 ;
        RECT 91.665 174.725 92.550 174.895 ;
        RECT 92.730 174.425 93.045 174.925 ;
        RECT 93.275 174.595 93.615 175.155 ;
        RECT 93.785 174.425 93.955 175.435 ;
        RECT 94.125 174.640 94.455 175.485 ;
        RECT 94.685 174.425 94.975 175.590 ;
        RECT 95.145 175.565 95.425 176.235 ;
        RECT 95.700 176.175 96.825 176.345 ;
        RECT 95.700 176.065 96.150 176.175 ;
        RECT 95.595 175.735 96.150 176.065 ;
        RECT 97.015 176.005 97.415 176.805 ;
        RECT 97.815 176.515 98.085 176.975 ;
        RECT 98.255 176.345 98.540 176.805 ;
        RECT 95.145 174.595 95.530 175.565 ;
        RECT 95.700 175.275 96.150 175.735 ;
        RECT 96.320 175.445 97.415 176.005 ;
        RECT 95.700 175.055 96.825 175.275 ;
        RECT 95.700 174.425 96.025 174.885 ;
        RECT 96.545 174.595 96.825 175.055 ;
        RECT 97.015 174.595 97.415 175.445 ;
        RECT 97.585 176.175 98.540 176.345 ;
        RECT 98.825 176.235 99.210 176.805 ;
        RECT 99.380 176.515 99.705 176.975 ;
        RECT 100.225 176.345 100.505 176.805 ;
        RECT 97.585 175.275 97.795 176.175 ;
        RECT 97.965 175.445 98.655 176.005 ;
        RECT 98.825 175.565 99.105 176.235 ;
        RECT 99.380 176.175 100.505 176.345 ;
        RECT 99.380 176.065 99.830 176.175 ;
        RECT 99.275 175.735 99.830 176.065 ;
        RECT 100.695 176.005 101.095 176.805 ;
        RECT 101.495 176.515 101.765 176.975 ;
        RECT 101.935 176.345 102.220 176.805 ;
        RECT 97.585 175.055 98.540 175.275 ;
        RECT 97.815 174.425 98.085 174.885 ;
        RECT 98.255 174.595 98.540 175.055 ;
        RECT 98.825 174.595 99.210 175.565 ;
        RECT 99.380 175.275 99.830 175.735 ;
        RECT 100.000 175.445 101.095 176.005 ;
        RECT 99.380 175.055 100.505 175.275 ;
        RECT 99.380 174.425 99.705 174.885 ;
        RECT 100.225 174.595 100.505 175.055 ;
        RECT 100.695 174.595 101.095 175.445 ;
        RECT 101.265 176.175 102.220 176.345 ;
        RECT 102.505 176.235 102.890 176.805 ;
        RECT 103.060 176.515 103.385 176.975 ;
        RECT 103.905 176.345 104.185 176.805 ;
        RECT 101.265 175.275 101.475 176.175 ;
        RECT 101.645 175.445 102.335 176.005 ;
        RECT 102.505 175.565 102.785 176.235 ;
        RECT 103.060 176.175 104.185 176.345 ;
        RECT 103.060 176.065 103.510 176.175 ;
        RECT 102.955 175.735 103.510 176.065 ;
        RECT 104.375 176.005 104.775 176.805 ;
        RECT 105.175 176.515 105.445 176.975 ;
        RECT 105.615 176.345 105.900 176.805 ;
        RECT 106.665 176.505 106.960 176.975 ;
        RECT 101.265 175.055 102.220 175.275 ;
        RECT 101.495 174.425 101.765 174.885 ;
        RECT 101.935 174.595 102.220 175.055 ;
        RECT 102.505 174.595 102.890 175.565 ;
        RECT 103.060 175.275 103.510 175.735 ;
        RECT 103.680 175.445 104.775 176.005 ;
        RECT 103.060 175.055 104.185 175.275 ;
        RECT 103.060 174.425 103.385 174.885 ;
        RECT 103.905 174.595 104.185 175.055 ;
        RECT 104.375 174.595 104.775 175.445 ;
        RECT 104.945 176.175 105.900 176.345 ;
        RECT 107.130 176.335 107.390 176.780 ;
        RECT 107.560 176.505 107.820 176.975 ;
        RECT 107.990 176.335 108.245 176.780 ;
        RECT 108.415 176.505 108.715 176.975 ;
        RECT 104.945 175.275 105.155 176.175 ;
        RECT 106.205 176.165 109.235 176.335 ;
        RECT 105.325 175.445 106.015 176.005 ;
        RECT 106.205 175.600 106.375 176.165 ;
        RECT 106.545 175.770 108.760 175.995 ;
        RECT 108.935 175.600 109.235 176.165 ;
        RECT 106.205 175.430 109.235 175.600 ;
        RECT 109.405 176.255 109.745 176.765 ;
        RECT 104.945 175.055 105.900 175.275 ;
        RECT 105.175 174.425 105.445 174.885 ;
        RECT 105.615 174.595 105.900 175.055 ;
        RECT 106.185 174.425 106.530 175.260 ;
        RECT 106.705 174.625 106.960 175.430 ;
        RECT 107.130 174.425 107.390 175.260 ;
        RECT 107.565 174.625 107.820 175.430 ;
        RECT 107.990 174.425 108.250 175.260 ;
        RECT 108.420 174.625 108.680 175.430 ;
        RECT 108.850 174.425 109.235 175.260 ;
        RECT 109.405 174.855 109.665 176.255 ;
        RECT 109.915 176.175 110.185 176.975 ;
        RECT 109.840 175.735 110.170 175.985 ;
        RECT 110.365 175.735 110.645 176.705 ;
        RECT 110.825 175.735 111.125 176.705 ;
        RECT 111.305 175.735 111.655 176.700 ;
        RECT 111.875 176.475 112.370 176.805 ;
        RECT 109.855 175.565 110.170 175.735 ;
        RECT 111.875 175.565 112.045 176.475 ;
        RECT 112.625 176.430 117.970 176.975 ;
        RECT 109.855 175.395 112.045 175.565 ;
        RECT 109.405 174.595 109.745 174.855 ;
        RECT 109.915 174.425 110.245 175.225 ;
        RECT 110.710 174.595 110.960 175.395 ;
        RECT 111.145 174.425 111.475 175.145 ;
        RECT 111.695 174.595 111.945 175.395 ;
        RECT 112.215 174.985 112.455 176.295 ;
        RECT 114.210 175.600 114.550 176.430 ;
        RECT 118.145 176.205 119.815 176.975 ;
        RECT 120.445 176.250 120.735 176.975 ;
        RECT 120.905 176.205 123.495 176.975 ;
        RECT 124.160 176.235 124.775 176.805 ;
        RECT 124.945 176.465 125.160 176.975 ;
        RECT 125.390 176.465 125.670 176.795 ;
        RECT 125.850 176.465 126.090 176.975 ;
        RECT 126.425 176.595 127.315 176.765 ;
        RECT 116.030 174.860 116.380 176.110 ;
        RECT 118.145 175.685 118.895 176.205 ;
        RECT 119.065 175.515 119.815 176.035 ;
        RECT 120.905 175.685 122.115 176.205 ;
        RECT 112.115 174.425 112.450 174.805 ;
        RECT 112.625 174.425 117.970 174.860 ;
        RECT 118.145 174.425 119.815 175.515 ;
        RECT 120.445 174.425 120.735 175.590 ;
        RECT 122.285 175.515 123.495 176.035 ;
        RECT 120.905 174.425 123.495 175.515 ;
        RECT 124.160 175.215 124.475 176.235 ;
        RECT 124.645 175.565 124.815 176.065 ;
        RECT 125.065 175.735 125.330 176.295 ;
        RECT 125.500 175.565 125.670 176.465 ;
        RECT 125.840 175.735 126.195 176.295 ;
        RECT 126.425 176.040 126.975 176.425 ;
        RECT 127.145 175.870 127.315 176.595 ;
        RECT 126.425 175.800 127.315 175.870 ;
        RECT 127.485 176.295 127.705 176.755 ;
        RECT 127.875 176.435 128.125 176.975 ;
        RECT 128.295 176.325 128.555 176.805 ;
        RECT 127.485 176.270 127.735 176.295 ;
        RECT 127.485 175.845 127.815 176.270 ;
        RECT 126.425 175.775 127.320 175.800 ;
        RECT 126.425 175.760 127.330 175.775 ;
        RECT 126.425 175.745 127.335 175.760 ;
        RECT 126.425 175.740 127.345 175.745 ;
        RECT 126.425 175.730 127.350 175.740 ;
        RECT 126.425 175.720 127.355 175.730 ;
        RECT 126.425 175.715 127.365 175.720 ;
        RECT 126.425 175.705 127.375 175.715 ;
        RECT 126.425 175.700 127.385 175.705 ;
        RECT 124.645 175.395 126.070 175.565 ;
        RECT 124.160 174.595 124.695 175.215 ;
        RECT 124.865 174.425 125.195 175.225 ;
        RECT 125.680 175.220 126.070 175.395 ;
        RECT 126.425 175.250 126.685 175.700 ;
        RECT 127.050 175.695 127.385 175.700 ;
        RECT 127.050 175.690 127.400 175.695 ;
        RECT 127.050 175.680 127.415 175.690 ;
        RECT 127.050 175.675 127.440 175.680 ;
        RECT 127.985 175.675 128.215 176.070 ;
        RECT 127.050 175.670 128.215 175.675 ;
        RECT 127.080 175.635 128.215 175.670 ;
        RECT 127.115 175.610 128.215 175.635 ;
        RECT 127.145 175.580 128.215 175.610 ;
        RECT 127.165 175.550 128.215 175.580 ;
        RECT 127.185 175.520 128.215 175.550 ;
        RECT 127.255 175.510 128.215 175.520 ;
        RECT 127.280 175.500 128.215 175.510 ;
        RECT 127.300 175.485 128.215 175.500 ;
        RECT 127.320 175.470 128.215 175.485 ;
        RECT 127.325 175.460 128.110 175.470 ;
        RECT 127.340 175.425 128.110 175.460 ;
        RECT 126.855 175.105 127.185 175.350 ;
        RECT 127.355 175.175 128.110 175.425 ;
        RECT 128.385 175.295 128.555 176.325 ;
        RECT 128.735 176.165 129.005 176.975 ;
        RECT 129.175 176.165 129.505 176.805 ;
        RECT 129.675 176.165 129.915 176.975 ;
        RECT 131.025 176.175 131.335 176.975 ;
        RECT 131.540 176.175 132.235 176.805 ;
        RECT 132.735 176.575 133.065 176.975 ;
        RECT 133.235 176.405 133.565 176.745 ;
        RECT 134.615 176.575 134.945 176.975 ;
        RECT 132.580 176.235 134.945 176.405 ;
        RECT 135.115 176.250 135.445 176.760 ;
        RECT 135.630 176.575 135.965 176.975 ;
        RECT 136.135 176.405 136.340 176.805 ;
        RECT 136.550 176.495 136.825 176.975 ;
        RECT 137.035 176.475 137.295 176.805 ;
        RECT 128.725 175.735 129.075 175.985 ;
        RECT 129.245 175.565 129.415 176.165 ;
        RECT 129.585 175.735 129.935 175.985 ;
        RECT 131.035 175.735 131.370 176.005 ;
        RECT 131.540 175.575 131.710 176.175 ;
        RECT 131.880 175.735 132.215 175.985 ;
        RECT 126.855 175.080 127.040 175.105 ;
        RECT 126.425 174.980 127.040 175.080 ;
        RECT 126.425 174.425 127.030 174.980 ;
        RECT 127.205 174.595 127.685 174.935 ;
        RECT 127.855 174.425 128.110 174.970 ;
        RECT 128.280 174.595 128.555 175.295 ;
        RECT 128.735 174.425 129.065 175.565 ;
        RECT 129.245 175.395 129.925 175.565 ;
        RECT 129.595 174.610 129.925 175.395 ;
        RECT 131.025 174.425 131.305 175.565 ;
        RECT 131.475 174.595 131.805 175.575 ;
        RECT 131.975 174.425 132.235 175.565 ;
        RECT 132.580 175.235 132.750 176.235 ;
        RECT 134.775 176.065 134.945 176.235 ;
        RECT 132.920 175.405 133.165 176.065 ;
        RECT 133.380 175.405 133.645 176.065 ;
        RECT 133.840 175.405 134.125 176.065 ;
        RECT 134.300 175.735 134.605 176.065 ;
        RECT 134.775 175.735 135.085 176.065 ;
        RECT 134.300 175.405 134.515 175.735 ;
        RECT 132.580 175.065 133.035 175.235 ;
        RECT 132.705 174.635 133.035 175.065 ;
        RECT 133.215 175.065 134.505 175.235 ;
        RECT 133.215 174.645 133.465 175.065 ;
        RECT 133.695 174.425 134.025 174.895 ;
        RECT 134.255 174.645 134.505 175.065 ;
        RECT 134.695 174.425 134.945 175.565 ;
        RECT 135.255 175.485 135.445 176.250 ;
        RECT 135.115 174.635 135.445 175.485 ;
        RECT 135.655 176.235 136.340 176.405 ;
        RECT 135.655 175.205 135.995 176.235 ;
        RECT 136.165 175.565 136.415 176.065 ;
        RECT 136.595 175.735 136.955 176.315 ;
        RECT 137.125 175.565 137.295 176.475 ;
        RECT 137.555 176.425 137.725 176.715 ;
        RECT 137.895 176.595 138.225 176.975 ;
        RECT 137.555 176.255 138.220 176.425 ;
        RECT 136.165 175.395 137.295 175.565 ;
        RECT 137.470 175.435 137.820 176.085 ;
        RECT 135.655 175.030 136.320 175.205 ;
        RECT 135.630 174.425 135.965 174.850 ;
        RECT 136.135 174.625 136.320 175.030 ;
        RECT 136.525 174.425 136.855 175.205 ;
        RECT 137.025 174.625 137.295 175.395 ;
        RECT 137.990 175.265 138.220 176.255 ;
        RECT 137.555 175.095 138.220 175.265 ;
        RECT 137.555 174.595 137.725 175.095 ;
        RECT 137.895 174.425 138.225 174.925 ;
        RECT 138.395 174.595 138.580 176.715 ;
        RECT 138.835 176.515 139.085 176.975 ;
        RECT 139.255 176.525 139.590 176.695 ;
        RECT 139.785 176.525 140.460 176.695 ;
        RECT 139.255 176.385 139.425 176.525 ;
        RECT 138.750 175.395 139.030 176.345 ;
        RECT 139.200 176.255 139.425 176.385 ;
        RECT 139.200 175.150 139.370 176.255 ;
        RECT 139.595 176.105 140.120 176.325 ;
        RECT 139.540 175.340 139.780 175.935 ;
        RECT 139.950 175.405 140.120 176.105 ;
        RECT 140.290 175.745 140.460 176.525 ;
        RECT 140.780 176.475 141.150 176.975 ;
        RECT 141.330 176.525 141.735 176.695 ;
        RECT 141.905 176.525 142.690 176.695 ;
        RECT 141.330 176.295 141.500 176.525 ;
        RECT 140.670 175.995 141.500 176.295 ;
        RECT 141.885 176.025 142.350 176.355 ;
        RECT 140.670 175.965 140.870 175.995 ;
        RECT 140.990 175.745 141.160 175.815 ;
        RECT 140.290 175.575 141.160 175.745 ;
        RECT 140.650 175.485 141.160 175.575 ;
        RECT 139.200 175.020 139.505 175.150 ;
        RECT 139.950 175.040 140.480 175.405 ;
        RECT 138.820 174.425 139.085 174.885 ;
        RECT 139.255 174.595 139.505 175.020 ;
        RECT 140.650 174.870 140.820 175.485 ;
        RECT 139.715 174.700 140.820 174.870 ;
        RECT 140.990 174.425 141.160 175.225 ;
        RECT 141.330 174.925 141.500 175.995 ;
        RECT 141.670 175.095 141.860 175.815 ;
        RECT 142.030 175.065 142.350 176.025 ;
        RECT 142.520 176.065 142.690 176.525 ;
        RECT 142.965 176.445 143.175 176.975 ;
        RECT 143.435 176.235 143.765 176.760 ;
        RECT 143.935 176.365 144.105 176.975 ;
        RECT 144.275 176.320 144.605 176.755 ;
        RECT 144.275 176.235 144.655 176.320 ;
        RECT 143.565 176.065 143.765 176.235 ;
        RECT 144.430 176.195 144.655 176.235 ;
        RECT 145.745 176.225 146.955 176.975 ;
        RECT 142.520 175.735 143.395 176.065 ;
        RECT 143.565 175.735 144.315 176.065 ;
        RECT 141.330 174.595 141.580 174.925 ;
        RECT 142.520 174.895 142.690 175.735 ;
        RECT 143.565 175.530 143.755 175.735 ;
        RECT 144.485 175.615 144.655 176.195 ;
        RECT 144.440 175.565 144.655 175.615 ;
        RECT 142.860 175.155 143.755 175.530 ;
        RECT 144.265 175.485 144.655 175.565 ;
        RECT 145.745 175.515 146.265 176.055 ;
        RECT 146.435 175.685 146.955 176.225 ;
        RECT 141.805 174.725 142.690 174.895 ;
        RECT 142.870 174.425 143.185 174.925 ;
        RECT 143.415 174.595 143.755 175.155 ;
        RECT 143.925 174.425 144.095 175.435 ;
        RECT 144.265 174.640 144.595 175.485 ;
        RECT 145.745 174.425 146.955 175.515 ;
        RECT 17.320 174.255 147.040 174.425 ;
        RECT 17.405 173.165 18.615 174.255 ;
        RECT 18.785 173.165 21.375 174.255 ;
        RECT 22.065 173.195 22.395 174.040 ;
        RECT 22.565 173.245 22.735 174.255 ;
        RECT 22.905 173.525 23.245 174.085 ;
        RECT 23.475 173.755 23.790 174.255 ;
        RECT 23.970 173.785 24.855 173.955 ;
        RECT 17.405 172.455 17.925 172.995 ;
        RECT 18.095 172.625 18.615 173.165 ;
        RECT 18.785 172.475 19.995 172.995 ;
        RECT 20.165 172.645 21.375 173.165 ;
        RECT 22.005 173.115 22.395 173.195 ;
        RECT 22.905 173.150 23.800 173.525 ;
        RECT 22.005 173.065 22.220 173.115 ;
        RECT 22.005 172.485 22.175 173.065 ;
        RECT 22.905 172.945 23.095 173.150 ;
        RECT 23.970 172.945 24.140 173.785 ;
        RECT 25.080 173.755 25.330 174.085 ;
        RECT 22.345 172.615 23.095 172.945 ;
        RECT 23.265 172.615 24.140 172.945 ;
        RECT 17.405 171.705 18.615 172.455 ;
        RECT 18.785 171.705 21.375 172.475 ;
        RECT 22.005 172.445 22.230 172.485 ;
        RECT 22.895 172.445 23.095 172.615 ;
        RECT 22.005 172.360 22.385 172.445 ;
        RECT 22.055 171.925 22.385 172.360 ;
        RECT 22.555 171.705 22.725 172.315 ;
        RECT 22.895 171.920 23.225 172.445 ;
        RECT 23.485 171.705 23.695 172.235 ;
        RECT 23.970 172.155 24.140 172.615 ;
        RECT 24.310 172.655 24.630 173.615 ;
        RECT 24.800 172.865 24.990 173.585 ;
        RECT 25.160 172.685 25.330 173.755 ;
        RECT 25.500 173.455 25.670 174.255 ;
        RECT 25.840 173.810 26.945 173.980 ;
        RECT 25.840 173.195 26.010 173.810 ;
        RECT 27.155 173.660 27.405 174.085 ;
        RECT 27.575 173.795 27.840 174.255 ;
        RECT 26.180 173.275 26.710 173.640 ;
        RECT 27.155 173.530 27.460 173.660 ;
        RECT 25.500 173.105 26.010 173.195 ;
        RECT 25.500 172.935 26.370 173.105 ;
        RECT 25.500 172.865 25.670 172.935 ;
        RECT 25.790 172.685 25.990 172.715 ;
        RECT 24.310 172.325 24.775 172.655 ;
        RECT 25.160 172.385 25.990 172.685 ;
        RECT 25.160 172.155 25.330 172.385 ;
        RECT 23.970 171.985 24.755 172.155 ;
        RECT 24.925 171.985 25.330 172.155 ;
        RECT 25.510 171.705 25.880 172.205 ;
        RECT 26.200 172.155 26.370 172.935 ;
        RECT 26.540 172.575 26.710 173.275 ;
        RECT 26.880 172.745 27.120 173.340 ;
        RECT 26.540 172.355 27.065 172.575 ;
        RECT 27.290 172.425 27.460 173.530 ;
        RECT 27.235 172.295 27.460 172.425 ;
        RECT 27.630 172.335 27.910 173.285 ;
        RECT 27.235 172.155 27.405 172.295 ;
        RECT 26.200 171.985 26.875 172.155 ;
        RECT 27.070 171.985 27.405 172.155 ;
        RECT 27.575 171.705 27.825 172.165 ;
        RECT 28.080 171.965 28.265 174.085 ;
        RECT 28.435 173.755 28.765 174.255 ;
        RECT 28.935 173.585 29.105 174.085 ;
        RECT 28.440 173.415 29.105 173.585 ;
        RECT 28.440 172.425 28.670 173.415 ;
        RECT 28.840 172.595 29.190 173.245 ;
        RECT 30.285 173.090 30.575 174.255 ;
        RECT 30.745 173.820 36.090 174.255 ;
        RECT 28.440 172.255 29.105 172.425 ;
        RECT 28.435 171.705 28.765 172.085 ;
        RECT 28.935 171.965 29.105 172.255 ;
        RECT 30.285 171.705 30.575 172.430 ;
        RECT 32.330 172.250 32.670 173.080 ;
        RECT 34.150 172.570 34.500 173.820 ;
        RECT 36.265 173.165 37.475 174.255 ;
        RECT 37.655 173.455 37.985 174.255 ;
        RECT 38.165 173.915 39.595 174.085 ;
        RECT 38.165 173.285 38.415 173.915 ;
        RECT 36.265 172.455 36.785 172.995 ;
        RECT 36.955 172.625 37.475 173.165 ;
        RECT 37.645 173.115 38.415 173.285 ;
        RECT 30.745 171.705 36.090 172.250 ;
        RECT 36.265 171.705 37.475 172.455 ;
        RECT 37.645 172.445 37.815 173.115 ;
        RECT 37.985 172.615 38.390 172.945 ;
        RECT 38.605 172.615 38.855 173.745 ;
        RECT 39.055 172.945 39.255 173.745 ;
        RECT 39.425 173.235 39.595 173.915 ;
        RECT 39.765 173.405 40.080 174.255 ;
        RECT 40.255 173.455 40.695 174.085 ;
        RECT 39.425 173.065 40.215 173.235 ;
        RECT 39.055 172.615 39.300 172.945 ;
        RECT 39.485 172.615 39.875 172.895 ;
        RECT 40.045 172.615 40.215 173.065 ;
        RECT 40.385 172.445 40.695 173.455 ;
        RECT 37.645 171.875 38.135 172.445 ;
        RECT 38.305 172.275 39.465 172.445 ;
        RECT 38.305 171.875 38.535 172.275 ;
        RECT 38.705 171.705 39.125 172.105 ;
        RECT 39.295 171.875 39.465 172.275 ;
        RECT 39.635 171.705 40.085 172.445 ;
        RECT 40.255 171.885 40.695 172.445 ;
        RECT 40.865 173.145 41.125 174.085 ;
        RECT 41.295 173.855 41.625 174.255 ;
        RECT 42.770 173.990 43.025 174.085 ;
        RECT 41.885 173.820 43.025 173.990 ;
        RECT 43.195 173.875 43.525 174.045 ;
        RECT 41.885 173.595 42.055 173.820 ;
        RECT 41.295 173.425 42.055 173.595 ;
        RECT 42.770 173.685 43.025 173.820 ;
        RECT 40.865 172.430 41.040 173.145 ;
        RECT 41.295 172.945 41.465 173.425 ;
        RECT 42.320 173.335 42.490 173.525 ;
        RECT 42.770 173.515 43.180 173.685 ;
        RECT 41.210 172.615 41.465 172.945 ;
        RECT 41.690 172.615 42.020 173.235 ;
        RECT 42.320 173.165 42.840 173.335 ;
        RECT 42.190 172.615 42.480 172.995 ;
        RECT 42.670 172.445 42.840 173.165 ;
        RECT 40.865 171.875 41.125 172.430 ;
        RECT 41.960 172.275 42.840 172.445 ;
        RECT 43.010 172.490 43.180 173.515 ;
        RECT 43.355 173.625 43.525 173.875 ;
        RECT 43.695 173.795 43.945 174.255 ;
        RECT 44.115 173.625 44.295 174.085 ;
        RECT 43.355 173.455 44.295 173.625 ;
        RECT 43.380 172.975 43.860 173.275 ;
        RECT 43.010 172.320 43.360 172.490 ;
        RECT 43.600 172.385 43.860 172.975 ;
        RECT 44.060 172.385 44.320 173.275 ;
        RECT 44.545 173.115 44.825 174.255 ;
        RECT 44.995 173.105 45.325 174.085 ;
        RECT 45.495 173.115 45.755 174.255 ;
        RECT 46.445 173.195 46.775 174.040 ;
        RECT 46.945 173.245 47.115 174.255 ;
        RECT 47.285 173.525 47.625 174.085 ;
        RECT 47.855 173.755 48.170 174.255 ;
        RECT 48.350 173.785 49.235 173.955 ;
        RECT 46.385 173.115 46.775 173.195 ;
        RECT 47.285 173.150 48.180 173.525 ;
        RECT 44.555 172.675 44.890 172.945 ;
        RECT 45.060 172.505 45.230 173.105 ;
        RECT 46.385 173.065 46.600 173.115 ;
        RECT 45.400 172.695 45.735 172.945 ;
        RECT 41.295 171.705 41.725 172.150 ;
        RECT 41.960 171.875 42.130 172.275 ;
        RECT 42.300 171.705 43.020 172.105 ;
        RECT 43.190 171.875 43.360 172.320 ;
        RECT 43.935 171.705 44.335 172.215 ;
        RECT 44.545 171.705 44.855 172.505 ;
        RECT 45.060 171.875 45.755 172.505 ;
        RECT 46.385 172.485 46.555 173.065 ;
        RECT 47.285 172.945 47.475 173.150 ;
        RECT 48.350 172.945 48.520 173.785 ;
        RECT 49.460 173.755 49.710 174.085 ;
        RECT 46.725 172.615 47.475 172.945 ;
        RECT 47.645 172.615 48.520 172.945 ;
        RECT 46.385 172.445 46.610 172.485 ;
        RECT 47.275 172.445 47.475 172.615 ;
        RECT 46.385 172.360 46.765 172.445 ;
        RECT 46.435 171.925 46.765 172.360 ;
        RECT 46.935 171.705 47.105 172.315 ;
        RECT 47.275 171.920 47.605 172.445 ;
        RECT 47.865 171.705 48.075 172.235 ;
        RECT 48.350 172.155 48.520 172.615 ;
        RECT 48.690 172.655 49.010 173.615 ;
        RECT 49.180 172.865 49.370 173.585 ;
        RECT 49.540 172.685 49.710 173.755 ;
        RECT 49.880 173.455 50.050 174.255 ;
        RECT 50.220 173.810 51.325 173.980 ;
        RECT 50.220 173.195 50.390 173.810 ;
        RECT 51.535 173.660 51.785 174.085 ;
        RECT 51.955 173.795 52.220 174.255 ;
        RECT 50.560 173.275 51.090 173.640 ;
        RECT 51.535 173.530 51.840 173.660 ;
        RECT 49.880 173.105 50.390 173.195 ;
        RECT 49.880 172.935 50.750 173.105 ;
        RECT 49.880 172.865 50.050 172.935 ;
        RECT 50.170 172.685 50.370 172.715 ;
        RECT 48.690 172.325 49.155 172.655 ;
        RECT 49.540 172.385 50.370 172.685 ;
        RECT 49.540 172.155 49.710 172.385 ;
        RECT 48.350 171.985 49.135 172.155 ;
        RECT 49.305 171.985 49.710 172.155 ;
        RECT 49.890 171.705 50.260 172.205 ;
        RECT 50.580 172.155 50.750 172.935 ;
        RECT 50.920 172.575 51.090 173.275 ;
        RECT 51.260 172.745 51.500 173.340 ;
        RECT 50.920 172.355 51.445 172.575 ;
        RECT 51.670 172.425 51.840 173.530 ;
        RECT 51.615 172.295 51.840 172.425 ;
        RECT 52.010 172.335 52.290 173.285 ;
        RECT 51.615 172.155 51.785 172.295 ;
        RECT 50.580 171.985 51.255 172.155 ;
        RECT 51.450 171.985 51.785 172.155 ;
        RECT 51.955 171.705 52.205 172.165 ;
        RECT 52.460 171.965 52.645 174.085 ;
        RECT 52.815 173.755 53.145 174.255 ;
        RECT 53.315 173.585 53.485 174.085 ;
        RECT 52.820 173.415 53.485 173.585 ;
        RECT 52.820 172.425 53.050 173.415 ;
        RECT 53.220 172.595 53.570 173.245 ;
        RECT 53.745 173.165 55.415 174.255 ;
        RECT 53.745 172.475 54.495 172.995 ;
        RECT 54.665 172.645 55.415 173.165 ;
        RECT 56.045 173.090 56.335 174.255 ;
        RECT 56.505 173.820 61.850 174.255 ;
        RECT 52.820 172.255 53.485 172.425 ;
        RECT 52.815 171.705 53.145 172.085 ;
        RECT 53.315 171.965 53.485 172.255 ;
        RECT 53.745 171.705 55.415 172.475 ;
        RECT 56.045 171.705 56.335 172.430 ;
        RECT 58.090 172.250 58.430 173.080 ;
        RECT 59.910 172.570 60.260 173.820 ;
        RECT 62.025 173.165 63.695 174.255 ;
        RECT 62.025 172.475 62.775 172.995 ;
        RECT 62.945 172.645 63.695 173.165 ;
        RECT 64.325 173.385 64.600 174.085 ;
        RECT 64.770 173.710 65.025 174.255 ;
        RECT 65.195 173.745 65.675 174.085 ;
        RECT 65.850 173.700 66.455 174.255 ;
        RECT 65.840 173.600 66.455 173.700 ;
        RECT 66.635 173.645 66.965 174.075 ;
        RECT 67.145 173.815 67.340 174.255 ;
        RECT 67.510 173.645 67.840 174.075 ;
        RECT 65.840 173.575 66.025 173.600 ;
        RECT 56.505 171.705 61.850 172.250 ;
        RECT 62.025 171.705 63.695 172.475 ;
        RECT 64.325 172.355 64.495 173.385 ;
        RECT 64.770 173.255 65.525 173.505 ;
        RECT 65.695 173.330 66.025 173.575 ;
        RECT 66.635 173.475 67.840 173.645 ;
        RECT 64.770 173.220 65.540 173.255 ;
        RECT 64.770 173.210 65.555 173.220 ;
        RECT 64.665 173.195 65.560 173.210 ;
        RECT 64.665 173.180 65.580 173.195 ;
        RECT 64.665 173.170 65.600 173.180 ;
        RECT 64.665 173.160 65.625 173.170 ;
        RECT 64.665 173.130 65.695 173.160 ;
        RECT 64.665 173.100 65.715 173.130 ;
        RECT 64.665 173.070 65.735 173.100 ;
        RECT 64.665 173.045 65.765 173.070 ;
        RECT 64.665 173.010 65.800 173.045 ;
        RECT 64.665 173.005 65.830 173.010 ;
        RECT 64.665 172.610 64.895 173.005 ;
        RECT 65.440 173.000 65.830 173.005 ;
        RECT 65.465 172.990 65.830 173.000 ;
        RECT 65.480 172.985 65.830 172.990 ;
        RECT 65.495 172.980 65.830 172.985 ;
        RECT 66.195 172.980 66.455 173.430 ;
        RECT 66.635 173.145 67.530 173.475 ;
        RECT 68.010 173.305 68.285 174.075 ;
        RECT 65.495 172.975 66.455 172.980 ;
        RECT 65.505 172.965 66.455 172.975 ;
        RECT 65.515 172.960 66.455 172.965 ;
        RECT 65.525 172.950 66.455 172.960 ;
        RECT 65.530 172.940 66.455 172.950 ;
        RECT 67.700 173.115 68.285 173.305 ;
        RECT 68.475 173.285 68.805 174.070 ;
        RECT 68.475 173.115 69.155 173.285 ;
        RECT 69.335 173.115 69.665 174.255 ;
        RECT 70.965 173.585 71.245 174.255 ;
        RECT 71.415 173.365 71.715 173.915 ;
        RECT 71.915 173.535 72.245 174.255 ;
        RECT 72.435 173.535 72.895 174.085 ;
        RECT 65.535 172.935 66.455 172.940 ;
        RECT 65.545 172.920 66.455 172.935 ;
        RECT 65.550 172.905 66.455 172.920 ;
        RECT 65.560 172.880 66.455 172.905 ;
        RECT 65.065 172.410 65.395 172.835 ;
        RECT 65.145 172.385 65.395 172.410 ;
        RECT 64.325 171.875 64.585 172.355 ;
        RECT 64.755 171.705 65.005 172.245 ;
        RECT 65.175 171.925 65.395 172.385 ;
        RECT 65.565 172.810 66.455 172.880 ;
        RECT 65.565 172.085 65.735 172.810 ;
        RECT 65.905 172.255 66.455 172.640 ;
        RECT 66.640 172.615 66.935 172.945 ;
        RECT 67.115 172.615 67.530 172.945 ;
        RECT 65.565 171.915 66.455 172.085 ;
        RECT 66.635 171.705 66.935 172.435 ;
        RECT 67.115 171.995 67.345 172.615 ;
        RECT 67.700 172.445 67.875 173.115 ;
        RECT 67.545 172.265 67.875 172.445 ;
        RECT 68.045 172.295 68.285 172.945 ;
        RECT 68.465 172.695 68.815 172.945 ;
        RECT 68.985 172.515 69.155 173.115 ;
        RECT 70.780 172.945 71.045 173.305 ;
        RECT 71.415 173.195 72.355 173.365 ;
        RECT 72.185 172.945 72.355 173.195 ;
        RECT 69.325 172.695 69.675 172.945 ;
        RECT 70.780 172.695 71.455 172.945 ;
        RECT 71.675 172.695 72.015 172.945 ;
        RECT 72.185 172.615 72.475 172.945 ;
        RECT 72.185 172.525 72.355 172.615 ;
        RECT 67.545 171.885 67.770 172.265 ;
        RECT 67.940 171.705 68.270 172.095 ;
        RECT 68.485 171.705 68.725 172.515 ;
        RECT 68.895 171.875 69.225 172.515 ;
        RECT 69.395 171.705 69.665 172.515 ;
        RECT 70.965 172.335 72.355 172.525 ;
        RECT 70.965 171.975 71.295 172.335 ;
        RECT 72.645 172.165 72.895 173.535 ;
        RECT 73.125 173.195 73.455 174.040 ;
        RECT 73.625 173.245 73.795 174.255 ;
        RECT 73.965 173.525 74.305 174.085 ;
        RECT 74.535 173.755 74.850 174.255 ;
        RECT 75.030 173.785 75.915 173.955 ;
        RECT 73.065 173.115 73.455 173.195 ;
        RECT 73.965 173.150 74.860 173.525 ;
        RECT 73.065 173.065 73.280 173.115 ;
        RECT 73.065 172.485 73.235 173.065 ;
        RECT 73.965 172.945 74.155 173.150 ;
        RECT 75.030 172.945 75.200 173.785 ;
        RECT 76.140 173.755 76.390 174.085 ;
        RECT 73.405 172.615 74.155 172.945 ;
        RECT 74.325 172.615 75.200 172.945 ;
        RECT 73.065 172.445 73.290 172.485 ;
        RECT 73.955 172.445 74.155 172.615 ;
        RECT 73.065 172.360 73.445 172.445 ;
        RECT 71.915 171.705 72.165 172.165 ;
        RECT 72.335 171.875 72.895 172.165 ;
        RECT 73.115 171.925 73.445 172.360 ;
        RECT 73.615 171.705 73.785 172.315 ;
        RECT 73.955 171.920 74.285 172.445 ;
        RECT 74.545 171.705 74.755 172.235 ;
        RECT 75.030 172.155 75.200 172.615 ;
        RECT 75.370 172.655 75.690 173.615 ;
        RECT 75.860 172.865 76.050 173.585 ;
        RECT 76.220 172.685 76.390 173.755 ;
        RECT 76.560 173.455 76.730 174.255 ;
        RECT 76.900 173.810 78.005 173.980 ;
        RECT 76.900 173.195 77.070 173.810 ;
        RECT 78.215 173.660 78.465 174.085 ;
        RECT 78.635 173.795 78.900 174.255 ;
        RECT 77.240 173.275 77.770 173.640 ;
        RECT 78.215 173.530 78.520 173.660 ;
        RECT 76.560 173.105 77.070 173.195 ;
        RECT 76.560 172.935 77.430 173.105 ;
        RECT 76.560 172.865 76.730 172.935 ;
        RECT 76.850 172.685 77.050 172.715 ;
        RECT 75.370 172.325 75.835 172.655 ;
        RECT 76.220 172.385 77.050 172.685 ;
        RECT 76.220 172.155 76.390 172.385 ;
        RECT 75.030 171.985 75.815 172.155 ;
        RECT 75.985 171.985 76.390 172.155 ;
        RECT 76.570 171.705 76.940 172.205 ;
        RECT 77.260 172.155 77.430 172.935 ;
        RECT 77.600 172.575 77.770 173.275 ;
        RECT 77.940 172.745 78.180 173.340 ;
        RECT 77.600 172.355 78.125 172.575 ;
        RECT 78.350 172.425 78.520 173.530 ;
        RECT 78.295 172.295 78.520 172.425 ;
        RECT 78.690 172.335 78.970 173.285 ;
        RECT 78.295 172.155 78.465 172.295 ;
        RECT 77.260 171.985 77.935 172.155 ;
        RECT 78.130 171.985 78.465 172.155 ;
        RECT 78.635 171.705 78.885 172.165 ;
        RECT 79.140 171.965 79.325 174.085 ;
        RECT 79.495 173.755 79.825 174.255 ;
        RECT 79.995 173.585 80.165 174.085 ;
        RECT 79.500 173.415 80.165 173.585 ;
        RECT 79.500 172.425 79.730 173.415 ;
        RECT 79.900 172.595 80.250 173.245 ;
        RECT 80.425 173.165 81.635 174.255 ;
        RECT 80.425 172.455 80.945 172.995 ;
        RECT 81.115 172.625 81.635 173.165 ;
        RECT 81.805 173.090 82.095 174.255 ;
        RECT 82.265 173.165 85.775 174.255 ;
        RECT 86.495 173.585 86.665 174.085 ;
        RECT 86.835 173.755 87.165 174.255 ;
        RECT 86.495 173.415 87.160 173.585 ;
        RECT 82.265 172.475 83.915 172.995 ;
        RECT 84.085 172.645 85.775 173.165 ;
        RECT 86.410 172.595 86.760 173.245 ;
        RECT 79.500 172.255 80.165 172.425 ;
        RECT 79.495 171.705 79.825 172.085 ;
        RECT 79.995 171.965 80.165 172.255 ;
        RECT 80.425 171.705 81.635 172.455 ;
        RECT 81.805 171.705 82.095 172.430 ;
        RECT 82.265 171.705 85.775 172.475 ;
        RECT 86.930 172.425 87.160 173.415 ;
        RECT 86.495 172.255 87.160 172.425 ;
        RECT 86.495 171.965 86.665 172.255 ;
        RECT 86.835 171.705 87.165 172.085 ;
        RECT 87.335 171.965 87.520 174.085 ;
        RECT 87.760 173.795 88.025 174.255 ;
        RECT 88.195 173.660 88.445 174.085 ;
        RECT 88.655 173.810 89.760 173.980 ;
        RECT 88.140 173.530 88.445 173.660 ;
        RECT 87.690 172.335 87.970 173.285 ;
        RECT 88.140 172.425 88.310 173.530 ;
        RECT 88.480 172.745 88.720 173.340 ;
        RECT 88.890 173.275 89.420 173.640 ;
        RECT 88.890 172.575 89.060 173.275 ;
        RECT 89.590 173.195 89.760 173.810 ;
        RECT 89.930 173.455 90.100 174.255 ;
        RECT 90.270 173.755 90.520 174.085 ;
        RECT 90.745 173.785 91.630 173.955 ;
        RECT 89.590 173.105 90.100 173.195 ;
        RECT 88.140 172.295 88.365 172.425 ;
        RECT 88.535 172.355 89.060 172.575 ;
        RECT 89.230 172.935 90.100 173.105 ;
        RECT 87.775 171.705 88.025 172.165 ;
        RECT 88.195 172.155 88.365 172.295 ;
        RECT 89.230 172.155 89.400 172.935 ;
        RECT 89.930 172.865 90.100 172.935 ;
        RECT 89.610 172.685 89.810 172.715 ;
        RECT 90.270 172.685 90.440 173.755 ;
        RECT 90.610 172.865 90.800 173.585 ;
        RECT 89.610 172.385 90.440 172.685 ;
        RECT 90.970 172.655 91.290 173.615 ;
        RECT 88.195 171.985 88.530 172.155 ;
        RECT 88.725 171.985 89.400 172.155 ;
        RECT 89.720 171.705 90.090 172.205 ;
        RECT 90.270 172.155 90.440 172.385 ;
        RECT 90.825 172.325 91.290 172.655 ;
        RECT 91.460 172.945 91.630 173.785 ;
        RECT 91.810 173.755 92.125 174.255 ;
        RECT 92.355 173.525 92.695 174.085 ;
        RECT 91.800 173.150 92.695 173.525 ;
        RECT 92.865 173.245 93.035 174.255 ;
        RECT 92.505 172.945 92.695 173.150 ;
        RECT 93.205 173.195 93.535 174.040 ;
        RECT 93.205 173.115 93.595 173.195 ;
        RECT 93.380 173.065 93.595 173.115 ;
        RECT 91.460 172.615 92.335 172.945 ;
        RECT 92.505 172.615 93.255 172.945 ;
        RECT 91.460 172.155 91.630 172.615 ;
        RECT 92.505 172.445 92.705 172.615 ;
        RECT 93.425 172.485 93.595 173.065 ;
        RECT 93.370 172.445 93.595 172.485 ;
        RECT 90.270 171.985 90.675 172.155 ;
        RECT 90.845 171.985 91.630 172.155 ;
        RECT 91.905 171.705 92.115 172.235 ;
        RECT 92.375 171.920 92.705 172.445 ;
        RECT 93.215 172.360 93.595 172.445 ;
        RECT 93.770 173.115 94.105 174.085 ;
        RECT 94.275 173.115 94.445 174.255 ;
        RECT 94.615 173.915 96.645 174.085 ;
        RECT 93.770 172.445 93.940 173.115 ;
        RECT 94.615 172.945 94.785 173.915 ;
        RECT 94.110 172.615 94.365 172.945 ;
        RECT 94.590 172.615 94.785 172.945 ;
        RECT 94.955 173.575 96.080 173.745 ;
        RECT 94.195 172.445 94.365 172.615 ;
        RECT 94.955 172.445 95.125 173.575 ;
        RECT 92.875 171.705 93.045 172.315 ;
        RECT 93.215 171.925 93.545 172.360 ;
        RECT 93.770 171.875 94.025 172.445 ;
        RECT 94.195 172.275 95.125 172.445 ;
        RECT 95.295 173.235 96.305 173.405 ;
        RECT 95.295 172.435 95.465 173.235 ;
        RECT 94.950 172.240 95.125 172.275 ;
        RECT 94.195 171.705 94.525 172.105 ;
        RECT 94.950 171.875 95.480 172.240 ;
        RECT 95.670 172.215 95.945 173.035 ;
        RECT 95.665 172.045 95.945 172.215 ;
        RECT 95.670 171.875 95.945 172.045 ;
        RECT 96.115 171.875 96.305 173.235 ;
        RECT 96.475 173.250 96.645 173.915 ;
        RECT 96.815 173.495 96.985 174.255 ;
        RECT 97.220 173.495 97.735 173.905 ;
        RECT 96.475 173.060 97.225 173.250 ;
        RECT 97.395 172.685 97.735 173.495 ;
        RECT 97.905 173.165 100.495 174.255 ;
        RECT 96.505 172.515 97.735 172.685 ;
        RECT 96.485 171.705 96.995 172.240 ;
        RECT 97.215 171.910 97.460 172.515 ;
        RECT 97.905 172.475 99.115 172.995 ;
        RECT 99.285 172.645 100.495 173.165 ;
        RECT 100.670 173.115 101.005 174.085 ;
        RECT 101.175 173.115 101.345 174.255 ;
        RECT 101.515 173.915 103.545 174.085 ;
        RECT 97.905 171.705 100.495 172.475 ;
        RECT 100.670 172.445 100.840 173.115 ;
        RECT 101.515 172.945 101.685 173.915 ;
        RECT 101.010 172.615 101.265 172.945 ;
        RECT 101.490 172.615 101.685 172.945 ;
        RECT 101.855 173.575 102.980 173.745 ;
        RECT 101.095 172.445 101.265 172.615 ;
        RECT 101.855 172.445 102.025 173.575 ;
        RECT 100.670 171.875 100.925 172.445 ;
        RECT 101.095 172.275 102.025 172.445 ;
        RECT 102.195 173.235 103.205 173.405 ;
        RECT 102.195 172.435 102.365 173.235 ;
        RECT 101.850 172.240 102.025 172.275 ;
        RECT 101.095 171.705 101.425 172.105 ;
        RECT 101.850 171.875 102.380 172.240 ;
        RECT 102.570 172.215 102.845 173.035 ;
        RECT 102.565 172.045 102.845 172.215 ;
        RECT 102.570 171.875 102.845 172.045 ;
        RECT 103.015 171.875 103.205 173.235 ;
        RECT 103.375 173.250 103.545 173.915 ;
        RECT 103.715 173.495 103.885 174.255 ;
        RECT 104.120 173.495 104.635 173.905 ;
        RECT 103.375 173.060 104.125 173.250 ;
        RECT 104.295 172.685 104.635 173.495 ;
        RECT 105.735 173.115 106.065 174.255 ;
        RECT 106.595 173.285 106.925 174.070 ;
        RECT 106.245 173.115 106.925 173.285 ;
        RECT 105.725 172.695 106.075 172.945 ;
        RECT 103.405 172.515 104.635 172.685 ;
        RECT 106.245 172.515 106.415 173.115 ;
        RECT 107.565 173.090 107.855 174.255 ;
        RECT 108.115 173.585 108.285 174.085 ;
        RECT 108.455 173.755 108.785 174.255 ;
        RECT 108.115 173.415 108.780 173.585 ;
        RECT 106.585 172.695 106.935 172.945 ;
        RECT 108.030 172.595 108.380 173.245 ;
        RECT 103.385 171.705 103.895 172.240 ;
        RECT 104.115 171.910 104.360 172.515 ;
        RECT 105.735 171.705 106.005 172.515 ;
        RECT 106.175 171.875 106.505 172.515 ;
        RECT 106.675 171.705 106.915 172.515 ;
        RECT 107.565 171.705 107.855 172.430 ;
        RECT 108.550 172.425 108.780 173.415 ;
        RECT 108.115 172.255 108.780 172.425 ;
        RECT 108.115 171.965 108.285 172.255 ;
        RECT 108.455 171.705 108.785 172.085 ;
        RECT 108.955 171.965 109.140 174.085 ;
        RECT 109.380 173.795 109.645 174.255 ;
        RECT 109.815 173.660 110.065 174.085 ;
        RECT 110.275 173.810 111.380 173.980 ;
        RECT 109.760 173.530 110.065 173.660 ;
        RECT 109.310 172.335 109.590 173.285 ;
        RECT 109.760 172.425 109.930 173.530 ;
        RECT 110.100 172.745 110.340 173.340 ;
        RECT 110.510 173.275 111.040 173.640 ;
        RECT 110.510 172.575 110.680 173.275 ;
        RECT 111.210 173.195 111.380 173.810 ;
        RECT 111.550 173.455 111.720 174.255 ;
        RECT 111.890 173.755 112.140 174.085 ;
        RECT 112.365 173.785 113.250 173.955 ;
        RECT 111.210 173.105 111.720 173.195 ;
        RECT 109.760 172.295 109.985 172.425 ;
        RECT 110.155 172.355 110.680 172.575 ;
        RECT 110.850 172.935 111.720 173.105 ;
        RECT 109.395 171.705 109.645 172.165 ;
        RECT 109.815 172.155 109.985 172.295 ;
        RECT 110.850 172.155 111.020 172.935 ;
        RECT 111.550 172.865 111.720 172.935 ;
        RECT 111.230 172.685 111.430 172.715 ;
        RECT 111.890 172.685 112.060 173.755 ;
        RECT 112.230 172.865 112.420 173.585 ;
        RECT 111.230 172.385 112.060 172.685 ;
        RECT 112.590 172.655 112.910 173.615 ;
        RECT 109.815 171.985 110.150 172.155 ;
        RECT 110.345 171.985 111.020 172.155 ;
        RECT 111.340 171.705 111.710 172.205 ;
        RECT 111.890 172.155 112.060 172.385 ;
        RECT 112.445 172.325 112.910 172.655 ;
        RECT 113.080 172.945 113.250 173.785 ;
        RECT 113.430 173.755 113.745 174.255 ;
        RECT 113.975 173.525 114.315 174.085 ;
        RECT 113.420 173.150 114.315 173.525 ;
        RECT 114.485 173.245 114.655 174.255 ;
        RECT 114.125 172.945 114.315 173.150 ;
        RECT 114.825 173.195 115.155 174.040 ;
        RECT 115.385 173.820 120.730 174.255 ;
        RECT 114.825 173.115 115.215 173.195 ;
        RECT 115.000 173.065 115.215 173.115 ;
        RECT 113.080 172.615 113.955 172.945 ;
        RECT 114.125 172.615 114.875 172.945 ;
        RECT 113.080 172.155 113.250 172.615 ;
        RECT 114.125 172.445 114.325 172.615 ;
        RECT 115.045 172.485 115.215 173.065 ;
        RECT 114.990 172.445 115.215 172.485 ;
        RECT 111.890 171.985 112.295 172.155 ;
        RECT 112.465 171.985 113.250 172.155 ;
        RECT 113.525 171.705 113.735 172.235 ;
        RECT 113.995 171.920 114.325 172.445 ;
        RECT 114.835 172.360 115.215 172.445 ;
        RECT 114.495 171.705 114.665 172.315 ;
        RECT 114.835 171.925 115.165 172.360 ;
        RECT 116.970 172.250 117.310 173.080 ;
        RECT 118.790 172.570 119.140 173.820 ;
        RECT 120.905 173.165 122.575 174.255 ;
        RECT 120.905 172.475 121.655 172.995 ;
        RECT 121.825 172.645 122.575 173.165 ;
        RECT 123.205 173.115 123.485 174.255 ;
        RECT 123.655 173.105 123.985 174.085 ;
        RECT 124.155 173.115 124.415 174.255 ;
        RECT 124.585 173.820 129.930 174.255 ;
        RECT 123.215 172.675 123.550 172.945 ;
        RECT 123.720 172.505 123.890 173.105 ;
        RECT 124.060 172.695 124.395 172.945 ;
        RECT 115.385 171.705 120.730 172.250 ;
        RECT 120.905 171.705 122.575 172.475 ;
        RECT 123.205 171.705 123.515 172.505 ;
        RECT 123.720 171.875 124.415 172.505 ;
        RECT 126.170 172.250 126.510 173.080 ;
        RECT 127.990 172.570 128.340 173.820 ;
        RECT 130.575 173.115 130.905 174.255 ;
        RECT 131.435 173.285 131.765 174.070 ;
        RECT 131.085 173.115 131.765 173.285 ;
        RECT 131.955 173.115 132.285 174.255 ;
        RECT 132.815 173.285 133.145 174.070 ;
        RECT 132.465 173.115 133.145 173.285 ;
        RECT 130.565 172.695 130.915 172.945 ;
        RECT 131.085 172.515 131.255 173.115 ;
        RECT 131.425 172.695 131.775 172.945 ;
        RECT 131.945 172.695 132.295 172.945 ;
        RECT 132.465 172.515 132.635 173.115 ;
        RECT 133.325 173.090 133.615 174.255 ;
        RECT 133.795 173.285 134.125 174.070 ;
        RECT 133.795 173.115 134.475 173.285 ;
        RECT 134.655 173.115 134.985 174.255 ;
        RECT 136.090 173.865 136.425 174.085 ;
        RECT 137.430 173.875 137.785 174.255 ;
        RECT 136.090 173.245 136.345 173.865 ;
        RECT 136.595 173.705 136.825 173.745 ;
        RECT 137.955 173.705 138.205 174.085 ;
        RECT 136.595 173.505 138.205 173.705 ;
        RECT 136.595 173.415 136.780 173.505 ;
        RECT 137.370 173.495 138.205 173.505 ;
        RECT 138.455 173.475 138.705 174.255 ;
        RECT 138.875 173.405 139.135 174.085 ;
        RECT 136.935 173.305 137.265 173.335 ;
        RECT 136.935 173.245 138.735 173.305 ;
        RECT 136.090 173.135 138.795 173.245 ;
        RECT 132.805 172.695 133.155 172.945 ;
        RECT 133.785 172.695 134.135 172.945 ;
        RECT 134.305 172.515 134.475 173.115 ;
        RECT 136.090 173.075 137.265 173.135 ;
        RECT 138.595 173.100 138.795 173.135 ;
        RECT 134.645 172.695 134.995 172.945 ;
        RECT 136.085 172.695 136.575 172.895 ;
        RECT 136.765 172.695 137.240 172.905 ;
        RECT 124.585 171.705 129.930 172.250 ;
        RECT 130.575 171.705 130.845 172.515 ;
        RECT 131.015 171.875 131.345 172.515 ;
        RECT 131.515 171.705 131.755 172.515 ;
        RECT 131.955 171.705 132.225 172.515 ;
        RECT 132.395 171.875 132.725 172.515 ;
        RECT 132.895 171.705 133.135 172.515 ;
        RECT 133.325 171.705 133.615 172.430 ;
        RECT 133.805 171.705 134.045 172.515 ;
        RECT 134.215 171.875 134.545 172.515 ;
        RECT 134.715 171.705 134.985 172.515 ;
        RECT 136.090 171.705 136.545 172.470 ;
        RECT 137.020 172.295 137.240 172.695 ;
        RECT 137.485 172.695 137.815 172.905 ;
        RECT 137.485 172.295 137.695 172.695 ;
        RECT 137.985 172.660 138.395 172.965 ;
        RECT 138.625 172.525 138.795 173.100 ;
        RECT 138.525 172.405 138.795 172.525 ;
        RECT 137.950 172.360 138.795 172.405 ;
        RECT 137.950 172.235 138.705 172.360 ;
        RECT 137.950 172.085 138.120 172.235 ;
        RECT 138.965 172.205 139.135 173.405 ;
        RECT 139.365 173.115 139.575 174.255 ;
        RECT 139.745 173.105 140.075 174.085 ;
        RECT 140.245 173.115 140.475 174.255 ;
        RECT 140.685 173.115 140.945 174.255 ;
        RECT 141.115 173.105 141.445 174.085 ;
        RECT 141.615 173.115 141.895 174.255 ;
        RECT 142.065 173.165 145.575 174.255 ;
        RECT 136.820 171.875 138.120 172.085 ;
        RECT 138.375 171.705 138.705 172.065 ;
        RECT 138.875 171.875 139.135 172.205 ;
        RECT 139.365 171.705 139.575 172.525 ;
        RECT 139.745 172.505 139.995 173.105 ;
        RECT 141.205 173.065 141.380 173.105 ;
        RECT 140.165 172.695 140.495 172.945 ;
        RECT 140.705 172.695 141.040 172.945 ;
        RECT 139.745 171.875 140.075 172.505 ;
        RECT 140.245 171.705 140.475 172.525 ;
        RECT 141.210 172.505 141.380 173.065 ;
        RECT 141.550 172.675 141.885 172.945 ;
        RECT 140.685 171.875 141.380 172.505 ;
        RECT 141.585 171.705 141.895 172.505 ;
        RECT 142.065 172.475 143.715 172.995 ;
        RECT 143.885 172.645 145.575 173.165 ;
        RECT 145.745 173.165 146.955 174.255 ;
        RECT 145.745 172.625 146.265 173.165 ;
        RECT 142.065 171.705 145.575 172.475 ;
        RECT 146.435 172.455 146.955 172.995 ;
        RECT 145.745 171.705 146.955 172.455 ;
        RECT 17.320 171.535 147.040 171.705 ;
        RECT 17.405 170.785 18.615 171.535 ;
        RECT 18.785 170.990 24.130 171.535 ;
        RECT 24.305 170.990 29.650 171.535 ;
        RECT 17.405 170.245 17.925 170.785 ;
        RECT 18.095 170.075 18.615 170.615 ;
        RECT 20.370 170.160 20.710 170.990 ;
        RECT 17.405 168.985 18.615 170.075 ;
        RECT 22.190 169.420 22.540 170.670 ;
        RECT 25.890 170.160 26.230 170.990 ;
        RECT 29.825 170.765 33.335 171.535 ;
        RECT 33.505 170.785 34.715 171.535 ;
        RECT 34.885 170.895 35.225 171.300 ;
        RECT 35.395 171.065 35.565 171.535 ;
        RECT 35.735 170.895 35.985 171.300 ;
        RECT 27.710 169.420 28.060 170.670 ;
        RECT 29.825 170.245 31.475 170.765 ;
        RECT 31.645 170.075 33.335 170.595 ;
        RECT 33.505 170.245 34.025 170.785 ;
        RECT 34.885 170.715 35.985 170.895 ;
        RECT 36.155 170.930 36.405 171.300 ;
        RECT 36.575 171.055 37.020 171.225 ;
        RECT 37.190 171.195 37.410 171.240 ;
        RECT 34.195 170.075 34.715 170.615 ;
        RECT 36.155 170.545 36.325 170.930 ;
        RECT 18.785 168.985 24.130 169.420 ;
        RECT 24.305 168.985 29.650 169.420 ;
        RECT 29.825 168.985 33.335 170.075 ;
        RECT 33.505 168.985 34.715 170.075 ;
        RECT 34.885 169.975 35.230 170.545 ;
        RECT 35.400 170.295 35.960 170.545 ;
        RECT 36.130 170.375 36.325 170.545 ;
        RECT 34.885 168.985 35.230 169.805 ;
        RECT 35.400 169.195 35.575 170.295 ;
        RECT 36.130 170.125 36.300 170.375 ;
        RECT 36.575 170.265 36.745 171.055 ;
        RECT 37.190 171.025 37.415 171.195 ;
        RECT 37.190 170.885 37.410 171.025 ;
        RECT 36.915 170.715 37.410 170.885 ;
        RECT 37.690 170.870 37.860 171.535 ;
        RECT 38.055 170.795 38.395 171.365 ;
        RECT 38.730 171.025 38.970 171.535 ;
        RECT 39.150 171.025 39.430 171.355 ;
        RECT 39.660 171.025 39.875 171.535 ;
        RECT 36.915 170.520 37.090 170.715 ;
        RECT 37.260 170.345 37.710 170.545 ;
        RECT 35.745 169.735 36.300 170.125 ;
        RECT 36.470 170.125 36.745 170.265 ;
        RECT 37.880 170.175 38.050 170.625 ;
        RECT 36.470 169.905 37.485 170.125 ;
        RECT 37.655 170.005 38.050 170.175 ;
        RECT 37.655 169.735 37.825 170.005 ;
        RECT 38.220 169.825 38.395 170.795 ;
        RECT 38.625 170.295 38.980 170.855 ;
        RECT 39.150 170.125 39.320 171.025 ;
        RECT 39.490 170.295 39.755 170.855 ;
        RECT 40.045 170.795 40.660 171.365 ;
        RECT 40.005 170.125 40.175 170.625 ;
        RECT 35.745 169.565 37.825 169.735 ;
        RECT 35.745 169.330 36.075 169.565 ;
        RECT 36.365 168.985 36.765 169.385 ;
        RECT 37.635 168.985 37.965 169.385 ;
        RECT 38.135 169.155 38.395 169.825 ;
        RECT 38.750 169.955 40.175 170.125 ;
        RECT 38.750 169.780 39.140 169.955 ;
        RECT 39.625 168.985 39.955 169.785 ;
        RECT 40.345 169.775 40.660 170.795 ;
        RECT 40.865 170.765 42.535 171.535 ;
        RECT 43.165 170.810 43.455 171.535 ;
        RECT 43.625 170.810 43.885 171.365 ;
        RECT 44.055 171.090 44.485 171.535 ;
        RECT 44.720 170.965 44.890 171.365 ;
        RECT 45.060 171.135 45.780 171.535 ;
        RECT 40.865 170.245 41.615 170.765 ;
        RECT 41.785 170.075 42.535 170.595 ;
        RECT 40.125 169.155 40.660 169.775 ;
        RECT 40.865 168.985 42.535 170.075 ;
        RECT 43.165 168.985 43.455 170.150 ;
        RECT 43.625 170.095 43.800 170.810 ;
        RECT 44.720 170.795 45.600 170.965 ;
        RECT 45.950 170.920 46.120 171.365 ;
        RECT 46.695 171.025 47.095 171.535 ;
        RECT 47.355 171.145 47.685 171.535 ;
        RECT 47.855 170.965 48.025 171.285 ;
        RECT 48.195 171.145 48.525 171.535 ;
        RECT 48.940 171.135 49.895 171.305 ;
        RECT 43.970 170.295 44.225 170.625 ;
        RECT 43.625 169.155 43.885 170.095 ;
        RECT 44.055 169.815 44.225 170.295 ;
        RECT 44.450 170.005 44.780 170.625 ;
        RECT 44.950 170.245 45.240 170.625 ;
        RECT 45.430 170.075 45.600 170.795 ;
        RECT 45.080 169.905 45.600 170.075 ;
        RECT 45.770 170.750 46.120 170.920 ;
        RECT 44.055 169.645 44.815 169.815 ;
        RECT 45.080 169.715 45.250 169.905 ;
        RECT 45.770 169.725 45.940 170.750 ;
        RECT 46.360 170.265 46.620 170.855 ;
        RECT 46.140 169.965 46.620 170.265 ;
        RECT 46.820 169.965 47.080 170.855 ;
        RECT 47.305 170.795 49.555 170.965 ;
        RECT 47.305 169.835 47.475 170.795 ;
        RECT 47.645 170.175 47.890 170.625 ;
        RECT 48.060 170.345 48.610 170.545 ;
        RECT 48.780 170.375 49.155 170.545 ;
        RECT 48.780 170.175 48.950 170.375 ;
        RECT 49.325 170.295 49.555 170.795 ;
        RECT 47.645 170.005 48.950 170.175 ;
        RECT 49.725 170.255 49.895 171.135 ;
        RECT 50.065 170.700 50.355 171.535 ;
        RECT 50.725 170.905 51.055 171.265 ;
        RECT 51.675 171.075 51.925 171.535 ;
        RECT 52.095 171.075 52.655 171.365 ;
        RECT 50.725 170.715 52.115 170.905 ;
        RECT 51.945 170.625 52.115 170.715 ;
        RECT 50.540 170.295 51.215 170.545 ;
        RECT 51.435 170.295 51.775 170.545 ;
        RECT 51.945 170.295 52.235 170.625 ;
        RECT 49.725 170.085 50.355 170.255 ;
        RECT 44.645 169.420 44.815 169.645 ;
        RECT 45.530 169.555 45.940 169.725 ;
        RECT 46.115 169.615 47.055 169.785 ;
        RECT 45.530 169.420 45.785 169.555 ;
        RECT 44.055 168.985 44.385 169.385 ;
        RECT 44.645 169.250 45.785 169.420 ;
        RECT 46.115 169.365 46.285 169.615 ;
        RECT 45.530 169.155 45.785 169.250 ;
        RECT 45.955 169.195 46.285 169.365 ;
        RECT 46.455 168.985 46.705 169.445 ;
        RECT 46.875 169.155 47.055 169.615 ;
        RECT 47.305 169.155 47.685 169.835 ;
        RECT 48.275 168.985 48.445 169.835 ;
        RECT 48.615 169.665 49.855 169.835 ;
        RECT 48.615 169.155 48.945 169.665 ;
        RECT 49.115 168.985 49.285 169.495 ;
        RECT 49.455 169.155 49.855 169.665 ;
        RECT 50.035 169.155 50.355 170.085 ;
        RECT 50.540 169.935 50.805 170.295 ;
        RECT 51.945 170.045 52.115 170.295 ;
        RECT 51.175 169.875 52.115 170.045 ;
        RECT 50.725 168.985 51.005 169.655 ;
        RECT 51.175 169.325 51.475 169.875 ;
        RECT 52.405 169.705 52.655 171.075 ;
        RECT 52.825 170.765 56.335 171.535 ;
        RECT 57.035 171.135 57.365 171.535 ;
        RECT 57.535 170.965 57.705 171.235 ;
        RECT 57.875 171.135 58.205 171.535 ;
        RECT 58.375 170.965 58.630 171.235 ;
        RECT 52.825 170.245 54.475 170.765 ;
        RECT 54.645 170.075 56.335 170.595 ;
        RECT 51.675 168.985 52.005 169.705 ;
        RECT 52.195 169.155 52.655 169.705 ;
        RECT 52.825 168.985 56.335 170.075 ;
        RECT 56.965 169.955 57.235 170.965 ;
        RECT 57.405 170.795 58.630 170.965 ;
        RECT 58.805 170.795 59.125 171.275 ;
        RECT 59.295 170.965 59.525 171.365 ;
        RECT 59.695 171.145 60.045 171.535 ;
        RECT 59.295 170.885 59.805 170.965 ;
        RECT 60.215 170.885 60.545 171.365 ;
        RECT 59.295 170.795 60.545 170.885 ;
        RECT 57.405 170.125 57.575 170.795 ;
        RECT 57.745 170.295 58.125 170.625 ;
        RECT 58.295 170.295 58.630 170.625 ;
        RECT 57.405 169.955 57.720 170.125 ;
        RECT 56.970 168.985 57.285 169.785 ;
        RECT 57.550 169.340 57.720 169.955 ;
        RECT 57.890 169.615 58.125 170.295 ;
        RECT 58.295 169.340 58.630 170.125 ;
        RECT 58.805 169.865 58.975 170.795 ;
        RECT 59.635 170.715 60.545 170.795 ;
        RECT 60.715 170.715 60.885 171.535 ;
        RECT 61.390 170.795 61.855 171.340 ;
        RECT 59.145 170.205 59.315 170.625 ;
        RECT 59.545 170.375 60.145 170.545 ;
        RECT 59.145 170.035 59.805 170.205 ;
        RECT 58.805 169.665 59.465 169.865 ;
        RECT 59.635 169.835 59.805 170.035 ;
        RECT 59.975 170.175 60.145 170.375 ;
        RECT 60.315 170.345 61.010 170.545 ;
        RECT 61.270 170.175 61.515 170.625 ;
        RECT 59.975 170.005 61.515 170.175 ;
        RECT 61.685 169.835 61.855 170.795 ;
        RECT 59.635 169.665 61.855 169.835 ;
        RECT 62.025 170.795 62.490 171.340 ;
        RECT 62.025 169.835 62.195 170.795 ;
        RECT 62.995 170.715 63.165 171.535 ;
        RECT 63.335 170.885 63.665 171.365 ;
        RECT 63.835 171.145 64.185 171.535 ;
        RECT 64.355 170.965 64.585 171.365 ;
        RECT 64.075 170.885 64.585 170.965 ;
        RECT 63.335 170.795 64.585 170.885 ;
        RECT 64.755 170.795 65.075 171.275 ;
        RECT 63.335 170.715 64.245 170.795 ;
        RECT 62.365 170.175 62.610 170.625 ;
        RECT 62.870 170.345 63.565 170.545 ;
        RECT 63.735 170.375 64.335 170.545 ;
        RECT 63.735 170.175 63.905 170.375 ;
        RECT 64.565 170.205 64.735 170.625 ;
        RECT 62.365 170.005 63.905 170.175 ;
        RECT 64.075 170.035 64.735 170.205 ;
        RECT 64.075 169.835 64.245 170.035 ;
        RECT 64.905 169.865 65.075 170.795 ;
        RECT 62.025 169.665 64.245 169.835 ;
        RECT 64.415 169.665 65.075 169.865 ;
        RECT 65.245 170.795 65.630 171.365 ;
        RECT 65.800 171.075 66.125 171.535 ;
        RECT 66.645 170.905 66.925 171.365 ;
        RECT 65.245 170.125 65.525 170.795 ;
        RECT 65.800 170.735 66.925 170.905 ;
        RECT 65.800 170.625 66.250 170.735 ;
        RECT 65.695 170.295 66.250 170.625 ;
        RECT 67.115 170.565 67.515 171.365 ;
        RECT 67.915 171.075 68.185 171.535 ;
        RECT 68.355 170.905 68.640 171.365 ;
        RECT 59.295 169.495 59.465 169.665 ;
        RECT 57.550 169.170 58.630 169.340 ;
        RECT 58.825 168.985 59.125 169.495 ;
        RECT 59.295 169.325 59.675 169.495 ;
        RECT 60.255 168.985 60.885 169.495 ;
        RECT 61.055 169.155 61.385 169.665 ;
        RECT 61.555 168.985 61.855 169.495 ;
        RECT 62.025 168.985 62.325 169.495 ;
        RECT 62.495 169.155 62.825 169.665 ;
        RECT 64.415 169.495 64.585 169.665 ;
        RECT 62.995 168.985 63.625 169.495 ;
        RECT 64.205 169.325 64.585 169.495 ;
        RECT 64.755 168.985 65.055 169.495 ;
        RECT 65.245 169.155 65.630 170.125 ;
        RECT 65.800 169.835 66.250 170.295 ;
        RECT 66.420 170.005 67.515 170.565 ;
        RECT 65.800 169.615 66.925 169.835 ;
        RECT 65.800 168.985 66.125 169.445 ;
        RECT 66.645 169.155 66.925 169.615 ;
        RECT 67.115 169.155 67.515 170.005 ;
        RECT 67.685 170.735 68.640 170.905 ;
        RECT 68.925 170.810 69.215 171.535 ;
        RECT 69.385 170.795 69.770 171.365 ;
        RECT 69.940 171.075 70.265 171.535 ;
        RECT 70.785 170.905 71.065 171.365 ;
        RECT 67.685 169.835 67.895 170.735 ;
        RECT 68.065 170.005 68.755 170.565 ;
        RECT 67.685 169.615 68.640 169.835 ;
        RECT 67.915 168.985 68.185 169.445 ;
        RECT 68.355 169.155 68.640 169.615 ;
        RECT 68.925 168.985 69.215 170.150 ;
        RECT 69.385 170.125 69.665 170.795 ;
        RECT 69.940 170.735 71.065 170.905 ;
        RECT 69.940 170.625 70.390 170.735 ;
        RECT 69.835 170.295 70.390 170.625 ;
        RECT 71.255 170.565 71.655 171.365 ;
        RECT 72.055 171.075 72.325 171.535 ;
        RECT 72.495 170.905 72.780 171.365 ;
        RECT 73.135 171.135 73.465 171.535 ;
        RECT 73.635 170.965 73.805 171.235 ;
        RECT 73.975 171.135 74.305 171.535 ;
        RECT 74.475 170.965 74.730 171.235 ;
        RECT 69.385 169.155 69.770 170.125 ;
        RECT 69.940 169.835 70.390 170.295 ;
        RECT 70.560 170.005 71.655 170.565 ;
        RECT 69.940 169.615 71.065 169.835 ;
        RECT 69.940 168.985 70.265 169.445 ;
        RECT 70.785 169.155 71.065 169.615 ;
        RECT 71.255 169.155 71.655 170.005 ;
        RECT 71.825 170.735 72.780 170.905 ;
        RECT 71.825 169.835 72.035 170.735 ;
        RECT 72.205 170.005 72.895 170.565 ;
        RECT 73.065 169.955 73.335 170.965 ;
        RECT 73.505 170.795 74.730 170.965 ;
        RECT 73.505 170.125 73.675 170.795 ;
        RECT 74.905 170.765 77.495 171.535 ;
        RECT 77.755 170.985 77.925 171.275 ;
        RECT 78.095 171.155 78.425 171.535 ;
        RECT 77.755 170.815 78.420 170.985 ;
        RECT 73.845 170.295 74.225 170.625 ;
        RECT 74.395 170.295 74.730 170.625 ;
        RECT 73.505 169.955 73.820 170.125 ;
        RECT 71.825 169.615 72.780 169.835 ;
        RECT 72.055 168.985 72.325 169.445 ;
        RECT 72.495 169.155 72.780 169.615 ;
        RECT 73.070 168.985 73.385 169.785 ;
        RECT 73.650 169.340 73.820 169.955 ;
        RECT 73.990 169.615 74.225 170.295 ;
        RECT 74.905 170.245 76.115 170.765 ;
        RECT 74.395 169.340 74.730 170.125 ;
        RECT 76.285 170.075 77.495 170.595 ;
        RECT 73.650 169.170 74.730 169.340 ;
        RECT 74.905 168.985 77.495 170.075 ;
        RECT 77.670 169.995 78.020 170.645 ;
        RECT 78.190 169.825 78.420 170.815 ;
        RECT 77.755 169.655 78.420 169.825 ;
        RECT 77.755 169.155 77.925 169.655 ;
        RECT 78.095 168.985 78.425 169.485 ;
        RECT 78.595 169.155 78.780 171.275 ;
        RECT 79.035 171.075 79.285 171.535 ;
        RECT 79.455 171.085 79.790 171.255 ;
        RECT 79.985 171.085 80.660 171.255 ;
        RECT 79.455 170.945 79.625 171.085 ;
        RECT 78.950 169.955 79.230 170.905 ;
        RECT 79.400 170.815 79.625 170.945 ;
        RECT 79.400 169.710 79.570 170.815 ;
        RECT 79.795 170.665 80.320 170.885 ;
        RECT 79.740 169.900 79.980 170.495 ;
        RECT 80.150 169.965 80.320 170.665 ;
        RECT 80.490 170.305 80.660 171.085 ;
        RECT 80.980 171.035 81.350 171.535 ;
        RECT 81.530 171.085 81.935 171.255 ;
        RECT 82.105 171.085 82.890 171.255 ;
        RECT 81.530 170.855 81.700 171.085 ;
        RECT 80.870 170.555 81.700 170.855 ;
        RECT 82.085 170.585 82.550 170.915 ;
        RECT 80.870 170.525 81.070 170.555 ;
        RECT 81.190 170.305 81.360 170.375 ;
        RECT 80.490 170.135 81.360 170.305 ;
        RECT 80.850 170.045 81.360 170.135 ;
        RECT 79.400 169.580 79.705 169.710 ;
        RECT 80.150 169.600 80.680 169.965 ;
        RECT 79.020 168.985 79.285 169.445 ;
        RECT 79.455 169.155 79.705 169.580 ;
        RECT 80.850 169.430 81.020 170.045 ;
        RECT 79.915 169.260 81.020 169.430 ;
        RECT 81.190 168.985 81.360 169.785 ;
        RECT 81.530 169.485 81.700 170.555 ;
        RECT 81.870 169.655 82.060 170.375 ;
        RECT 82.230 169.625 82.550 170.585 ;
        RECT 82.720 170.625 82.890 171.085 ;
        RECT 83.165 171.005 83.375 171.535 ;
        RECT 83.635 170.795 83.965 171.320 ;
        RECT 84.135 170.925 84.305 171.535 ;
        RECT 84.475 170.880 84.805 171.315 ;
        RECT 85.025 170.990 90.370 171.535 ;
        RECT 84.475 170.795 84.855 170.880 ;
        RECT 83.765 170.625 83.965 170.795 ;
        RECT 84.630 170.755 84.855 170.795 ;
        RECT 82.720 170.295 83.595 170.625 ;
        RECT 83.765 170.295 84.515 170.625 ;
        RECT 81.530 169.155 81.780 169.485 ;
        RECT 82.720 169.455 82.890 170.295 ;
        RECT 83.765 170.090 83.955 170.295 ;
        RECT 84.685 170.175 84.855 170.755 ;
        RECT 84.640 170.125 84.855 170.175 ;
        RECT 86.610 170.160 86.950 170.990 ;
        RECT 90.545 170.765 94.055 171.535 ;
        RECT 94.685 170.810 94.975 171.535 ;
        RECT 95.150 170.795 95.405 171.365 ;
        RECT 95.575 171.135 95.905 171.535 ;
        RECT 96.330 171.000 96.860 171.365 ;
        RECT 96.330 170.965 96.505 171.000 ;
        RECT 95.575 170.795 96.505 170.965 ;
        RECT 83.060 169.715 83.955 170.090 ;
        RECT 84.465 170.045 84.855 170.125 ;
        RECT 82.005 169.285 82.890 169.455 ;
        RECT 83.070 168.985 83.385 169.485 ;
        RECT 83.615 169.155 83.955 169.715 ;
        RECT 84.125 168.985 84.295 169.995 ;
        RECT 84.465 169.200 84.795 170.045 ;
        RECT 88.430 169.420 88.780 170.670 ;
        RECT 90.545 170.245 92.195 170.765 ;
        RECT 92.365 170.075 94.055 170.595 ;
        RECT 85.025 168.985 90.370 169.420 ;
        RECT 90.545 168.985 94.055 170.075 ;
        RECT 94.685 168.985 94.975 170.150 ;
        RECT 95.150 170.125 95.320 170.795 ;
        RECT 95.575 170.625 95.745 170.795 ;
        RECT 95.490 170.295 95.745 170.625 ;
        RECT 95.970 170.295 96.165 170.625 ;
        RECT 95.150 169.155 95.485 170.125 ;
        RECT 95.655 168.985 95.825 170.125 ;
        RECT 95.995 169.325 96.165 170.295 ;
        RECT 96.335 169.665 96.505 170.795 ;
        RECT 96.675 170.005 96.845 170.805 ;
        RECT 97.050 170.515 97.325 171.365 ;
        RECT 97.045 170.345 97.325 170.515 ;
        RECT 97.050 170.205 97.325 170.345 ;
        RECT 97.495 170.005 97.685 171.365 ;
        RECT 97.865 171.000 98.375 171.535 ;
        RECT 98.595 170.725 98.840 171.330 ;
        RECT 99.285 170.765 100.955 171.535 ;
        RECT 101.185 171.075 101.430 171.535 ;
        RECT 97.885 170.555 99.115 170.725 ;
        RECT 96.675 169.835 97.685 170.005 ;
        RECT 97.855 169.990 98.605 170.180 ;
        RECT 96.335 169.495 97.460 169.665 ;
        RECT 97.855 169.325 98.025 169.990 ;
        RECT 98.775 169.745 99.115 170.555 ;
        RECT 99.285 170.245 100.035 170.765 ;
        RECT 100.205 170.075 100.955 170.595 ;
        RECT 101.125 170.295 101.440 170.905 ;
        RECT 101.610 170.545 101.860 171.355 ;
        RECT 102.030 171.010 102.290 171.535 ;
        RECT 102.460 170.885 102.720 171.340 ;
        RECT 102.890 171.055 103.150 171.535 ;
        RECT 103.320 170.885 103.580 171.340 ;
        RECT 103.750 171.055 104.010 171.535 ;
        RECT 104.180 170.885 104.440 171.340 ;
        RECT 104.610 171.055 104.870 171.535 ;
        RECT 105.040 170.885 105.300 171.340 ;
        RECT 105.470 171.055 105.770 171.535 ;
        RECT 102.460 170.715 105.770 170.885 ;
        RECT 101.610 170.295 104.630 170.545 ;
        RECT 95.995 169.155 98.025 169.325 ;
        RECT 98.195 168.985 98.365 169.745 ;
        RECT 98.600 169.335 99.115 169.745 ;
        RECT 99.285 168.985 100.955 170.075 ;
        RECT 101.135 168.985 101.430 170.095 ;
        RECT 101.610 169.160 101.860 170.295 ;
        RECT 104.800 170.125 105.770 170.715 ;
        RECT 106.185 170.765 107.855 171.535 ;
        RECT 108.115 170.985 108.285 171.275 ;
        RECT 108.455 171.155 108.785 171.535 ;
        RECT 108.115 170.815 108.780 170.985 ;
        RECT 106.185 170.245 106.935 170.765 ;
        RECT 102.030 168.985 102.290 170.095 ;
        RECT 102.460 169.885 105.770 170.125 ;
        RECT 107.105 170.075 107.855 170.595 ;
        RECT 102.460 169.160 102.720 169.885 ;
        RECT 102.890 168.985 103.150 169.715 ;
        RECT 103.320 169.160 103.580 169.885 ;
        RECT 103.750 168.985 104.010 169.715 ;
        RECT 104.180 169.160 104.440 169.885 ;
        RECT 104.610 168.985 104.870 169.715 ;
        RECT 105.040 169.160 105.300 169.885 ;
        RECT 105.470 168.985 105.765 169.715 ;
        RECT 106.185 168.985 107.855 170.075 ;
        RECT 108.030 169.995 108.380 170.645 ;
        RECT 108.550 169.825 108.780 170.815 ;
        RECT 108.115 169.655 108.780 169.825 ;
        RECT 108.115 169.155 108.285 169.655 ;
        RECT 108.455 168.985 108.785 169.485 ;
        RECT 108.955 169.155 109.140 171.275 ;
        RECT 109.395 171.075 109.645 171.535 ;
        RECT 109.815 171.085 110.150 171.255 ;
        RECT 110.345 171.085 111.020 171.255 ;
        RECT 109.815 170.945 109.985 171.085 ;
        RECT 109.310 169.955 109.590 170.905 ;
        RECT 109.760 170.815 109.985 170.945 ;
        RECT 109.760 169.710 109.930 170.815 ;
        RECT 110.155 170.665 110.680 170.885 ;
        RECT 110.100 169.900 110.340 170.495 ;
        RECT 110.510 169.965 110.680 170.665 ;
        RECT 110.850 170.305 111.020 171.085 ;
        RECT 111.340 171.035 111.710 171.535 ;
        RECT 111.890 171.085 112.295 171.255 ;
        RECT 112.465 171.085 113.250 171.255 ;
        RECT 111.890 170.855 112.060 171.085 ;
        RECT 111.230 170.555 112.060 170.855 ;
        RECT 112.445 170.585 112.910 170.915 ;
        RECT 111.230 170.525 111.430 170.555 ;
        RECT 111.550 170.305 111.720 170.375 ;
        RECT 110.850 170.135 111.720 170.305 ;
        RECT 111.210 170.045 111.720 170.135 ;
        RECT 109.760 169.580 110.065 169.710 ;
        RECT 110.510 169.600 111.040 169.965 ;
        RECT 109.380 168.985 109.645 169.445 ;
        RECT 109.815 169.155 110.065 169.580 ;
        RECT 111.210 169.430 111.380 170.045 ;
        RECT 110.275 169.260 111.380 169.430 ;
        RECT 111.550 168.985 111.720 169.785 ;
        RECT 111.890 169.485 112.060 170.555 ;
        RECT 112.230 169.655 112.420 170.375 ;
        RECT 112.590 169.625 112.910 170.585 ;
        RECT 113.080 170.625 113.250 171.085 ;
        RECT 113.525 171.005 113.735 171.535 ;
        RECT 113.995 170.795 114.325 171.320 ;
        RECT 114.495 170.925 114.665 171.535 ;
        RECT 114.835 170.880 115.165 171.315 ;
        RECT 114.835 170.795 115.215 170.880 ;
        RECT 114.125 170.625 114.325 170.795 ;
        RECT 114.990 170.755 115.215 170.795 ;
        RECT 113.080 170.295 113.955 170.625 ;
        RECT 114.125 170.295 114.875 170.625 ;
        RECT 111.890 169.155 112.140 169.485 ;
        RECT 113.080 169.455 113.250 170.295 ;
        RECT 114.125 170.090 114.315 170.295 ;
        RECT 115.045 170.175 115.215 170.755 ;
        RECT 115.000 170.125 115.215 170.175 ;
        RECT 113.420 169.715 114.315 170.090 ;
        RECT 114.825 170.045 115.215 170.125 ;
        RECT 112.365 169.285 113.250 169.455 ;
        RECT 113.430 168.985 113.745 169.485 ;
        RECT 113.975 169.155 114.315 169.715 ;
        RECT 114.485 168.985 114.655 169.995 ;
        RECT 114.825 169.200 115.155 170.045 ;
        RECT 116.325 169.955 116.555 171.295 ;
        RECT 116.735 170.455 116.965 171.355 ;
        RECT 117.165 170.755 117.410 171.535 ;
        RECT 117.580 170.995 118.010 171.355 ;
        RECT 118.590 171.165 119.320 171.535 ;
        RECT 117.580 170.805 119.320 170.995 ;
        RECT 117.580 170.575 117.800 170.805 ;
        RECT 116.735 169.775 117.075 170.455 ;
        RECT 116.325 169.575 117.075 169.775 ;
        RECT 117.255 170.275 117.800 170.575 ;
        RECT 116.325 169.185 116.565 169.575 ;
        RECT 116.735 168.985 117.085 169.395 ;
        RECT 117.255 169.165 117.585 170.275 ;
        RECT 117.970 170.005 118.395 170.625 ;
        RECT 118.590 170.005 118.850 170.625 ;
        RECT 119.060 170.295 119.320 170.805 ;
        RECT 117.755 169.635 118.780 169.835 ;
        RECT 117.755 169.165 117.935 169.635 ;
        RECT 118.105 168.985 118.435 169.465 ;
        RECT 118.610 169.165 118.780 169.635 ;
        RECT 119.045 168.985 119.330 170.125 ;
        RECT 119.520 169.165 119.800 171.355 ;
        RECT 120.445 170.810 120.735 171.535 ;
        RECT 120.905 170.990 126.250 171.535 ;
        RECT 126.450 171.145 126.780 171.535 ;
        RECT 122.490 170.160 122.830 170.990 ;
        RECT 126.950 170.975 127.175 171.355 ;
        RECT 120.445 168.985 120.735 170.150 ;
        RECT 124.310 169.420 124.660 170.670 ;
        RECT 126.435 170.295 126.675 170.945 ;
        RECT 126.845 170.795 127.175 170.975 ;
        RECT 126.845 170.125 127.020 170.795 ;
        RECT 127.375 170.625 127.605 171.245 ;
        RECT 127.785 170.805 128.085 171.535 ;
        RECT 128.285 170.725 128.525 171.535 ;
        RECT 128.695 170.725 129.025 171.365 ;
        RECT 129.195 170.725 129.465 171.535 ;
        RECT 129.645 170.765 132.235 171.535 ;
        RECT 132.405 170.795 132.990 171.365 ;
        RECT 133.240 170.965 133.570 171.310 ;
        RECT 133.785 171.135 134.160 171.535 ;
        RECT 134.340 170.965 134.635 171.310 ;
        RECT 133.240 170.795 134.635 170.965 ;
        RECT 134.805 170.795 135.475 171.535 ;
        RECT 127.190 170.295 127.605 170.625 ;
        RECT 127.785 170.295 128.080 170.625 ;
        RECT 128.265 170.295 128.615 170.545 ;
        RECT 128.785 170.125 128.955 170.725 ;
        RECT 129.125 170.295 129.475 170.545 ;
        RECT 129.645 170.245 130.855 170.765 ;
        RECT 126.435 169.935 127.020 170.125 ;
        RECT 120.905 168.985 126.250 169.420 ;
        RECT 126.435 169.165 126.710 169.935 ;
        RECT 127.190 169.765 128.085 170.095 ;
        RECT 126.880 169.595 128.085 169.765 ;
        RECT 126.880 169.165 127.210 169.595 ;
        RECT 127.380 168.985 127.575 169.425 ;
        RECT 127.755 169.165 128.085 169.595 ;
        RECT 128.275 169.955 128.955 170.125 ;
        RECT 128.275 169.170 128.605 169.955 ;
        RECT 129.135 168.985 129.465 170.125 ;
        RECT 131.025 170.075 132.235 170.595 ;
        RECT 132.405 170.295 132.650 170.625 ;
        RECT 132.820 170.125 132.990 170.795 ;
        RECT 133.160 170.295 133.560 170.625 ;
        RECT 133.730 170.295 134.020 170.625 ;
        RECT 129.645 168.985 132.235 170.075 ;
        RECT 132.405 169.955 133.615 170.125 ;
        RECT 132.405 169.155 132.695 169.955 ;
        RECT 132.865 168.985 133.100 169.785 ;
        RECT 133.285 169.325 133.615 169.955 ;
        RECT 133.785 169.550 134.020 170.295 ;
        RECT 134.210 170.295 134.550 170.625 ;
        RECT 134.720 170.295 135.055 170.625 ;
        RECT 134.210 169.550 134.480 170.295 ;
        RECT 135.225 170.125 135.395 170.625 ;
        RECT 135.645 170.550 135.915 171.365 ;
        RECT 134.650 169.955 135.395 170.125 ;
        RECT 134.650 169.325 134.820 169.955 ;
        RECT 133.285 169.155 134.820 169.325 ;
        RECT 134.990 168.985 135.395 169.785 ;
        RECT 135.565 169.155 135.915 170.550 ;
        RECT 136.085 171.075 136.645 171.365 ;
        RECT 136.815 171.075 137.065 171.535 ;
        RECT 136.085 169.705 136.335 171.075 ;
        RECT 137.685 170.905 138.015 171.265 ;
        RECT 136.625 170.715 138.015 170.905 ;
        RECT 138.405 170.725 138.645 171.535 ;
        RECT 138.815 170.725 139.145 171.365 ;
        RECT 139.315 170.725 139.585 171.535 ;
        RECT 139.765 170.990 145.110 171.535 ;
        RECT 136.625 170.625 136.795 170.715 ;
        RECT 136.505 170.295 136.795 170.625 ;
        RECT 136.965 170.295 137.305 170.545 ;
        RECT 137.525 170.295 138.200 170.545 ;
        RECT 138.385 170.295 138.735 170.545 ;
        RECT 136.625 170.045 136.795 170.295 ;
        RECT 136.625 169.875 137.565 170.045 ;
        RECT 137.935 169.935 138.200 170.295 ;
        RECT 138.905 170.125 139.075 170.725 ;
        RECT 139.245 170.295 139.595 170.545 ;
        RECT 141.350 170.160 141.690 170.990 ;
        RECT 145.745 170.785 146.955 171.535 ;
        RECT 138.395 169.955 139.075 170.125 ;
        RECT 136.085 169.155 136.545 169.705 ;
        RECT 136.735 168.985 137.065 169.705 ;
        RECT 137.265 169.325 137.565 169.875 ;
        RECT 137.735 168.985 138.015 169.655 ;
        RECT 138.395 169.170 138.725 169.955 ;
        RECT 139.255 168.985 139.585 170.125 ;
        RECT 143.170 169.420 143.520 170.670 ;
        RECT 145.745 170.075 146.265 170.615 ;
        RECT 146.435 170.245 146.955 170.785 ;
        RECT 139.765 168.985 145.110 169.420 ;
        RECT 145.745 168.985 146.955 170.075 ;
        RECT 17.320 168.815 147.040 168.985 ;
        RECT 17.405 167.725 18.615 168.815 ;
        RECT 18.785 167.725 22.295 168.815 ;
        RECT 22.465 167.725 23.675 168.815 ;
        RECT 17.405 167.015 17.925 167.555 ;
        RECT 18.095 167.185 18.615 167.725 ;
        RECT 18.785 167.035 20.435 167.555 ;
        RECT 20.605 167.205 22.295 167.725 ;
        RECT 17.405 166.265 18.615 167.015 ;
        RECT 18.785 166.265 22.295 167.035 ;
        RECT 22.465 167.015 22.985 167.555 ;
        RECT 23.155 167.185 23.675 167.725 ;
        RECT 23.905 167.675 24.115 168.815 ;
        RECT 24.285 167.665 24.615 168.645 ;
        RECT 24.785 167.675 25.015 168.815 ;
        RECT 25.685 168.095 26.145 168.645 ;
        RECT 26.335 168.095 26.665 168.815 ;
        RECT 22.465 166.265 23.675 167.015 ;
        RECT 23.905 166.265 24.115 167.085 ;
        RECT 24.285 167.065 24.535 167.665 ;
        RECT 24.705 167.255 25.035 167.505 ;
        RECT 24.285 166.435 24.615 167.065 ;
        RECT 24.785 166.265 25.015 167.085 ;
        RECT 25.685 166.725 25.935 168.095 ;
        RECT 26.865 167.925 27.165 168.475 ;
        RECT 27.335 168.145 27.615 168.815 ;
        RECT 26.225 167.755 27.165 167.925 ;
        RECT 26.225 167.505 26.395 167.755 ;
        RECT 27.535 167.505 27.800 167.865 ;
        RECT 27.985 167.725 29.655 168.815 ;
        RECT 26.105 167.175 26.395 167.505 ;
        RECT 26.565 167.255 26.905 167.505 ;
        RECT 27.125 167.255 27.800 167.505 ;
        RECT 26.225 167.085 26.395 167.175 ;
        RECT 26.225 166.895 27.615 167.085 ;
        RECT 25.685 166.435 26.245 166.725 ;
        RECT 26.415 166.265 26.665 166.725 ;
        RECT 27.285 166.535 27.615 166.895 ;
        RECT 27.985 167.035 28.735 167.555 ;
        RECT 28.905 167.205 29.655 167.725 ;
        RECT 30.285 167.650 30.575 168.815 ;
        RECT 30.750 168.425 31.085 168.645 ;
        RECT 32.090 168.435 32.445 168.815 ;
        RECT 30.750 167.805 31.005 168.425 ;
        RECT 31.255 168.265 31.485 168.305 ;
        RECT 32.615 168.265 32.865 168.645 ;
        RECT 31.255 168.065 32.865 168.265 ;
        RECT 31.255 167.975 31.440 168.065 ;
        RECT 32.030 168.055 32.865 168.065 ;
        RECT 33.115 168.035 33.365 168.815 ;
        RECT 33.535 167.965 33.795 168.645 ;
        RECT 31.595 167.865 31.925 167.895 ;
        RECT 31.595 167.805 33.395 167.865 ;
        RECT 30.750 167.695 33.455 167.805 ;
        RECT 30.750 167.635 31.925 167.695 ;
        RECT 33.255 167.660 33.455 167.695 ;
        RECT 30.745 167.255 31.235 167.455 ;
        RECT 31.425 167.255 31.900 167.465 ;
        RECT 27.985 166.265 29.655 167.035 ;
        RECT 30.285 166.265 30.575 166.990 ;
        RECT 30.750 166.265 31.205 167.030 ;
        RECT 31.680 166.855 31.900 167.255 ;
        RECT 32.145 167.255 32.475 167.465 ;
        RECT 32.145 166.855 32.355 167.255 ;
        RECT 32.645 167.220 33.055 167.525 ;
        RECT 33.285 167.085 33.455 167.660 ;
        RECT 33.185 166.965 33.455 167.085 ;
        RECT 32.610 166.920 33.455 166.965 ;
        RECT 32.610 166.795 33.365 166.920 ;
        RECT 32.610 166.645 32.780 166.795 ;
        RECT 33.625 166.765 33.795 167.965 ;
        RECT 33.965 167.635 34.285 168.815 ;
        RECT 34.455 167.795 34.655 168.585 ;
        RECT 34.845 168.225 35.345 168.645 ;
        RECT 35.835 168.355 36.045 168.815 ;
        RECT 34.845 168.015 35.685 168.225 ;
        RECT 34.455 167.625 34.775 167.795 ;
        RECT 33.965 167.255 34.425 167.455 ;
        RECT 34.595 167.425 34.775 167.625 ;
        RECT 34.945 167.595 35.345 167.845 ;
        RECT 34.595 167.255 34.960 167.425 ;
        RECT 35.175 167.175 35.345 167.595 ;
        RECT 31.480 166.435 32.780 166.645 ;
        RECT 33.035 166.265 33.365 166.625 ;
        RECT 33.535 166.435 33.795 166.765 ;
        RECT 33.965 167.005 34.995 167.045 ;
        RECT 35.515 167.005 35.685 168.015 ;
        RECT 33.965 166.875 35.165 167.005 ;
        RECT 33.965 166.460 34.305 166.875 ;
        RECT 34.475 166.265 34.645 166.705 ;
        RECT 34.835 166.655 35.165 166.875 ;
        RECT 35.335 166.825 35.685 167.005 ;
        RECT 35.855 166.845 36.095 168.170 ;
        RECT 36.265 167.675 36.525 168.815 ;
        RECT 36.695 167.665 37.025 168.645 ;
        RECT 37.195 167.675 37.475 168.815 ;
        RECT 37.645 168.380 42.990 168.815 ;
        RECT 36.285 167.255 36.620 167.505 ;
        RECT 36.790 167.065 36.960 167.665 ;
        RECT 37.130 167.235 37.465 167.505 ;
        RECT 34.835 166.475 36.095 166.655 ;
        RECT 36.265 166.435 36.960 167.065 ;
        RECT 37.165 166.265 37.475 167.065 ;
        RECT 39.230 166.810 39.570 167.640 ;
        RECT 41.050 167.130 41.400 168.380 ;
        RECT 43.630 168.305 45.285 168.595 ;
        RECT 43.630 167.965 45.220 168.135 ;
        RECT 45.455 168.015 45.735 168.815 ;
        RECT 43.630 167.675 43.950 167.965 ;
        RECT 45.050 167.845 45.220 167.965 ;
        RECT 43.630 166.935 43.980 167.505 ;
        RECT 44.150 167.175 44.860 167.795 ;
        RECT 45.050 167.675 45.775 167.845 ;
        RECT 45.945 167.675 46.215 168.645 ;
        RECT 46.385 168.260 46.990 168.815 ;
        RECT 47.165 168.305 47.645 168.645 ;
        RECT 47.815 168.270 48.070 168.815 ;
        RECT 46.385 168.160 47.000 168.260 ;
        RECT 46.815 168.135 47.000 168.160 ;
        RECT 45.605 167.505 45.775 167.675 ;
        RECT 45.030 167.175 45.435 167.505 ;
        RECT 45.605 167.175 45.875 167.505 ;
        RECT 45.605 167.005 45.775 167.175 ;
        RECT 44.165 166.835 45.775 167.005 ;
        RECT 46.045 166.940 46.215 167.675 ;
        RECT 46.385 167.540 46.645 167.990 ;
        RECT 46.815 167.890 47.145 168.135 ;
        RECT 47.315 167.815 48.070 168.065 ;
        RECT 48.240 167.945 48.515 168.645 ;
        RECT 47.300 167.780 48.070 167.815 ;
        RECT 47.285 167.770 48.070 167.780 ;
        RECT 47.280 167.755 48.175 167.770 ;
        RECT 47.260 167.740 48.175 167.755 ;
        RECT 47.240 167.730 48.175 167.740 ;
        RECT 47.215 167.720 48.175 167.730 ;
        RECT 47.145 167.690 48.175 167.720 ;
        RECT 47.125 167.660 48.175 167.690 ;
        RECT 47.105 167.630 48.175 167.660 ;
        RECT 47.075 167.605 48.175 167.630 ;
        RECT 47.040 167.570 48.175 167.605 ;
        RECT 47.010 167.565 48.175 167.570 ;
        RECT 47.010 167.560 47.400 167.565 ;
        RECT 47.010 167.550 47.375 167.560 ;
        RECT 47.010 167.545 47.360 167.550 ;
        RECT 47.010 167.540 47.345 167.545 ;
        RECT 46.385 167.535 47.345 167.540 ;
        RECT 46.385 167.525 47.335 167.535 ;
        RECT 46.385 167.520 47.325 167.525 ;
        RECT 46.385 167.510 47.315 167.520 ;
        RECT 46.385 167.500 47.310 167.510 ;
        RECT 46.385 167.495 47.305 167.500 ;
        RECT 46.385 167.480 47.295 167.495 ;
        RECT 46.385 167.465 47.290 167.480 ;
        RECT 46.385 167.440 47.280 167.465 ;
        RECT 46.385 167.370 47.275 167.440 ;
        RECT 37.645 166.265 42.990 166.810 ;
        RECT 43.635 166.265 43.965 166.765 ;
        RECT 44.165 166.485 44.335 166.835 ;
        RECT 44.535 166.265 44.865 166.665 ;
        RECT 45.035 166.485 45.205 166.835 ;
        RECT 45.375 166.265 45.755 166.665 ;
        RECT 45.945 166.595 46.215 166.940 ;
        RECT 46.385 166.815 46.935 167.200 ;
        RECT 47.105 166.645 47.275 167.370 ;
        RECT 46.385 166.475 47.275 166.645 ;
        RECT 47.445 166.970 47.775 167.395 ;
        RECT 47.945 167.170 48.175 167.565 ;
        RECT 47.445 166.485 47.665 166.970 ;
        RECT 48.345 166.915 48.515 167.945 ;
        RECT 48.725 167.675 48.955 168.815 ;
        RECT 49.125 167.665 49.455 168.645 ;
        RECT 49.625 167.675 49.835 168.815 ;
        RECT 50.065 167.725 52.655 168.815 ;
        RECT 48.705 167.255 49.035 167.505 ;
        RECT 47.835 166.265 48.085 166.805 ;
        RECT 48.255 166.435 48.515 166.915 ;
        RECT 48.725 166.265 48.955 167.085 ;
        RECT 49.205 167.065 49.455 167.665 ;
        RECT 49.125 166.435 49.455 167.065 ;
        RECT 49.625 166.265 49.835 167.085 ;
        RECT 50.065 167.035 51.275 167.555 ;
        RECT 51.445 167.205 52.655 167.725 ;
        RECT 53.325 167.675 53.555 168.815 ;
        RECT 53.725 167.665 54.055 168.645 ;
        RECT 54.225 167.675 54.435 168.815 ;
        RECT 54.665 167.725 55.875 168.815 ;
        RECT 53.305 167.255 53.635 167.505 ;
        RECT 50.065 166.265 52.655 167.035 ;
        RECT 53.325 166.265 53.555 167.085 ;
        RECT 53.805 167.065 54.055 167.665 ;
        RECT 53.725 166.435 54.055 167.065 ;
        RECT 54.225 166.265 54.435 167.085 ;
        RECT 54.665 167.015 55.185 167.555 ;
        RECT 55.355 167.185 55.875 167.725 ;
        RECT 56.045 167.650 56.335 168.815 ;
        RECT 56.975 167.675 57.305 168.815 ;
        RECT 57.835 167.845 58.165 168.630 ;
        RECT 58.435 168.145 58.605 168.645 ;
        RECT 58.775 168.315 59.105 168.815 ;
        RECT 58.435 167.975 59.100 168.145 ;
        RECT 57.485 167.675 58.165 167.845 ;
        RECT 56.965 167.255 57.315 167.505 ;
        RECT 57.485 167.075 57.655 167.675 ;
        RECT 57.825 167.255 58.175 167.505 ;
        RECT 58.350 167.155 58.700 167.805 ;
        RECT 54.665 166.265 55.875 167.015 ;
        RECT 56.045 166.265 56.335 166.990 ;
        RECT 56.975 166.265 57.245 167.075 ;
        RECT 57.415 166.435 57.745 167.075 ;
        RECT 57.915 166.265 58.155 167.075 ;
        RECT 58.870 166.985 59.100 167.975 ;
        RECT 58.435 166.815 59.100 166.985 ;
        RECT 58.435 166.525 58.605 166.815 ;
        RECT 58.775 166.265 59.105 166.645 ;
        RECT 59.275 166.525 59.460 168.645 ;
        RECT 59.700 168.355 59.965 168.815 ;
        RECT 60.135 168.220 60.385 168.645 ;
        RECT 60.595 168.370 61.700 168.540 ;
        RECT 60.080 168.090 60.385 168.220 ;
        RECT 59.630 166.895 59.910 167.845 ;
        RECT 60.080 166.985 60.250 168.090 ;
        RECT 60.420 167.305 60.660 167.900 ;
        RECT 60.830 167.835 61.360 168.200 ;
        RECT 60.830 167.135 61.000 167.835 ;
        RECT 61.530 167.755 61.700 168.370 ;
        RECT 61.870 168.015 62.040 168.815 ;
        RECT 62.210 168.315 62.460 168.645 ;
        RECT 62.685 168.345 63.570 168.515 ;
        RECT 61.530 167.665 62.040 167.755 ;
        RECT 60.080 166.855 60.305 166.985 ;
        RECT 60.475 166.915 61.000 167.135 ;
        RECT 61.170 167.495 62.040 167.665 ;
        RECT 59.715 166.265 59.965 166.725 ;
        RECT 60.135 166.715 60.305 166.855 ;
        RECT 61.170 166.715 61.340 167.495 ;
        RECT 61.870 167.425 62.040 167.495 ;
        RECT 61.550 167.245 61.750 167.275 ;
        RECT 62.210 167.245 62.380 168.315 ;
        RECT 62.550 167.425 62.740 168.145 ;
        RECT 61.550 166.945 62.380 167.245 ;
        RECT 62.910 167.215 63.230 168.175 ;
        RECT 60.135 166.545 60.470 166.715 ;
        RECT 60.665 166.545 61.340 166.715 ;
        RECT 61.660 166.265 62.030 166.765 ;
        RECT 62.210 166.715 62.380 166.945 ;
        RECT 62.765 166.885 63.230 167.215 ;
        RECT 63.400 167.505 63.570 168.345 ;
        RECT 63.750 168.315 64.065 168.815 ;
        RECT 64.295 168.085 64.635 168.645 ;
        RECT 63.740 167.710 64.635 168.085 ;
        RECT 64.805 167.805 64.975 168.815 ;
        RECT 64.445 167.505 64.635 167.710 ;
        RECT 65.145 167.755 65.475 168.600 ;
        RECT 65.765 167.755 66.095 168.600 ;
        RECT 66.265 167.805 66.435 168.815 ;
        RECT 66.605 168.085 66.945 168.645 ;
        RECT 67.175 168.315 67.490 168.815 ;
        RECT 67.670 168.345 68.555 168.515 ;
        RECT 65.145 167.675 65.535 167.755 ;
        RECT 65.320 167.625 65.535 167.675 ;
        RECT 63.400 167.175 64.275 167.505 ;
        RECT 64.445 167.175 65.195 167.505 ;
        RECT 63.400 166.715 63.570 167.175 ;
        RECT 64.445 167.005 64.645 167.175 ;
        RECT 65.365 167.045 65.535 167.625 ;
        RECT 65.310 167.005 65.535 167.045 ;
        RECT 62.210 166.545 62.615 166.715 ;
        RECT 62.785 166.545 63.570 166.715 ;
        RECT 63.845 166.265 64.055 166.795 ;
        RECT 64.315 166.480 64.645 167.005 ;
        RECT 65.155 166.920 65.535 167.005 ;
        RECT 65.705 167.675 66.095 167.755 ;
        RECT 66.605 167.710 67.500 168.085 ;
        RECT 65.705 167.625 65.920 167.675 ;
        RECT 65.705 167.045 65.875 167.625 ;
        RECT 66.605 167.505 66.795 167.710 ;
        RECT 67.670 167.505 67.840 168.345 ;
        RECT 68.780 168.315 69.030 168.645 ;
        RECT 66.045 167.175 66.795 167.505 ;
        RECT 66.965 167.175 67.840 167.505 ;
        RECT 65.705 167.005 65.930 167.045 ;
        RECT 66.595 167.005 66.795 167.175 ;
        RECT 65.705 166.920 66.085 167.005 ;
        RECT 64.815 166.265 64.985 166.875 ;
        RECT 65.155 166.485 65.485 166.920 ;
        RECT 65.755 166.485 66.085 166.920 ;
        RECT 66.255 166.265 66.425 166.875 ;
        RECT 66.595 166.480 66.925 167.005 ;
        RECT 67.185 166.265 67.395 166.795 ;
        RECT 67.670 166.715 67.840 167.175 ;
        RECT 68.010 167.215 68.330 168.175 ;
        RECT 68.500 167.425 68.690 168.145 ;
        RECT 68.860 167.245 69.030 168.315 ;
        RECT 69.200 168.015 69.370 168.815 ;
        RECT 69.540 168.370 70.645 168.540 ;
        RECT 69.540 167.755 69.710 168.370 ;
        RECT 70.855 168.220 71.105 168.645 ;
        RECT 71.275 168.355 71.540 168.815 ;
        RECT 69.880 167.835 70.410 168.200 ;
        RECT 70.855 168.090 71.160 168.220 ;
        RECT 69.200 167.665 69.710 167.755 ;
        RECT 69.200 167.495 70.070 167.665 ;
        RECT 69.200 167.425 69.370 167.495 ;
        RECT 69.490 167.245 69.690 167.275 ;
        RECT 68.010 166.885 68.475 167.215 ;
        RECT 68.860 166.945 69.690 167.245 ;
        RECT 68.860 166.715 69.030 166.945 ;
        RECT 67.670 166.545 68.455 166.715 ;
        RECT 68.625 166.545 69.030 166.715 ;
        RECT 69.210 166.265 69.580 166.765 ;
        RECT 69.900 166.715 70.070 167.495 ;
        RECT 70.240 167.135 70.410 167.835 ;
        RECT 70.580 167.305 70.820 167.900 ;
        RECT 70.240 166.915 70.765 167.135 ;
        RECT 70.990 166.985 71.160 168.090 ;
        RECT 70.935 166.855 71.160 166.985 ;
        RECT 71.330 166.895 71.610 167.845 ;
        RECT 70.935 166.715 71.105 166.855 ;
        RECT 69.900 166.545 70.575 166.715 ;
        RECT 70.770 166.545 71.105 166.715 ;
        RECT 71.275 166.265 71.525 166.725 ;
        RECT 71.780 166.525 71.965 168.645 ;
        RECT 72.135 168.315 72.465 168.815 ;
        RECT 72.635 168.145 72.805 168.645 ;
        RECT 73.065 168.380 78.410 168.815 ;
        RECT 72.140 167.975 72.805 168.145 ;
        RECT 72.140 166.985 72.370 167.975 ;
        RECT 72.540 167.155 72.890 167.805 ;
        RECT 72.140 166.815 72.805 166.985 ;
        RECT 72.135 166.265 72.465 166.645 ;
        RECT 72.635 166.525 72.805 166.815 ;
        RECT 74.650 166.810 74.990 167.640 ;
        RECT 76.470 167.130 76.820 168.380 ;
        RECT 78.585 167.725 81.175 168.815 ;
        RECT 78.585 167.035 79.795 167.555 ;
        RECT 79.965 167.205 81.175 167.725 ;
        RECT 81.805 167.650 82.095 168.815 ;
        RECT 82.265 167.725 83.935 168.815 ;
        RECT 84.680 168.185 84.965 168.645 ;
        RECT 85.135 168.355 85.405 168.815 ;
        RECT 84.680 167.965 85.635 168.185 ;
        RECT 82.265 167.035 83.015 167.555 ;
        RECT 83.185 167.205 83.935 167.725 ;
        RECT 84.565 167.235 85.255 167.795 ;
        RECT 85.425 167.065 85.635 167.965 ;
        RECT 73.065 166.265 78.410 166.810 ;
        RECT 78.585 166.265 81.175 167.035 ;
        RECT 81.805 166.265 82.095 166.990 ;
        RECT 82.265 166.265 83.935 167.035 ;
        RECT 84.680 166.895 85.635 167.065 ;
        RECT 85.805 167.795 86.205 168.645 ;
        RECT 86.395 168.185 86.675 168.645 ;
        RECT 87.195 168.355 87.520 168.815 ;
        RECT 86.395 167.965 87.520 168.185 ;
        RECT 85.805 167.235 86.900 167.795 ;
        RECT 87.070 167.505 87.520 167.965 ;
        RECT 87.690 167.675 88.075 168.645 ;
        RECT 88.245 167.725 91.755 168.815 ;
        RECT 91.925 167.725 93.135 168.815 ;
        RECT 93.395 168.145 93.565 168.645 ;
        RECT 93.735 168.315 94.065 168.815 ;
        RECT 93.395 167.975 94.060 168.145 ;
        RECT 84.680 166.435 84.965 166.895 ;
        RECT 85.135 166.265 85.405 166.725 ;
        RECT 85.805 166.435 86.205 167.235 ;
        RECT 87.070 167.175 87.625 167.505 ;
        RECT 87.070 167.065 87.520 167.175 ;
        RECT 86.395 166.895 87.520 167.065 ;
        RECT 87.795 167.005 88.075 167.675 ;
        RECT 86.395 166.435 86.675 166.895 ;
        RECT 87.195 166.265 87.520 166.725 ;
        RECT 87.690 166.435 88.075 167.005 ;
        RECT 88.245 167.035 89.895 167.555 ;
        RECT 90.065 167.205 91.755 167.725 ;
        RECT 88.245 166.265 91.755 167.035 ;
        RECT 91.925 167.015 92.445 167.555 ;
        RECT 92.615 167.185 93.135 167.725 ;
        RECT 93.310 167.155 93.660 167.805 ;
        RECT 91.925 166.265 93.135 167.015 ;
        RECT 93.830 166.985 94.060 167.975 ;
        RECT 93.395 166.815 94.060 166.985 ;
        RECT 93.395 166.525 93.565 166.815 ;
        RECT 93.735 166.265 94.065 166.645 ;
        RECT 94.235 166.525 94.420 168.645 ;
        RECT 94.660 168.355 94.925 168.815 ;
        RECT 95.095 168.220 95.345 168.645 ;
        RECT 95.555 168.370 96.660 168.540 ;
        RECT 95.040 168.090 95.345 168.220 ;
        RECT 94.590 166.895 94.870 167.845 ;
        RECT 95.040 166.985 95.210 168.090 ;
        RECT 95.380 167.305 95.620 167.900 ;
        RECT 95.790 167.835 96.320 168.200 ;
        RECT 95.790 167.135 95.960 167.835 ;
        RECT 96.490 167.755 96.660 168.370 ;
        RECT 96.830 168.015 97.000 168.815 ;
        RECT 97.170 168.315 97.420 168.645 ;
        RECT 97.645 168.345 98.530 168.515 ;
        RECT 96.490 167.665 97.000 167.755 ;
        RECT 95.040 166.855 95.265 166.985 ;
        RECT 95.435 166.915 95.960 167.135 ;
        RECT 96.130 167.495 97.000 167.665 ;
        RECT 94.675 166.265 94.925 166.725 ;
        RECT 95.095 166.715 95.265 166.855 ;
        RECT 96.130 166.715 96.300 167.495 ;
        RECT 96.830 167.425 97.000 167.495 ;
        RECT 96.510 167.245 96.710 167.275 ;
        RECT 97.170 167.245 97.340 168.315 ;
        RECT 97.510 167.425 97.700 168.145 ;
        RECT 96.510 166.945 97.340 167.245 ;
        RECT 97.870 167.215 98.190 168.175 ;
        RECT 95.095 166.545 95.430 166.715 ;
        RECT 95.625 166.545 96.300 166.715 ;
        RECT 96.620 166.265 96.990 166.765 ;
        RECT 97.170 166.715 97.340 166.945 ;
        RECT 97.725 166.885 98.190 167.215 ;
        RECT 98.360 167.505 98.530 168.345 ;
        RECT 98.710 168.315 99.025 168.815 ;
        RECT 99.255 168.085 99.595 168.645 ;
        RECT 98.700 167.710 99.595 168.085 ;
        RECT 99.765 167.805 99.935 168.815 ;
        RECT 99.405 167.505 99.595 167.710 ;
        RECT 100.105 167.755 100.435 168.600 ;
        RECT 100.105 167.675 100.495 167.755 ;
        RECT 100.280 167.625 100.495 167.675 ;
        RECT 98.360 167.175 99.235 167.505 ;
        RECT 99.405 167.175 100.155 167.505 ;
        RECT 98.360 166.715 98.530 167.175 ;
        RECT 99.405 167.005 99.605 167.175 ;
        RECT 100.325 167.045 100.495 167.625 ;
        RECT 100.270 167.005 100.495 167.045 ;
        RECT 97.170 166.545 97.575 166.715 ;
        RECT 97.745 166.545 98.530 166.715 ;
        RECT 98.805 166.265 99.015 166.795 ;
        RECT 99.275 166.480 99.605 167.005 ;
        RECT 100.115 166.920 100.495 167.005 ;
        RECT 100.670 167.675 101.005 168.645 ;
        RECT 101.175 167.675 101.345 168.815 ;
        RECT 101.515 168.475 103.545 168.645 ;
        RECT 100.670 167.005 100.840 167.675 ;
        RECT 101.515 167.505 101.685 168.475 ;
        RECT 101.010 167.175 101.265 167.505 ;
        RECT 101.490 167.175 101.685 167.505 ;
        RECT 101.855 168.135 102.980 168.305 ;
        RECT 101.095 167.005 101.265 167.175 ;
        RECT 101.855 167.005 102.025 168.135 ;
        RECT 99.775 166.265 99.945 166.875 ;
        RECT 100.115 166.485 100.445 166.920 ;
        RECT 100.670 166.435 100.925 167.005 ;
        RECT 101.095 166.835 102.025 167.005 ;
        RECT 102.195 167.795 103.205 167.965 ;
        RECT 102.195 166.995 102.365 167.795 ;
        RECT 102.570 167.115 102.845 167.595 ;
        RECT 102.565 166.945 102.845 167.115 ;
        RECT 101.850 166.800 102.025 166.835 ;
        RECT 101.095 166.265 101.425 166.665 ;
        RECT 101.850 166.435 102.380 166.800 ;
        RECT 102.570 166.435 102.845 166.945 ;
        RECT 103.015 166.435 103.205 167.795 ;
        RECT 103.375 167.810 103.545 168.475 ;
        RECT 103.715 168.055 103.885 168.815 ;
        RECT 104.120 168.055 104.635 168.465 ;
        RECT 103.375 167.620 104.125 167.810 ;
        RECT 104.295 167.245 104.635 168.055 ;
        RECT 105.735 168.205 106.065 168.635 ;
        RECT 106.245 168.375 106.440 168.815 ;
        RECT 106.610 168.205 106.940 168.635 ;
        RECT 105.735 168.035 106.940 168.205 ;
        RECT 105.735 167.705 106.630 168.035 ;
        RECT 107.110 167.865 107.385 168.635 ;
        RECT 106.800 167.675 107.385 167.865 ;
        RECT 103.405 167.075 104.635 167.245 ;
        RECT 105.740 167.175 106.035 167.505 ;
        RECT 106.215 167.175 106.630 167.505 ;
        RECT 103.385 166.265 103.895 166.800 ;
        RECT 104.115 166.470 104.360 167.075 ;
        RECT 105.735 166.265 106.035 166.995 ;
        RECT 106.215 166.555 106.445 167.175 ;
        RECT 106.800 167.005 106.975 167.675 ;
        RECT 107.565 167.650 107.855 168.815 ;
        RECT 108.065 167.675 108.295 168.815 ;
        RECT 108.465 167.665 108.795 168.645 ;
        RECT 108.965 167.675 109.175 168.815 ;
        RECT 109.405 167.675 109.665 168.645 ;
        RECT 109.835 168.390 110.220 168.815 ;
        RECT 110.390 168.220 110.645 168.645 ;
        RECT 109.835 168.025 110.645 168.220 ;
        RECT 106.645 166.825 106.975 167.005 ;
        RECT 107.145 166.855 107.385 167.505 ;
        RECT 108.045 167.255 108.375 167.505 ;
        RECT 106.645 166.445 106.870 166.825 ;
        RECT 107.040 166.265 107.370 166.655 ;
        RECT 107.565 166.265 107.855 166.990 ;
        RECT 108.065 166.265 108.295 167.085 ;
        RECT 108.545 167.065 108.795 167.665 ;
        RECT 108.465 166.435 108.795 167.065 ;
        RECT 108.965 166.265 109.175 167.085 ;
        RECT 109.405 167.005 109.590 167.675 ;
        RECT 109.835 167.505 110.185 168.025 ;
        RECT 110.835 167.855 111.080 168.645 ;
        RECT 111.250 168.390 111.635 168.815 ;
        RECT 111.805 168.220 112.080 168.645 ;
        RECT 109.760 167.175 110.185 167.505 ;
        RECT 110.355 167.675 111.080 167.855 ;
        RECT 111.250 168.025 112.080 168.220 ;
        RECT 110.355 167.175 111.005 167.675 ;
        RECT 111.250 167.505 111.600 168.025 ;
        RECT 112.250 167.855 112.675 168.645 ;
        RECT 112.845 168.390 113.230 168.815 ;
        RECT 113.400 168.220 113.835 168.645 ;
        RECT 111.175 167.175 111.600 167.505 ;
        RECT 111.770 167.675 112.675 167.855 ;
        RECT 112.845 168.050 113.835 168.220 ;
        RECT 111.770 167.175 112.600 167.675 ;
        RECT 112.845 167.505 113.180 168.050 ;
        RECT 112.770 167.175 113.180 167.505 ;
        RECT 113.350 167.175 113.835 167.880 ;
        RECT 114.005 167.675 114.280 168.645 ;
        RECT 114.490 168.015 114.770 168.815 ;
        RECT 114.940 168.305 116.990 168.595 ;
        RECT 114.940 167.965 116.570 168.135 ;
        RECT 114.940 167.845 115.110 167.965 ;
        RECT 114.450 167.675 115.110 167.845 ;
        RECT 109.835 167.005 110.185 167.175 ;
        RECT 110.835 167.005 111.005 167.175 ;
        RECT 111.250 167.005 111.600 167.175 ;
        RECT 112.250 167.005 112.600 167.175 ;
        RECT 112.845 167.005 113.180 167.175 ;
        RECT 109.405 166.435 109.665 167.005 ;
        RECT 109.835 166.835 110.645 167.005 ;
        RECT 109.835 166.265 110.220 166.665 ;
        RECT 110.390 166.435 110.645 166.835 ;
        RECT 110.835 166.435 111.080 167.005 ;
        RECT 111.250 166.835 112.060 167.005 ;
        RECT 111.250 166.265 111.635 166.665 ;
        RECT 111.805 166.435 112.060 166.835 ;
        RECT 112.250 166.435 112.675 167.005 ;
        RECT 112.845 166.835 113.835 167.005 ;
        RECT 112.845 166.265 113.230 166.665 ;
        RECT 113.400 166.435 113.835 166.835 ;
        RECT 114.005 166.940 114.175 167.675 ;
        RECT 114.450 167.505 114.620 167.675 ;
        RECT 114.345 167.175 114.620 167.505 ;
        RECT 114.790 167.175 115.170 167.505 ;
        RECT 115.340 167.175 116.080 167.795 ;
        RECT 116.250 167.675 116.570 167.965 ;
        RECT 116.765 167.505 117.005 168.100 ;
        RECT 117.175 167.740 117.515 168.815 ;
        RECT 117.885 168.145 118.165 168.815 ;
        RECT 118.335 167.925 118.635 168.475 ;
        RECT 118.835 168.095 119.165 168.815 ;
        RECT 119.355 168.095 119.815 168.645 ;
        RECT 117.700 167.505 117.965 167.865 ;
        RECT 118.335 167.755 119.275 167.925 ;
        RECT 119.105 167.505 119.275 167.755 ;
        RECT 116.350 167.175 117.005 167.505 ;
        RECT 114.450 167.005 114.620 167.175 ;
        RECT 114.005 166.595 114.280 166.940 ;
        RECT 114.450 166.835 116.035 167.005 ;
        RECT 114.470 166.265 114.850 166.665 ;
        RECT 115.020 166.485 115.190 166.835 ;
        RECT 115.360 166.265 115.690 166.665 ;
        RECT 115.865 166.485 116.035 166.835 ;
        RECT 116.235 166.265 116.565 166.765 ;
        RECT 116.760 166.485 117.005 167.175 ;
        RECT 117.175 166.935 117.515 167.505 ;
        RECT 117.700 167.255 118.375 167.505 ;
        RECT 118.595 167.255 118.935 167.505 ;
        RECT 119.105 167.175 119.395 167.505 ;
        RECT 119.105 167.085 119.275 167.175 ;
        RECT 117.885 166.895 119.275 167.085 ;
        RECT 117.175 166.265 117.515 166.765 ;
        RECT 117.885 166.535 118.215 166.895 ;
        RECT 119.565 166.725 119.815 168.095 ;
        RECT 119.985 167.675 120.265 168.815 ;
        RECT 120.435 167.665 120.765 168.645 ;
        RECT 120.935 167.675 121.195 168.815 ;
        RECT 121.365 167.725 122.575 168.815 ;
        RECT 119.995 167.235 120.330 167.505 ;
        RECT 120.500 167.065 120.670 167.665 ;
        RECT 120.840 167.255 121.175 167.505 ;
        RECT 118.835 166.265 119.085 166.725 ;
        RECT 119.255 166.435 119.815 166.725 ;
        RECT 119.985 166.265 120.295 167.065 ;
        RECT 120.500 166.435 121.195 167.065 ;
        RECT 121.365 167.015 121.885 167.555 ;
        RECT 122.055 167.185 122.575 167.725 ;
        RECT 122.745 167.675 123.020 168.645 ;
        RECT 123.230 168.015 123.510 168.815 ;
        RECT 123.680 168.305 125.295 168.635 ;
        RECT 123.680 167.965 124.855 168.135 ;
        RECT 123.680 167.845 123.850 167.965 ;
        RECT 123.190 167.675 123.850 167.845 ;
        RECT 121.365 166.265 122.575 167.015 ;
        RECT 122.745 166.940 122.915 167.675 ;
        RECT 123.190 167.505 123.360 167.675 ;
        RECT 124.110 167.505 124.355 167.795 ;
        RECT 124.525 167.675 124.855 167.965 ;
        RECT 125.115 167.505 125.285 168.065 ;
        RECT 125.535 167.675 125.795 168.815 ;
        RECT 126.055 168.195 126.225 168.625 ;
        RECT 126.395 168.365 126.725 168.815 ;
        RECT 126.055 167.965 126.730 168.195 ;
        RECT 123.085 167.175 123.360 167.505 ;
        RECT 123.530 167.175 124.355 167.505 ;
        RECT 124.570 167.175 125.285 167.505 ;
        RECT 125.455 167.255 125.790 167.505 ;
        RECT 123.190 167.005 123.360 167.175 ;
        RECT 125.035 167.085 125.285 167.175 ;
        RECT 122.745 166.595 123.020 166.940 ;
        RECT 123.190 166.835 124.855 167.005 ;
        RECT 123.210 166.265 123.585 166.665 ;
        RECT 123.755 166.485 123.925 166.835 ;
        RECT 124.095 166.265 124.425 166.665 ;
        RECT 124.595 166.435 124.855 166.835 ;
        RECT 125.035 166.665 125.365 167.085 ;
        RECT 125.535 166.265 125.795 167.085 ;
        RECT 126.025 166.945 126.325 167.795 ;
        RECT 126.495 167.315 126.730 167.965 ;
        RECT 126.900 167.655 127.185 168.600 ;
        RECT 127.365 168.345 128.050 168.815 ;
        RECT 127.360 167.825 128.055 168.135 ;
        RECT 128.230 167.760 128.535 168.545 ;
        RECT 126.900 167.505 127.760 167.655 ;
        RECT 126.900 167.485 128.185 167.505 ;
        RECT 126.495 166.985 127.030 167.315 ;
        RECT 127.200 167.125 128.185 167.485 ;
        RECT 126.495 166.835 126.715 166.985 ;
        RECT 125.970 166.265 126.305 166.770 ;
        RECT 126.475 166.460 126.715 166.835 ;
        RECT 127.200 166.790 127.370 167.125 ;
        RECT 128.360 166.955 128.535 167.760 ;
        RECT 128.735 168.205 129.065 168.635 ;
        RECT 129.245 168.375 129.440 168.815 ;
        RECT 129.610 168.205 129.940 168.635 ;
        RECT 128.735 168.035 129.940 168.205 ;
        RECT 128.735 167.705 129.630 168.035 ;
        RECT 130.110 167.865 130.385 168.635 ;
        RECT 129.800 167.675 130.385 167.865 ;
        RECT 130.575 167.675 130.905 168.815 ;
        RECT 131.435 167.845 131.765 168.630 ;
        RECT 131.085 167.675 131.765 167.845 ;
        RECT 131.945 167.725 133.155 168.815 ;
        RECT 128.740 167.175 129.035 167.505 ;
        RECT 129.215 167.175 129.630 167.505 ;
        RECT 126.995 166.595 127.370 166.790 ;
        RECT 126.995 166.450 127.165 166.595 ;
        RECT 127.730 166.265 128.125 166.760 ;
        RECT 128.295 166.435 128.535 166.955 ;
        RECT 128.735 166.265 129.035 166.995 ;
        RECT 129.215 166.555 129.445 167.175 ;
        RECT 129.800 167.005 129.975 167.675 ;
        RECT 129.645 166.825 129.975 167.005 ;
        RECT 130.145 166.855 130.385 167.505 ;
        RECT 130.565 167.255 130.915 167.505 ;
        RECT 131.085 167.075 131.255 167.675 ;
        RECT 131.425 167.255 131.775 167.505 ;
        RECT 129.645 166.445 129.870 166.825 ;
        RECT 130.040 166.265 130.370 166.655 ;
        RECT 130.575 166.265 130.845 167.075 ;
        RECT 131.015 166.435 131.345 167.075 ;
        RECT 131.515 166.265 131.755 167.075 ;
        RECT 131.945 167.015 132.465 167.555 ;
        RECT 132.635 167.185 133.155 167.725 ;
        RECT 133.325 167.650 133.615 168.815 ;
        RECT 133.785 168.305 134.975 168.595 ;
        RECT 133.805 167.965 134.975 168.135 ;
        RECT 135.145 168.015 135.425 168.815 ;
        RECT 133.805 167.675 134.130 167.965 ;
        RECT 134.805 167.845 134.975 167.965 ;
        RECT 134.300 167.505 134.495 167.795 ;
        RECT 134.805 167.675 135.465 167.845 ;
        RECT 135.635 167.675 135.910 168.645 ;
        RECT 136.085 167.675 136.345 168.815 ;
        RECT 135.295 167.505 135.465 167.675 ;
        RECT 133.785 167.175 134.130 167.505 ;
        RECT 134.300 167.175 135.125 167.505 ;
        RECT 135.295 167.175 135.570 167.505 ;
        RECT 131.945 166.265 133.155 167.015 ;
        RECT 135.295 167.005 135.465 167.175 ;
        RECT 133.325 166.265 133.615 166.990 ;
        RECT 133.800 166.835 135.465 167.005 ;
        RECT 135.740 166.940 135.910 167.675 ;
        RECT 136.515 167.665 136.845 168.645 ;
        RECT 137.015 167.675 137.295 168.815 ;
        RECT 137.465 168.380 142.810 168.815 ;
        RECT 136.105 167.255 136.440 167.505 ;
        RECT 136.610 167.065 136.780 167.665 ;
        RECT 136.950 167.235 137.285 167.505 ;
        RECT 133.800 166.485 134.055 166.835 ;
        RECT 134.225 166.265 134.555 166.665 ;
        RECT 134.725 166.485 134.895 166.835 ;
        RECT 135.065 166.265 135.445 166.665 ;
        RECT 135.635 166.595 135.910 166.940 ;
        RECT 136.085 166.435 136.780 167.065 ;
        RECT 136.985 166.265 137.295 167.065 ;
        RECT 139.050 166.810 139.390 167.640 ;
        RECT 140.870 167.130 141.220 168.380 ;
        RECT 143.910 167.665 144.170 168.815 ;
        RECT 144.345 167.740 144.600 168.645 ;
        RECT 144.770 168.055 145.100 168.815 ;
        RECT 145.315 167.885 145.485 168.645 ;
        RECT 137.465 166.265 142.810 166.810 ;
        RECT 143.910 166.265 144.170 167.105 ;
        RECT 144.345 167.010 144.515 167.740 ;
        RECT 144.770 167.715 145.485 167.885 ;
        RECT 145.745 167.725 146.955 168.815 ;
        RECT 144.770 167.505 144.940 167.715 ;
        RECT 144.685 167.175 144.940 167.505 ;
        RECT 144.345 166.435 144.600 167.010 ;
        RECT 144.770 166.985 144.940 167.175 ;
        RECT 145.220 167.165 145.575 167.535 ;
        RECT 145.745 167.185 146.265 167.725 ;
        RECT 146.435 167.015 146.955 167.555 ;
        RECT 144.770 166.815 145.485 166.985 ;
        RECT 144.770 166.265 145.100 166.645 ;
        RECT 145.315 166.435 145.485 166.815 ;
        RECT 145.745 166.265 146.955 167.015 ;
        RECT 17.320 166.095 147.040 166.265 ;
        RECT 17.405 165.345 18.615 166.095 ;
        RECT 17.405 164.805 17.925 165.345 ;
        RECT 18.785 165.325 20.455 166.095 ;
        RECT 20.660 165.355 21.275 165.925 ;
        RECT 21.445 165.585 21.660 166.095 ;
        RECT 21.890 165.585 22.170 165.915 ;
        RECT 22.350 165.585 22.590 166.095 ;
        RECT 18.095 164.635 18.615 165.175 ;
        RECT 18.785 164.805 19.535 165.325 ;
        RECT 19.705 164.635 20.455 165.155 ;
        RECT 17.405 163.545 18.615 164.635 ;
        RECT 18.785 163.545 20.455 164.635 ;
        RECT 20.660 164.335 20.975 165.355 ;
        RECT 21.145 164.685 21.315 165.185 ;
        RECT 21.565 164.855 21.830 165.415 ;
        RECT 22.000 164.685 22.170 165.585 ;
        RECT 22.925 165.445 23.185 165.925 ;
        RECT 23.355 165.555 23.605 166.095 ;
        RECT 22.340 164.855 22.695 165.415 ;
        RECT 21.145 164.515 22.570 164.685 ;
        RECT 20.660 163.715 21.195 164.335 ;
        RECT 21.365 163.545 21.695 164.345 ;
        RECT 22.180 164.340 22.570 164.515 ;
        RECT 22.925 164.415 23.095 165.445 ;
        RECT 23.775 165.390 23.995 165.875 ;
        RECT 23.265 164.795 23.495 165.190 ;
        RECT 23.665 164.965 23.995 165.390 ;
        RECT 24.165 165.715 25.055 165.885 ;
        RECT 24.165 164.990 24.335 165.715 ;
        RECT 24.505 165.160 25.055 165.545 ;
        RECT 25.260 165.355 25.875 165.925 ;
        RECT 26.045 165.585 26.260 166.095 ;
        RECT 26.490 165.585 26.770 165.915 ;
        RECT 26.950 165.585 27.190 166.095 ;
        RECT 28.315 165.695 28.645 166.095 ;
        RECT 24.165 164.920 25.055 164.990 ;
        RECT 24.160 164.895 25.055 164.920 ;
        RECT 24.150 164.880 25.055 164.895 ;
        RECT 24.145 164.865 25.055 164.880 ;
        RECT 24.135 164.860 25.055 164.865 ;
        RECT 24.130 164.850 25.055 164.860 ;
        RECT 24.125 164.840 25.055 164.850 ;
        RECT 24.115 164.835 25.055 164.840 ;
        RECT 24.105 164.825 25.055 164.835 ;
        RECT 24.095 164.820 25.055 164.825 ;
        RECT 24.095 164.815 24.430 164.820 ;
        RECT 24.080 164.810 24.430 164.815 ;
        RECT 24.065 164.800 24.430 164.810 ;
        RECT 24.040 164.795 24.430 164.800 ;
        RECT 23.265 164.790 24.430 164.795 ;
        RECT 23.265 164.755 24.400 164.790 ;
        RECT 23.265 164.730 24.365 164.755 ;
        RECT 23.265 164.700 24.335 164.730 ;
        RECT 23.265 164.670 24.315 164.700 ;
        RECT 23.265 164.640 24.295 164.670 ;
        RECT 23.265 164.630 24.225 164.640 ;
        RECT 23.265 164.620 24.200 164.630 ;
        RECT 23.265 164.605 24.180 164.620 ;
        RECT 23.265 164.590 24.160 164.605 ;
        RECT 23.370 164.580 24.155 164.590 ;
        RECT 23.370 164.545 24.140 164.580 ;
        RECT 22.925 163.715 23.200 164.415 ;
        RECT 23.370 164.295 24.125 164.545 ;
        RECT 24.295 164.225 24.625 164.470 ;
        RECT 24.795 164.370 25.055 164.820 ;
        RECT 24.440 164.200 24.625 164.225 ;
        RECT 25.260 164.335 25.575 165.355 ;
        RECT 25.745 164.685 25.915 165.185 ;
        RECT 26.165 164.855 26.430 165.415 ;
        RECT 26.600 164.685 26.770 165.585 ;
        RECT 28.815 165.525 29.145 165.865 ;
        RECT 30.195 165.695 30.525 166.095 ;
        RECT 26.940 164.855 27.295 165.415 ;
        RECT 28.160 165.355 30.525 165.525 ;
        RECT 30.695 165.370 31.025 165.880 ;
        RECT 25.745 164.515 27.170 164.685 ;
        RECT 24.440 164.100 25.055 164.200 ;
        RECT 23.370 163.545 23.625 164.090 ;
        RECT 23.795 163.715 24.275 164.055 ;
        RECT 24.450 163.545 25.055 164.100 ;
        RECT 25.260 163.715 25.795 164.335 ;
        RECT 25.965 163.545 26.295 164.345 ;
        RECT 26.780 164.340 27.170 164.515 ;
        RECT 28.160 164.355 28.330 165.355 ;
        RECT 30.355 165.185 30.525 165.355 ;
        RECT 28.500 164.525 28.745 165.185 ;
        RECT 28.960 164.525 29.225 165.185 ;
        RECT 29.420 164.525 29.705 165.185 ;
        RECT 29.880 164.855 30.185 165.185 ;
        RECT 30.355 164.855 30.665 165.185 ;
        RECT 29.880 164.525 30.095 164.855 ;
        RECT 28.160 164.185 28.615 164.355 ;
        RECT 28.285 163.755 28.615 164.185 ;
        RECT 28.795 164.185 30.085 164.355 ;
        RECT 28.795 163.765 29.045 164.185 ;
        RECT 29.275 163.545 29.605 164.015 ;
        RECT 29.835 163.765 30.085 164.185 ;
        RECT 30.275 163.545 30.525 164.685 ;
        RECT 30.835 164.605 31.025 165.370 ;
        RECT 31.265 165.275 31.475 166.095 ;
        RECT 31.645 165.295 31.975 165.925 ;
        RECT 31.645 164.695 31.895 165.295 ;
        RECT 32.145 165.275 32.375 166.095 ;
        RECT 32.585 165.325 36.095 166.095 ;
        RECT 36.760 165.355 37.375 165.925 ;
        RECT 37.545 165.585 37.760 166.095 ;
        RECT 37.990 165.585 38.270 165.915 ;
        RECT 38.450 165.585 38.690 166.095 ;
        RECT 32.065 164.855 32.395 165.105 ;
        RECT 32.585 164.805 34.235 165.325 ;
        RECT 30.695 163.755 31.025 164.605 ;
        RECT 31.265 163.545 31.475 164.685 ;
        RECT 31.645 163.715 31.975 164.695 ;
        RECT 32.145 163.545 32.375 164.685 ;
        RECT 34.405 164.635 36.095 165.155 ;
        RECT 32.585 163.545 36.095 164.635 ;
        RECT 36.760 164.335 37.075 165.355 ;
        RECT 37.245 164.685 37.415 165.185 ;
        RECT 37.665 164.855 37.930 165.415 ;
        RECT 38.100 164.685 38.270 165.585 ;
        RECT 38.440 164.855 38.795 165.415 ;
        RECT 39.085 165.275 39.295 166.095 ;
        RECT 39.465 165.295 39.795 165.925 ;
        RECT 39.465 164.695 39.715 165.295 ;
        RECT 39.965 165.275 40.195 166.095 ;
        RECT 40.405 165.345 41.615 166.095 ;
        RECT 39.885 164.855 40.215 165.105 ;
        RECT 40.405 164.805 40.925 165.345 ;
        RECT 41.795 165.285 42.065 166.095 ;
        RECT 42.235 165.285 42.565 165.925 ;
        RECT 42.735 165.285 42.975 166.095 ;
        RECT 43.165 165.370 43.455 166.095 ;
        RECT 43.625 165.595 43.885 165.925 ;
        RECT 44.055 165.735 44.385 166.095 ;
        RECT 44.640 165.715 45.940 165.925 ;
        RECT 43.625 165.585 43.855 165.595 ;
        RECT 37.245 164.515 38.670 164.685 ;
        RECT 36.760 163.715 37.295 164.335 ;
        RECT 37.465 163.545 37.795 164.345 ;
        RECT 38.280 164.340 38.670 164.515 ;
        RECT 39.085 163.545 39.295 164.685 ;
        RECT 39.465 163.715 39.795 164.695 ;
        RECT 39.965 163.545 40.195 164.685 ;
        RECT 41.095 164.635 41.615 165.175 ;
        RECT 41.785 164.855 42.135 165.105 ;
        RECT 42.305 164.685 42.475 165.285 ;
        RECT 42.645 164.855 42.995 165.105 ;
        RECT 40.405 163.545 41.615 164.635 ;
        RECT 41.795 163.545 42.125 164.685 ;
        RECT 42.305 164.515 42.985 164.685 ;
        RECT 42.655 163.730 42.985 164.515 ;
        RECT 43.165 163.545 43.455 164.710 ;
        RECT 43.625 164.395 43.795 165.585 ;
        RECT 44.640 165.565 44.810 165.715 ;
        RECT 44.055 165.440 44.810 165.565 ;
        RECT 43.965 165.395 44.810 165.440 ;
        RECT 43.965 165.275 44.235 165.395 ;
        RECT 43.965 164.700 44.135 165.275 ;
        RECT 44.365 164.835 44.775 165.140 ;
        RECT 45.065 165.105 45.275 165.505 ;
        RECT 44.945 164.895 45.275 165.105 ;
        RECT 45.520 165.105 45.740 165.505 ;
        RECT 46.215 165.330 46.670 166.095 ;
        RECT 46.845 165.295 47.540 165.925 ;
        RECT 47.745 165.295 48.055 166.095 ;
        RECT 48.735 165.440 49.065 165.875 ;
        RECT 49.235 165.485 49.405 166.095 ;
        RECT 48.685 165.355 49.065 165.440 ;
        RECT 49.575 165.355 49.905 165.880 ;
        RECT 50.165 165.565 50.375 166.095 ;
        RECT 50.650 165.645 51.435 165.815 ;
        RECT 51.605 165.645 52.010 165.815 ;
        RECT 48.685 165.315 48.910 165.355 ;
        RECT 45.520 164.895 45.995 165.105 ;
        RECT 46.185 164.905 46.675 165.105 ;
        RECT 46.865 164.855 47.200 165.105 ;
        RECT 43.965 164.665 44.165 164.700 ;
        RECT 45.495 164.665 46.670 164.725 ;
        RECT 47.370 164.695 47.540 165.295 ;
        RECT 47.710 164.855 48.045 165.125 ;
        RECT 48.685 164.735 48.855 165.315 ;
        RECT 49.575 165.185 49.775 165.355 ;
        RECT 50.650 165.185 50.820 165.645 ;
        RECT 49.025 164.855 49.775 165.185 ;
        RECT 49.945 164.855 50.820 165.185 ;
        RECT 43.965 164.555 46.670 164.665 ;
        RECT 44.025 164.495 45.825 164.555 ;
        RECT 45.495 164.465 45.825 164.495 ;
        RECT 43.625 163.715 43.885 164.395 ;
        RECT 44.055 163.545 44.305 164.325 ;
        RECT 44.555 164.295 45.390 164.305 ;
        RECT 45.980 164.295 46.165 164.385 ;
        RECT 44.555 164.095 46.165 164.295 ;
        RECT 44.555 163.715 44.805 164.095 ;
        RECT 45.935 164.055 46.165 164.095 ;
        RECT 46.415 163.935 46.670 164.555 ;
        RECT 44.975 163.545 45.330 163.925 ;
        RECT 46.335 163.715 46.670 163.935 ;
        RECT 46.845 163.545 47.105 164.685 ;
        RECT 47.275 163.715 47.605 164.695 ;
        RECT 48.685 164.685 48.900 164.735 ;
        RECT 47.775 163.545 48.055 164.685 ;
        RECT 48.685 164.605 49.075 164.685 ;
        RECT 48.745 163.760 49.075 164.605 ;
        RECT 49.585 164.650 49.775 164.855 ;
        RECT 49.245 163.545 49.415 164.555 ;
        RECT 49.585 164.275 50.480 164.650 ;
        RECT 49.585 163.715 49.925 164.275 ;
        RECT 50.155 163.545 50.470 164.045 ;
        RECT 50.650 164.015 50.820 164.855 ;
        RECT 50.990 165.145 51.455 165.475 ;
        RECT 51.840 165.415 52.010 165.645 ;
        RECT 52.190 165.595 52.560 166.095 ;
        RECT 52.880 165.645 53.555 165.815 ;
        RECT 53.750 165.645 54.085 165.815 ;
        RECT 50.990 164.185 51.310 165.145 ;
        RECT 51.840 165.115 52.670 165.415 ;
        RECT 51.480 164.215 51.670 164.935 ;
        RECT 51.840 164.045 52.010 165.115 ;
        RECT 52.470 165.085 52.670 165.115 ;
        RECT 52.180 164.865 52.350 164.935 ;
        RECT 52.880 164.865 53.050 165.645 ;
        RECT 53.915 165.505 54.085 165.645 ;
        RECT 54.255 165.635 54.505 166.095 ;
        RECT 52.180 164.695 53.050 164.865 ;
        RECT 53.220 165.225 53.745 165.445 ;
        RECT 53.915 165.375 54.140 165.505 ;
        RECT 52.180 164.605 52.690 164.695 ;
        RECT 50.650 163.845 51.535 164.015 ;
        RECT 51.760 163.715 52.010 164.045 ;
        RECT 52.180 163.545 52.350 164.345 ;
        RECT 52.520 163.990 52.690 164.605 ;
        RECT 53.220 164.525 53.390 165.225 ;
        RECT 52.860 164.160 53.390 164.525 ;
        RECT 53.560 164.460 53.800 165.055 ;
        RECT 53.970 164.270 54.140 165.375 ;
        RECT 54.310 164.515 54.590 165.465 ;
        RECT 53.835 164.140 54.140 164.270 ;
        RECT 52.520 163.820 53.625 163.990 ;
        RECT 53.835 163.715 54.085 164.140 ;
        RECT 54.255 163.545 54.520 164.005 ;
        RECT 54.760 163.715 54.945 165.835 ;
        RECT 55.115 165.715 55.445 166.095 ;
        RECT 55.615 165.545 55.785 165.835 ;
        RECT 56.045 165.550 61.390 166.095 ;
        RECT 55.120 165.375 55.785 165.545 ;
        RECT 55.120 164.385 55.350 165.375 ;
        RECT 55.520 164.555 55.870 165.205 ;
        RECT 57.630 164.720 57.970 165.550 ;
        RECT 61.655 165.545 61.825 165.835 ;
        RECT 61.995 165.715 62.325 166.095 ;
        RECT 61.655 165.375 62.320 165.545 ;
        RECT 55.120 164.215 55.785 164.385 ;
        RECT 55.115 163.545 55.445 164.045 ;
        RECT 55.615 163.715 55.785 164.215 ;
        RECT 59.450 163.980 59.800 165.230 ;
        RECT 61.570 164.555 61.920 165.205 ;
        RECT 62.090 164.385 62.320 165.375 ;
        RECT 61.655 164.215 62.320 164.385 ;
        RECT 56.045 163.545 61.390 163.980 ;
        RECT 61.655 163.715 61.825 164.215 ;
        RECT 61.995 163.545 62.325 164.045 ;
        RECT 62.495 163.715 62.680 165.835 ;
        RECT 62.935 165.635 63.185 166.095 ;
        RECT 63.355 165.645 63.690 165.815 ;
        RECT 63.885 165.645 64.560 165.815 ;
        RECT 63.355 165.505 63.525 165.645 ;
        RECT 62.850 164.515 63.130 165.465 ;
        RECT 63.300 165.375 63.525 165.505 ;
        RECT 63.300 164.270 63.470 165.375 ;
        RECT 63.695 165.225 64.220 165.445 ;
        RECT 63.640 164.460 63.880 165.055 ;
        RECT 64.050 164.525 64.220 165.225 ;
        RECT 64.390 164.865 64.560 165.645 ;
        RECT 64.880 165.595 65.250 166.095 ;
        RECT 65.430 165.645 65.835 165.815 ;
        RECT 66.005 165.645 66.790 165.815 ;
        RECT 65.430 165.415 65.600 165.645 ;
        RECT 64.770 165.115 65.600 165.415 ;
        RECT 65.985 165.145 66.450 165.475 ;
        RECT 64.770 165.085 64.970 165.115 ;
        RECT 65.090 164.865 65.260 164.935 ;
        RECT 64.390 164.695 65.260 164.865 ;
        RECT 64.750 164.605 65.260 164.695 ;
        RECT 63.300 164.140 63.605 164.270 ;
        RECT 64.050 164.160 64.580 164.525 ;
        RECT 62.920 163.545 63.185 164.005 ;
        RECT 63.355 163.715 63.605 164.140 ;
        RECT 64.750 163.990 64.920 164.605 ;
        RECT 63.815 163.820 64.920 163.990 ;
        RECT 65.090 163.545 65.260 164.345 ;
        RECT 65.430 164.045 65.600 165.115 ;
        RECT 65.770 164.215 65.960 164.935 ;
        RECT 66.130 164.185 66.450 165.145 ;
        RECT 66.620 165.185 66.790 165.645 ;
        RECT 67.065 165.565 67.275 166.095 ;
        RECT 67.535 165.355 67.865 165.880 ;
        RECT 68.035 165.485 68.205 166.095 ;
        RECT 68.375 165.440 68.705 165.875 ;
        RECT 68.375 165.355 68.755 165.440 ;
        RECT 68.925 165.370 69.215 166.095 ;
        RECT 69.385 165.550 74.730 166.095 ;
        RECT 67.665 165.185 67.865 165.355 ;
        RECT 68.530 165.315 68.755 165.355 ;
        RECT 66.620 164.855 67.495 165.185 ;
        RECT 67.665 164.855 68.415 165.185 ;
        RECT 65.430 163.715 65.680 164.045 ;
        RECT 66.620 164.015 66.790 164.855 ;
        RECT 67.665 164.650 67.855 164.855 ;
        RECT 68.585 164.735 68.755 165.315 ;
        RECT 68.540 164.685 68.755 164.735 ;
        RECT 70.970 164.720 71.310 165.550 ;
        RECT 74.905 165.325 76.575 166.095 ;
        RECT 76.795 165.440 77.125 165.875 ;
        RECT 77.295 165.485 77.465 166.095 ;
        RECT 76.745 165.355 77.125 165.440 ;
        RECT 77.635 165.355 77.965 165.880 ;
        RECT 78.225 165.565 78.435 166.095 ;
        RECT 78.710 165.645 79.495 165.815 ;
        RECT 79.665 165.645 80.070 165.815 ;
        RECT 66.960 164.275 67.855 164.650 ;
        RECT 68.365 164.605 68.755 164.685 ;
        RECT 65.905 163.845 66.790 164.015 ;
        RECT 66.970 163.545 67.285 164.045 ;
        RECT 67.515 163.715 67.855 164.275 ;
        RECT 68.025 163.545 68.195 164.555 ;
        RECT 68.365 163.760 68.695 164.605 ;
        RECT 68.925 163.545 69.215 164.710 ;
        RECT 72.790 163.980 73.140 165.230 ;
        RECT 74.905 164.805 75.655 165.325 ;
        RECT 76.745 165.315 76.970 165.355 ;
        RECT 75.825 164.635 76.575 165.155 ;
        RECT 69.385 163.545 74.730 163.980 ;
        RECT 74.905 163.545 76.575 164.635 ;
        RECT 76.745 164.735 76.915 165.315 ;
        RECT 77.635 165.185 77.835 165.355 ;
        RECT 78.710 165.185 78.880 165.645 ;
        RECT 77.085 164.855 77.835 165.185 ;
        RECT 78.005 164.855 78.880 165.185 ;
        RECT 76.745 164.685 76.960 164.735 ;
        RECT 76.745 164.605 77.135 164.685 ;
        RECT 76.805 163.760 77.135 164.605 ;
        RECT 77.645 164.650 77.835 164.855 ;
        RECT 77.305 163.545 77.475 164.555 ;
        RECT 77.645 164.275 78.540 164.650 ;
        RECT 77.645 163.715 77.985 164.275 ;
        RECT 78.215 163.545 78.530 164.045 ;
        RECT 78.710 164.015 78.880 164.855 ;
        RECT 79.050 165.145 79.515 165.475 ;
        RECT 79.900 165.415 80.070 165.645 ;
        RECT 80.250 165.595 80.620 166.095 ;
        RECT 80.940 165.645 81.615 165.815 ;
        RECT 81.810 165.645 82.145 165.815 ;
        RECT 79.050 164.185 79.370 165.145 ;
        RECT 79.900 165.115 80.730 165.415 ;
        RECT 79.540 164.215 79.730 164.935 ;
        RECT 79.900 164.045 80.070 165.115 ;
        RECT 80.530 165.085 80.730 165.115 ;
        RECT 80.240 164.865 80.410 164.935 ;
        RECT 80.940 164.865 81.110 165.645 ;
        RECT 81.975 165.505 82.145 165.645 ;
        RECT 82.315 165.635 82.565 166.095 ;
        RECT 80.240 164.695 81.110 164.865 ;
        RECT 81.280 165.225 81.805 165.445 ;
        RECT 81.975 165.375 82.200 165.505 ;
        RECT 80.240 164.605 80.750 164.695 ;
        RECT 78.710 163.845 79.595 164.015 ;
        RECT 79.820 163.715 80.070 164.045 ;
        RECT 80.240 163.545 80.410 164.345 ;
        RECT 80.580 163.990 80.750 164.605 ;
        RECT 81.280 164.525 81.450 165.225 ;
        RECT 80.920 164.160 81.450 164.525 ;
        RECT 81.620 164.460 81.860 165.055 ;
        RECT 82.030 164.270 82.200 165.375 ;
        RECT 82.370 164.515 82.650 165.465 ;
        RECT 81.895 164.140 82.200 164.270 ;
        RECT 80.580 163.820 81.685 163.990 ;
        RECT 81.895 163.715 82.145 164.140 ;
        RECT 82.315 163.545 82.580 164.005 ;
        RECT 82.820 163.715 83.005 165.835 ;
        RECT 83.175 165.715 83.505 166.095 ;
        RECT 83.675 165.545 83.845 165.835 ;
        RECT 83.180 165.375 83.845 165.545 ;
        RECT 83.180 164.385 83.410 165.375 ;
        RECT 84.105 165.370 84.365 165.925 ;
        RECT 84.535 165.650 84.965 166.095 ;
        RECT 85.200 165.525 85.370 165.925 ;
        RECT 85.540 165.695 86.260 166.095 ;
        RECT 83.580 164.555 83.930 165.205 ;
        RECT 84.105 164.655 84.280 165.370 ;
        RECT 85.200 165.355 86.080 165.525 ;
        RECT 86.430 165.480 86.600 165.925 ;
        RECT 87.175 165.585 87.575 166.095 ;
        RECT 87.805 165.585 88.045 166.095 ;
        RECT 84.450 164.855 84.705 165.185 ;
        RECT 83.180 164.215 83.845 164.385 ;
        RECT 83.175 163.545 83.505 164.045 ;
        RECT 83.675 163.715 83.845 164.215 ;
        RECT 84.105 163.715 84.365 164.655 ;
        RECT 84.535 164.375 84.705 164.855 ;
        RECT 84.930 164.565 85.260 165.185 ;
        RECT 85.430 164.805 85.720 165.185 ;
        RECT 85.910 164.635 86.080 165.355 ;
        RECT 85.560 164.465 86.080 164.635 ;
        RECT 86.250 165.310 86.600 165.480 ;
        RECT 84.535 164.205 85.295 164.375 ;
        RECT 85.560 164.275 85.730 164.465 ;
        RECT 86.250 164.285 86.420 165.310 ;
        RECT 86.840 164.825 87.100 165.415 ;
        RECT 86.620 164.525 87.100 164.825 ;
        RECT 87.300 164.525 87.560 165.415 ;
        RECT 87.790 164.855 88.045 165.415 ;
        RECT 88.215 165.355 88.545 165.890 ;
        RECT 88.760 165.355 88.930 166.095 ;
        RECT 89.140 165.445 89.470 165.915 ;
        RECT 89.640 165.615 89.810 166.095 ;
        RECT 89.980 165.445 90.310 165.915 ;
        RECT 90.480 165.615 90.650 166.095 ;
        RECT 88.215 164.685 88.395 165.355 ;
        RECT 89.140 165.275 90.835 165.445 ;
        RECT 88.565 164.855 88.940 165.185 ;
        RECT 89.110 164.935 90.320 165.105 ;
        RECT 89.110 164.685 89.315 164.935 ;
        RECT 90.490 164.685 90.835 165.275 ;
        RECT 91.005 165.325 94.515 166.095 ;
        RECT 94.685 165.370 94.975 166.095 ;
        RECT 95.145 165.325 98.655 166.095 ;
        RECT 91.005 164.805 92.655 165.325 ;
        RECT 87.855 164.515 89.315 164.685 ;
        RECT 89.980 164.515 90.835 164.685 ;
        RECT 92.825 164.635 94.515 165.155 ;
        RECT 95.145 164.805 96.795 165.325 ;
        RECT 98.825 165.295 99.135 166.095 ;
        RECT 99.340 165.295 100.035 165.925 ;
        RECT 100.255 165.440 100.585 165.875 ;
        RECT 100.755 165.485 100.925 166.095 ;
        RECT 100.205 165.355 100.585 165.440 ;
        RECT 101.095 165.355 101.425 165.880 ;
        RECT 101.685 165.565 101.895 166.095 ;
        RECT 102.170 165.645 102.955 165.815 ;
        RECT 103.125 165.645 103.530 165.815 ;
        RECT 100.205 165.315 100.430 165.355 ;
        RECT 85.125 163.980 85.295 164.205 ;
        RECT 86.010 164.115 86.420 164.285 ;
        RECT 86.595 164.175 87.535 164.345 ;
        RECT 86.010 163.980 86.265 164.115 ;
        RECT 84.535 163.545 84.865 163.945 ;
        RECT 85.125 163.810 86.265 163.980 ;
        RECT 86.595 163.925 86.765 164.175 ;
        RECT 86.010 163.715 86.265 163.810 ;
        RECT 86.435 163.755 86.765 163.925 ;
        RECT 86.935 163.545 87.185 164.005 ;
        RECT 87.355 163.715 87.535 164.175 ;
        RECT 87.855 163.715 88.215 164.515 ;
        RECT 89.980 164.345 90.310 164.515 ;
        RECT 88.760 163.545 88.930 164.345 ;
        RECT 89.140 164.175 90.310 164.345 ;
        RECT 89.140 163.715 89.470 164.175 ;
        RECT 89.640 163.545 89.810 164.005 ;
        RECT 89.980 163.715 90.310 164.175 ;
        RECT 90.480 163.545 90.650 164.345 ;
        RECT 91.005 163.545 94.515 164.635 ;
        RECT 94.685 163.545 94.975 164.710 ;
        RECT 96.965 164.635 98.655 165.155 ;
        RECT 98.835 164.855 99.170 165.125 ;
        RECT 99.340 164.695 99.510 165.295 ;
        RECT 99.680 164.855 100.015 165.105 ;
        RECT 100.205 164.735 100.375 165.315 ;
        RECT 101.095 165.185 101.295 165.355 ;
        RECT 102.170 165.185 102.340 165.645 ;
        RECT 100.545 164.855 101.295 165.185 ;
        RECT 101.465 164.855 102.340 165.185 ;
        RECT 95.145 163.545 98.655 164.635 ;
        RECT 98.825 163.545 99.105 164.685 ;
        RECT 99.275 163.715 99.605 164.695 ;
        RECT 100.205 164.685 100.420 164.735 ;
        RECT 99.775 163.545 100.035 164.685 ;
        RECT 100.205 164.605 100.595 164.685 ;
        RECT 100.265 163.760 100.595 164.605 ;
        RECT 101.105 164.650 101.295 164.855 ;
        RECT 100.765 163.545 100.935 164.555 ;
        RECT 101.105 164.275 102.000 164.650 ;
        RECT 101.105 163.715 101.445 164.275 ;
        RECT 101.675 163.545 101.990 164.045 ;
        RECT 102.170 164.015 102.340 164.855 ;
        RECT 102.510 165.145 102.975 165.475 ;
        RECT 103.360 165.415 103.530 165.645 ;
        RECT 103.710 165.595 104.080 166.095 ;
        RECT 104.400 165.645 105.075 165.815 ;
        RECT 105.270 165.645 105.605 165.815 ;
        RECT 102.510 164.185 102.830 165.145 ;
        RECT 103.360 165.115 104.190 165.415 ;
        RECT 103.000 164.215 103.190 164.935 ;
        RECT 103.360 164.045 103.530 165.115 ;
        RECT 103.990 165.085 104.190 165.115 ;
        RECT 103.700 164.865 103.870 164.935 ;
        RECT 104.400 164.865 104.570 165.645 ;
        RECT 105.435 165.505 105.605 165.645 ;
        RECT 105.775 165.635 106.025 166.095 ;
        RECT 103.700 164.695 104.570 164.865 ;
        RECT 104.740 165.225 105.265 165.445 ;
        RECT 105.435 165.375 105.660 165.505 ;
        RECT 103.700 164.605 104.210 164.695 ;
        RECT 102.170 163.845 103.055 164.015 ;
        RECT 103.280 163.715 103.530 164.045 ;
        RECT 103.700 163.545 103.870 164.345 ;
        RECT 104.040 163.990 104.210 164.605 ;
        RECT 104.740 164.525 104.910 165.225 ;
        RECT 104.380 164.160 104.910 164.525 ;
        RECT 105.080 164.460 105.320 165.055 ;
        RECT 105.490 164.270 105.660 165.375 ;
        RECT 105.830 164.515 106.110 165.465 ;
        RECT 105.355 164.140 105.660 164.270 ;
        RECT 104.040 163.820 105.145 163.990 ;
        RECT 105.355 163.715 105.605 164.140 ;
        RECT 105.775 163.545 106.040 164.005 ;
        RECT 106.280 163.715 106.465 165.835 ;
        RECT 106.635 165.715 106.965 166.095 ;
        RECT 107.135 165.545 107.305 165.835 ;
        RECT 106.640 165.375 107.305 165.545 ;
        RECT 106.640 164.385 106.870 165.375 ;
        RECT 107.565 165.355 107.950 165.925 ;
        RECT 108.120 165.635 108.445 166.095 ;
        RECT 108.965 165.465 109.245 165.925 ;
        RECT 107.040 164.555 107.390 165.205 ;
        RECT 107.565 164.685 107.845 165.355 ;
        RECT 108.120 165.295 109.245 165.465 ;
        RECT 108.120 165.185 108.570 165.295 ;
        RECT 108.015 164.855 108.570 165.185 ;
        RECT 109.435 165.125 109.835 165.925 ;
        RECT 110.235 165.635 110.505 166.095 ;
        RECT 110.675 165.465 110.960 165.925 ;
        RECT 106.640 164.215 107.305 164.385 ;
        RECT 106.635 163.545 106.965 164.045 ;
        RECT 107.135 163.715 107.305 164.215 ;
        RECT 107.565 163.715 107.950 164.685 ;
        RECT 108.120 164.395 108.570 164.855 ;
        RECT 108.740 164.565 109.835 165.125 ;
        RECT 108.120 164.175 109.245 164.395 ;
        RECT 108.120 163.545 108.445 164.005 ;
        RECT 108.965 163.715 109.245 164.175 ;
        RECT 109.435 163.715 109.835 164.565 ;
        RECT 110.005 165.295 110.960 165.465 ;
        RECT 110.005 164.395 110.215 165.295 ;
        RECT 110.385 164.565 111.075 165.125 ;
        RECT 111.265 164.515 111.495 165.855 ;
        RECT 111.675 165.015 111.905 165.915 ;
        RECT 112.105 165.315 112.350 166.095 ;
        RECT 112.520 165.555 112.950 165.915 ;
        RECT 113.530 165.725 114.260 166.095 ;
        RECT 112.520 165.365 114.260 165.555 ;
        RECT 112.520 165.135 112.740 165.365 ;
        RECT 110.005 164.175 110.960 164.395 ;
        RECT 111.675 164.335 112.015 165.015 ;
        RECT 110.235 163.545 110.505 164.005 ;
        RECT 110.675 163.715 110.960 164.175 ;
        RECT 111.265 164.135 112.015 164.335 ;
        RECT 112.195 164.835 112.740 165.135 ;
        RECT 111.265 163.745 111.505 164.135 ;
        RECT 111.675 163.545 112.025 163.955 ;
        RECT 112.195 163.725 112.525 164.835 ;
        RECT 112.910 164.565 113.335 165.185 ;
        RECT 113.530 164.565 113.790 165.185 ;
        RECT 114.000 164.855 114.260 165.365 ;
        RECT 112.695 164.195 113.720 164.395 ;
        RECT 112.695 163.725 112.875 164.195 ;
        RECT 113.045 163.545 113.375 164.025 ;
        RECT 113.550 163.725 113.720 164.195 ;
        RECT 113.985 163.545 114.270 164.685 ;
        RECT 114.460 163.725 114.740 165.915 ;
        RECT 114.925 165.595 115.265 166.095 ;
        RECT 114.925 164.855 115.265 165.425 ;
        RECT 115.435 165.185 115.680 165.875 ;
        RECT 115.875 165.595 116.205 166.095 ;
        RECT 116.405 165.525 116.575 165.875 ;
        RECT 116.750 165.695 117.080 166.095 ;
        RECT 117.250 165.525 117.420 165.875 ;
        RECT 117.590 165.695 117.970 166.095 ;
        RECT 116.405 165.355 117.990 165.525 ;
        RECT 118.160 165.420 118.435 165.765 ;
        RECT 117.820 165.185 117.990 165.355 ;
        RECT 115.435 164.855 116.090 165.185 ;
        RECT 114.925 163.545 115.265 164.620 ;
        RECT 115.435 164.260 115.675 164.855 ;
        RECT 115.870 164.395 116.190 164.685 ;
        RECT 116.360 164.565 117.100 165.185 ;
        RECT 117.270 164.855 117.650 165.185 ;
        RECT 117.820 164.855 118.095 165.185 ;
        RECT 117.820 164.685 117.990 164.855 ;
        RECT 118.265 164.685 118.435 165.420 ;
        RECT 118.605 165.325 120.275 166.095 ;
        RECT 120.445 165.370 120.735 166.095 ;
        RECT 120.905 165.445 121.165 165.925 ;
        RECT 121.335 165.555 121.585 166.095 ;
        RECT 118.605 164.805 119.355 165.325 ;
        RECT 117.330 164.515 117.990 164.685 ;
        RECT 117.330 164.395 117.500 164.515 ;
        RECT 115.870 164.225 117.500 164.395 ;
        RECT 115.445 163.885 117.500 164.055 ;
        RECT 115.450 163.765 117.500 163.885 ;
        RECT 117.670 163.545 117.950 164.345 ;
        RECT 118.160 163.715 118.435 164.685 ;
        RECT 119.525 164.635 120.275 165.155 ;
        RECT 118.605 163.545 120.275 164.635 ;
        RECT 120.445 163.545 120.735 164.710 ;
        RECT 120.905 164.415 121.075 165.445 ;
        RECT 121.755 165.390 121.975 165.875 ;
        RECT 121.245 164.795 121.475 165.190 ;
        RECT 121.645 164.965 121.975 165.390 ;
        RECT 122.145 165.715 123.035 165.885 ;
        RECT 122.145 164.990 122.315 165.715 ;
        RECT 123.265 165.635 123.510 166.095 ;
        RECT 122.485 165.160 123.035 165.545 ;
        RECT 122.145 164.920 123.035 164.990 ;
        RECT 122.140 164.895 123.035 164.920 ;
        RECT 122.130 164.880 123.035 164.895 ;
        RECT 122.125 164.865 123.035 164.880 ;
        RECT 122.115 164.860 123.035 164.865 ;
        RECT 122.110 164.850 123.035 164.860 ;
        RECT 123.205 164.855 123.520 165.465 ;
        RECT 123.690 165.105 123.940 165.915 ;
        RECT 124.110 165.570 124.370 166.095 ;
        RECT 124.540 165.445 124.800 165.900 ;
        RECT 124.970 165.615 125.230 166.095 ;
        RECT 125.400 165.445 125.660 165.900 ;
        RECT 125.830 165.615 126.090 166.095 ;
        RECT 126.260 165.445 126.520 165.900 ;
        RECT 126.690 165.615 126.950 166.095 ;
        RECT 127.120 165.445 127.380 165.900 ;
        RECT 127.550 165.615 127.850 166.095 ;
        RECT 129.345 165.535 129.675 165.925 ;
        RECT 129.845 165.705 131.030 165.875 ;
        RECT 131.290 165.625 131.460 166.095 ;
        RECT 124.540 165.275 127.850 165.445 ;
        RECT 129.345 165.355 129.855 165.535 ;
        RECT 123.690 164.855 126.710 165.105 ;
        RECT 122.105 164.840 123.035 164.850 ;
        RECT 122.095 164.835 123.035 164.840 ;
        RECT 122.085 164.825 123.035 164.835 ;
        RECT 122.075 164.820 123.035 164.825 ;
        RECT 122.075 164.815 122.410 164.820 ;
        RECT 122.060 164.810 122.410 164.815 ;
        RECT 122.045 164.800 122.410 164.810 ;
        RECT 122.020 164.795 122.410 164.800 ;
        RECT 121.245 164.790 122.410 164.795 ;
        RECT 121.245 164.755 122.380 164.790 ;
        RECT 121.245 164.730 122.345 164.755 ;
        RECT 121.245 164.700 122.315 164.730 ;
        RECT 121.245 164.670 122.295 164.700 ;
        RECT 121.245 164.640 122.275 164.670 ;
        RECT 121.245 164.630 122.205 164.640 ;
        RECT 121.245 164.620 122.180 164.630 ;
        RECT 121.245 164.605 122.160 164.620 ;
        RECT 121.245 164.590 122.140 164.605 ;
        RECT 121.350 164.580 122.135 164.590 ;
        RECT 121.350 164.545 122.120 164.580 ;
        RECT 120.905 163.715 121.180 164.415 ;
        RECT 121.350 164.295 122.105 164.545 ;
        RECT 122.275 164.225 122.605 164.470 ;
        RECT 122.775 164.370 123.035 164.820 ;
        RECT 122.420 164.200 122.605 164.225 ;
        RECT 122.420 164.100 123.035 164.200 ;
        RECT 121.350 163.545 121.605 164.090 ;
        RECT 121.775 163.715 122.255 164.055 ;
        RECT 122.430 163.545 123.035 164.100 ;
        RECT 123.215 163.545 123.510 164.655 ;
        RECT 123.690 163.720 123.940 164.855 ;
        RECT 126.880 164.685 127.850 165.275 ;
        RECT 129.185 164.895 129.515 165.185 ;
        RECT 129.685 164.725 129.855 165.355 ;
        RECT 130.260 165.445 130.645 165.535 ;
        RECT 131.630 165.445 131.960 165.910 ;
        RECT 130.260 165.275 131.960 165.445 ;
        RECT 132.130 165.275 132.300 166.095 ;
        RECT 132.470 165.275 133.155 165.915 ;
        RECT 130.025 164.895 130.355 165.105 ;
        RECT 130.535 164.855 130.915 165.105 ;
        RECT 131.105 165.075 131.590 165.105 ;
        RECT 131.085 164.905 131.590 165.075 ;
        RECT 124.110 163.545 124.370 164.655 ;
        RECT 124.540 164.445 127.850 164.685 ;
        RECT 129.340 164.555 130.425 164.725 ;
        RECT 124.540 163.720 124.800 164.445 ;
        RECT 124.970 163.545 125.230 164.275 ;
        RECT 125.400 163.720 125.660 164.445 ;
        RECT 125.830 163.545 126.090 164.275 ;
        RECT 126.260 163.720 126.520 164.445 ;
        RECT 126.690 163.545 126.950 164.275 ;
        RECT 127.120 163.720 127.380 164.445 ;
        RECT 127.550 163.545 127.845 164.275 ;
        RECT 129.340 163.715 129.640 164.555 ;
        RECT 129.835 163.545 130.085 164.385 ;
        RECT 130.255 164.305 130.425 164.555 ;
        RECT 130.595 164.475 130.915 164.855 ;
        RECT 131.105 164.895 131.590 164.905 ;
        RECT 131.780 164.895 132.230 165.105 ;
        RECT 132.400 164.895 132.735 165.105 ;
        RECT 131.105 164.475 131.480 164.895 ;
        RECT 132.400 164.725 132.570 164.895 ;
        RECT 131.650 164.555 132.570 164.725 ;
        RECT 131.650 164.305 131.820 164.555 ;
        RECT 130.255 164.135 131.820 164.305 ;
        RECT 130.675 163.715 131.480 164.135 ;
        RECT 131.990 163.545 132.320 164.385 ;
        RECT 132.905 164.305 133.155 165.275 ;
        RECT 132.490 163.715 133.155 164.305 ;
        RECT 133.820 165.355 134.435 165.925 ;
        RECT 134.605 165.585 134.820 166.095 ;
        RECT 135.050 165.585 135.330 165.915 ;
        RECT 135.510 165.585 135.750 166.095 ;
        RECT 133.820 164.335 134.135 165.355 ;
        RECT 134.305 164.685 134.475 165.185 ;
        RECT 134.725 164.855 134.990 165.415 ;
        RECT 135.160 164.685 135.330 165.585 ;
        RECT 136.635 165.545 136.805 165.835 ;
        RECT 136.975 165.715 137.305 166.095 ;
        RECT 135.500 164.855 135.855 165.415 ;
        RECT 136.635 165.375 137.300 165.545 ;
        RECT 134.305 164.515 135.730 164.685 ;
        RECT 136.550 164.555 136.900 165.205 ;
        RECT 133.820 163.715 134.355 164.335 ;
        RECT 134.525 163.545 134.855 164.345 ;
        RECT 135.340 164.340 135.730 164.515 ;
        RECT 137.070 164.385 137.300 165.375 ;
        RECT 136.635 164.215 137.300 164.385 ;
        RECT 136.635 163.715 136.805 164.215 ;
        RECT 136.975 163.545 137.305 164.045 ;
        RECT 137.475 163.715 137.660 165.835 ;
        RECT 137.915 165.635 138.165 166.095 ;
        RECT 138.335 165.645 138.670 165.815 ;
        RECT 138.865 165.645 139.540 165.815 ;
        RECT 138.335 165.505 138.505 165.645 ;
        RECT 137.830 164.515 138.110 165.465 ;
        RECT 138.280 165.375 138.505 165.505 ;
        RECT 138.280 164.270 138.450 165.375 ;
        RECT 138.675 165.225 139.200 165.445 ;
        RECT 138.620 164.460 138.860 165.055 ;
        RECT 139.030 164.525 139.200 165.225 ;
        RECT 139.370 164.865 139.540 165.645 ;
        RECT 139.860 165.595 140.230 166.095 ;
        RECT 140.410 165.645 140.815 165.815 ;
        RECT 140.985 165.645 141.770 165.815 ;
        RECT 140.410 165.415 140.580 165.645 ;
        RECT 139.750 165.115 140.580 165.415 ;
        RECT 140.965 165.145 141.430 165.475 ;
        RECT 139.750 165.085 139.950 165.115 ;
        RECT 140.070 164.865 140.240 164.935 ;
        RECT 139.370 164.695 140.240 164.865 ;
        RECT 139.730 164.605 140.240 164.695 ;
        RECT 138.280 164.140 138.585 164.270 ;
        RECT 139.030 164.160 139.560 164.525 ;
        RECT 137.900 163.545 138.165 164.005 ;
        RECT 138.335 163.715 138.585 164.140 ;
        RECT 139.730 163.990 139.900 164.605 ;
        RECT 138.795 163.820 139.900 163.990 ;
        RECT 140.070 163.545 140.240 164.345 ;
        RECT 140.410 164.045 140.580 165.115 ;
        RECT 140.750 164.215 140.940 164.935 ;
        RECT 141.110 164.185 141.430 165.145 ;
        RECT 141.600 165.185 141.770 165.645 ;
        RECT 142.045 165.565 142.255 166.095 ;
        RECT 142.515 165.355 142.845 165.880 ;
        RECT 143.015 165.485 143.185 166.095 ;
        RECT 143.355 165.440 143.685 165.875 ;
        RECT 143.995 165.545 144.165 165.925 ;
        RECT 144.380 165.715 144.710 166.095 ;
        RECT 143.355 165.355 143.735 165.440 ;
        RECT 143.995 165.375 144.710 165.545 ;
        RECT 142.645 165.185 142.845 165.355 ;
        RECT 143.510 165.315 143.735 165.355 ;
        RECT 141.600 164.855 142.475 165.185 ;
        RECT 142.645 164.855 143.395 165.185 ;
        RECT 140.410 163.715 140.660 164.045 ;
        RECT 141.600 164.015 141.770 164.855 ;
        RECT 142.645 164.650 142.835 164.855 ;
        RECT 143.565 164.735 143.735 165.315 ;
        RECT 143.905 164.825 144.260 165.195 ;
        RECT 144.540 165.185 144.710 165.375 ;
        RECT 144.880 165.350 145.135 165.925 ;
        RECT 144.540 164.855 144.795 165.185 ;
        RECT 143.520 164.685 143.735 164.735 ;
        RECT 141.940 164.275 142.835 164.650 ;
        RECT 143.345 164.605 143.735 164.685 ;
        RECT 144.540 164.645 144.710 164.855 ;
        RECT 140.885 163.845 141.770 164.015 ;
        RECT 141.950 163.545 142.265 164.045 ;
        RECT 142.495 163.715 142.835 164.275 ;
        RECT 143.005 163.545 143.175 164.555 ;
        RECT 143.345 163.760 143.675 164.605 ;
        RECT 143.995 164.475 144.710 164.645 ;
        RECT 144.965 164.620 145.135 165.350 ;
        RECT 145.310 165.255 145.570 166.095 ;
        RECT 145.745 165.345 146.955 166.095 ;
        RECT 143.995 163.715 144.165 164.475 ;
        RECT 144.380 163.545 144.710 164.305 ;
        RECT 144.880 163.715 145.135 164.620 ;
        RECT 145.310 163.545 145.570 164.695 ;
        RECT 145.745 164.635 146.265 165.175 ;
        RECT 146.435 164.805 146.955 165.345 ;
        RECT 145.745 163.545 146.955 164.635 ;
        RECT 17.320 163.375 147.040 163.545 ;
        RECT 17.405 162.285 18.615 163.375 ;
        RECT 19.335 162.705 19.505 163.205 ;
        RECT 19.675 162.875 20.005 163.375 ;
        RECT 19.335 162.535 20.000 162.705 ;
        RECT 17.405 161.575 17.925 162.115 ;
        RECT 18.095 161.745 18.615 162.285 ;
        RECT 19.250 161.715 19.600 162.365 ;
        RECT 17.405 160.825 18.615 161.575 ;
        RECT 19.770 161.545 20.000 162.535 ;
        RECT 19.335 161.375 20.000 161.545 ;
        RECT 19.335 161.085 19.505 161.375 ;
        RECT 19.675 160.825 20.005 161.205 ;
        RECT 20.175 161.085 20.360 163.205 ;
        RECT 20.600 162.915 20.865 163.375 ;
        RECT 21.035 162.780 21.285 163.205 ;
        RECT 21.495 162.930 22.600 163.100 ;
        RECT 20.980 162.650 21.285 162.780 ;
        RECT 20.530 161.455 20.810 162.405 ;
        RECT 20.980 161.545 21.150 162.650 ;
        RECT 21.320 161.865 21.560 162.460 ;
        RECT 21.730 162.395 22.260 162.760 ;
        RECT 21.730 161.695 21.900 162.395 ;
        RECT 22.430 162.315 22.600 162.930 ;
        RECT 22.770 162.575 22.940 163.375 ;
        RECT 23.110 162.875 23.360 163.205 ;
        RECT 23.585 162.905 24.470 163.075 ;
        RECT 22.430 162.225 22.940 162.315 ;
        RECT 20.980 161.415 21.205 161.545 ;
        RECT 21.375 161.475 21.900 161.695 ;
        RECT 22.070 162.055 22.940 162.225 ;
        RECT 20.615 160.825 20.865 161.285 ;
        RECT 21.035 161.275 21.205 161.415 ;
        RECT 22.070 161.275 22.240 162.055 ;
        RECT 22.770 161.985 22.940 162.055 ;
        RECT 22.450 161.805 22.650 161.835 ;
        RECT 23.110 161.805 23.280 162.875 ;
        RECT 23.450 161.985 23.640 162.705 ;
        RECT 22.450 161.505 23.280 161.805 ;
        RECT 23.810 161.775 24.130 162.735 ;
        RECT 21.035 161.105 21.370 161.275 ;
        RECT 21.565 161.105 22.240 161.275 ;
        RECT 22.560 160.825 22.930 161.325 ;
        RECT 23.110 161.275 23.280 161.505 ;
        RECT 23.665 161.445 24.130 161.775 ;
        RECT 24.300 162.065 24.470 162.905 ;
        RECT 24.650 162.875 24.965 163.375 ;
        RECT 25.195 162.645 25.535 163.205 ;
        RECT 24.640 162.270 25.535 162.645 ;
        RECT 25.705 162.365 25.875 163.375 ;
        RECT 25.345 162.065 25.535 162.270 ;
        RECT 26.045 162.315 26.375 163.160 ;
        RECT 26.045 162.235 26.435 162.315 ;
        RECT 26.605 162.235 26.865 163.375 ;
        RECT 26.220 162.185 26.435 162.235 ;
        RECT 27.035 162.225 27.365 163.205 ;
        RECT 27.535 162.235 27.815 163.375 ;
        RECT 27.985 162.820 28.590 163.375 ;
        RECT 28.765 162.865 29.245 163.205 ;
        RECT 29.415 162.830 29.670 163.375 ;
        RECT 27.985 162.720 28.600 162.820 ;
        RECT 28.415 162.695 28.600 162.720 ;
        RECT 24.300 161.735 25.175 162.065 ;
        RECT 25.345 161.735 26.095 162.065 ;
        RECT 24.300 161.275 24.470 161.735 ;
        RECT 25.345 161.565 25.545 161.735 ;
        RECT 26.265 161.605 26.435 162.185 ;
        RECT 26.625 161.815 26.960 162.065 ;
        RECT 27.130 161.625 27.300 162.225 ;
        RECT 27.985 162.100 28.245 162.550 ;
        RECT 28.415 162.450 28.745 162.695 ;
        RECT 28.915 162.375 29.670 162.625 ;
        RECT 29.840 162.505 30.115 163.205 ;
        RECT 28.900 162.340 29.670 162.375 ;
        RECT 28.885 162.330 29.670 162.340 ;
        RECT 28.880 162.315 29.775 162.330 ;
        RECT 28.860 162.300 29.775 162.315 ;
        RECT 28.840 162.290 29.775 162.300 ;
        RECT 28.815 162.280 29.775 162.290 ;
        RECT 28.745 162.250 29.775 162.280 ;
        RECT 28.725 162.220 29.775 162.250 ;
        RECT 28.705 162.190 29.775 162.220 ;
        RECT 28.675 162.165 29.775 162.190 ;
        RECT 28.640 162.130 29.775 162.165 ;
        RECT 28.610 162.125 29.775 162.130 ;
        RECT 28.610 162.120 29.000 162.125 ;
        RECT 28.610 162.110 28.975 162.120 ;
        RECT 28.610 162.105 28.960 162.110 ;
        RECT 28.610 162.100 28.945 162.105 ;
        RECT 27.985 162.095 28.945 162.100 ;
        RECT 27.985 162.085 28.935 162.095 ;
        RECT 27.985 162.080 28.925 162.085 ;
        RECT 27.985 162.070 28.915 162.080 ;
        RECT 27.470 161.795 27.805 162.065 ;
        RECT 27.985 162.060 28.910 162.070 ;
        RECT 27.985 162.055 28.905 162.060 ;
        RECT 27.985 162.040 28.895 162.055 ;
        RECT 27.985 162.025 28.890 162.040 ;
        RECT 27.985 162.000 28.880 162.025 ;
        RECT 27.985 161.930 28.875 162.000 ;
        RECT 26.210 161.565 26.435 161.605 ;
        RECT 23.110 161.105 23.515 161.275 ;
        RECT 23.685 161.105 24.470 161.275 ;
        RECT 24.745 160.825 24.955 161.355 ;
        RECT 25.215 161.040 25.545 161.565 ;
        RECT 26.055 161.480 26.435 161.565 ;
        RECT 25.715 160.825 25.885 161.435 ;
        RECT 26.055 161.045 26.385 161.480 ;
        RECT 26.605 160.995 27.300 161.625 ;
        RECT 27.505 160.825 27.815 161.625 ;
        RECT 27.985 161.375 28.535 161.760 ;
        RECT 28.705 161.205 28.875 161.930 ;
        RECT 27.985 161.035 28.875 161.205 ;
        RECT 29.045 161.530 29.375 161.955 ;
        RECT 29.545 161.730 29.775 162.125 ;
        RECT 29.045 161.045 29.265 161.530 ;
        RECT 29.945 161.475 30.115 162.505 ;
        RECT 30.285 162.210 30.575 163.375 ;
        RECT 30.835 162.705 31.005 163.205 ;
        RECT 31.175 162.875 31.505 163.375 ;
        RECT 30.835 162.535 31.500 162.705 ;
        RECT 30.750 161.715 31.100 162.365 ;
        RECT 29.435 160.825 29.685 161.365 ;
        RECT 29.855 160.995 30.115 161.475 ;
        RECT 30.285 160.825 30.575 161.550 ;
        RECT 31.270 161.545 31.500 162.535 ;
        RECT 30.835 161.375 31.500 161.545 ;
        RECT 30.835 161.085 31.005 161.375 ;
        RECT 31.175 160.825 31.505 161.205 ;
        RECT 31.675 161.085 31.860 163.205 ;
        RECT 32.100 162.915 32.365 163.375 ;
        RECT 32.535 162.780 32.785 163.205 ;
        RECT 32.995 162.930 34.100 163.100 ;
        RECT 32.480 162.650 32.785 162.780 ;
        RECT 32.030 161.455 32.310 162.405 ;
        RECT 32.480 161.545 32.650 162.650 ;
        RECT 32.820 161.865 33.060 162.460 ;
        RECT 33.230 162.395 33.760 162.760 ;
        RECT 33.230 161.695 33.400 162.395 ;
        RECT 33.930 162.315 34.100 162.930 ;
        RECT 34.270 162.575 34.440 163.375 ;
        RECT 34.610 162.875 34.860 163.205 ;
        RECT 35.085 162.905 35.970 163.075 ;
        RECT 33.930 162.225 34.440 162.315 ;
        RECT 32.480 161.415 32.705 161.545 ;
        RECT 32.875 161.475 33.400 161.695 ;
        RECT 33.570 162.055 34.440 162.225 ;
        RECT 32.115 160.825 32.365 161.285 ;
        RECT 32.535 161.275 32.705 161.415 ;
        RECT 33.570 161.275 33.740 162.055 ;
        RECT 34.270 161.985 34.440 162.055 ;
        RECT 33.950 161.805 34.150 161.835 ;
        RECT 34.610 161.805 34.780 162.875 ;
        RECT 34.950 161.985 35.140 162.705 ;
        RECT 33.950 161.505 34.780 161.805 ;
        RECT 35.310 161.775 35.630 162.735 ;
        RECT 32.535 161.105 32.870 161.275 ;
        RECT 33.065 161.105 33.740 161.275 ;
        RECT 34.060 160.825 34.430 161.325 ;
        RECT 34.610 161.275 34.780 161.505 ;
        RECT 35.165 161.445 35.630 161.775 ;
        RECT 35.800 162.065 35.970 162.905 ;
        RECT 36.150 162.875 36.465 163.375 ;
        RECT 36.695 162.645 37.035 163.205 ;
        RECT 36.140 162.270 37.035 162.645 ;
        RECT 37.205 162.365 37.375 163.375 ;
        RECT 36.845 162.065 37.035 162.270 ;
        RECT 37.545 162.315 37.875 163.160 ;
        RECT 38.305 162.705 38.585 163.375 ;
        RECT 38.755 162.485 39.055 163.035 ;
        RECT 39.255 162.655 39.585 163.375 ;
        RECT 39.775 162.655 40.235 163.205 ;
        RECT 40.410 162.950 40.745 163.375 ;
        RECT 40.915 162.770 41.100 163.175 ;
        RECT 37.545 162.235 37.935 162.315 ;
        RECT 37.720 162.185 37.935 162.235 ;
        RECT 35.800 161.735 36.675 162.065 ;
        RECT 36.845 161.735 37.595 162.065 ;
        RECT 35.800 161.275 35.970 161.735 ;
        RECT 36.845 161.565 37.045 161.735 ;
        RECT 37.765 161.605 37.935 162.185 ;
        RECT 38.120 162.065 38.385 162.425 ;
        RECT 38.755 162.315 39.695 162.485 ;
        RECT 39.525 162.065 39.695 162.315 ;
        RECT 38.120 161.815 38.795 162.065 ;
        RECT 39.015 161.815 39.355 162.065 ;
        RECT 39.525 161.735 39.815 162.065 ;
        RECT 39.525 161.645 39.695 161.735 ;
        RECT 37.710 161.565 37.935 161.605 ;
        RECT 34.610 161.105 35.015 161.275 ;
        RECT 35.185 161.105 35.970 161.275 ;
        RECT 36.245 160.825 36.455 161.355 ;
        RECT 36.715 161.040 37.045 161.565 ;
        RECT 37.555 161.480 37.935 161.565 ;
        RECT 37.215 160.825 37.385 161.435 ;
        RECT 37.555 161.045 37.885 161.480 ;
        RECT 38.305 161.455 39.695 161.645 ;
        RECT 38.305 161.095 38.635 161.455 ;
        RECT 39.985 161.285 40.235 162.655 ;
        RECT 40.435 162.595 41.100 162.770 ;
        RECT 41.305 162.595 41.635 163.375 ;
        RECT 40.435 161.565 40.775 162.595 ;
        RECT 41.805 162.405 42.075 163.175 ;
        RECT 40.945 162.235 42.075 162.405 ;
        RECT 42.430 162.405 42.820 162.580 ;
        RECT 43.305 162.575 43.635 163.375 ;
        RECT 43.805 162.585 44.340 163.205 ;
        RECT 44.545 162.820 45.150 163.375 ;
        RECT 45.325 162.865 45.805 163.205 ;
        RECT 45.975 162.830 46.230 163.375 ;
        RECT 44.545 162.720 45.160 162.820 ;
        RECT 42.430 162.235 43.855 162.405 ;
        RECT 40.945 161.735 41.195 162.235 ;
        RECT 40.435 161.395 41.120 161.565 ;
        RECT 41.375 161.485 41.735 162.065 ;
        RECT 39.255 160.825 39.505 161.285 ;
        RECT 39.675 160.995 40.235 161.285 ;
        RECT 40.410 160.825 40.745 161.225 ;
        RECT 40.915 160.995 41.120 161.395 ;
        RECT 41.905 161.325 42.075 162.235 ;
        RECT 42.305 161.505 42.660 162.065 ;
        RECT 42.830 161.335 43.000 162.235 ;
        RECT 43.170 161.505 43.435 162.065 ;
        RECT 43.685 161.735 43.855 162.235 ;
        RECT 44.025 161.565 44.340 162.585 ;
        RECT 44.975 162.695 45.160 162.720 ;
        RECT 44.545 162.100 44.805 162.550 ;
        RECT 44.975 162.450 45.305 162.695 ;
        RECT 45.475 162.375 46.230 162.625 ;
        RECT 46.400 162.505 46.675 163.205 ;
        RECT 46.845 162.865 47.145 163.375 ;
        RECT 47.315 162.695 47.645 163.205 ;
        RECT 47.815 162.865 48.445 163.375 ;
        RECT 49.025 162.865 49.405 163.035 ;
        RECT 49.575 162.865 49.875 163.375 ;
        RECT 49.235 162.695 49.405 162.865 ;
        RECT 50.265 162.705 50.545 163.375 ;
        RECT 45.460 162.340 46.230 162.375 ;
        RECT 45.445 162.330 46.230 162.340 ;
        RECT 45.440 162.315 46.335 162.330 ;
        RECT 45.420 162.300 46.335 162.315 ;
        RECT 45.400 162.290 46.335 162.300 ;
        RECT 45.375 162.280 46.335 162.290 ;
        RECT 45.305 162.250 46.335 162.280 ;
        RECT 45.285 162.220 46.335 162.250 ;
        RECT 45.265 162.190 46.335 162.220 ;
        RECT 45.235 162.165 46.335 162.190 ;
        RECT 45.200 162.130 46.335 162.165 ;
        RECT 45.170 162.125 46.335 162.130 ;
        RECT 45.170 162.120 45.560 162.125 ;
        RECT 45.170 162.110 45.535 162.120 ;
        RECT 45.170 162.105 45.520 162.110 ;
        RECT 45.170 162.100 45.505 162.105 ;
        RECT 44.545 162.095 45.505 162.100 ;
        RECT 44.545 162.085 45.495 162.095 ;
        RECT 44.545 162.080 45.485 162.085 ;
        RECT 44.545 162.070 45.475 162.080 ;
        RECT 44.545 162.060 45.470 162.070 ;
        RECT 44.545 162.055 45.465 162.060 ;
        RECT 44.545 162.040 45.455 162.055 ;
        RECT 44.545 162.025 45.450 162.040 ;
        RECT 44.545 162.000 45.440 162.025 ;
        RECT 44.545 161.930 45.435 162.000 ;
        RECT 41.330 160.825 41.605 161.305 ;
        RECT 41.815 160.995 42.075 161.325 ;
        RECT 42.410 160.825 42.650 161.335 ;
        RECT 42.830 161.005 43.110 161.335 ;
        RECT 43.340 160.825 43.555 161.335 ;
        RECT 43.725 160.995 44.340 161.565 ;
        RECT 44.545 161.375 45.095 161.760 ;
        RECT 45.265 161.205 45.435 161.930 ;
        RECT 44.545 161.035 45.435 161.205 ;
        RECT 45.605 161.530 45.935 161.955 ;
        RECT 46.105 161.730 46.335 162.125 ;
        RECT 45.605 161.045 45.825 161.530 ;
        RECT 46.505 161.475 46.675 162.505 ;
        RECT 45.995 160.825 46.245 161.365 ;
        RECT 46.415 160.995 46.675 161.475 ;
        RECT 46.845 162.525 49.065 162.695 ;
        RECT 46.845 161.565 47.015 162.525 ;
        RECT 47.185 162.185 48.725 162.355 ;
        RECT 47.185 161.735 47.430 162.185 ;
        RECT 47.690 161.815 48.385 162.015 ;
        RECT 48.555 161.985 48.725 162.185 ;
        RECT 48.895 162.325 49.065 162.525 ;
        RECT 49.235 162.495 49.895 162.695 ;
        RECT 48.895 162.155 49.555 162.325 ;
        RECT 48.555 161.815 49.155 161.985 ;
        RECT 49.385 161.735 49.555 162.155 ;
        RECT 46.845 161.020 47.310 161.565 ;
        RECT 47.815 160.825 47.985 161.645 ;
        RECT 48.155 161.565 49.065 161.645 ;
        RECT 49.725 161.565 49.895 162.495 ;
        RECT 50.715 162.485 51.015 163.035 ;
        RECT 51.215 162.655 51.545 163.375 ;
        RECT 51.735 162.655 52.195 163.205 ;
        RECT 50.080 162.065 50.345 162.425 ;
        RECT 50.715 162.315 51.655 162.485 ;
        RECT 51.485 162.065 51.655 162.315 ;
        RECT 50.080 161.815 50.755 162.065 ;
        RECT 50.975 161.815 51.315 162.065 ;
        RECT 51.485 161.735 51.775 162.065 ;
        RECT 51.485 161.645 51.655 161.735 ;
        RECT 48.155 161.475 49.405 161.565 ;
        RECT 48.155 160.995 48.485 161.475 ;
        RECT 48.895 161.395 49.405 161.475 ;
        RECT 48.655 160.825 49.005 161.215 ;
        RECT 49.175 160.995 49.405 161.395 ;
        RECT 49.575 161.085 49.895 161.565 ;
        RECT 50.265 161.455 51.655 161.645 ;
        RECT 50.265 161.095 50.595 161.455 ;
        RECT 51.945 161.285 52.195 162.655 ;
        RECT 52.365 162.285 55.875 163.375 ;
        RECT 51.215 160.825 51.465 161.285 ;
        RECT 51.635 160.995 52.195 161.285 ;
        RECT 52.365 161.595 54.015 162.115 ;
        RECT 54.185 161.765 55.875 162.285 ;
        RECT 56.045 162.210 56.335 163.375 ;
        RECT 56.505 162.940 61.850 163.375 ;
        RECT 62.025 162.940 67.370 163.375 ;
        RECT 67.545 162.940 72.890 163.375 ;
        RECT 73.065 162.940 78.410 163.375 ;
        RECT 52.365 160.825 55.875 161.595 ;
        RECT 56.045 160.825 56.335 161.550 ;
        RECT 58.090 161.370 58.430 162.200 ;
        RECT 59.910 161.690 60.260 162.940 ;
        RECT 63.610 161.370 63.950 162.200 ;
        RECT 65.430 161.690 65.780 162.940 ;
        RECT 69.130 161.370 69.470 162.200 ;
        RECT 70.950 161.690 71.300 162.940 ;
        RECT 74.650 161.370 74.990 162.200 ;
        RECT 76.470 161.690 76.820 162.940 ;
        RECT 78.585 162.285 81.175 163.375 ;
        RECT 78.585 161.595 79.795 162.115 ;
        RECT 79.965 161.765 81.175 162.285 ;
        RECT 81.805 162.210 82.095 163.375 ;
        RECT 82.725 162.085 82.995 163.185 ;
        RECT 83.165 162.445 83.440 162.950 ;
        RECT 83.610 162.615 83.940 163.375 ;
        RECT 83.165 162.275 83.655 162.445 ;
        RECT 84.110 162.365 84.435 163.205 ;
        RECT 82.725 161.735 83.175 162.085 ;
        RECT 83.360 161.735 83.655 162.275 ;
        RECT 83.825 162.195 84.435 162.365 ;
        RECT 84.910 162.275 85.285 163.375 ;
        RECT 85.485 162.865 85.745 163.375 ;
        RECT 56.505 160.825 61.850 161.370 ;
        RECT 62.025 160.825 67.370 161.370 ;
        RECT 67.545 160.825 72.890 161.370 ;
        RECT 73.065 160.825 78.410 161.370 ;
        RECT 78.585 160.825 81.175 161.595 ;
        RECT 83.360 161.565 83.530 161.735 ;
        RECT 83.825 161.565 83.995 162.195 ;
        RECT 84.165 161.815 84.665 162.025 ;
        RECT 84.835 161.815 85.315 162.025 ;
        RECT 85.485 161.815 85.825 162.695 ;
        RECT 85.995 161.985 86.165 163.205 ;
        RECT 86.405 162.870 87.020 163.375 ;
        RECT 86.405 162.335 86.655 162.700 ;
        RECT 86.825 162.695 87.020 162.870 ;
        RECT 87.190 162.865 87.665 163.205 ;
        RECT 87.835 162.830 88.050 163.375 ;
        RECT 86.825 162.505 87.155 162.695 ;
        RECT 87.375 162.335 88.090 162.630 ;
        RECT 88.260 162.505 88.535 163.205 ;
        RECT 86.405 162.165 88.195 162.335 ;
        RECT 85.995 161.735 86.790 161.985 ;
        RECT 85.995 161.645 86.245 161.735 ;
        RECT 81.805 160.825 82.095 161.550 ;
        RECT 82.725 160.825 83.000 161.565 ;
        RECT 83.220 161.395 83.530 161.565 ;
        RECT 83.220 161.235 83.410 161.395 ;
        RECT 83.755 161.385 83.995 161.565 ;
        RECT 84.210 161.475 85.305 161.645 ;
        RECT 83.755 160.995 83.925 161.385 ;
        RECT 84.210 161.225 84.380 161.475 ;
        RECT 84.130 160.995 84.460 161.225 ;
        RECT 84.635 160.825 84.805 161.295 ;
        RECT 84.975 161.010 85.305 161.475 ;
        RECT 85.485 160.825 85.745 161.645 ;
        RECT 85.915 161.225 86.245 161.645 ;
        RECT 86.960 161.310 87.215 162.165 ;
        RECT 86.425 161.045 87.215 161.310 ;
        RECT 87.385 161.465 87.795 161.985 ;
        RECT 87.965 161.735 88.195 162.165 ;
        RECT 88.365 161.475 88.535 162.505 ;
        RECT 88.705 162.235 88.965 163.375 ;
        RECT 89.135 162.225 89.465 163.205 ;
        RECT 89.635 162.235 89.915 163.375 ;
        RECT 90.635 162.705 90.805 163.205 ;
        RECT 90.975 162.875 91.305 163.375 ;
        RECT 90.635 162.535 91.300 162.705 ;
        RECT 88.725 161.815 89.060 162.065 ;
        RECT 89.230 161.625 89.400 162.225 ;
        RECT 89.570 161.795 89.905 162.065 ;
        RECT 90.550 161.715 90.900 162.365 ;
        RECT 87.385 161.045 87.585 161.465 ;
        RECT 87.775 160.825 88.105 161.285 ;
        RECT 88.275 160.995 88.535 161.475 ;
        RECT 88.705 160.995 89.400 161.625 ;
        RECT 89.605 160.825 89.915 161.625 ;
        RECT 91.070 161.545 91.300 162.535 ;
        RECT 90.635 161.375 91.300 161.545 ;
        RECT 90.635 161.085 90.805 161.375 ;
        RECT 90.975 160.825 91.305 161.205 ;
        RECT 91.475 161.085 91.660 163.205 ;
        RECT 91.900 162.915 92.165 163.375 ;
        RECT 92.335 162.780 92.585 163.205 ;
        RECT 92.795 162.930 93.900 163.100 ;
        RECT 92.280 162.650 92.585 162.780 ;
        RECT 91.830 161.455 92.110 162.405 ;
        RECT 92.280 161.545 92.450 162.650 ;
        RECT 92.620 161.865 92.860 162.460 ;
        RECT 93.030 162.395 93.560 162.760 ;
        RECT 93.030 161.695 93.200 162.395 ;
        RECT 93.730 162.315 93.900 162.930 ;
        RECT 94.070 162.575 94.240 163.375 ;
        RECT 94.410 162.875 94.660 163.205 ;
        RECT 94.885 162.905 95.770 163.075 ;
        RECT 93.730 162.225 94.240 162.315 ;
        RECT 92.280 161.415 92.505 161.545 ;
        RECT 92.675 161.475 93.200 161.695 ;
        RECT 93.370 162.055 94.240 162.225 ;
        RECT 91.915 160.825 92.165 161.285 ;
        RECT 92.335 161.275 92.505 161.415 ;
        RECT 93.370 161.275 93.540 162.055 ;
        RECT 94.070 161.985 94.240 162.055 ;
        RECT 93.750 161.805 93.950 161.835 ;
        RECT 94.410 161.805 94.580 162.875 ;
        RECT 94.750 161.985 94.940 162.705 ;
        RECT 93.750 161.505 94.580 161.805 ;
        RECT 95.110 161.775 95.430 162.735 ;
        RECT 92.335 161.105 92.670 161.275 ;
        RECT 92.865 161.105 93.540 161.275 ;
        RECT 93.860 160.825 94.230 161.325 ;
        RECT 94.410 161.275 94.580 161.505 ;
        RECT 94.965 161.445 95.430 161.775 ;
        RECT 95.600 162.065 95.770 162.905 ;
        RECT 95.950 162.875 96.265 163.375 ;
        RECT 96.495 162.645 96.835 163.205 ;
        RECT 95.940 162.270 96.835 162.645 ;
        RECT 97.005 162.365 97.175 163.375 ;
        RECT 96.645 162.065 96.835 162.270 ;
        RECT 97.345 162.315 97.675 163.160 ;
        RECT 98.155 162.645 98.450 163.375 ;
        RECT 98.620 162.475 98.880 163.200 ;
        RECT 99.050 162.645 99.310 163.375 ;
        RECT 99.480 162.475 99.740 163.200 ;
        RECT 99.910 162.645 100.170 163.375 ;
        RECT 100.340 162.475 100.600 163.200 ;
        RECT 100.770 162.645 101.030 163.375 ;
        RECT 101.200 162.475 101.460 163.200 ;
        RECT 97.345 162.235 97.735 162.315 ;
        RECT 97.520 162.185 97.735 162.235 ;
        RECT 95.600 161.735 96.475 162.065 ;
        RECT 96.645 161.735 97.395 162.065 ;
        RECT 95.600 161.275 95.770 161.735 ;
        RECT 96.645 161.565 96.845 161.735 ;
        RECT 97.565 161.605 97.735 162.185 ;
        RECT 97.510 161.565 97.735 161.605 ;
        RECT 94.410 161.105 94.815 161.275 ;
        RECT 94.985 161.105 95.770 161.275 ;
        RECT 96.045 160.825 96.255 161.355 ;
        RECT 96.515 161.040 96.845 161.565 ;
        RECT 97.355 161.480 97.735 161.565 ;
        RECT 98.150 162.235 101.460 162.475 ;
        RECT 101.630 162.265 101.890 163.375 ;
        RECT 98.150 161.645 99.120 162.235 ;
        RECT 102.060 162.065 102.310 163.200 ;
        RECT 102.490 162.265 102.785 163.375 ;
        RECT 102.965 162.235 103.350 163.205 ;
        RECT 103.520 162.915 103.845 163.375 ;
        RECT 104.365 162.745 104.645 163.205 ;
        RECT 103.520 162.525 104.645 162.745 ;
        RECT 99.290 161.815 102.310 162.065 ;
        RECT 97.015 160.825 97.185 161.435 ;
        RECT 97.355 161.045 97.685 161.480 ;
        RECT 98.150 161.475 101.460 161.645 ;
        RECT 98.150 160.825 98.450 161.305 ;
        RECT 98.620 161.020 98.880 161.475 ;
        RECT 99.050 160.825 99.310 161.305 ;
        RECT 99.480 161.020 99.740 161.475 ;
        RECT 99.910 160.825 100.170 161.305 ;
        RECT 100.340 161.020 100.600 161.475 ;
        RECT 100.770 160.825 101.030 161.305 ;
        RECT 101.200 161.020 101.460 161.475 ;
        RECT 101.630 160.825 101.890 161.350 ;
        RECT 102.060 161.005 102.310 161.815 ;
        RECT 102.480 161.455 102.795 162.065 ;
        RECT 102.965 161.565 103.245 162.235 ;
        RECT 103.520 162.065 103.970 162.525 ;
        RECT 104.835 162.355 105.235 163.205 ;
        RECT 105.635 162.915 105.905 163.375 ;
        RECT 106.075 162.745 106.360 163.205 ;
        RECT 103.415 161.735 103.970 162.065 ;
        RECT 104.140 161.795 105.235 162.355 ;
        RECT 103.520 161.625 103.970 161.735 ;
        RECT 102.490 160.825 102.735 161.285 ;
        RECT 102.965 160.995 103.350 161.565 ;
        RECT 103.520 161.455 104.645 161.625 ;
        RECT 103.520 160.825 103.845 161.285 ;
        RECT 104.365 160.995 104.645 161.455 ;
        RECT 104.835 160.995 105.235 161.795 ;
        RECT 105.405 162.525 106.360 162.745 ;
        RECT 105.405 161.625 105.615 162.525 ;
        RECT 105.785 161.795 106.475 162.355 ;
        RECT 107.565 162.210 107.855 163.375 ;
        RECT 108.070 162.235 108.365 163.375 ;
        RECT 108.625 162.405 108.955 163.205 ;
        RECT 109.125 162.575 109.295 163.375 ;
        RECT 109.465 162.405 109.795 163.205 ;
        RECT 109.965 162.575 110.135 163.375 ;
        RECT 110.305 162.425 110.635 163.205 ;
        RECT 110.805 162.915 110.975 163.375 ;
        RECT 111.245 162.865 111.505 163.375 ;
        RECT 110.305 162.405 111.075 162.425 ;
        RECT 108.625 162.235 111.075 162.405 ;
        RECT 108.045 161.815 110.555 162.065 ;
        RECT 110.725 161.645 111.075 162.235 ;
        RECT 111.245 161.815 111.585 162.695 ;
        RECT 111.755 161.985 111.925 163.205 ;
        RECT 112.165 162.870 112.780 163.375 ;
        RECT 112.165 162.335 112.415 162.700 ;
        RECT 112.585 162.695 112.780 162.870 ;
        RECT 112.950 162.865 113.425 163.205 ;
        RECT 113.595 162.830 113.810 163.375 ;
        RECT 112.585 162.505 112.915 162.695 ;
        RECT 113.135 162.335 113.850 162.630 ;
        RECT 114.020 162.505 114.295 163.205 ;
        RECT 114.505 163.035 115.645 163.205 ;
        RECT 114.505 162.575 114.805 163.035 ;
        RECT 112.165 162.165 113.955 162.335 ;
        RECT 111.755 161.735 112.550 161.985 ;
        RECT 111.755 161.645 112.005 161.735 ;
        RECT 105.405 161.455 106.360 161.625 ;
        RECT 105.635 160.825 105.905 161.285 ;
        RECT 106.075 160.995 106.360 161.455 ;
        RECT 107.565 160.825 107.855 161.550 ;
        RECT 108.705 161.465 111.075 161.645 ;
        RECT 108.070 160.825 108.335 161.285 ;
        RECT 108.705 160.995 108.875 161.465 ;
        RECT 109.125 160.825 109.295 161.285 ;
        RECT 109.545 160.995 109.715 161.465 ;
        RECT 109.965 160.825 110.135 161.285 ;
        RECT 110.385 160.995 110.555 161.465 ;
        RECT 110.725 160.825 110.975 161.290 ;
        RECT 111.245 160.825 111.505 161.645 ;
        RECT 111.675 161.225 112.005 161.645 ;
        RECT 112.720 161.310 112.975 162.165 ;
        RECT 112.185 161.045 112.975 161.310 ;
        RECT 113.145 161.465 113.555 161.985 ;
        RECT 113.725 161.735 113.955 162.165 ;
        RECT 114.125 161.475 114.295 162.505 ;
        RECT 114.975 162.405 115.305 162.865 ;
        RECT 114.545 162.355 115.305 162.405 ;
        RECT 114.525 162.185 115.305 162.355 ;
        RECT 115.475 162.405 115.645 163.035 ;
        RECT 115.815 162.575 116.145 163.375 ;
        RECT 116.315 162.405 116.590 163.205 ;
        RECT 115.475 162.195 116.590 162.405 ;
        RECT 114.545 161.645 114.760 162.185 ;
        RECT 114.930 161.815 115.700 162.015 ;
        RECT 115.870 161.815 116.590 162.015 ;
        RECT 114.545 161.475 116.145 161.645 ;
        RECT 113.145 161.045 113.345 161.465 ;
        RECT 113.535 160.825 113.865 161.285 ;
        RECT 114.035 160.995 114.295 161.475 ;
        RECT 114.975 161.465 116.145 161.475 ;
        RECT 114.515 160.825 114.805 161.295 ;
        RECT 114.975 160.995 115.305 161.465 ;
        RECT 115.475 160.825 115.645 161.295 ;
        RECT 115.815 160.995 116.145 161.465 ;
        RECT 116.315 160.825 116.590 161.645 ;
        RECT 117.695 161.005 117.955 163.195 ;
        RECT 118.125 162.645 118.465 163.375 ;
        RECT 118.645 162.465 118.915 163.195 ;
        RECT 118.145 162.245 118.915 162.465 ;
        RECT 119.095 162.485 119.325 163.195 ;
        RECT 119.495 162.665 119.825 163.375 ;
        RECT 119.995 162.485 120.255 163.195 ;
        RECT 119.095 162.245 120.255 162.485 ;
        RECT 118.145 161.575 118.435 162.245 ;
        RECT 118.615 161.755 119.080 162.065 ;
        RECT 119.260 161.755 119.785 162.065 ;
        RECT 118.145 161.375 119.375 161.575 ;
        RECT 118.215 160.825 118.885 161.195 ;
        RECT 119.065 161.005 119.375 161.375 ;
        RECT 119.555 161.115 119.785 161.755 ;
        RECT 119.965 161.735 120.265 162.065 ;
        RECT 119.965 160.825 120.255 161.555 ;
        RECT 120.915 161.005 121.175 163.195 ;
        RECT 121.345 162.645 121.685 163.375 ;
        RECT 121.865 162.465 122.135 163.195 ;
        RECT 121.365 162.245 122.135 162.465 ;
        RECT 122.315 162.485 122.545 163.195 ;
        RECT 122.715 162.665 123.045 163.375 ;
        RECT 123.215 162.485 123.475 163.195 ;
        RECT 122.315 162.245 123.475 162.485 ;
        RECT 121.365 161.575 121.655 162.245 ;
        RECT 123.795 162.205 124.125 163.375 ;
        RECT 121.835 161.755 122.300 162.065 ;
        RECT 122.480 161.755 123.005 162.065 ;
        RECT 121.365 161.375 122.595 161.575 ;
        RECT 121.435 160.825 122.105 161.195 ;
        RECT 122.285 161.005 122.595 161.375 ;
        RECT 122.775 161.115 123.005 161.755 ;
        RECT 123.185 161.735 123.485 162.065 ;
        RECT 124.325 162.035 124.655 163.205 ;
        RECT 124.855 162.205 125.185 163.375 ;
        RECT 125.385 162.035 125.745 163.205 ;
        RECT 125.915 162.235 126.245 163.375 ;
        RECT 126.580 162.365 126.880 163.205 ;
        RECT 127.075 162.535 127.325 163.375 ;
        RECT 127.915 162.785 128.720 163.205 ;
        RECT 127.495 162.615 129.060 162.785 ;
        RECT 127.495 162.365 127.665 162.615 ;
        RECT 126.580 162.195 127.665 162.365 ;
        RECT 124.325 161.755 125.745 162.035 ;
        RECT 123.185 160.825 123.475 161.555 ;
        RECT 124.335 160.825 124.665 161.515 ;
        RECT 125.385 161.420 125.745 161.755 ;
        RECT 125.915 161.485 126.255 162.065 ;
        RECT 126.425 161.735 126.755 162.025 ;
        RECT 126.925 161.565 127.095 162.195 ;
        RECT 127.835 162.065 128.155 162.445 ;
        RECT 128.345 162.355 128.720 162.445 ;
        RECT 128.325 162.185 128.720 162.355 ;
        RECT 128.890 162.365 129.060 162.615 ;
        RECT 129.230 162.535 129.560 163.375 ;
        RECT 129.730 162.615 130.395 163.205 ;
        RECT 128.890 162.195 129.810 162.365 ;
        RECT 127.265 161.815 127.595 162.025 ;
        RECT 127.775 161.815 128.155 162.065 ;
        RECT 128.345 162.025 128.720 162.185 ;
        RECT 129.640 162.025 129.810 162.195 ;
        RECT 128.345 161.815 128.830 162.025 ;
        RECT 129.020 161.815 129.470 162.025 ;
        RECT 129.640 161.815 129.975 162.025 ;
        RECT 130.145 161.645 130.395 162.615 ;
        RECT 125.125 160.995 125.745 161.420 ;
        RECT 126.585 161.385 127.095 161.565 ;
        RECT 127.500 161.475 129.200 161.645 ;
        RECT 127.500 161.385 127.885 161.475 ;
        RECT 125.915 160.825 126.245 161.315 ;
        RECT 126.585 160.995 126.915 161.385 ;
        RECT 127.085 161.045 128.270 161.215 ;
        RECT 128.530 160.825 128.700 161.295 ;
        RECT 128.870 161.010 129.200 161.475 ;
        RECT 129.370 160.825 129.540 161.645 ;
        RECT 129.710 161.005 130.395 161.645 ;
        RECT 130.600 162.585 131.135 163.205 ;
        RECT 130.600 161.565 130.915 162.585 ;
        RECT 131.305 162.575 131.635 163.375 ;
        RECT 132.120 162.405 132.510 162.580 ;
        RECT 131.085 162.235 132.510 162.405 ;
        RECT 131.085 161.735 131.255 162.235 ;
        RECT 130.600 160.995 131.215 161.565 ;
        RECT 131.505 161.505 131.770 162.065 ;
        RECT 131.940 161.335 132.110 162.235 ;
        RECT 133.325 162.210 133.615 163.375 ;
        RECT 133.785 162.865 134.975 163.155 ;
        RECT 133.805 162.525 134.975 162.695 ;
        RECT 135.145 162.575 135.425 163.375 ;
        RECT 133.805 162.235 134.130 162.525 ;
        RECT 134.805 162.405 134.975 162.525 ;
        RECT 134.300 162.065 134.495 162.355 ;
        RECT 134.805 162.235 135.465 162.405 ;
        RECT 135.635 162.235 135.910 163.205 ;
        RECT 136.085 162.285 137.295 163.375 ;
        RECT 135.295 162.065 135.465 162.235 ;
        RECT 132.280 161.505 132.635 162.065 ;
        RECT 133.785 161.735 134.130 162.065 ;
        RECT 134.300 161.735 135.125 162.065 ;
        RECT 135.295 161.735 135.570 162.065 ;
        RECT 135.295 161.565 135.465 161.735 ;
        RECT 131.385 160.825 131.600 161.335 ;
        RECT 131.830 161.005 132.110 161.335 ;
        RECT 132.290 160.825 132.530 161.335 ;
        RECT 133.325 160.825 133.615 161.550 ;
        RECT 133.800 161.395 135.465 161.565 ;
        RECT 135.740 161.500 135.910 162.235 ;
        RECT 133.800 161.045 134.055 161.395 ;
        RECT 134.225 160.825 134.555 161.225 ;
        RECT 134.725 161.045 134.895 161.395 ;
        RECT 135.065 160.825 135.445 161.225 ;
        RECT 135.635 161.155 135.910 161.500 ;
        RECT 136.085 161.575 136.605 162.115 ;
        RECT 136.775 161.745 137.295 162.285 ;
        RECT 137.470 162.235 137.805 163.205 ;
        RECT 137.975 162.235 138.145 163.375 ;
        RECT 138.315 163.035 140.345 163.205 ;
        RECT 136.085 160.825 137.295 161.575 ;
        RECT 137.470 161.565 137.640 162.235 ;
        RECT 138.315 162.065 138.485 163.035 ;
        RECT 137.810 161.735 138.065 162.065 ;
        RECT 138.290 161.735 138.485 162.065 ;
        RECT 138.655 162.695 139.780 162.865 ;
        RECT 137.895 161.565 138.065 161.735 ;
        RECT 138.655 161.565 138.825 162.695 ;
        RECT 137.470 160.995 137.725 161.565 ;
        RECT 137.895 161.395 138.825 161.565 ;
        RECT 138.995 162.355 140.005 162.525 ;
        RECT 138.995 161.555 139.165 162.355 ;
        RECT 139.370 161.675 139.645 162.155 ;
        RECT 139.365 161.505 139.645 161.675 ;
        RECT 138.650 161.360 138.825 161.395 ;
        RECT 137.895 160.825 138.225 161.225 ;
        RECT 138.650 160.995 139.180 161.360 ;
        RECT 139.370 160.995 139.645 161.505 ;
        RECT 139.815 160.995 140.005 162.355 ;
        RECT 140.175 162.370 140.345 163.035 ;
        RECT 140.515 162.615 140.685 163.375 ;
        RECT 140.920 162.615 141.435 163.025 ;
        RECT 140.175 162.180 140.925 162.370 ;
        RECT 141.095 161.805 141.435 162.615 ;
        RECT 140.205 161.635 141.435 161.805 ;
        RECT 141.605 162.235 141.990 163.205 ;
        RECT 142.160 162.915 142.485 163.375 ;
        RECT 143.005 162.745 143.285 163.205 ;
        RECT 142.160 162.525 143.285 162.745 ;
        RECT 140.185 160.825 140.695 161.360 ;
        RECT 140.915 161.030 141.160 161.635 ;
        RECT 141.605 161.565 141.885 162.235 ;
        RECT 142.160 162.065 142.610 162.525 ;
        RECT 143.475 162.355 143.875 163.205 ;
        RECT 144.275 162.915 144.545 163.375 ;
        RECT 144.715 162.745 145.000 163.205 ;
        RECT 142.055 161.735 142.610 162.065 ;
        RECT 142.780 161.795 143.875 162.355 ;
        RECT 142.160 161.625 142.610 161.735 ;
        RECT 141.605 160.995 141.990 161.565 ;
        RECT 142.160 161.455 143.285 161.625 ;
        RECT 142.160 160.825 142.485 161.285 ;
        RECT 143.005 160.995 143.285 161.455 ;
        RECT 143.475 160.995 143.875 161.795 ;
        RECT 144.045 162.525 145.000 162.745 ;
        RECT 144.045 161.625 144.255 162.525 ;
        RECT 144.425 161.795 145.115 162.355 ;
        RECT 145.745 162.285 146.955 163.375 ;
        RECT 145.745 161.745 146.265 162.285 ;
        RECT 144.045 161.455 145.000 161.625 ;
        RECT 146.435 161.575 146.955 162.115 ;
        RECT 144.275 160.825 144.545 161.285 ;
        RECT 144.715 160.995 145.000 161.455 ;
        RECT 145.745 160.825 146.955 161.575 ;
        RECT 17.320 160.655 147.040 160.825 ;
        RECT 17.405 159.905 18.615 160.655 ;
        RECT 18.785 159.905 19.995 160.655 ;
        RECT 20.165 160.005 20.425 160.485 ;
        RECT 20.595 160.115 20.845 160.655 ;
        RECT 17.405 159.365 17.925 159.905 ;
        RECT 18.095 159.195 18.615 159.735 ;
        RECT 18.785 159.365 19.305 159.905 ;
        RECT 19.475 159.195 19.995 159.735 ;
        RECT 17.405 158.105 18.615 159.195 ;
        RECT 18.785 158.105 19.995 159.195 ;
        RECT 20.165 158.975 20.335 160.005 ;
        RECT 21.015 159.950 21.235 160.435 ;
        RECT 20.505 159.355 20.735 159.750 ;
        RECT 20.905 159.525 21.235 159.950 ;
        RECT 21.405 160.275 22.295 160.445 ;
        RECT 21.405 159.550 21.575 160.275 ;
        RECT 22.555 160.105 22.725 160.395 ;
        RECT 22.895 160.275 23.225 160.655 ;
        RECT 21.745 159.720 22.295 160.105 ;
        RECT 22.555 159.935 23.220 160.105 ;
        RECT 21.405 159.480 22.295 159.550 ;
        RECT 21.400 159.455 22.295 159.480 ;
        RECT 21.390 159.440 22.295 159.455 ;
        RECT 21.385 159.425 22.295 159.440 ;
        RECT 21.375 159.420 22.295 159.425 ;
        RECT 21.370 159.410 22.295 159.420 ;
        RECT 21.365 159.400 22.295 159.410 ;
        RECT 21.355 159.395 22.295 159.400 ;
        RECT 21.345 159.385 22.295 159.395 ;
        RECT 21.335 159.380 22.295 159.385 ;
        RECT 21.335 159.375 21.670 159.380 ;
        RECT 21.320 159.370 21.670 159.375 ;
        RECT 21.305 159.360 21.670 159.370 ;
        RECT 21.280 159.355 21.670 159.360 ;
        RECT 20.505 159.350 21.670 159.355 ;
        RECT 20.505 159.315 21.640 159.350 ;
        RECT 20.505 159.290 21.605 159.315 ;
        RECT 20.505 159.260 21.575 159.290 ;
        RECT 20.505 159.230 21.555 159.260 ;
        RECT 20.505 159.200 21.535 159.230 ;
        RECT 20.505 159.190 21.465 159.200 ;
        RECT 20.505 159.180 21.440 159.190 ;
        RECT 20.505 159.165 21.420 159.180 ;
        RECT 20.505 159.150 21.400 159.165 ;
        RECT 20.610 159.140 21.395 159.150 ;
        RECT 20.610 159.105 21.380 159.140 ;
        RECT 20.165 158.275 20.440 158.975 ;
        RECT 20.610 158.855 21.365 159.105 ;
        RECT 21.535 158.785 21.865 159.030 ;
        RECT 22.035 158.930 22.295 159.380 ;
        RECT 22.470 159.115 22.820 159.765 ;
        RECT 22.990 158.945 23.220 159.935 ;
        RECT 21.680 158.760 21.865 158.785 ;
        RECT 22.555 158.775 23.220 158.945 ;
        RECT 21.680 158.660 22.295 158.760 ;
        RECT 20.610 158.105 20.865 158.650 ;
        RECT 21.035 158.275 21.515 158.615 ;
        RECT 21.690 158.105 22.295 158.660 ;
        RECT 22.555 158.275 22.725 158.775 ;
        RECT 22.895 158.105 23.225 158.605 ;
        RECT 23.395 158.275 23.580 160.395 ;
        RECT 23.835 160.195 24.085 160.655 ;
        RECT 24.255 160.205 24.590 160.375 ;
        RECT 24.785 160.205 25.460 160.375 ;
        RECT 24.255 160.065 24.425 160.205 ;
        RECT 23.750 159.075 24.030 160.025 ;
        RECT 24.200 159.935 24.425 160.065 ;
        RECT 24.200 158.830 24.370 159.935 ;
        RECT 24.595 159.785 25.120 160.005 ;
        RECT 24.540 159.020 24.780 159.615 ;
        RECT 24.950 159.085 25.120 159.785 ;
        RECT 25.290 159.425 25.460 160.205 ;
        RECT 25.780 160.155 26.150 160.655 ;
        RECT 26.330 160.205 26.735 160.375 ;
        RECT 26.905 160.205 27.690 160.375 ;
        RECT 26.330 159.975 26.500 160.205 ;
        RECT 25.670 159.675 26.500 159.975 ;
        RECT 26.885 159.705 27.350 160.035 ;
        RECT 25.670 159.645 25.870 159.675 ;
        RECT 25.990 159.425 26.160 159.495 ;
        RECT 25.290 159.255 26.160 159.425 ;
        RECT 25.650 159.165 26.160 159.255 ;
        RECT 24.200 158.700 24.505 158.830 ;
        RECT 24.950 158.720 25.480 159.085 ;
        RECT 23.820 158.105 24.085 158.565 ;
        RECT 24.255 158.275 24.505 158.700 ;
        RECT 25.650 158.550 25.820 159.165 ;
        RECT 24.715 158.380 25.820 158.550 ;
        RECT 25.990 158.105 26.160 158.905 ;
        RECT 26.330 158.605 26.500 159.675 ;
        RECT 26.670 158.775 26.860 159.495 ;
        RECT 27.030 158.745 27.350 159.705 ;
        RECT 27.520 159.745 27.690 160.205 ;
        RECT 27.965 160.125 28.175 160.655 ;
        RECT 28.435 159.915 28.765 160.440 ;
        RECT 28.935 160.045 29.105 160.655 ;
        RECT 29.275 160.000 29.605 160.435 ;
        RECT 29.825 160.275 30.715 160.445 ;
        RECT 29.275 159.915 29.655 160.000 ;
        RECT 28.565 159.745 28.765 159.915 ;
        RECT 29.430 159.875 29.655 159.915 ;
        RECT 27.520 159.415 28.395 159.745 ;
        RECT 28.565 159.415 29.315 159.745 ;
        RECT 26.330 158.275 26.580 158.605 ;
        RECT 27.520 158.575 27.690 159.415 ;
        RECT 28.565 159.210 28.755 159.415 ;
        RECT 29.485 159.295 29.655 159.875 ;
        RECT 29.825 159.720 30.375 160.105 ;
        RECT 30.545 159.550 30.715 160.275 ;
        RECT 29.440 159.245 29.655 159.295 ;
        RECT 27.860 158.835 28.755 159.210 ;
        RECT 29.265 159.165 29.655 159.245 ;
        RECT 29.825 159.480 30.715 159.550 ;
        RECT 30.885 159.950 31.105 160.435 ;
        RECT 31.275 160.115 31.525 160.655 ;
        RECT 31.695 160.005 31.955 160.485 ;
        RECT 30.885 159.525 31.215 159.950 ;
        RECT 29.825 159.455 30.720 159.480 ;
        RECT 29.825 159.440 30.730 159.455 ;
        RECT 29.825 159.425 30.735 159.440 ;
        RECT 29.825 159.420 30.745 159.425 ;
        RECT 29.825 159.410 30.750 159.420 ;
        RECT 29.825 159.400 30.755 159.410 ;
        RECT 29.825 159.395 30.765 159.400 ;
        RECT 29.825 159.385 30.775 159.395 ;
        RECT 29.825 159.380 30.785 159.385 ;
        RECT 26.805 158.405 27.690 158.575 ;
        RECT 27.870 158.105 28.185 158.605 ;
        RECT 28.415 158.275 28.755 158.835 ;
        RECT 28.925 158.105 29.095 159.115 ;
        RECT 29.265 158.320 29.595 159.165 ;
        RECT 29.825 158.930 30.085 159.380 ;
        RECT 30.450 159.375 30.785 159.380 ;
        RECT 30.450 159.370 30.800 159.375 ;
        RECT 30.450 159.360 30.815 159.370 ;
        RECT 30.450 159.355 30.840 159.360 ;
        RECT 31.385 159.355 31.615 159.750 ;
        RECT 30.450 159.350 31.615 159.355 ;
        RECT 30.480 159.315 31.615 159.350 ;
        RECT 30.515 159.290 31.615 159.315 ;
        RECT 30.545 159.260 31.615 159.290 ;
        RECT 30.565 159.230 31.615 159.260 ;
        RECT 30.585 159.200 31.615 159.230 ;
        RECT 30.655 159.190 31.615 159.200 ;
        RECT 30.680 159.180 31.615 159.190 ;
        RECT 30.700 159.165 31.615 159.180 ;
        RECT 30.720 159.150 31.615 159.165 ;
        RECT 30.725 159.140 31.510 159.150 ;
        RECT 30.740 159.105 31.510 159.140 ;
        RECT 30.255 158.785 30.585 159.030 ;
        RECT 30.755 158.855 31.510 159.105 ;
        RECT 31.785 158.975 31.955 160.005 ;
        RECT 32.125 159.885 34.715 160.655 ;
        RECT 35.435 160.105 35.605 160.395 ;
        RECT 35.775 160.275 36.105 160.655 ;
        RECT 35.435 159.935 36.100 160.105 ;
        RECT 32.125 159.365 33.335 159.885 ;
        RECT 33.505 159.195 34.715 159.715 ;
        RECT 30.255 158.760 30.440 158.785 ;
        RECT 29.825 158.660 30.440 158.760 ;
        RECT 29.825 158.105 30.430 158.660 ;
        RECT 30.605 158.275 31.085 158.615 ;
        RECT 31.255 158.105 31.510 158.650 ;
        RECT 31.680 158.275 31.955 158.975 ;
        RECT 32.125 158.105 34.715 159.195 ;
        RECT 35.350 159.115 35.700 159.765 ;
        RECT 35.870 158.945 36.100 159.935 ;
        RECT 35.435 158.775 36.100 158.945 ;
        RECT 35.435 158.275 35.605 158.775 ;
        RECT 35.775 158.105 36.105 158.605 ;
        RECT 36.275 158.275 36.460 160.395 ;
        RECT 36.715 160.195 36.965 160.655 ;
        RECT 37.135 160.205 37.470 160.375 ;
        RECT 37.665 160.205 38.340 160.375 ;
        RECT 37.135 160.065 37.305 160.205 ;
        RECT 36.630 159.075 36.910 160.025 ;
        RECT 37.080 159.935 37.305 160.065 ;
        RECT 37.080 158.830 37.250 159.935 ;
        RECT 37.475 159.785 38.000 160.005 ;
        RECT 37.420 159.020 37.660 159.615 ;
        RECT 37.830 159.085 38.000 159.785 ;
        RECT 38.170 159.425 38.340 160.205 ;
        RECT 38.660 160.155 39.030 160.655 ;
        RECT 39.210 160.205 39.615 160.375 ;
        RECT 39.785 160.205 40.570 160.375 ;
        RECT 39.210 159.975 39.380 160.205 ;
        RECT 38.550 159.675 39.380 159.975 ;
        RECT 39.765 159.705 40.230 160.035 ;
        RECT 38.550 159.645 38.750 159.675 ;
        RECT 38.870 159.425 39.040 159.495 ;
        RECT 38.170 159.255 39.040 159.425 ;
        RECT 38.530 159.165 39.040 159.255 ;
        RECT 37.080 158.700 37.385 158.830 ;
        RECT 37.830 158.720 38.360 159.085 ;
        RECT 36.700 158.105 36.965 158.565 ;
        RECT 37.135 158.275 37.385 158.700 ;
        RECT 38.530 158.550 38.700 159.165 ;
        RECT 37.595 158.380 38.700 158.550 ;
        RECT 38.870 158.105 39.040 158.905 ;
        RECT 39.210 158.605 39.380 159.675 ;
        RECT 39.550 158.775 39.740 159.495 ;
        RECT 39.910 158.745 40.230 159.705 ;
        RECT 40.400 159.745 40.570 160.205 ;
        RECT 40.845 160.125 41.055 160.655 ;
        RECT 41.315 159.915 41.645 160.440 ;
        RECT 41.815 160.045 41.985 160.655 ;
        RECT 42.155 160.000 42.485 160.435 ;
        RECT 42.155 159.915 42.535 160.000 ;
        RECT 43.165 159.930 43.455 160.655 ;
        RECT 41.445 159.745 41.645 159.915 ;
        RECT 42.310 159.875 42.535 159.915 ;
        RECT 40.400 159.415 41.275 159.745 ;
        RECT 41.445 159.415 42.195 159.745 ;
        RECT 39.210 158.275 39.460 158.605 ;
        RECT 40.400 158.575 40.570 159.415 ;
        RECT 41.445 159.210 41.635 159.415 ;
        RECT 42.365 159.295 42.535 159.875 ;
        RECT 43.625 159.905 44.835 160.655 ;
        RECT 45.055 160.000 45.385 160.435 ;
        RECT 45.555 160.045 45.725 160.655 ;
        RECT 45.005 159.915 45.385 160.000 ;
        RECT 45.895 159.915 46.225 160.440 ;
        RECT 46.485 160.125 46.695 160.655 ;
        RECT 46.970 160.205 47.755 160.375 ;
        RECT 47.925 160.205 48.330 160.375 ;
        RECT 43.625 159.365 44.145 159.905 ;
        RECT 45.005 159.875 45.230 159.915 ;
        RECT 42.320 159.245 42.535 159.295 ;
        RECT 40.740 158.835 41.635 159.210 ;
        RECT 42.145 159.165 42.535 159.245 ;
        RECT 39.685 158.405 40.570 158.575 ;
        RECT 40.750 158.105 41.065 158.605 ;
        RECT 41.295 158.275 41.635 158.835 ;
        RECT 41.805 158.105 41.975 159.115 ;
        RECT 42.145 158.320 42.475 159.165 ;
        RECT 43.165 158.105 43.455 159.270 ;
        RECT 44.315 159.195 44.835 159.735 ;
        RECT 43.625 158.105 44.835 159.195 ;
        RECT 45.005 159.295 45.175 159.875 ;
        RECT 45.895 159.745 46.095 159.915 ;
        RECT 46.970 159.745 47.140 160.205 ;
        RECT 45.345 159.415 46.095 159.745 ;
        RECT 46.265 159.415 47.140 159.745 ;
        RECT 45.005 159.245 45.220 159.295 ;
        RECT 45.005 159.165 45.395 159.245 ;
        RECT 45.065 158.320 45.395 159.165 ;
        RECT 45.905 159.210 46.095 159.415 ;
        RECT 45.565 158.105 45.735 159.115 ;
        RECT 45.905 158.835 46.800 159.210 ;
        RECT 45.905 158.275 46.245 158.835 ;
        RECT 46.475 158.105 46.790 158.605 ;
        RECT 46.970 158.575 47.140 159.415 ;
        RECT 47.310 159.705 47.775 160.035 ;
        RECT 48.160 159.975 48.330 160.205 ;
        RECT 48.510 160.155 48.880 160.655 ;
        RECT 49.200 160.205 49.875 160.375 ;
        RECT 50.070 160.205 50.405 160.375 ;
        RECT 47.310 158.745 47.630 159.705 ;
        RECT 48.160 159.675 48.990 159.975 ;
        RECT 47.800 158.775 47.990 159.495 ;
        RECT 48.160 158.605 48.330 159.675 ;
        RECT 48.790 159.645 48.990 159.675 ;
        RECT 48.500 159.425 48.670 159.495 ;
        RECT 49.200 159.425 49.370 160.205 ;
        RECT 50.235 160.065 50.405 160.205 ;
        RECT 50.575 160.195 50.825 160.655 ;
        RECT 48.500 159.255 49.370 159.425 ;
        RECT 49.540 159.785 50.065 160.005 ;
        RECT 50.235 159.935 50.460 160.065 ;
        RECT 48.500 159.165 49.010 159.255 ;
        RECT 46.970 158.405 47.855 158.575 ;
        RECT 48.080 158.275 48.330 158.605 ;
        RECT 48.500 158.105 48.670 158.905 ;
        RECT 48.840 158.550 49.010 159.165 ;
        RECT 49.540 159.085 49.710 159.785 ;
        RECT 49.180 158.720 49.710 159.085 ;
        RECT 49.880 159.020 50.120 159.615 ;
        RECT 50.290 158.830 50.460 159.935 ;
        RECT 50.630 159.075 50.910 160.025 ;
        RECT 50.155 158.700 50.460 158.830 ;
        RECT 48.840 158.380 49.945 158.550 ;
        RECT 50.155 158.275 50.405 158.700 ;
        RECT 50.575 158.105 50.840 158.565 ;
        RECT 51.080 158.275 51.265 160.395 ;
        RECT 51.435 160.275 51.765 160.655 ;
        RECT 51.935 160.105 52.105 160.395 ;
        RECT 52.365 160.110 57.710 160.655 ;
        RECT 51.440 159.935 52.105 160.105 ;
        RECT 51.440 158.945 51.670 159.935 ;
        RECT 51.840 159.115 52.190 159.765 ;
        RECT 53.950 159.280 54.290 160.110 ;
        RECT 57.885 159.885 61.395 160.655 ;
        RECT 51.440 158.775 52.105 158.945 ;
        RECT 51.435 158.105 51.765 158.605 ;
        RECT 51.935 158.275 52.105 158.775 ;
        RECT 55.770 158.540 56.120 159.790 ;
        RECT 57.885 159.365 59.535 159.885 ;
        RECT 62.085 159.835 62.295 160.655 ;
        RECT 62.465 159.855 62.795 160.485 ;
        RECT 59.705 159.195 61.395 159.715 ;
        RECT 62.465 159.255 62.715 159.855 ;
        RECT 62.965 159.835 63.195 160.655 ;
        RECT 64.325 159.915 64.710 160.485 ;
        RECT 64.880 160.195 65.205 160.655 ;
        RECT 65.725 160.025 66.005 160.485 ;
        RECT 62.885 159.415 63.215 159.665 ;
        RECT 52.365 158.105 57.710 158.540 ;
        RECT 57.885 158.105 61.395 159.195 ;
        RECT 62.085 158.105 62.295 159.245 ;
        RECT 62.465 158.275 62.795 159.255 ;
        RECT 64.325 159.245 64.605 159.915 ;
        RECT 64.880 159.855 66.005 160.025 ;
        RECT 64.880 159.745 65.330 159.855 ;
        RECT 64.775 159.415 65.330 159.745 ;
        RECT 66.195 159.685 66.595 160.485 ;
        RECT 66.995 160.195 67.265 160.655 ;
        RECT 67.435 160.025 67.720 160.485 ;
        RECT 62.965 158.105 63.195 159.245 ;
        RECT 64.325 158.275 64.710 159.245 ;
        RECT 64.880 158.955 65.330 159.415 ;
        RECT 65.500 159.125 66.595 159.685 ;
        RECT 64.880 158.735 66.005 158.955 ;
        RECT 64.880 158.105 65.205 158.565 ;
        RECT 65.725 158.275 66.005 158.735 ;
        RECT 66.195 158.275 66.595 159.125 ;
        RECT 66.765 159.855 67.720 160.025 ;
        RECT 68.925 159.930 69.215 160.655 ;
        RECT 69.385 160.110 74.730 160.655 ;
        RECT 66.765 158.955 66.975 159.855 ;
        RECT 67.145 159.125 67.835 159.685 ;
        RECT 70.970 159.280 71.310 160.110 ;
        RECT 74.905 159.885 78.415 160.655 ;
        RECT 79.620 160.025 79.905 160.485 ;
        RECT 80.075 160.195 80.345 160.655 ;
        RECT 66.765 158.735 67.720 158.955 ;
        RECT 66.995 158.105 67.265 158.565 ;
        RECT 67.435 158.275 67.720 158.735 ;
        RECT 68.925 158.105 69.215 159.270 ;
        RECT 72.790 158.540 73.140 159.790 ;
        RECT 74.905 159.365 76.555 159.885 ;
        RECT 79.620 159.855 80.575 160.025 ;
        RECT 76.725 159.195 78.415 159.715 ;
        RECT 69.385 158.105 74.730 158.540 ;
        RECT 74.905 158.105 78.415 159.195 ;
        RECT 79.505 159.125 80.195 159.685 ;
        RECT 80.365 158.955 80.575 159.855 ;
        RECT 79.620 158.735 80.575 158.955 ;
        RECT 80.745 159.685 81.145 160.485 ;
        RECT 81.335 160.025 81.615 160.485 ;
        RECT 82.135 160.195 82.460 160.655 ;
        RECT 81.335 159.855 82.460 160.025 ;
        RECT 82.630 159.915 83.015 160.485 ;
        RECT 82.010 159.745 82.460 159.855 ;
        RECT 80.745 159.125 81.840 159.685 ;
        RECT 82.010 159.415 82.565 159.745 ;
        RECT 79.620 158.275 79.905 158.735 ;
        RECT 80.075 158.105 80.345 158.565 ;
        RECT 80.745 158.275 81.145 159.125 ;
        RECT 82.010 158.955 82.460 159.415 ;
        RECT 82.735 159.245 83.015 159.915 ;
        RECT 83.185 159.885 86.695 160.655 ;
        RECT 86.915 160.135 87.170 160.435 ;
        RECT 87.340 160.255 87.670 160.655 ;
        RECT 86.865 160.085 87.170 160.135 ;
        RECT 87.840 160.085 88.010 160.435 ;
        RECT 88.310 160.175 88.480 160.655 ;
        RECT 88.715 160.145 89.065 160.475 ;
        RECT 89.235 160.175 89.405 160.655 ;
        RECT 86.865 160.005 88.010 160.085 ;
        RECT 86.865 159.975 88.575 160.005 ;
        RECT 86.865 159.915 88.725 159.975 ;
        RECT 83.185 159.365 84.835 159.885 ;
        RECT 81.335 158.735 82.460 158.955 ;
        RECT 81.335 158.275 81.615 158.735 ;
        RECT 82.135 158.105 82.460 158.565 ;
        RECT 82.630 158.275 83.015 159.245 ;
        RECT 85.005 159.195 86.695 159.715 ;
        RECT 83.185 158.105 86.695 159.195 ;
        RECT 86.865 159.245 87.035 159.915 ;
        RECT 87.840 159.835 88.725 159.915 ;
        RECT 88.405 159.805 88.725 159.835 ;
        RECT 87.210 159.415 87.510 159.745 ;
        RECT 86.865 158.815 87.170 159.245 ;
        RECT 87.340 158.955 87.510 159.415 ;
        RECT 87.770 159.125 88.305 159.665 ;
        RECT 88.555 159.415 88.725 159.805 ;
        RECT 88.895 159.245 89.065 160.145 ;
        RECT 89.655 160.005 89.915 160.450 ;
        RECT 88.670 159.040 89.065 159.245 ;
        RECT 89.235 159.835 89.915 160.005 ;
        RECT 90.550 159.835 90.825 160.655 ;
        RECT 90.995 160.015 91.325 160.485 ;
        RECT 91.495 160.185 91.665 160.655 ;
        RECT 91.835 160.015 92.165 160.485 ;
        RECT 92.335 160.185 92.505 160.655 ;
        RECT 92.675 160.015 93.005 160.485 ;
        RECT 93.175 160.185 93.345 160.655 ;
        RECT 93.515 160.015 93.845 160.485 ;
        RECT 94.015 160.185 94.300 160.655 ;
        RECT 90.995 159.835 94.515 160.015 ;
        RECT 94.685 159.930 94.975 160.655 ;
        RECT 95.310 160.145 95.550 160.655 ;
        RECT 95.730 160.145 96.010 160.475 ;
        RECT 96.240 160.145 96.455 160.655 ;
        RECT 87.340 158.870 88.450 158.955 ;
        RECT 89.235 158.930 89.405 159.835 ;
        RECT 89.575 159.100 89.915 159.665 ;
        RECT 90.600 159.465 92.260 159.665 ;
        RECT 92.580 159.465 93.945 159.665 ;
        RECT 94.115 159.295 94.515 159.835 ;
        RECT 95.205 159.415 95.560 159.975 ;
        RECT 90.550 159.075 92.585 159.285 ;
        RECT 89.235 158.870 89.915 158.930 ;
        RECT 87.340 158.785 89.915 158.870 ;
        RECT 88.280 158.700 89.915 158.785 ;
        RECT 86.865 158.375 88.065 158.615 ;
        RECT 88.245 158.105 88.575 158.530 ;
        RECT 89.090 158.105 89.450 158.530 ;
        RECT 89.655 158.520 89.915 158.700 ;
        RECT 90.550 158.275 90.825 159.075 ;
        RECT 90.995 158.105 91.325 158.905 ;
        RECT 91.495 158.275 91.665 159.075 ;
        RECT 91.835 158.105 92.085 158.905 ;
        RECT 92.255 158.445 92.585 159.075 ;
        RECT 92.755 158.995 94.515 159.295 ;
        RECT 92.755 158.615 92.925 158.995 ;
        RECT 93.095 158.445 93.425 158.805 ;
        RECT 93.595 158.615 93.765 158.995 ;
        RECT 93.935 158.445 94.350 158.825 ;
        RECT 92.255 158.275 94.350 158.445 ;
        RECT 94.685 158.105 94.975 159.270 ;
        RECT 95.730 159.245 95.900 160.145 ;
        RECT 96.070 159.415 96.335 159.975 ;
        RECT 96.625 159.915 97.240 160.485 ;
        RECT 96.585 159.245 96.755 159.745 ;
        RECT 95.330 159.075 96.755 159.245 ;
        RECT 95.330 158.900 95.720 159.075 ;
        RECT 96.205 158.105 96.535 158.905 ;
        RECT 96.925 158.895 97.240 159.915 ;
        RECT 97.905 160.035 98.170 160.485 ;
        RECT 98.340 160.205 98.630 160.655 ;
        RECT 98.800 160.035 99.090 160.485 ;
        RECT 97.905 159.865 99.090 160.035 ;
        RECT 99.270 159.745 99.515 160.350 ;
        RECT 97.925 159.080 98.255 159.665 ;
        RECT 98.425 159.415 98.910 159.665 ;
        RECT 99.255 159.415 99.515 159.745 ;
        RECT 99.765 159.415 100.035 160.350 ;
        RECT 100.215 159.665 100.425 160.350 ;
        RECT 100.595 160.005 100.935 160.485 ;
        RECT 101.115 160.175 101.425 160.655 ;
        RECT 100.595 159.835 101.265 160.005 ;
        RECT 101.095 159.745 101.265 159.835 ;
        RECT 100.215 159.415 100.695 159.665 ;
        RECT 101.095 159.415 101.435 159.745 ;
        RECT 96.705 158.275 97.240 158.895 ;
        RECT 97.905 158.105 98.230 158.905 ;
        RECT 98.425 158.325 98.610 159.415 ;
        RECT 101.095 159.245 101.265 159.415 ;
        RECT 98.780 159.075 101.265 159.245 ;
        RECT 98.780 158.275 99.030 159.075 ;
        RECT 99.200 158.105 99.940 158.905 ;
        RECT 100.125 158.275 100.455 159.075 ;
        RECT 100.625 158.105 101.435 158.905 ;
        RECT 101.605 158.275 101.865 160.485 ;
        RECT 102.045 159.915 102.430 160.485 ;
        RECT 102.600 160.195 102.925 160.655 ;
        RECT 103.445 160.025 103.725 160.485 ;
        RECT 102.045 159.245 102.325 159.915 ;
        RECT 102.600 159.855 103.725 160.025 ;
        RECT 102.600 159.745 103.050 159.855 ;
        RECT 102.495 159.415 103.050 159.745 ;
        RECT 103.915 159.685 104.315 160.485 ;
        RECT 104.715 160.195 104.985 160.655 ;
        RECT 105.155 160.025 105.440 160.485 ;
        RECT 102.045 158.275 102.430 159.245 ;
        RECT 102.600 158.955 103.050 159.415 ;
        RECT 103.220 159.125 104.315 159.685 ;
        RECT 102.600 158.735 103.725 158.955 ;
        RECT 102.600 158.105 102.925 158.565 ;
        RECT 103.445 158.275 103.725 158.735 ;
        RECT 103.915 158.275 104.315 159.125 ;
        RECT 104.485 159.855 105.440 160.025 ;
        RECT 105.725 160.155 105.985 160.485 ;
        RECT 106.155 160.295 106.485 160.655 ;
        RECT 106.740 160.275 108.040 160.485 ;
        RECT 105.725 160.145 105.955 160.155 ;
        RECT 104.485 158.955 104.695 159.855 ;
        RECT 104.865 159.125 105.555 159.685 ;
        RECT 105.725 158.955 105.895 160.145 ;
        RECT 106.740 160.125 106.910 160.275 ;
        RECT 106.155 160.000 106.910 160.125 ;
        RECT 106.065 159.955 106.910 160.000 ;
        RECT 106.065 159.835 106.335 159.955 ;
        RECT 106.065 159.260 106.235 159.835 ;
        RECT 106.465 159.395 106.875 159.700 ;
        RECT 107.165 159.665 107.375 160.065 ;
        RECT 107.045 159.455 107.375 159.665 ;
        RECT 107.620 159.665 107.840 160.065 ;
        RECT 108.315 159.890 108.770 160.655 ;
        RECT 110.135 159.855 110.395 160.655 ;
        RECT 110.565 160.005 110.895 160.485 ;
        RECT 111.065 160.175 111.255 160.655 ;
        RECT 111.425 160.235 113.475 160.485 ;
        RECT 111.425 160.005 111.685 160.235 ;
        RECT 113.645 160.215 113.925 160.655 ;
        RECT 114.115 160.125 114.305 160.485 ;
        RECT 114.475 160.295 114.805 160.655 ;
        RECT 114.975 160.125 115.165 160.370 ;
        RECT 110.565 159.835 111.685 160.005 ;
        RECT 111.855 160.045 113.485 160.065 ;
        RECT 114.115 160.045 115.165 160.125 ;
        RECT 111.855 159.875 115.165 160.045 ;
        RECT 115.335 159.935 115.670 160.655 ;
        RECT 111.855 159.845 114.160 159.875 ;
        RECT 107.620 159.455 108.095 159.665 ;
        RECT 108.285 159.465 108.775 159.665 ;
        RECT 106.065 159.225 106.265 159.260 ;
        RECT 107.595 159.225 108.770 159.285 ;
        RECT 106.065 159.115 108.770 159.225 ;
        RECT 106.125 159.055 107.925 159.115 ;
        RECT 107.595 159.025 107.925 159.055 ;
        RECT 104.485 158.735 105.440 158.955 ;
        RECT 104.715 158.105 104.985 158.565 ;
        RECT 105.155 158.275 105.440 158.735 ;
        RECT 105.725 158.275 105.985 158.955 ;
        RECT 106.155 158.105 106.405 158.885 ;
        RECT 106.655 158.855 107.490 158.865 ;
        RECT 108.080 158.855 108.265 158.945 ;
        RECT 106.655 158.655 108.265 158.855 ;
        RECT 106.655 158.275 106.905 158.655 ;
        RECT 108.035 158.615 108.265 158.655 ;
        RECT 108.515 158.495 108.770 159.115 ;
        RECT 110.290 159.260 111.535 159.665 ;
        RECT 111.760 159.430 113.195 159.675 ;
        RECT 113.365 159.260 113.710 159.675 ;
        RECT 110.290 159.035 113.710 159.260 ;
        RECT 113.880 159.155 114.160 159.845 ;
        RECT 115.885 159.835 116.115 160.655 ;
        RECT 116.285 159.855 116.615 160.485 ;
        RECT 115.360 159.705 115.670 159.745 ;
        RECT 114.330 159.325 115.670 159.705 ;
        RECT 115.865 159.415 116.195 159.665 ;
        RECT 116.365 159.255 116.615 159.855 ;
        RECT 116.785 159.835 116.995 160.655 ;
        RECT 117.225 159.855 117.920 160.485 ;
        RECT 118.125 159.855 118.435 160.655 ;
        RECT 119.065 159.855 119.375 160.655 ;
        RECT 119.580 159.855 120.275 160.485 ;
        RECT 120.445 159.930 120.735 160.655 ;
        RECT 120.920 160.085 121.175 160.435 ;
        RECT 121.345 160.255 121.675 160.655 ;
        RECT 121.845 160.085 122.015 160.435 ;
        RECT 122.185 160.255 122.565 160.655 ;
        RECT 120.920 159.915 122.585 160.085 ;
        RECT 122.755 159.980 123.030 160.325 ;
        RECT 123.265 160.195 123.510 160.655 ;
        RECT 117.245 159.415 117.580 159.665 ;
        RECT 117.750 159.255 117.920 159.855 ;
        RECT 118.090 159.415 118.425 159.685 ;
        RECT 119.075 159.415 119.410 159.685 ;
        RECT 119.580 159.255 119.750 159.855 ;
        RECT 122.415 159.745 122.585 159.915 ;
        RECT 119.920 159.415 120.255 159.665 ;
        RECT 120.905 159.415 121.250 159.745 ;
        RECT 121.420 159.415 122.245 159.745 ;
        RECT 122.415 159.415 122.690 159.745 ;
        RECT 113.880 159.035 115.180 159.155 ;
        RECT 107.075 158.105 107.430 158.485 ;
        RECT 108.435 158.275 108.770 158.495 ;
        RECT 110.135 158.635 113.845 158.865 ;
        RECT 114.015 158.705 115.180 159.035 ;
        RECT 110.135 158.275 110.395 158.635 ;
        RECT 110.565 158.105 110.895 158.465 ;
        RECT 111.075 158.275 111.255 158.635 ;
        RECT 111.425 158.105 111.755 158.465 ;
        RECT 111.925 158.275 112.115 158.635 ;
        RECT 112.285 158.105 112.615 158.465 ;
        RECT 112.785 158.275 112.975 158.635 ;
        RECT 113.645 158.535 113.845 158.635 ;
        RECT 113.645 158.525 114.805 158.535 ;
        RECT 115.385 158.525 115.580 158.945 ;
        RECT 113.145 158.105 113.475 158.465 ;
        RECT 113.645 158.275 115.580 158.525 ;
        RECT 115.885 158.105 116.115 159.245 ;
        RECT 116.285 158.275 116.615 159.255 ;
        RECT 116.785 158.105 116.995 159.245 ;
        RECT 117.225 158.105 117.485 159.245 ;
        RECT 117.655 158.275 117.985 159.255 ;
        RECT 118.155 158.105 118.435 159.245 ;
        RECT 119.065 158.105 119.345 159.245 ;
        RECT 119.515 158.275 119.845 159.255 ;
        RECT 120.015 158.105 120.275 159.245 ;
        RECT 120.445 158.105 120.735 159.270 ;
        RECT 120.925 158.955 121.250 159.245 ;
        RECT 121.420 159.125 121.615 159.415 ;
        RECT 122.415 159.245 122.585 159.415 ;
        RECT 122.860 159.245 123.030 159.980 ;
        RECT 123.205 159.415 123.520 160.025 ;
        RECT 123.690 159.665 123.940 160.475 ;
        RECT 124.110 160.130 124.370 160.655 ;
        RECT 124.540 160.005 124.800 160.460 ;
        RECT 124.970 160.175 125.230 160.655 ;
        RECT 125.400 160.005 125.660 160.460 ;
        RECT 125.830 160.175 126.090 160.655 ;
        RECT 126.260 160.005 126.520 160.460 ;
        RECT 126.690 160.175 126.950 160.655 ;
        RECT 127.120 160.005 127.380 160.460 ;
        RECT 127.550 160.175 127.850 160.655 ;
        RECT 124.540 159.835 127.850 160.005 ;
        RECT 128.470 159.875 128.970 160.485 ;
        RECT 123.690 159.415 126.710 159.665 ;
        RECT 121.925 159.075 122.585 159.245 ;
        RECT 121.925 158.955 122.095 159.075 ;
        RECT 120.925 158.785 122.095 158.955 ;
        RECT 120.905 158.325 122.095 158.615 ;
        RECT 122.265 158.105 122.545 158.905 ;
        RECT 122.755 158.275 123.030 159.245 ;
        RECT 123.215 158.105 123.510 159.215 ;
        RECT 123.690 158.280 123.940 159.415 ;
        RECT 126.880 159.245 127.850 159.835 ;
        RECT 128.265 159.415 128.615 159.665 ;
        RECT 128.800 159.245 128.970 159.875 ;
        RECT 129.600 160.005 129.930 160.485 ;
        RECT 130.100 160.195 130.325 160.655 ;
        RECT 130.495 160.005 130.825 160.485 ;
        RECT 129.600 159.835 130.825 160.005 ;
        RECT 131.015 159.855 131.265 160.655 ;
        RECT 131.435 159.855 131.775 160.485 ;
        RECT 131.950 159.890 132.405 160.655 ;
        RECT 132.680 160.275 133.980 160.485 ;
        RECT 134.235 160.295 134.565 160.655 ;
        RECT 133.810 160.125 133.980 160.275 ;
        RECT 134.735 160.155 134.995 160.485 ;
        RECT 134.765 160.145 134.995 160.155 ;
        RECT 131.545 159.805 131.775 159.855 ;
        RECT 129.140 159.465 129.470 159.665 ;
        RECT 129.640 159.465 129.970 159.665 ;
        RECT 130.140 159.465 130.560 159.665 ;
        RECT 130.735 159.495 131.430 159.665 ;
        RECT 130.735 159.245 130.905 159.495 ;
        RECT 131.600 159.245 131.775 159.805 ;
        RECT 132.880 159.665 133.100 160.065 ;
        RECT 131.945 159.465 132.435 159.665 ;
        RECT 132.625 159.455 133.100 159.665 ;
        RECT 133.345 159.665 133.555 160.065 ;
        RECT 133.810 160.000 134.565 160.125 ;
        RECT 133.810 159.955 134.655 160.000 ;
        RECT 134.385 159.835 134.655 159.955 ;
        RECT 133.345 159.455 133.675 159.665 ;
        RECT 133.845 159.395 134.255 159.700 ;
        RECT 124.110 158.105 124.370 159.215 ;
        RECT 124.540 159.005 127.850 159.245 ;
        RECT 128.470 159.075 130.905 159.245 ;
        RECT 124.540 158.280 124.800 159.005 ;
        RECT 124.970 158.105 125.230 158.835 ;
        RECT 125.400 158.280 125.660 159.005 ;
        RECT 125.830 158.105 126.090 158.835 ;
        RECT 126.260 158.280 126.520 159.005 ;
        RECT 126.690 158.105 126.950 158.835 ;
        RECT 127.120 158.280 127.380 159.005 ;
        RECT 127.550 158.105 127.845 158.835 ;
        RECT 128.470 158.275 128.800 159.075 ;
        RECT 128.970 158.105 129.300 158.905 ;
        RECT 129.600 158.275 129.930 159.075 ;
        RECT 130.575 158.105 130.825 158.905 ;
        RECT 131.095 158.105 131.265 159.245 ;
        RECT 131.435 158.275 131.775 159.245 ;
        RECT 131.950 159.225 133.125 159.285 ;
        RECT 134.485 159.260 134.655 159.835 ;
        RECT 134.455 159.225 134.655 159.260 ;
        RECT 131.950 159.115 134.655 159.225 ;
        RECT 131.950 158.495 132.205 159.115 ;
        RECT 132.795 159.055 134.595 159.115 ;
        RECT 132.795 159.025 133.125 159.055 ;
        RECT 134.825 158.955 134.995 160.145 ;
        RECT 135.715 160.105 135.885 160.395 ;
        RECT 136.055 160.275 136.385 160.655 ;
        RECT 135.715 159.935 136.380 160.105 ;
        RECT 135.630 159.115 135.980 159.765 ;
        RECT 132.455 158.855 132.640 158.945 ;
        RECT 133.230 158.855 134.065 158.865 ;
        RECT 132.455 158.655 134.065 158.855 ;
        RECT 132.455 158.615 132.685 158.655 ;
        RECT 131.950 158.275 132.285 158.495 ;
        RECT 133.290 158.105 133.645 158.485 ;
        RECT 133.815 158.275 134.065 158.655 ;
        RECT 134.315 158.105 134.565 158.885 ;
        RECT 134.735 158.275 134.995 158.955 ;
        RECT 136.150 158.945 136.380 159.935 ;
        RECT 135.715 158.775 136.380 158.945 ;
        RECT 135.715 158.275 135.885 158.775 ;
        RECT 136.055 158.105 136.385 158.605 ;
        RECT 136.555 158.275 136.740 160.395 ;
        RECT 136.995 160.195 137.245 160.655 ;
        RECT 137.415 160.205 137.750 160.375 ;
        RECT 137.945 160.205 138.620 160.375 ;
        RECT 137.415 160.065 137.585 160.205 ;
        RECT 136.910 159.075 137.190 160.025 ;
        RECT 137.360 159.935 137.585 160.065 ;
        RECT 137.360 158.830 137.530 159.935 ;
        RECT 137.755 159.785 138.280 160.005 ;
        RECT 137.700 159.020 137.940 159.615 ;
        RECT 138.110 159.085 138.280 159.785 ;
        RECT 138.450 159.425 138.620 160.205 ;
        RECT 138.940 160.155 139.310 160.655 ;
        RECT 139.490 160.205 139.895 160.375 ;
        RECT 140.065 160.205 140.850 160.375 ;
        RECT 139.490 159.975 139.660 160.205 ;
        RECT 138.830 159.675 139.660 159.975 ;
        RECT 140.045 159.705 140.510 160.035 ;
        RECT 138.830 159.645 139.030 159.675 ;
        RECT 139.150 159.425 139.320 159.495 ;
        RECT 138.450 159.255 139.320 159.425 ;
        RECT 138.810 159.165 139.320 159.255 ;
        RECT 137.360 158.700 137.665 158.830 ;
        RECT 138.110 158.720 138.640 159.085 ;
        RECT 136.980 158.105 137.245 158.565 ;
        RECT 137.415 158.275 137.665 158.700 ;
        RECT 138.810 158.550 138.980 159.165 ;
        RECT 137.875 158.380 138.980 158.550 ;
        RECT 139.150 158.105 139.320 158.905 ;
        RECT 139.490 158.605 139.660 159.675 ;
        RECT 139.830 158.775 140.020 159.495 ;
        RECT 140.190 158.745 140.510 159.705 ;
        RECT 140.680 159.745 140.850 160.205 ;
        RECT 141.125 160.125 141.335 160.655 ;
        RECT 141.595 159.915 141.925 160.440 ;
        RECT 142.095 160.045 142.265 160.655 ;
        RECT 142.435 160.000 142.765 160.435 ;
        RECT 143.995 160.105 144.165 160.485 ;
        RECT 144.380 160.275 144.710 160.655 ;
        RECT 142.435 159.915 142.815 160.000 ;
        RECT 143.995 159.935 144.710 160.105 ;
        RECT 141.725 159.745 141.925 159.915 ;
        RECT 142.590 159.875 142.815 159.915 ;
        RECT 140.680 159.415 141.555 159.745 ;
        RECT 141.725 159.415 142.475 159.745 ;
        RECT 139.490 158.275 139.740 158.605 ;
        RECT 140.680 158.575 140.850 159.415 ;
        RECT 141.725 159.210 141.915 159.415 ;
        RECT 142.645 159.295 142.815 159.875 ;
        RECT 143.905 159.385 144.260 159.755 ;
        RECT 144.540 159.745 144.710 159.935 ;
        RECT 144.880 159.910 145.135 160.485 ;
        RECT 144.540 159.415 144.795 159.745 ;
        RECT 142.600 159.245 142.815 159.295 ;
        RECT 141.020 158.835 141.915 159.210 ;
        RECT 142.425 159.165 142.815 159.245 ;
        RECT 144.540 159.205 144.710 159.415 ;
        RECT 139.965 158.405 140.850 158.575 ;
        RECT 141.030 158.105 141.345 158.605 ;
        RECT 141.575 158.275 141.915 158.835 ;
        RECT 142.085 158.105 142.255 159.115 ;
        RECT 142.425 158.320 142.755 159.165 ;
        RECT 143.995 159.035 144.710 159.205 ;
        RECT 144.965 159.180 145.135 159.910 ;
        RECT 145.310 159.815 145.570 160.655 ;
        RECT 145.745 159.905 146.955 160.655 ;
        RECT 143.995 158.275 144.165 159.035 ;
        RECT 144.380 158.105 144.710 158.865 ;
        RECT 144.880 158.275 145.135 159.180 ;
        RECT 145.310 158.105 145.570 159.255 ;
        RECT 145.745 159.195 146.265 159.735 ;
        RECT 146.435 159.365 146.955 159.905 ;
        RECT 145.745 158.105 146.955 159.195 ;
        RECT 17.320 157.935 147.040 158.105 ;
        RECT 17.405 156.845 18.615 157.935 ;
        RECT 18.785 157.500 24.130 157.935 ;
        RECT 24.305 157.500 29.650 157.935 ;
        RECT 17.405 156.135 17.925 156.675 ;
        RECT 18.095 156.305 18.615 156.845 ;
        RECT 17.405 155.385 18.615 156.135 ;
        RECT 20.370 155.930 20.710 156.760 ;
        RECT 22.190 156.250 22.540 157.500 ;
        RECT 25.890 155.930 26.230 156.760 ;
        RECT 27.710 156.250 28.060 157.500 ;
        RECT 30.285 156.770 30.575 157.935 ;
        RECT 30.745 157.500 36.090 157.935 ;
        RECT 18.785 155.385 24.130 155.930 ;
        RECT 24.305 155.385 29.650 155.930 ;
        RECT 30.285 155.385 30.575 156.110 ;
        RECT 32.330 155.930 32.670 156.760 ;
        RECT 34.150 156.250 34.500 157.500 ;
        RECT 36.725 157.065 37.000 157.765 ;
        RECT 37.170 157.390 37.425 157.935 ;
        RECT 37.595 157.425 38.075 157.765 ;
        RECT 38.250 157.380 38.855 157.935 ;
        RECT 39.025 157.500 44.370 157.935 ;
        RECT 44.545 157.500 49.890 157.935 ;
        RECT 50.065 157.500 55.410 157.935 ;
        RECT 38.240 157.280 38.855 157.380 ;
        RECT 38.240 157.255 38.425 157.280 ;
        RECT 36.725 156.035 36.895 157.065 ;
        RECT 37.170 156.935 37.925 157.185 ;
        RECT 38.095 157.010 38.425 157.255 ;
        RECT 37.170 156.900 37.940 156.935 ;
        RECT 37.170 156.890 37.955 156.900 ;
        RECT 37.065 156.875 37.960 156.890 ;
        RECT 37.065 156.860 37.980 156.875 ;
        RECT 37.065 156.850 38.000 156.860 ;
        RECT 37.065 156.840 38.025 156.850 ;
        RECT 37.065 156.810 38.095 156.840 ;
        RECT 37.065 156.780 38.115 156.810 ;
        RECT 37.065 156.750 38.135 156.780 ;
        RECT 37.065 156.725 38.165 156.750 ;
        RECT 37.065 156.690 38.200 156.725 ;
        RECT 37.065 156.685 38.230 156.690 ;
        RECT 37.065 156.290 37.295 156.685 ;
        RECT 37.840 156.680 38.230 156.685 ;
        RECT 37.865 156.670 38.230 156.680 ;
        RECT 37.880 156.665 38.230 156.670 ;
        RECT 37.895 156.660 38.230 156.665 ;
        RECT 38.595 156.660 38.855 157.110 ;
        RECT 37.895 156.655 38.855 156.660 ;
        RECT 37.905 156.645 38.855 156.655 ;
        RECT 37.915 156.640 38.855 156.645 ;
        RECT 37.925 156.630 38.855 156.640 ;
        RECT 37.930 156.620 38.855 156.630 ;
        RECT 37.935 156.615 38.855 156.620 ;
        RECT 37.945 156.600 38.855 156.615 ;
        RECT 37.950 156.585 38.855 156.600 ;
        RECT 37.960 156.560 38.855 156.585 ;
        RECT 37.465 156.090 37.795 156.515 ;
        RECT 30.745 155.385 36.090 155.930 ;
        RECT 36.725 155.555 36.985 156.035 ;
        RECT 37.155 155.385 37.405 155.925 ;
        RECT 37.575 155.605 37.795 156.090 ;
        RECT 37.965 156.490 38.855 156.560 ;
        RECT 37.965 155.765 38.135 156.490 ;
        RECT 38.305 155.935 38.855 156.320 ;
        RECT 40.610 155.930 40.950 156.760 ;
        RECT 42.430 156.250 42.780 157.500 ;
        RECT 46.130 155.930 46.470 156.760 ;
        RECT 47.950 156.250 48.300 157.500 ;
        RECT 51.650 155.930 51.990 156.760 ;
        RECT 53.470 156.250 53.820 157.500 ;
        RECT 56.045 156.770 56.335 157.935 ;
        RECT 56.505 156.845 58.175 157.935 ;
        RECT 58.920 157.305 59.205 157.765 ;
        RECT 59.375 157.475 59.645 157.935 ;
        RECT 58.920 157.085 59.875 157.305 ;
        RECT 56.505 156.155 57.255 156.675 ;
        RECT 57.425 156.325 58.175 156.845 ;
        RECT 58.805 156.355 59.495 156.915 ;
        RECT 59.665 156.185 59.875 157.085 ;
        RECT 37.965 155.595 38.855 155.765 ;
        RECT 39.025 155.385 44.370 155.930 ;
        RECT 44.545 155.385 49.890 155.930 ;
        RECT 50.065 155.385 55.410 155.930 ;
        RECT 56.045 155.385 56.335 156.110 ;
        RECT 56.505 155.385 58.175 156.155 ;
        RECT 58.920 156.015 59.875 156.185 ;
        RECT 60.045 156.915 60.445 157.765 ;
        RECT 60.635 157.305 60.915 157.765 ;
        RECT 61.435 157.475 61.760 157.935 ;
        RECT 60.635 157.085 61.760 157.305 ;
        RECT 60.045 156.355 61.140 156.915 ;
        RECT 61.310 156.625 61.760 157.085 ;
        RECT 61.930 156.795 62.315 157.765 ;
        RECT 58.920 155.555 59.205 156.015 ;
        RECT 59.375 155.385 59.645 155.845 ;
        RECT 60.045 155.555 60.445 156.355 ;
        RECT 61.310 156.295 61.865 156.625 ;
        RECT 61.310 156.185 61.760 156.295 ;
        RECT 60.635 156.015 61.760 156.185 ;
        RECT 62.035 156.125 62.315 156.795 ;
        RECT 60.635 155.555 60.915 156.015 ;
        RECT 61.435 155.385 61.760 155.845 ;
        RECT 61.930 155.555 62.315 156.125 ;
        RECT 62.495 155.565 62.755 157.755 ;
        RECT 62.925 157.205 63.265 157.935 ;
        RECT 63.445 157.025 63.715 157.755 ;
        RECT 62.945 156.805 63.715 157.025 ;
        RECT 63.895 157.045 64.125 157.755 ;
        RECT 64.295 157.225 64.625 157.935 ;
        RECT 64.795 157.045 65.055 157.755 ;
        RECT 63.895 156.805 65.055 157.045 ;
        RECT 66.200 157.145 66.735 157.765 ;
        RECT 62.945 156.135 63.235 156.805 ;
        RECT 63.415 156.315 63.880 156.625 ;
        RECT 64.060 156.315 64.585 156.625 ;
        RECT 62.945 155.935 64.175 156.135 ;
        RECT 63.015 155.385 63.685 155.755 ;
        RECT 63.865 155.565 64.175 155.935 ;
        RECT 64.355 155.675 64.585 156.315 ;
        RECT 64.765 156.295 65.065 156.625 ;
        RECT 66.200 156.125 66.515 157.145 ;
        RECT 66.905 157.135 67.235 157.935 ;
        RECT 68.470 157.510 68.805 157.935 ;
        RECT 68.975 157.330 69.160 157.735 ;
        RECT 68.495 157.155 69.160 157.330 ;
        RECT 69.365 157.155 69.695 157.935 ;
        RECT 67.720 156.965 68.110 157.140 ;
        RECT 66.685 156.795 68.110 156.965 ;
        RECT 66.685 156.295 66.855 156.795 ;
        RECT 64.765 155.385 65.055 156.115 ;
        RECT 66.200 155.555 66.815 156.125 ;
        RECT 67.105 156.065 67.370 156.625 ;
        RECT 67.540 155.895 67.710 156.795 ;
        RECT 67.880 156.065 68.235 156.625 ;
        RECT 68.495 156.125 68.835 157.155 ;
        RECT 69.865 156.965 70.135 157.735 ;
        RECT 69.005 156.795 70.135 156.965 ;
        RECT 70.315 156.965 70.645 157.750 ;
        RECT 70.315 156.795 70.995 156.965 ;
        RECT 71.175 156.795 71.505 157.935 ;
        RECT 71.775 157.265 71.945 157.765 ;
        RECT 72.115 157.435 72.445 157.935 ;
        RECT 71.775 157.095 72.440 157.265 ;
        RECT 69.005 156.295 69.255 156.795 ;
        RECT 68.495 155.955 69.180 156.125 ;
        RECT 69.435 156.045 69.795 156.625 ;
        RECT 66.985 155.385 67.200 155.895 ;
        RECT 67.430 155.565 67.710 155.895 ;
        RECT 67.890 155.385 68.130 155.895 ;
        RECT 68.470 155.385 68.805 155.785 ;
        RECT 68.975 155.555 69.180 155.955 ;
        RECT 69.965 155.885 70.135 156.795 ;
        RECT 70.305 156.375 70.655 156.625 ;
        RECT 70.825 156.195 70.995 156.795 ;
        RECT 71.165 156.375 71.515 156.625 ;
        RECT 71.690 156.275 72.040 156.925 ;
        RECT 69.390 155.385 69.665 155.865 ;
        RECT 69.875 155.555 70.135 155.885 ;
        RECT 70.325 155.385 70.565 156.195 ;
        RECT 70.735 155.555 71.065 156.195 ;
        RECT 71.235 155.385 71.505 156.195 ;
        RECT 72.210 156.105 72.440 157.095 ;
        RECT 71.775 155.935 72.440 156.105 ;
        RECT 71.775 155.645 71.945 155.935 ;
        RECT 72.115 155.385 72.445 155.765 ;
        RECT 72.615 155.645 72.800 157.765 ;
        RECT 73.040 157.475 73.305 157.935 ;
        RECT 73.475 157.340 73.725 157.765 ;
        RECT 73.935 157.490 75.040 157.660 ;
        RECT 73.420 157.210 73.725 157.340 ;
        RECT 72.970 156.015 73.250 156.965 ;
        RECT 73.420 156.105 73.590 157.210 ;
        RECT 73.760 156.425 74.000 157.020 ;
        RECT 74.170 156.955 74.700 157.320 ;
        RECT 74.170 156.255 74.340 156.955 ;
        RECT 74.870 156.875 75.040 157.490 ;
        RECT 75.210 157.135 75.380 157.935 ;
        RECT 75.550 157.435 75.800 157.765 ;
        RECT 76.025 157.465 76.910 157.635 ;
        RECT 74.870 156.785 75.380 156.875 ;
        RECT 73.420 155.975 73.645 156.105 ;
        RECT 73.815 156.035 74.340 156.255 ;
        RECT 74.510 156.615 75.380 156.785 ;
        RECT 73.055 155.385 73.305 155.845 ;
        RECT 73.475 155.835 73.645 155.975 ;
        RECT 74.510 155.835 74.680 156.615 ;
        RECT 75.210 156.545 75.380 156.615 ;
        RECT 74.890 156.365 75.090 156.395 ;
        RECT 75.550 156.365 75.720 157.435 ;
        RECT 75.890 156.545 76.080 157.265 ;
        RECT 74.890 156.065 75.720 156.365 ;
        RECT 76.250 156.335 76.570 157.295 ;
        RECT 73.475 155.665 73.810 155.835 ;
        RECT 74.005 155.665 74.680 155.835 ;
        RECT 75.000 155.385 75.370 155.885 ;
        RECT 75.550 155.835 75.720 156.065 ;
        RECT 76.105 156.005 76.570 156.335 ;
        RECT 76.740 156.625 76.910 157.465 ;
        RECT 77.090 157.435 77.405 157.935 ;
        RECT 77.635 157.205 77.975 157.765 ;
        RECT 77.080 156.830 77.975 157.205 ;
        RECT 78.145 156.925 78.315 157.935 ;
        RECT 77.785 156.625 77.975 156.830 ;
        RECT 78.485 156.875 78.815 157.720 ;
        RECT 79.045 157.065 79.320 157.765 ;
        RECT 79.490 157.390 79.745 157.935 ;
        RECT 79.915 157.425 80.395 157.765 ;
        RECT 80.570 157.380 81.175 157.935 ;
        RECT 80.560 157.280 81.175 157.380 ;
        RECT 80.560 157.255 80.745 157.280 ;
        RECT 78.485 156.795 78.875 156.875 ;
        RECT 78.660 156.745 78.875 156.795 ;
        RECT 76.740 156.295 77.615 156.625 ;
        RECT 77.785 156.295 78.535 156.625 ;
        RECT 76.740 155.835 76.910 156.295 ;
        RECT 77.785 156.125 77.985 156.295 ;
        RECT 78.705 156.165 78.875 156.745 ;
        RECT 78.650 156.125 78.875 156.165 ;
        RECT 75.550 155.665 75.955 155.835 ;
        RECT 76.125 155.665 76.910 155.835 ;
        RECT 77.185 155.385 77.395 155.915 ;
        RECT 77.655 155.600 77.985 156.125 ;
        RECT 78.495 156.040 78.875 156.125 ;
        RECT 78.155 155.385 78.325 155.995 ;
        RECT 78.495 155.605 78.825 156.040 ;
        RECT 79.045 156.035 79.215 157.065 ;
        RECT 79.490 156.935 80.245 157.185 ;
        RECT 80.415 157.010 80.745 157.255 ;
        RECT 79.490 156.900 80.260 156.935 ;
        RECT 79.490 156.890 80.275 156.900 ;
        RECT 79.385 156.875 80.280 156.890 ;
        RECT 79.385 156.860 80.300 156.875 ;
        RECT 79.385 156.850 80.320 156.860 ;
        RECT 79.385 156.840 80.345 156.850 ;
        RECT 79.385 156.810 80.415 156.840 ;
        RECT 79.385 156.780 80.435 156.810 ;
        RECT 79.385 156.750 80.455 156.780 ;
        RECT 79.385 156.725 80.485 156.750 ;
        RECT 79.385 156.690 80.520 156.725 ;
        RECT 79.385 156.685 80.550 156.690 ;
        RECT 79.385 156.290 79.615 156.685 ;
        RECT 80.160 156.680 80.550 156.685 ;
        RECT 80.185 156.670 80.550 156.680 ;
        RECT 80.200 156.665 80.550 156.670 ;
        RECT 80.215 156.660 80.550 156.665 ;
        RECT 80.915 156.660 81.175 157.110 ;
        RECT 81.805 156.770 82.095 157.935 ;
        RECT 82.265 157.500 87.610 157.935 ;
        RECT 87.785 157.500 93.130 157.935 ;
        RECT 80.215 156.655 81.175 156.660 ;
        RECT 80.225 156.645 81.175 156.655 ;
        RECT 80.235 156.640 81.175 156.645 ;
        RECT 80.245 156.630 81.175 156.640 ;
        RECT 80.250 156.620 81.175 156.630 ;
        RECT 80.255 156.615 81.175 156.620 ;
        RECT 80.265 156.600 81.175 156.615 ;
        RECT 80.270 156.585 81.175 156.600 ;
        RECT 80.280 156.560 81.175 156.585 ;
        RECT 79.785 156.090 80.115 156.515 ;
        RECT 79.865 156.065 80.115 156.090 ;
        RECT 79.045 155.555 79.305 156.035 ;
        RECT 79.475 155.385 79.725 155.925 ;
        RECT 79.895 155.605 80.115 156.065 ;
        RECT 80.285 156.490 81.175 156.560 ;
        RECT 80.285 155.765 80.455 156.490 ;
        RECT 80.625 155.935 81.175 156.320 ;
        RECT 80.285 155.595 81.175 155.765 ;
        RECT 81.805 155.385 82.095 156.110 ;
        RECT 83.850 155.930 84.190 156.760 ;
        RECT 85.670 156.250 86.020 157.500 ;
        RECT 89.370 155.930 89.710 156.760 ;
        RECT 91.190 156.250 91.540 157.500 ;
        RECT 93.305 156.845 96.815 157.935 ;
        RECT 93.305 156.155 94.955 156.675 ;
        RECT 95.125 156.325 96.815 156.845 ;
        RECT 97.455 156.965 97.785 157.750 ;
        RECT 97.455 156.795 98.135 156.965 ;
        RECT 98.315 156.795 98.645 157.935 ;
        RECT 98.825 157.500 104.170 157.935 ;
        RECT 97.445 156.375 97.795 156.625 ;
        RECT 97.965 156.195 98.135 156.795 ;
        RECT 98.305 156.375 98.655 156.625 ;
        RECT 82.265 155.385 87.610 155.930 ;
        RECT 87.785 155.385 93.130 155.930 ;
        RECT 93.305 155.385 96.815 156.155 ;
        RECT 97.465 155.385 97.705 156.195 ;
        RECT 97.875 155.555 98.205 156.195 ;
        RECT 98.375 155.385 98.645 156.195 ;
        RECT 100.410 155.930 100.750 156.760 ;
        RECT 102.230 156.250 102.580 157.500 ;
        RECT 104.345 156.845 106.935 157.935 ;
        RECT 104.345 156.155 105.555 156.675 ;
        RECT 105.725 156.325 106.935 156.845 ;
        RECT 107.565 156.770 107.855 157.935 ;
        RECT 108.025 156.845 111.535 157.935 ;
        RECT 112.280 157.305 112.565 157.765 ;
        RECT 112.735 157.475 113.005 157.935 ;
        RECT 112.280 157.085 113.235 157.305 ;
        RECT 108.025 156.155 109.675 156.675 ;
        RECT 109.845 156.325 111.535 156.845 ;
        RECT 112.165 156.355 112.855 156.915 ;
        RECT 113.025 156.185 113.235 157.085 ;
        RECT 98.825 155.385 104.170 155.930 ;
        RECT 104.345 155.385 106.935 156.155 ;
        RECT 107.565 155.385 107.855 156.110 ;
        RECT 108.025 155.385 111.535 156.155 ;
        RECT 112.280 156.015 113.235 156.185 ;
        RECT 113.405 156.915 113.805 157.765 ;
        RECT 113.995 157.305 114.275 157.765 ;
        RECT 114.795 157.475 115.120 157.935 ;
        RECT 113.995 157.085 115.120 157.305 ;
        RECT 113.405 156.355 114.500 156.915 ;
        RECT 114.670 156.625 115.120 157.085 ;
        RECT 115.290 156.795 115.675 157.765 ;
        RECT 115.845 156.795 116.135 157.935 ;
        RECT 116.930 157.595 118.295 157.765 ;
        RECT 116.930 157.385 117.260 157.595 ;
        RECT 116.305 157.135 117.260 157.385 ;
        RECT 112.280 155.555 112.565 156.015 ;
        RECT 112.735 155.385 113.005 155.845 ;
        RECT 113.405 155.555 113.805 156.355 ;
        RECT 114.670 156.295 115.225 156.625 ;
        RECT 114.670 156.185 115.120 156.295 ;
        RECT 113.995 156.015 115.120 156.185 ;
        RECT 115.395 156.125 115.675 156.795 ;
        RECT 115.845 156.295 116.120 156.625 ;
        RECT 113.995 155.555 114.275 156.015 ;
        RECT 114.795 155.385 115.120 155.845 ;
        RECT 115.290 155.555 115.675 156.125 ;
        RECT 116.305 156.125 116.475 157.135 ;
        RECT 116.645 156.295 117.000 156.960 ;
        RECT 117.185 156.295 117.460 156.960 ;
        RECT 117.630 156.625 117.955 157.425 ;
        RECT 118.125 156.965 118.295 157.595 ;
        RECT 118.465 157.135 118.755 157.935 ;
        RECT 118.125 156.795 118.800 156.965 ;
        RECT 118.970 156.795 119.355 157.755 ;
        RECT 119.525 156.845 121.195 157.935 ;
        RECT 118.630 156.625 118.800 156.795 ;
        RECT 117.630 156.295 117.975 156.625 ;
        RECT 118.185 156.375 118.435 156.625 ;
        RECT 118.630 156.375 118.995 156.625 ;
        RECT 118.265 156.295 118.435 156.375 ;
        RECT 118.805 156.295 118.995 156.375 ;
        RECT 119.180 156.125 119.355 156.795 ;
        RECT 115.845 155.765 116.135 156.035 ;
        RECT 116.305 155.935 116.730 156.125 ;
        RECT 116.900 155.955 118.300 156.125 ;
        RECT 116.900 155.765 117.230 155.955 ;
        RECT 115.845 155.555 117.230 155.765 ;
        RECT 117.465 155.385 117.795 155.785 ;
        RECT 117.970 155.555 118.300 155.955 ;
        RECT 118.505 155.385 118.675 155.945 ;
        RECT 118.845 155.555 119.355 156.125 ;
        RECT 119.525 156.155 120.275 156.675 ;
        RECT 120.445 156.325 121.195 156.845 ;
        RECT 121.835 156.795 122.165 157.935 ;
        RECT 122.695 156.965 123.025 157.750 ;
        RECT 123.205 157.100 123.550 157.935 ;
        RECT 122.345 156.795 123.025 156.965 ;
        RECT 123.725 156.930 123.980 157.735 ;
        RECT 124.150 157.100 124.410 157.935 ;
        RECT 124.585 156.930 124.840 157.735 ;
        RECT 125.010 157.100 125.270 157.935 ;
        RECT 125.440 156.930 125.700 157.735 ;
        RECT 125.870 157.100 126.255 157.935 ;
        RECT 127.070 156.965 127.460 157.140 ;
        RECT 127.945 157.135 128.275 157.935 ;
        RECT 128.445 157.145 128.980 157.765 ;
        RECT 129.195 157.215 129.525 157.935 ;
        RECT 121.825 156.375 122.175 156.625 ;
        RECT 122.345 156.195 122.515 156.795 ;
        RECT 123.225 156.760 126.255 156.930 ;
        RECT 127.070 156.795 128.495 156.965 ;
        RECT 122.685 156.375 123.035 156.625 ;
        RECT 123.225 156.195 123.395 156.760 ;
        RECT 123.565 156.365 125.780 156.590 ;
        RECT 125.955 156.195 126.255 156.760 ;
        RECT 119.525 155.385 121.195 156.155 ;
        RECT 121.835 155.385 122.105 156.195 ;
        RECT 122.275 155.555 122.605 156.195 ;
        RECT 122.775 155.385 123.015 156.195 ;
        RECT 123.225 156.025 126.255 156.195 ;
        RECT 126.945 156.065 127.300 156.625 ;
        RECT 123.685 155.385 123.980 155.855 ;
        RECT 124.150 155.580 124.410 156.025 ;
        RECT 124.580 155.385 124.840 155.855 ;
        RECT 125.010 155.580 125.265 156.025 ;
        RECT 127.470 155.895 127.640 156.795 ;
        RECT 127.810 156.065 128.075 156.625 ;
        RECT 128.325 156.295 128.495 156.795 ;
        RECT 128.665 156.125 128.980 157.145 ;
        RECT 129.185 156.575 129.415 156.915 ;
        RECT 129.705 156.575 129.920 157.690 ;
        RECT 130.115 156.990 130.445 157.765 ;
        RECT 130.615 157.160 131.325 157.935 ;
        RECT 130.115 156.775 131.265 156.990 ;
        RECT 129.185 156.375 129.515 156.575 ;
        RECT 129.705 156.395 130.155 156.575 ;
        RECT 129.825 156.375 130.155 156.395 ;
        RECT 130.325 156.375 130.795 156.605 ;
        RECT 130.980 156.205 131.265 156.775 ;
        RECT 131.495 156.330 131.775 157.765 ;
        RECT 131.945 156.845 133.155 157.935 ;
        RECT 125.435 155.385 125.735 155.855 ;
        RECT 127.050 155.385 127.290 155.895 ;
        RECT 127.470 155.565 127.750 155.895 ;
        RECT 127.980 155.385 128.195 155.895 ;
        RECT 128.365 155.555 128.980 156.125 ;
        RECT 129.185 156.015 130.365 156.205 ;
        RECT 129.185 155.555 129.525 156.015 ;
        RECT 130.035 155.935 130.365 156.015 ;
        RECT 130.555 156.015 131.265 156.205 ;
        RECT 130.555 155.875 130.855 156.015 ;
        RECT 130.540 155.865 130.855 155.875 ;
        RECT 130.530 155.855 130.855 155.865 ;
        RECT 130.520 155.850 130.855 155.855 ;
        RECT 129.695 155.385 129.865 155.845 ;
        RECT 130.515 155.840 130.855 155.850 ;
        RECT 130.510 155.835 130.855 155.840 ;
        RECT 130.505 155.825 130.855 155.835 ;
        RECT 130.500 155.820 130.855 155.825 ;
        RECT 130.495 155.555 130.855 155.820 ;
        RECT 131.095 155.385 131.265 155.845 ;
        RECT 131.435 155.555 131.775 156.330 ;
        RECT 131.945 156.135 132.465 156.675 ;
        RECT 132.635 156.305 133.155 156.845 ;
        RECT 133.325 156.770 133.615 157.935 ;
        RECT 133.790 157.135 134.045 157.935 ;
        RECT 134.245 157.085 134.575 157.765 ;
        RECT 133.790 156.595 134.035 156.955 ;
        RECT 134.225 156.805 134.575 157.085 ;
        RECT 134.225 156.425 134.395 156.805 ;
        RECT 134.755 156.625 134.950 157.675 ;
        RECT 135.130 156.795 135.450 157.935 ;
        RECT 135.715 157.005 135.885 157.765 ;
        RECT 136.065 157.175 136.395 157.935 ;
        RECT 135.715 156.835 136.380 157.005 ;
        RECT 136.565 156.860 136.835 157.765 ;
        RECT 136.210 156.690 136.380 156.835 ;
        RECT 133.875 156.255 134.395 156.425 ;
        RECT 134.565 156.295 134.950 156.625 ;
        RECT 135.130 156.575 135.390 156.625 ;
        RECT 135.130 156.405 135.395 156.575 ;
        RECT 135.130 156.295 135.390 156.405 ;
        RECT 135.645 156.285 135.975 156.655 ;
        RECT 136.210 156.360 136.495 156.690 ;
        RECT 131.945 155.385 133.155 156.135 ;
        RECT 133.325 155.385 133.615 156.110 ;
        RECT 133.875 155.690 134.045 156.255 ;
        RECT 136.210 156.105 136.380 156.360 ;
        RECT 134.235 155.915 135.450 156.085 ;
        RECT 134.235 155.610 134.465 155.915 ;
        RECT 134.635 155.385 134.965 155.745 ;
        RECT 135.160 155.565 135.450 155.915 ;
        RECT 135.715 155.935 136.380 156.105 ;
        RECT 136.665 156.060 136.835 156.860 ;
        RECT 135.715 155.555 135.885 155.935 ;
        RECT 136.065 155.385 136.395 155.765 ;
        RECT 136.575 155.555 136.835 156.060 ;
        RECT 137.010 156.795 137.345 157.765 ;
        RECT 137.515 156.795 137.685 157.935 ;
        RECT 137.855 157.595 139.885 157.765 ;
        RECT 137.010 156.125 137.180 156.795 ;
        RECT 137.855 156.625 138.025 157.595 ;
        RECT 137.350 156.295 137.605 156.625 ;
        RECT 137.830 156.295 138.025 156.625 ;
        RECT 138.195 157.255 139.320 157.425 ;
        RECT 137.435 156.125 137.605 156.295 ;
        RECT 138.195 156.125 138.365 157.255 ;
        RECT 137.010 155.555 137.265 156.125 ;
        RECT 137.435 155.955 138.365 156.125 ;
        RECT 138.535 156.915 139.545 157.085 ;
        RECT 138.535 156.115 138.705 156.915 ;
        RECT 138.910 156.235 139.185 156.715 ;
        RECT 138.905 156.065 139.185 156.235 ;
        RECT 138.190 155.920 138.365 155.955 ;
        RECT 137.435 155.385 137.765 155.785 ;
        RECT 138.190 155.555 138.720 155.920 ;
        RECT 138.910 155.555 139.185 156.065 ;
        RECT 139.355 155.555 139.545 156.915 ;
        RECT 139.715 156.930 139.885 157.595 ;
        RECT 140.055 157.175 140.225 157.935 ;
        RECT 140.460 157.175 140.975 157.585 ;
        RECT 139.715 156.740 140.465 156.930 ;
        RECT 140.635 156.365 140.975 157.175 ;
        RECT 139.745 156.195 140.975 156.365 ;
        RECT 141.145 156.795 141.530 157.765 ;
        RECT 141.700 157.475 142.025 157.935 ;
        RECT 142.545 157.305 142.825 157.765 ;
        RECT 141.700 157.085 142.825 157.305 ;
        RECT 139.725 155.385 140.235 155.920 ;
        RECT 140.455 155.590 140.700 156.195 ;
        RECT 141.145 156.125 141.425 156.795 ;
        RECT 141.700 156.625 142.150 157.085 ;
        RECT 143.015 156.915 143.415 157.765 ;
        RECT 143.815 157.475 144.085 157.935 ;
        RECT 144.255 157.305 144.540 157.765 ;
        RECT 141.595 156.295 142.150 156.625 ;
        RECT 142.320 156.355 143.415 156.915 ;
        RECT 141.700 156.185 142.150 156.295 ;
        RECT 141.145 155.555 141.530 156.125 ;
        RECT 141.700 156.015 142.825 156.185 ;
        RECT 141.700 155.385 142.025 155.845 ;
        RECT 142.545 155.555 142.825 156.015 ;
        RECT 143.015 155.555 143.415 156.355 ;
        RECT 143.585 157.085 144.540 157.305 ;
        RECT 143.585 156.185 143.795 157.085 ;
        RECT 143.965 156.355 144.655 156.915 ;
        RECT 145.745 156.845 146.955 157.935 ;
        RECT 145.745 156.305 146.265 156.845 ;
        RECT 143.585 156.015 144.540 156.185 ;
        RECT 146.435 156.135 146.955 156.675 ;
        RECT 143.815 155.385 144.085 155.845 ;
        RECT 144.255 155.555 144.540 156.015 ;
        RECT 145.745 155.385 146.955 156.135 ;
        RECT 17.320 155.215 147.040 155.385 ;
        RECT 17.405 154.465 18.615 155.215 ;
        RECT 18.875 154.665 19.045 155.045 ;
        RECT 19.260 154.835 19.590 155.215 ;
        RECT 18.875 154.495 19.590 154.665 ;
        RECT 17.405 153.925 17.925 154.465 ;
        RECT 18.095 153.755 18.615 154.295 ;
        RECT 18.785 153.945 19.140 154.315 ;
        RECT 19.420 154.305 19.590 154.495 ;
        RECT 19.760 154.470 20.015 155.045 ;
        RECT 19.420 153.975 19.675 154.305 ;
        RECT 19.420 153.765 19.590 153.975 ;
        RECT 17.405 152.665 18.615 153.755 ;
        RECT 18.875 153.595 19.590 153.765 ;
        RECT 19.845 153.740 20.015 154.470 ;
        RECT 20.190 154.375 20.450 155.215 ;
        RECT 20.625 154.670 25.970 155.215 ;
        RECT 26.145 154.670 31.490 155.215 ;
        RECT 31.665 154.670 37.010 155.215 ;
        RECT 37.185 154.670 42.530 155.215 ;
        RECT 22.210 153.840 22.550 154.670 ;
        RECT 18.875 152.835 19.045 153.595 ;
        RECT 19.260 152.665 19.590 153.425 ;
        RECT 19.760 152.835 20.015 153.740 ;
        RECT 20.190 152.665 20.450 153.815 ;
        RECT 24.030 153.100 24.380 154.350 ;
        RECT 27.730 153.840 28.070 154.670 ;
        RECT 29.550 153.100 29.900 154.350 ;
        RECT 33.250 153.840 33.590 154.670 ;
        RECT 35.070 153.100 35.420 154.350 ;
        RECT 38.770 153.840 39.110 154.670 ;
        RECT 43.165 154.490 43.455 155.215 ;
        RECT 43.625 154.670 48.970 155.215 ;
        RECT 49.145 154.670 54.490 155.215 ;
        RECT 40.590 153.100 40.940 154.350 ;
        RECT 45.210 153.840 45.550 154.670 ;
        RECT 20.625 152.665 25.970 153.100 ;
        RECT 26.145 152.665 31.490 153.100 ;
        RECT 31.665 152.665 37.010 153.100 ;
        RECT 37.185 152.665 42.530 153.100 ;
        RECT 43.165 152.665 43.455 153.830 ;
        RECT 47.030 153.100 47.380 154.350 ;
        RECT 50.730 153.840 51.070 154.670 ;
        RECT 54.665 154.465 55.875 155.215 ;
        RECT 56.325 154.585 56.705 155.035 ;
        RECT 52.550 153.100 52.900 154.350 ;
        RECT 54.665 153.925 55.185 154.465 ;
        RECT 55.355 153.755 55.875 154.295 ;
        RECT 43.625 152.665 48.970 153.100 ;
        RECT 49.145 152.665 54.490 153.100 ;
        RECT 54.665 152.665 55.875 153.755 ;
        RECT 56.065 153.635 56.295 154.325 ;
        RECT 56.475 154.135 56.705 154.585 ;
        RECT 56.885 154.435 57.115 155.215 ;
        RECT 57.295 154.505 57.725 155.035 ;
        RECT 57.295 154.255 57.540 154.505 ;
        RECT 57.905 154.305 58.115 154.925 ;
        RECT 58.285 154.485 58.615 155.215 ;
        RECT 58.895 154.665 59.065 154.955 ;
        RECT 59.235 154.835 59.565 155.215 ;
        RECT 58.895 154.495 59.560 154.665 ;
        RECT 56.475 153.455 56.815 154.135 ;
        RECT 56.055 153.255 56.815 153.455 ;
        RECT 57.005 153.955 57.540 154.255 ;
        RECT 57.720 153.955 58.115 154.305 ;
        RECT 58.310 153.955 58.600 154.305 ;
        RECT 56.055 152.865 56.315 153.255 ;
        RECT 56.485 152.665 56.815 153.075 ;
        RECT 57.005 152.845 57.335 153.955 ;
        RECT 57.505 153.575 58.545 153.775 ;
        RECT 58.810 153.675 59.160 154.325 ;
        RECT 57.505 152.845 57.695 153.575 ;
        RECT 57.865 152.665 58.195 153.395 ;
        RECT 58.375 152.845 58.545 153.575 ;
        RECT 59.330 153.505 59.560 154.495 ;
        RECT 58.895 153.335 59.560 153.505 ;
        RECT 58.895 152.835 59.065 153.335 ;
        RECT 59.235 152.665 59.565 153.165 ;
        RECT 59.735 152.835 59.920 154.955 ;
        RECT 60.175 154.755 60.425 155.215 ;
        RECT 60.595 154.765 60.930 154.935 ;
        RECT 61.125 154.765 61.800 154.935 ;
        RECT 60.595 154.625 60.765 154.765 ;
        RECT 60.090 153.635 60.370 154.585 ;
        RECT 60.540 154.495 60.765 154.625 ;
        RECT 60.540 153.390 60.710 154.495 ;
        RECT 60.935 154.345 61.460 154.565 ;
        RECT 60.880 153.580 61.120 154.175 ;
        RECT 61.290 153.645 61.460 154.345 ;
        RECT 61.630 153.985 61.800 154.765 ;
        RECT 62.120 154.715 62.490 155.215 ;
        RECT 62.670 154.765 63.075 154.935 ;
        RECT 63.245 154.765 64.030 154.935 ;
        RECT 62.670 154.535 62.840 154.765 ;
        RECT 62.010 154.235 62.840 154.535 ;
        RECT 63.225 154.265 63.690 154.595 ;
        RECT 62.010 154.205 62.210 154.235 ;
        RECT 62.330 153.985 62.500 154.055 ;
        RECT 61.630 153.815 62.500 153.985 ;
        RECT 61.990 153.725 62.500 153.815 ;
        RECT 60.540 153.260 60.845 153.390 ;
        RECT 61.290 153.280 61.820 153.645 ;
        RECT 60.160 152.665 60.425 153.125 ;
        RECT 60.595 152.835 60.845 153.260 ;
        RECT 61.990 153.110 62.160 153.725 ;
        RECT 61.055 152.940 62.160 153.110 ;
        RECT 62.330 152.665 62.500 153.465 ;
        RECT 62.670 153.165 62.840 154.235 ;
        RECT 63.010 153.335 63.200 154.055 ;
        RECT 63.370 153.305 63.690 154.265 ;
        RECT 63.860 154.305 64.030 154.765 ;
        RECT 64.305 154.685 64.515 155.215 ;
        RECT 64.775 154.475 65.105 155.000 ;
        RECT 65.275 154.605 65.445 155.215 ;
        RECT 65.615 154.560 65.945 154.995 ;
        RECT 66.170 154.710 66.505 155.215 ;
        RECT 66.675 154.645 66.915 155.020 ;
        RECT 67.195 154.885 67.365 155.030 ;
        RECT 67.195 154.690 67.570 154.885 ;
        RECT 67.930 154.720 68.325 155.215 ;
        RECT 65.615 154.475 65.995 154.560 ;
        RECT 64.905 154.305 65.105 154.475 ;
        RECT 65.770 154.435 65.995 154.475 ;
        RECT 63.860 153.975 64.735 154.305 ;
        RECT 64.905 153.975 65.655 154.305 ;
        RECT 62.670 152.835 62.920 153.165 ;
        RECT 63.860 153.135 64.030 153.975 ;
        RECT 64.905 153.770 65.095 153.975 ;
        RECT 65.825 153.855 65.995 154.435 ;
        RECT 65.780 153.805 65.995 153.855 ;
        RECT 64.200 153.395 65.095 153.770 ;
        RECT 65.605 153.725 65.995 153.805 ;
        RECT 63.145 152.965 64.030 153.135 ;
        RECT 64.210 152.665 64.525 153.165 ;
        RECT 64.755 152.835 65.095 153.395 ;
        RECT 65.265 152.665 65.435 153.675 ;
        RECT 65.605 152.880 65.935 153.725 ;
        RECT 66.225 153.685 66.525 154.535 ;
        RECT 66.695 154.495 66.915 154.645 ;
        RECT 66.695 154.165 67.230 154.495 ;
        RECT 67.400 154.355 67.570 154.690 ;
        RECT 68.495 154.525 68.735 155.045 ;
        RECT 66.695 153.515 66.930 154.165 ;
        RECT 67.400 153.995 68.385 154.355 ;
        RECT 66.255 153.285 66.930 153.515 ;
        RECT 67.100 153.975 68.385 153.995 ;
        RECT 67.100 153.825 67.960 153.975 ;
        RECT 66.255 152.855 66.425 153.285 ;
        RECT 66.595 152.665 66.925 153.115 ;
        RECT 67.100 152.880 67.385 153.825 ;
        RECT 68.560 153.720 68.735 154.525 ;
        RECT 68.925 154.490 69.215 155.215 ;
        RECT 69.385 154.585 69.725 155.045 ;
        RECT 69.895 154.755 70.065 155.215 ;
        RECT 70.695 154.780 71.055 155.045 ;
        RECT 70.700 154.775 71.055 154.780 ;
        RECT 70.705 154.765 71.055 154.775 ;
        RECT 70.710 154.760 71.055 154.765 ;
        RECT 70.715 154.750 71.055 154.760 ;
        RECT 71.295 154.755 71.465 155.215 ;
        RECT 70.720 154.745 71.055 154.750 ;
        RECT 70.730 154.735 71.055 154.745 ;
        RECT 70.740 154.725 71.055 154.735 ;
        RECT 70.235 154.585 70.565 154.665 ;
        RECT 69.385 154.395 70.565 154.585 ;
        RECT 70.755 154.585 71.055 154.725 ;
        RECT 70.755 154.395 71.465 154.585 ;
        RECT 69.385 154.025 69.715 154.225 ;
        RECT 70.025 154.205 70.355 154.225 ;
        RECT 69.905 154.025 70.355 154.205 ;
        RECT 67.560 153.345 68.255 153.655 ;
        RECT 67.565 152.665 68.250 153.135 ;
        RECT 68.430 152.935 68.735 153.720 ;
        RECT 68.925 152.665 69.215 153.830 ;
        RECT 69.385 153.685 69.615 154.025 ;
        RECT 69.395 152.665 69.725 153.385 ;
        RECT 69.905 152.910 70.120 154.025 ;
        RECT 70.525 153.995 70.995 154.225 ;
        RECT 71.180 153.825 71.465 154.395 ;
        RECT 71.635 154.270 71.975 155.045 ;
        RECT 72.260 154.585 72.545 155.045 ;
        RECT 72.715 154.755 72.985 155.215 ;
        RECT 72.260 154.415 73.215 154.585 ;
        RECT 70.315 153.610 71.465 153.825 ;
        RECT 70.315 152.835 70.645 153.610 ;
        RECT 70.815 152.665 71.525 153.440 ;
        RECT 71.695 152.835 71.975 154.270 ;
        RECT 72.145 153.685 72.835 154.245 ;
        RECT 73.005 153.515 73.215 154.415 ;
        RECT 72.260 153.295 73.215 153.515 ;
        RECT 73.385 154.245 73.785 155.045 ;
        RECT 73.975 154.585 74.255 155.045 ;
        RECT 74.775 154.755 75.100 155.215 ;
        RECT 73.975 154.415 75.100 154.585 ;
        RECT 75.270 154.475 75.655 155.045 ;
        RECT 75.915 154.665 76.085 154.955 ;
        RECT 76.255 154.835 76.585 155.215 ;
        RECT 75.915 154.495 76.580 154.665 ;
        RECT 74.650 154.305 75.100 154.415 ;
        RECT 73.385 153.685 74.480 154.245 ;
        RECT 74.650 153.975 75.205 154.305 ;
        RECT 72.260 152.835 72.545 153.295 ;
        RECT 72.715 152.665 72.985 153.125 ;
        RECT 73.385 152.835 73.785 153.685 ;
        RECT 74.650 153.515 75.100 153.975 ;
        RECT 75.375 153.805 75.655 154.475 ;
        RECT 73.975 153.295 75.100 153.515 ;
        RECT 73.975 152.835 74.255 153.295 ;
        RECT 74.775 152.665 75.100 153.125 ;
        RECT 75.270 152.835 75.655 153.805 ;
        RECT 75.830 153.675 76.180 154.325 ;
        RECT 76.350 153.505 76.580 154.495 ;
        RECT 75.915 153.335 76.580 153.505 ;
        RECT 75.915 152.835 76.085 153.335 ;
        RECT 76.255 152.665 76.585 153.165 ;
        RECT 76.755 152.835 76.940 154.955 ;
        RECT 77.195 154.755 77.445 155.215 ;
        RECT 77.615 154.765 77.950 154.935 ;
        RECT 78.145 154.765 78.820 154.935 ;
        RECT 77.615 154.625 77.785 154.765 ;
        RECT 77.110 153.635 77.390 154.585 ;
        RECT 77.560 154.495 77.785 154.625 ;
        RECT 77.560 153.390 77.730 154.495 ;
        RECT 77.955 154.345 78.480 154.565 ;
        RECT 77.900 153.580 78.140 154.175 ;
        RECT 78.310 153.645 78.480 154.345 ;
        RECT 78.650 153.985 78.820 154.765 ;
        RECT 79.140 154.715 79.510 155.215 ;
        RECT 79.690 154.765 80.095 154.935 ;
        RECT 80.265 154.765 81.050 154.935 ;
        RECT 79.690 154.535 79.860 154.765 ;
        RECT 79.030 154.235 79.860 154.535 ;
        RECT 80.245 154.265 80.710 154.595 ;
        RECT 79.030 154.205 79.230 154.235 ;
        RECT 79.350 153.985 79.520 154.055 ;
        RECT 78.650 153.815 79.520 153.985 ;
        RECT 79.010 153.725 79.520 153.815 ;
        RECT 77.560 153.260 77.865 153.390 ;
        RECT 78.310 153.280 78.840 153.645 ;
        RECT 77.180 152.665 77.445 153.125 ;
        RECT 77.615 152.835 77.865 153.260 ;
        RECT 79.010 153.110 79.180 153.725 ;
        RECT 78.075 152.940 79.180 153.110 ;
        RECT 79.350 152.665 79.520 153.465 ;
        RECT 79.690 153.165 79.860 154.235 ;
        RECT 80.030 153.335 80.220 154.055 ;
        RECT 80.390 153.305 80.710 154.265 ;
        RECT 80.880 154.305 81.050 154.765 ;
        RECT 81.325 154.685 81.535 155.215 ;
        RECT 81.795 154.475 82.125 155.000 ;
        RECT 82.295 154.605 82.465 155.215 ;
        RECT 82.635 154.560 82.965 154.995 ;
        RECT 82.635 154.475 83.015 154.560 ;
        RECT 81.925 154.305 82.125 154.475 ;
        RECT 82.790 154.435 83.015 154.475 ;
        RECT 80.880 153.975 81.755 154.305 ;
        RECT 81.925 153.975 82.675 154.305 ;
        RECT 79.690 152.835 79.940 153.165 ;
        RECT 80.880 153.135 81.050 153.975 ;
        RECT 81.925 153.770 82.115 153.975 ;
        RECT 82.845 153.855 83.015 154.435 ;
        RECT 82.800 153.805 83.015 153.855 ;
        RECT 81.220 153.395 82.115 153.770 ;
        RECT 82.625 153.725 83.015 153.805 ;
        RECT 83.185 154.475 83.570 155.045 ;
        RECT 83.740 154.755 84.065 155.215 ;
        RECT 84.585 154.585 84.865 155.045 ;
        RECT 83.185 153.805 83.465 154.475 ;
        RECT 83.740 154.415 84.865 154.585 ;
        RECT 83.740 154.305 84.190 154.415 ;
        RECT 83.635 153.975 84.190 154.305 ;
        RECT 85.055 154.245 85.455 155.045 ;
        RECT 85.855 154.755 86.125 155.215 ;
        RECT 86.295 154.585 86.580 155.045 ;
        RECT 86.885 154.705 87.125 155.215 ;
        RECT 87.295 154.705 87.585 155.045 ;
        RECT 87.815 154.705 88.130 155.215 ;
        RECT 80.165 152.965 81.050 153.135 ;
        RECT 81.230 152.665 81.545 153.165 ;
        RECT 81.775 152.835 82.115 153.395 ;
        RECT 82.285 152.665 82.455 153.675 ;
        RECT 82.625 152.880 82.955 153.725 ;
        RECT 83.185 152.835 83.570 153.805 ;
        RECT 83.740 153.515 84.190 153.975 ;
        RECT 84.360 153.685 85.455 154.245 ;
        RECT 83.740 153.295 84.865 153.515 ;
        RECT 83.740 152.665 84.065 153.125 ;
        RECT 84.585 152.835 84.865 153.295 ;
        RECT 85.055 152.835 85.455 153.685 ;
        RECT 85.625 154.415 86.580 154.585 ;
        RECT 85.625 153.515 85.835 154.415 ;
        RECT 86.005 153.685 86.695 154.245 ;
        RECT 86.930 154.195 87.125 154.535 ;
        RECT 86.925 154.025 87.125 154.195 ;
        RECT 86.930 153.975 87.125 154.025 ;
        RECT 87.295 153.805 87.475 154.705 ;
        RECT 88.300 154.645 88.470 154.915 ;
        RECT 88.640 154.815 88.970 155.215 ;
        RECT 90.565 154.745 90.860 155.215 ;
        RECT 87.645 153.975 88.055 154.535 ;
        RECT 88.300 154.475 88.995 154.645 ;
        RECT 91.030 154.575 91.290 155.020 ;
        RECT 91.460 154.745 91.720 155.215 ;
        RECT 91.890 154.575 92.145 155.020 ;
        RECT 92.315 154.745 92.615 155.215 ;
        RECT 88.225 153.805 88.395 154.305 ;
        RECT 86.935 153.635 88.395 153.805 ;
        RECT 85.625 153.295 86.580 153.515 ;
        RECT 86.935 153.460 87.295 153.635 ;
        RECT 88.565 153.465 88.995 154.475 ;
        RECT 90.105 154.405 93.135 154.575 ;
        RECT 90.105 153.840 90.275 154.405 ;
        RECT 90.445 154.010 92.660 154.235 ;
        RECT 92.835 153.840 93.135 154.405 ;
        RECT 93.305 154.465 94.515 155.215 ;
        RECT 94.685 154.490 94.975 155.215 ;
        RECT 95.145 154.670 100.490 155.215 ;
        RECT 93.305 153.925 93.825 154.465 ;
        RECT 90.105 153.670 93.135 153.840 ;
        RECT 93.995 153.755 94.515 154.295 ;
        RECT 96.730 153.840 97.070 154.670 ;
        RECT 100.665 154.445 102.335 155.215 ;
        RECT 103.055 154.665 103.225 154.955 ;
        RECT 103.395 154.835 103.725 155.215 ;
        RECT 103.055 154.495 103.720 154.665 ;
        RECT 85.855 152.665 86.125 153.125 ;
        RECT 86.295 152.835 86.580 153.295 ;
        RECT 87.880 152.665 88.050 153.465 ;
        RECT 88.220 153.295 88.995 153.465 ;
        RECT 88.220 152.835 88.550 153.295 ;
        RECT 88.720 152.665 88.890 153.125 ;
        RECT 90.085 152.665 90.430 153.500 ;
        RECT 90.605 152.865 90.860 153.670 ;
        RECT 91.030 152.665 91.290 153.500 ;
        RECT 91.465 152.865 91.720 153.670 ;
        RECT 91.890 152.665 92.150 153.500 ;
        RECT 92.320 152.865 92.580 153.670 ;
        RECT 92.750 152.665 93.135 153.500 ;
        RECT 93.305 152.665 94.515 153.755 ;
        RECT 94.685 152.665 94.975 153.830 ;
        RECT 98.550 153.100 98.900 154.350 ;
        RECT 100.665 153.925 101.415 154.445 ;
        RECT 101.585 153.755 102.335 154.275 ;
        RECT 95.145 152.665 100.490 153.100 ;
        RECT 100.665 152.665 102.335 153.755 ;
        RECT 102.970 153.675 103.320 154.325 ;
        RECT 103.490 153.505 103.720 154.495 ;
        RECT 103.055 153.335 103.720 153.505 ;
        RECT 103.055 152.835 103.225 153.335 ;
        RECT 103.395 152.665 103.725 153.165 ;
        RECT 103.895 152.835 104.080 154.955 ;
        RECT 104.335 154.755 104.585 155.215 ;
        RECT 104.755 154.765 105.090 154.935 ;
        RECT 105.285 154.765 105.960 154.935 ;
        RECT 104.755 154.625 104.925 154.765 ;
        RECT 104.250 153.635 104.530 154.585 ;
        RECT 104.700 154.495 104.925 154.625 ;
        RECT 104.700 153.390 104.870 154.495 ;
        RECT 105.095 154.345 105.620 154.565 ;
        RECT 105.040 153.580 105.280 154.175 ;
        RECT 105.450 153.645 105.620 154.345 ;
        RECT 105.790 153.985 105.960 154.765 ;
        RECT 106.280 154.715 106.650 155.215 ;
        RECT 106.830 154.765 107.235 154.935 ;
        RECT 107.405 154.765 108.190 154.935 ;
        RECT 106.830 154.535 107.000 154.765 ;
        RECT 106.170 154.235 107.000 154.535 ;
        RECT 107.385 154.265 107.850 154.595 ;
        RECT 106.170 154.205 106.370 154.235 ;
        RECT 106.490 153.985 106.660 154.055 ;
        RECT 105.790 153.815 106.660 153.985 ;
        RECT 106.150 153.725 106.660 153.815 ;
        RECT 104.700 153.260 105.005 153.390 ;
        RECT 105.450 153.280 105.980 153.645 ;
        RECT 104.320 152.665 104.585 153.125 ;
        RECT 104.755 152.835 105.005 153.260 ;
        RECT 106.150 153.110 106.320 153.725 ;
        RECT 105.215 152.940 106.320 153.110 ;
        RECT 106.490 152.665 106.660 153.465 ;
        RECT 106.830 153.165 107.000 154.235 ;
        RECT 107.170 153.335 107.360 154.055 ;
        RECT 107.530 153.305 107.850 154.265 ;
        RECT 108.020 154.305 108.190 154.765 ;
        RECT 108.465 154.685 108.675 155.215 ;
        RECT 108.935 154.475 109.265 155.000 ;
        RECT 109.435 154.605 109.605 155.215 ;
        RECT 109.775 154.560 110.105 154.995 ;
        RECT 111.245 154.715 111.505 155.045 ;
        RECT 111.675 154.855 112.005 155.215 ;
        RECT 112.260 154.835 113.560 155.045 ;
        RECT 111.245 154.705 111.475 154.715 ;
        RECT 109.775 154.475 110.155 154.560 ;
        RECT 109.065 154.305 109.265 154.475 ;
        RECT 109.930 154.435 110.155 154.475 ;
        RECT 108.020 153.975 108.895 154.305 ;
        RECT 109.065 153.975 109.815 154.305 ;
        RECT 106.830 152.835 107.080 153.165 ;
        RECT 108.020 153.135 108.190 153.975 ;
        RECT 109.065 153.770 109.255 153.975 ;
        RECT 109.985 153.855 110.155 154.435 ;
        RECT 109.940 153.805 110.155 153.855 ;
        RECT 108.360 153.395 109.255 153.770 ;
        RECT 109.765 153.725 110.155 153.805 ;
        RECT 107.305 152.965 108.190 153.135 ;
        RECT 108.370 152.665 108.685 153.165 ;
        RECT 108.915 152.835 109.255 153.395 ;
        RECT 109.425 152.665 109.595 153.675 ;
        RECT 109.765 152.880 110.095 153.725 ;
        RECT 111.245 153.515 111.415 154.705 ;
        RECT 112.260 154.685 112.430 154.835 ;
        RECT 111.675 154.560 112.430 154.685 ;
        RECT 111.585 154.515 112.430 154.560 ;
        RECT 111.585 154.395 111.855 154.515 ;
        RECT 111.585 153.820 111.755 154.395 ;
        RECT 111.985 153.955 112.395 154.260 ;
        RECT 112.685 154.225 112.895 154.625 ;
        RECT 112.565 154.015 112.895 154.225 ;
        RECT 113.140 154.225 113.360 154.625 ;
        RECT 113.835 154.450 114.290 155.215 ;
        RECT 114.470 154.540 114.745 154.885 ;
        RECT 114.935 154.815 115.315 155.215 ;
        RECT 115.485 154.645 115.655 154.995 ;
        RECT 115.825 154.815 116.155 155.215 ;
        RECT 116.325 154.645 116.580 154.995 ;
        RECT 113.140 154.015 113.615 154.225 ;
        RECT 113.805 154.025 114.295 154.225 ;
        RECT 111.585 153.785 111.785 153.820 ;
        RECT 113.115 153.785 114.290 153.845 ;
        RECT 111.585 153.675 114.290 153.785 ;
        RECT 111.645 153.615 113.445 153.675 ;
        RECT 113.115 153.585 113.445 153.615 ;
        RECT 111.245 152.835 111.505 153.515 ;
        RECT 111.675 152.665 111.925 153.445 ;
        RECT 112.175 153.415 113.010 153.425 ;
        RECT 113.600 153.415 113.785 153.505 ;
        RECT 112.175 153.215 113.785 153.415 ;
        RECT 112.175 152.835 112.425 153.215 ;
        RECT 113.555 153.175 113.785 153.215 ;
        RECT 114.035 153.055 114.290 153.675 ;
        RECT 112.595 152.665 112.950 153.045 ;
        RECT 113.955 152.835 114.290 153.055 ;
        RECT 114.470 153.805 114.640 154.540 ;
        RECT 114.915 154.475 116.580 154.645 ;
        RECT 114.915 154.305 115.085 154.475 ;
        RECT 116.805 154.395 117.035 155.215 ;
        RECT 117.205 154.415 117.535 155.045 ;
        RECT 114.810 153.975 115.085 154.305 ;
        RECT 115.255 153.975 116.080 154.305 ;
        RECT 116.250 153.975 116.595 154.305 ;
        RECT 116.785 153.975 117.115 154.225 ;
        RECT 114.915 153.805 115.085 153.975 ;
        RECT 114.470 152.835 114.745 153.805 ;
        RECT 114.915 153.635 115.575 153.805 ;
        RECT 115.885 153.685 116.080 153.975 ;
        RECT 117.285 153.815 117.535 154.415 ;
        RECT 117.705 154.395 117.915 155.215 ;
        RECT 118.310 154.705 118.550 155.215 ;
        RECT 118.730 154.705 119.010 155.035 ;
        RECT 119.240 154.705 119.455 155.215 ;
        RECT 118.205 153.975 118.560 154.535 ;
        RECT 115.405 153.515 115.575 153.635 ;
        RECT 116.250 153.515 116.575 153.805 ;
        RECT 114.955 152.665 115.235 153.465 ;
        RECT 115.405 153.345 116.575 153.515 ;
        RECT 115.405 152.885 116.595 153.175 ;
        RECT 116.805 152.665 117.035 153.805 ;
        RECT 117.205 152.835 117.535 153.815 ;
        RECT 118.730 153.805 118.900 154.705 ;
        RECT 119.070 153.975 119.335 154.535 ;
        RECT 119.625 154.475 120.240 155.045 ;
        RECT 120.445 154.490 120.735 155.215 ;
        RECT 119.585 153.805 119.755 154.305 ;
        RECT 117.705 152.665 117.915 153.805 ;
        RECT 118.330 153.635 119.755 153.805 ;
        RECT 118.330 153.460 118.720 153.635 ;
        RECT 119.205 152.665 119.535 153.465 ;
        RECT 119.925 153.455 120.240 154.475 ;
        RECT 120.910 154.450 121.365 155.215 ;
        RECT 121.640 154.835 122.940 155.045 ;
        RECT 123.195 154.855 123.525 155.215 ;
        RECT 122.770 154.685 122.940 154.835 ;
        RECT 123.695 154.715 123.955 155.045 ;
        RECT 123.725 154.705 123.955 154.715 ;
        RECT 121.840 154.225 122.060 154.625 ;
        RECT 120.905 154.025 121.395 154.225 ;
        RECT 121.585 154.015 122.060 154.225 ;
        RECT 122.305 154.225 122.515 154.625 ;
        RECT 122.770 154.560 123.525 154.685 ;
        RECT 122.770 154.515 123.615 154.560 ;
        RECT 123.345 154.395 123.615 154.515 ;
        RECT 122.305 154.015 122.635 154.225 ;
        RECT 122.805 153.955 123.215 154.260 ;
        RECT 119.705 152.835 120.240 153.455 ;
        RECT 120.445 152.665 120.735 153.830 ;
        RECT 120.910 153.785 122.085 153.845 ;
        RECT 123.445 153.820 123.615 154.395 ;
        RECT 123.415 153.785 123.615 153.820 ;
        RECT 120.910 153.675 123.615 153.785 ;
        RECT 120.910 153.055 121.165 153.675 ;
        RECT 121.755 153.615 123.555 153.675 ;
        RECT 121.755 153.585 122.085 153.615 ;
        RECT 123.785 153.515 123.955 154.705 ;
        RECT 124.125 154.670 129.470 155.215 ;
        RECT 125.710 153.840 126.050 154.670 ;
        RECT 129.735 154.665 129.905 155.045 ;
        RECT 130.085 154.835 130.415 155.215 ;
        RECT 129.735 154.495 130.400 154.665 ;
        RECT 130.595 154.540 130.855 155.045 ;
        RECT 121.415 153.415 121.600 153.505 ;
        RECT 122.190 153.415 123.025 153.425 ;
        RECT 121.415 153.215 123.025 153.415 ;
        RECT 121.415 153.175 121.645 153.215 ;
        RECT 120.910 152.835 121.245 153.055 ;
        RECT 122.250 152.665 122.605 153.045 ;
        RECT 122.775 152.835 123.025 153.215 ;
        RECT 123.275 152.665 123.525 153.445 ;
        RECT 123.695 152.835 123.955 153.515 ;
        RECT 127.530 153.100 127.880 154.350 ;
        RECT 129.665 153.945 129.995 154.315 ;
        RECT 130.230 154.240 130.400 154.495 ;
        RECT 130.230 153.910 130.515 154.240 ;
        RECT 130.230 153.765 130.400 153.910 ;
        RECT 129.735 153.595 130.400 153.765 ;
        RECT 130.685 153.740 130.855 154.540 ;
        RECT 131.030 154.375 131.290 155.215 ;
        RECT 131.465 154.470 131.720 155.045 ;
        RECT 131.890 154.835 132.220 155.215 ;
        RECT 132.435 154.665 132.605 155.045 ;
        RECT 131.890 154.495 132.605 154.665 ;
        RECT 124.125 152.665 129.470 153.100 ;
        RECT 129.735 152.835 129.905 153.595 ;
        RECT 130.085 152.665 130.415 153.425 ;
        RECT 130.585 152.835 130.855 153.740 ;
        RECT 131.030 152.665 131.290 153.815 ;
        RECT 131.465 153.740 131.635 154.470 ;
        RECT 131.890 154.305 132.060 154.495 ;
        RECT 132.870 154.375 133.130 155.215 ;
        RECT 133.305 154.470 133.560 155.045 ;
        RECT 133.730 154.835 134.060 155.215 ;
        RECT 134.275 154.665 134.445 155.045 ;
        RECT 133.730 154.495 134.445 154.665 ;
        RECT 131.805 153.975 132.060 154.305 ;
        RECT 131.890 153.765 132.060 153.975 ;
        RECT 132.340 153.945 132.695 154.315 ;
        RECT 131.465 152.835 131.720 153.740 ;
        RECT 131.890 153.595 132.605 153.765 ;
        RECT 131.890 152.665 132.220 153.425 ;
        RECT 132.435 152.835 132.605 153.595 ;
        RECT 132.870 152.665 133.130 153.815 ;
        RECT 133.305 153.740 133.475 154.470 ;
        RECT 133.730 154.305 133.900 154.495 ;
        RECT 134.710 154.475 134.965 155.045 ;
        RECT 135.135 154.815 135.465 155.215 ;
        RECT 135.890 154.680 136.420 155.045 ;
        RECT 135.890 154.645 136.065 154.680 ;
        RECT 135.135 154.475 136.065 154.645 ;
        RECT 133.645 153.975 133.900 154.305 ;
        RECT 133.730 153.765 133.900 153.975 ;
        RECT 134.180 153.945 134.535 154.315 ;
        RECT 134.710 153.805 134.880 154.475 ;
        RECT 135.135 154.305 135.305 154.475 ;
        RECT 135.050 153.975 135.305 154.305 ;
        RECT 135.530 153.975 135.725 154.305 ;
        RECT 133.305 152.835 133.560 153.740 ;
        RECT 133.730 153.595 134.445 153.765 ;
        RECT 133.730 152.665 134.060 153.425 ;
        RECT 134.275 152.835 134.445 153.595 ;
        RECT 134.710 152.835 135.045 153.805 ;
        RECT 135.215 152.665 135.385 153.805 ;
        RECT 135.555 153.005 135.725 153.975 ;
        RECT 135.895 153.345 136.065 154.475 ;
        RECT 136.235 153.685 136.405 154.485 ;
        RECT 136.610 154.195 136.885 155.045 ;
        RECT 136.605 154.025 136.885 154.195 ;
        RECT 136.610 153.885 136.885 154.025 ;
        RECT 137.055 153.685 137.245 155.045 ;
        RECT 137.425 154.680 137.935 155.215 ;
        RECT 138.155 154.405 138.400 155.010 ;
        RECT 138.845 154.475 139.230 155.045 ;
        RECT 139.400 154.755 139.725 155.215 ;
        RECT 140.245 154.585 140.525 155.045 ;
        RECT 137.445 154.235 138.675 154.405 ;
        RECT 136.235 153.515 137.245 153.685 ;
        RECT 137.415 153.670 138.165 153.860 ;
        RECT 135.895 153.175 137.020 153.345 ;
        RECT 137.415 153.005 137.585 153.670 ;
        RECT 138.335 153.425 138.675 154.235 ;
        RECT 135.555 152.835 137.585 153.005 ;
        RECT 137.755 152.665 137.925 153.425 ;
        RECT 138.160 153.015 138.675 153.425 ;
        RECT 138.845 153.805 139.125 154.475 ;
        RECT 139.400 154.415 140.525 154.585 ;
        RECT 139.400 154.305 139.850 154.415 ;
        RECT 139.295 153.975 139.850 154.305 ;
        RECT 140.715 154.245 141.115 155.045 ;
        RECT 141.515 154.755 141.785 155.215 ;
        RECT 141.955 154.585 142.240 155.045 ;
        RECT 138.845 152.835 139.230 153.805 ;
        RECT 139.400 153.515 139.850 153.975 ;
        RECT 140.020 153.685 141.115 154.245 ;
        RECT 139.400 153.295 140.525 153.515 ;
        RECT 139.400 152.665 139.725 153.125 ;
        RECT 140.245 152.835 140.525 153.295 ;
        RECT 140.715 152.835 141.115 153.685 ;
        RECT 141.285 154.415 142.240 154.585 ;
        RECT 142.615 154.665 142.785 155.045 ;
        RECT 142.965 154.835 143.295 155.215 ;
        RECT 142.615 154.495 143.280 154.665 ;
        RECT 143.475 154.540 143.735 155.045 ;
        RECT 141.285 153.515 141.495 154.415 ;
        RECT 141.665 153.685 142.355 154.245 ;
        RECT 142.545 153.945 142.875 154.315 ;
        RECT 143.110 154.240 143.280 154.495 ;
        RECT 143.110 153.910 143.395 154.240 ;
        RECT 143.110 153.765 143.280 153.910 ;
        RECT 142.615 153.595 143.280 153.765 ;
        RECT 143.565 153.740 143.735 154.540 ;
        RECT 143.995 154.665 144.165 155.045 ;
        RECT 144.380 154.835 144.710 155.215 ;
        RECT 143.995 154.495 144.710 154.665 ;
        RECT 143.905 153.945 144.260 154.315 ;
        RECT 144.540 154.305 144.710 154.495 ;
        RECT 144.880 154.470 145.135 155.045 ;
        RECT 144.540 153.975 144.795 154.305 ;
        RECT 144.540 153.765 144.710 153.975 ;
        RECT 141.285 153.295 142.240 153.515 ;
        RECT 141.515 152.665 141.785 153.125 ;
        RECT 141.955 152.835 142.240 153.295 ;
        RECT 142.615 152.835 142.785 153.595 ;
        RECT 142.965 152.665 143.295 153.425 ;
        RECT 143.465 152.835 143.735 153.740 ;
        RECT 143.995 153.595 144.710 153.765 ;
        RECT 144.965 153.740 145.135 154.470 ;
        RECT 145.310 154.375 145.570 155.215 ;
        RECT 145.745 154.465 146.955 155.215 ;
        RECT 143.995 152.835 144.165 153.595 ;
        RECT 144.380 152.665 144.710 153.425 ;
        RECT 144.880 152.835 145.135 153.740 ;
        RECT 145.310 152.665 145.570 153.815 ;
        RECT 145.745 153.755 146.265 154.295 ;
        RECT 146.435 153.925 146.955 154.465 ;
        RECT 145.745 152.665 146.955 153.755 ;
        RECT 17.320 152.495 147.040 152.665 ;
        RECT 17.405 151.405 18.615 152.495 ;
        RECT 18.785 152.060 24.130 152.495 ;
        RECT 24.305 152.060 29.650 152.495 ;
        RECT 17.405 150.695 17.925 151.235 ;
        RECT 18.095 150.865 18.615 151.405 ;
        RECT 17.405 149.945 18.615 150.695 ;
        RECT 20.370 150.490 20.710 151.320 ;
        RECT 22.190 150.810 22.540 152.060 ;
        RECT 25.890 150.490 26.230 151.320 ;
        RECT 27.710 150.810 28.060 152.060 ;
        RECT 30.285 151.330 30.575 152.495 ;
        RECT 30.745 151.405 33.335 152.495 ;
        RECT 30.745 150.715 31.955 151.235 ;
        RECT 32.125 150.885 33.335 151.405 ;
        RECT 34.000 151.705 34.535 152.325 ;
        RECT 18.785 149.945 24.130 150.490 ;
        RECT 24.305 149.945 29.650 150.490 ;
        RECT 30.285 149.945 30.575 150.670 ;
        RECT 30.745 149.945 33.335 150.715 ;
        RECT 34.000 150.685 34.315 151.705 ;
        RECT 34.705 151.695 35.035 152.495 ;
        RECT 35.520 151.525 35.910 151.700 ;
        RECT 34.485 151.355 35.910 151.525 ;
        RECT 36.265 151.625 36.540 152.325 ;
        RECT 36.710 151.950 36.965 152.495 ;
        RECT 37.135 151.985 37.615 152.325 ;
        RECT 37.790 151.940 38.395 152.495 ;
        RECT 37.780 151.840 38.395 151.940 ;
        RECT 37.780 151.815 37.965 151.840 ;
        RECT 34.485 150.855 34.655 151.355 ;
        RECT 34.000 150.115 34.615 150.685 ;
        RECT 34.905 150.625 35.170 151.185 ;
        RECT 35.340 150.455 35.510 151.355 ;
        RECT 35.680 150.625 36.035 151.185 ;
        RECT 36.265 150.595 36.435 151.625 ;
        RECT 36.710 151.495 37.465 151.745 ;
        RECT 37.635 151.570 37.965 151.815 ;
        RECT 36.710 151.460 37.480 151.495 ;
        RECT 36.710 151.450 37.495 151.460 ;
        RECT 36.605 151.435 37.500 151.450 ;
        RECT 36.605 151.420 37.520 151.435 ;
        RECT 36.605 151.410 37.540 151.420 ;
        RECT 36.605 151.400 37.565 151.410 ;
        RECT 36.605 151.370 37.635 151.400 ;
        RECT 36.605 151.340 37.655 151.370 ;
        RECT 36.605 151.310 37.675 151.340 ;
        RECT 36.605 151.285 37.705 151.310 ;
        RECT 36.605 151.250 37.740 151.285 ;
        RECT 36.605 151.245 37.770 151.250 ;
        RECT 36.605 150.850 36.835 151.245 ;
        RECT 37.380 151.240 37.770 151.245 ;
        RECT 37.405 151.230 37.770 151.240 ;
        RECT 37.420 151.225 37.770 151.230 ;
        RECT 37.435 151.220 37.770 151.225 ;
        RECT 38.135 151.220 38.395 151.670 ;
        RECT 38.575 151.525 38.905 152.325 ;
        RECT 39.075 151.695 39.305 152.495 ;
        RECT 39.475 151.525 39.805 152.325 ;
        RECT 38.575 151.355 39.805 151.525 ;
        RECT 39.975 151.355 40.230 152.495 ;
        RECT 40.415 151.775 40.745 152.495 ;
        RECT 37.435 151.215 38.395 151.220 ;
        RECT 37.445 151.205 38.395 151.215 ;
        RECT 37.455 151.200 38.395 151.205 ;
        RECT 37.465 151.190 38.395 151.200 ;
        RECT 37.470 151.180 38.395 151.190 ;
        RECT 37.475 151.175 38.395 151.180 ;
        RECT 37.485 151.160 38.395 151.175 ;
        RECT 37.490 151.145 38.395 151.160 ;
        RECT 37.500 151.120 38.395 151.145 ;
        RECT 37.005 150.650 37.335 151.075 ;
        RECT 34.785 149.945 35.000 150.455 ;
        RECT 35.230 150.125 35.510 150.455 ;
        RECT 35.690 149.945 35.930 150.455 ;
        RECT 36.265 150.115 36.525 150.595 ;
        RECT 36.695 149.945 36.945 150.485 ;
        RECT 37.115 150.165 37.335 150.650 ;
        RECT 37.505 151.050 38.395 151.120 ;
        RECT 37.505 150.325 37.675 151.050 ;
        RECT 37.845 150.495 38.395 150.880 ;
        RECT 38.565 150.855 38.875 151.185 ;
        RECT 38.575 150.455 38.905 150.685 ;
        RECT 39.080 150.625 39.455 151.185 ;
        RECT 39.625 150.455 39.805 151.355 ;
        RECT 39.990 150.605 40.210 151.185 ;
        RECT 40.405 151.135 40.635 151.475 ;
        RECT 40.925 151.135 41.140 152.250 ;
        RECT 41.335 151.550 41.665 152.325 ;
        RECT 41.835 151.720 42.545 152.495 ;
        RECT 41.335 151.335 42.485 151.550 ;
        RECT 40.405 150.935 40.735 151.135 ;
        RECT 40.925 150.955 41.375 151.135 ;
        RECT 41.045 150.935 41.375 150.955 ;
        RECT 41.545 150.935 42.015 151.165 ;
        RECT 42.200 150.765 42.485 151.335 ;
        RECT 42.715 150.890 42.995 152.325 ;
        RECT 43.165 151.405 46.675 152.495 ;
        RECT 46.845 151.940 47.450 152.495 ;
        RECT 47.625 151.985 48.105 152.325 ;
        RECT 48.275 151.950 48.530 152.495 ;
        RECT 46.845 151.840 47.460 151.940 ;
        RECT 47.275 151.815 47.460 151.840 ;
        RECT 37.505 150.155 38.395 150.325 ;
        RECT 38.575 150.115 39.805 150.455 ;
        RECT 40.405 150.575 41.585 150.765 ;
        RECT 39.975 149.945 40.230 150.435 ;
        RECT 40.405 150.115 40.745 150.575 ;
        RECT 41.255 150.495 41.585 150.575 ;
        RECT 41.775 150.575 42.485 150.765 ;
        RECT 41.775 150.435 42.075 150.575 ;
        RECT 41.760 150.425 42.075 150.435 ;
        RECT 41.750 150.415 42.075 150.425 ;
        RECT 41.740 150.410 42.075 150.415 ;
        RECT 40.915 149.945 41.085 150.405 ;
        RECT 41.735 150.400 42.075 150.410 ;
        RECT 41.730 150.395 42.075 150.400 ;
        RECT 41.725 150.385 42.075 150.395 ;
        RECT 41.720 150.380 42.075 150.385 ;
        RECT 41.715 150.115 42.075 150.380 ;
        RECT 42.315 149.945 42.485 150.405 ;
        RECT 42.655 150.115 42.995 150.890 ;
        RECT 43.165 150.715 44.815 151.235 ;
        RECT 44.985 150.885 46.675 151.405 ;
        RECT 46.845 151.220 47.105 151.670 ;
        RECT 47.275 151.570 47.605 151.815 ;
        RECT 47.775 151.495 48.530 151.745 ;
        RECT 48.700 151.625 48.975 152.325 ;
        RECT 49.145 152.060 54.490 152.495 ;
        RECT 47.760 151.460 48.530 151.495 ;
        RECT 47.745 151.450 48.530 151.460 ;
        RECT 47.740 151.435 48.635 151.450 ;
        RECT 47.720 151.420 48.635 151.435 ;
        RECT 47.700 151.410 48.635 151.420 ;
        RECT 47.675 151.400 48.635 151.410 ;
        RECT 47.605 151.370 48.635 151.400 ;
        RECT 47.585 151.340 48.635 151.370 ;
        RECT 47.565 151.310 48.635 151.340 ;
        RECT 47.535 151.285 48.635 151.310 ;
        RECT 47.500 151.250 48.635 151.285 ;
        RECT 47.470 151.245 48.635 151.250 ;
        RECT 47.470 151.240 47.860 151.245 ;
        RECT 47.470 151.230 47.835 151.240 ;
        RECT 47.470 151.225 47.820 151.230 ;
        RECT 47.470 151.220 47.805 151.225 ;
        RECT 46.845 151.215 47.805 151.220 ;
        RECT 46.845 151.205 47.795 151.215 ;
        RECT 46.845 151.200 47.785 151.205 ;
        RECT 46.845 151.190 47.775 151.200 ;
        RECT 46.845 151.180 47.770 151.190 ;
        RECT 46.845 151.175 47.765 151.180 ;
        RECT 46.845 151.160 47.755 151.175 ;
        RECT 46.845 151.145 47.750 151.160 ;
        RECT 46.845 151.120 47.740 151.145 ;
        RECT 46.845 151.050 47.735 151.120 ;
        RECT 43.165 149.945 46.675 150.715 ;
        RECT 46.845 150.495 47.395 150.880 ;
        RECT 47.565 150.325 47.735 151.050 ;
        RECT 46.845 150.155 47.735 150.325 ;
        RECT 47.905 150.650 48.235 151.075 ;
        RECT 48.405 150.850 48.635 151.245 ;
        RECT 47.905 150.165 48.125 150.650 ;
        RECT 48.805 150.595 48.975 151.625 ;
        RECT 48.295 149.945 48.545 150.485 ;
        RECT 48.715 150.115 48.975 150.595 ;
        RECT 50.730 150.490 51.070 151.320 ;
        RECT 52.550 150.810 52.900 152.060 ;
        RECT 54.675 151.525 55.005 152.310 ;
        RECT 54.675 151.355 55.355 151.525 ;
        RECT 55.535 151.355 55.865 152.495 ;
        RECT 54.665 150.935 55.015 151.185 ;
        RECT 55.185 150.755 55.355 151.355 ;
        RECT 56.045 151.330 56.335 152.495 ;
        RECT 56.505 151.940 57.110 152.495 ;
        RECT 57.285 151.985 57.765 152.325 ;
        RECT 57.935 151.950 58.190 152.495 ;
        RECT 56.505 151.840 57.120 151.940 ;
        RECT 56.935 151.815 57.120 151.840 ;
        RECT 56.505 151.220 56.765 151.670 ;
        RECT 56.935 151.570 57.265 151.815 ;
        RECT 57.435 151.495 58.190 151.745 ;
        RECT 58.360 151.625 58.635 152.325 ;
        RECT 58.895 151.825 59.065 152.325 ;
        RECT 59.235 151.995 59.565 152.495 ;
        RECT 58.895 151.655 59.560 151.825 ;
        RECT 57.420 151.460 58.190 151.495 ;
        RECT 57.405 151.450 58.190 151.460 ;
        RECT 57.400 151.435 58.295 151.450 ;
        RECT 57.380 151.420 58.295 151.435 ;
        RECT 57.360 151.410 58.295 151.420 ;
        RECT 57.335 151.400 58.295 151.410 ;
        RECT 57.265 151.370 58.295 151.400 ;
        RECT 57.245 151.340 58.295 151.370 ;
        RECT 57.225 151.310 58.295 151.340 ;
        RECT 57.195 151.285 58.295 151.310 ;
        RECT 57.160 151.250 58.295 151.285 ;
        RECT 57.130 151.245 58.295 151.250 ;
        RECT 57.130 151.240 57.520 151.245 ;
        RECT 57.130 151.230 57.495 151.240 ;
        RECT 57.130 151.225 57.480 151.230 ;
        RECT 57.130 151.220 57.465 151.225 ;
        RECT 56.505 151.215 57.465 151.220 ;
        RECT 56.505 151.205 57.455 151.215 ;
        RECT 56.505 151.200 57.445 151.205 ;
        RECT 56.505 151.190 57.435 151.200 ;
        RECT 55.525 150.935 55.875 151.185 ;
        RECT 56.505 151.180 57.430 151.190 ;
        RECT 56.505 151.175 57.425 151.180 ;
        RECT 56.505 151.160 57.415 151.175 ;
        RECT 56.505 151.145 57.410 151.160 ;
        RECT 56.505 151.120 57.400 151.145 ;
        RECT 56.505 151.050 57.395 151.120 ;
        RECT 49.145 149.945 54.490 150.490 ;
        RECT 54.685 149.945 54.925 150.755 ;
        RECT 55.095 150.115 55.425 150.755 ;
        RECT 55.595 149.945 55.865 150.755 ;
        RECT 56.045 149.945 56.335 150.670 ;
        RECT 56.505 150.495 57.055 150.880 ;
        RECT 57.225 150.325 57.395 151.050 ;
        RECT 56.505 150.155 57.395 150.325 ;
        RECT 57.565 150.650 57.895 151.075 ;
        RECT 58.065 150.850 58.295 151.245 ;
        RECT 57.565 150.165 57.785 150.650 ;
        RECT 58.465 150.595 58.635 151.625 ;
        RECT 58.810 150.835 59.160 151.485 ;
        RECT 59.330 150.665 59.560 151.655 ;
        RECT 57.955 149.945 58.205 150.485 ;
        RECT 58.375 150.115 58.635 150.595 ;
        RECT 58.895 150.495 59.560 150.665 ;
        RECT 58.895 150.205 59.065 150.495 ;
        RECT 59.235 149.945 59.565 150.325 ;
        RECT 59.735 150.205 59.920 152.325 ;
        RECT 60.160 152.035 60.425 152.495 ;
        RECT 60.595 151.900 60.845 152.325 ;
        RECT 61.055 152.050 62.160 152.220 ;
        RECT 60.540 151.770 60.845 151.900 ;
        RECT 60.090 150.575 60.370 151.525 ;
        RECT 60.540 150.665 60.710 151.770 ;
        RECT 60.880 150.985 61.120 151.580 ;
        RECT 61.290 151.515 61.820 151.880 ;
        RECT 61.290 150.815 61.460 151.515 ;
        RECT 61.990 151.435 62.160 152.050 ;
        RECT 62.330 151.695 62.500 152.495 ;
        RECT 62.670 151.995 62.920 152.325 ;
        RECT 63.145 152.025 64.030 152.195 ;
        RECT 61.990 151.345 62.500 151.435 ;
        RECT 60.540 150.535 60.765 150.665 ;
        RECT 60.935 150.595 61.460 150.815 ;
        RECT 61.630 151.175 62.500 151.345 ;
        RECT 60.175 149.945 60.425 150.405 ;
        RECT 60.595 150.395 60.765 150.535 ;
        RECT 61.630 150.395 61.800 151.175 ;
        RECT 62.330 151.105 62.500 151.175 ;
        RECT 62.010 150.925 62.210 150.955 ;
        RECT 62.670 150.925 62.840 151.995 ;
        RECT 63.010 151.105 63.200 151.825 ;
        RECT 62.010 150.625 62.840 150.925 ;
        RECT 63.370 150.895 63.690 151.855 ;
        RECT 60.595 150.225 60.930 150.395 ;
        RECT 61.125 150.225 61.800 150.395 ;
        RECT 62.120 149.945 62.490 150.445 ;
        RECT 62.670 150.395 62.840 150.625 ;
        RECT 63.225 150.565 63.690 150.895 ;
        RECT 63.860 151.185 64.030 152.025 ;
        RECT 64.210 151.995 64.525 152.495 ;
        RECT 64.755 151.765 65.095 152.325 ;
        RECT 64.200 151.390 65.095 151.765 ;
        RECT 65.265 151.485 65.435 152.495 ;
        RECT 64.905 151.185 65.095 151.390 ;
        RECT 65.605 151.435 65.935 152.280 ;
        RECT 65.605 151.355 65.995 151.435 ;
        RECT 65.780 151.305 65.995 151.355 ;
        RECT 63.860 150.855 64.735 151.185 ;
        RECT 64.905 150.855 65.655 151.185 ;
        RECT 63.860 150.395 64.030 150.855 ;
        RECT 64.905 150.685 65.105 150.855 ;
        RECT 65.825 150.725 65.995 151.305 ;
        RECT 65.770 150.685 65.995 150.725 ;
        RECT 62.670 150.225 63.075 150.395 ;
        RECT 63.245 150.225 64.030 150.395 ;
        RECT 64.305 149.945 64.515 150.475 ;
        RECT 64.775 150.160 65.105 150.685 ;
        RECT 65.615 150.600 65.995 150.685 ;
        RECT 65.275 149.945 65.445 150.555 ;
        RECT 65.615 150.165 65.945 150.600 ;
        RECT 66.175 150.125 66.435 152.315 ;
        RECT 66.605 151.765 66.945 152.495 ;
        RECT 67.125 151.585 67.395 152.315 ;
        RECT 66.625 151.365 67.395 151.585 ;
        RECT 67.575 151.605 67.805 152.315 ;
        RECT 67.975 151.785 68.305 152.495 ;
        RECT 68.475 151.605 68.735 152.315 ;
        RECT 67.575 151.365 68.735 151.605 ;
        RECT 66.625 150.695 66.915 151.365 ;
        RECT 68.925 151.355 69.185 152.495 ;
        RECT 69.355 151.345 69.685 152.325 ;
        RECT 69.855 151.355 70.135 152.495 ;
        RECT 70.765 151.355 71.150 152.325 ;
        RECT 71.320 152.035 71.645 152.495 ;
        RECT 72.165 151.865 72.445 152.325 ;
        RECT 71.320 151.645 72.445 151.865 ;
        RECT 67.095 150.875 67.560 151.185 ;
        RECT 67.740 150.875 68.265 151.185 ;
        RECT 66.625 150.495 67.855 150.695 ;
        RECT 66.695 149.945 67.365 150.315 ;
        RECT 67.545 150.125 67.855 150.495 ;
        RECT 68.035 150.235 68.265 150.875 ;
        RECT 68.445 150.855 68.745 151.185 ;
        RECT 68.945 150.935 69.280 151.185 ;
        RECT 69.450 150.745 69.620 151.345 ;
        RECT 69.790 150.915 70.125 151.185 ;
        RECT 68.445 149.945 68.735 150.675 ;
        RECT 68.925 150.115 69.620 150.745 ;
        RECT 69.825 149.945 70.135 150.745 ;
        RECT 70.765 150.685 71.045 151.355 ;
        RECT 71.320 151.185 71.770 151.645 ;
        RECT 72.635 151.475 73.035 152.325 ;
        RECT 73.435 152.035 73.705 152.495 ;
        RECT 73.875 151.865 74.160 152.325 ;
        RECT 71.215 150.855 71.770 151.185 ;
        RECT 71.940 150.915 73.035 151.475 ;
        RECT 71.320 150.745 71.770 150.855 ;
        RECT 70.765 150.115 71.150 150.685 ;
        RECT 71.320 150.575 72.445 150.745 ;
        RECT 71.320 149.945 71.645 150.405 ;
        RECT 72.165 150.115 72.445 150.575 ;
        RECT 72.635 150.115 73.035 150.915 ;
        RECT 73.205 151.645 74.160 151.865 ;
        RECT 74.535 151.825 74.705 152.325 ;
        RECT 74.875 151.995 75.205 152.495 ;
        RECT 74.535 151.655 75.200 151.825 ;
        RECT 73.205 150.745 73.415 151.645 ;
        RECT 73.585 150.915 74.275 151.475 ;
        RECT 74.450 150.835 74.800 151.485 ;
        RECT 73.205 150.575 74.160 150.745 ;
        RECT 74.970 150.665 75.200 151.655 ;
        RECT 73.435 149.945 73.705 150.405 ;
        RECT 73.875 150.115 74.160 150.575 ;
        RECT 74.535 150.495 75.200 150.665 ;
        RECT 74.535 150.205 74.705 150.495 ;
        RECT 74.875 149.945 75.205 150.325 ;
        RECT 75.375 150.205 75.560 152.325 ;
        RECT 75.800 152.035 76.065 152.495 ;
        RECT 76.235 151.900 76.485 152.325 ;
        RECT 76.695 152.050 77.800 152.220 ;
        RECT 76.180 151.770 76.485 151.900 ;
        RECT 75.730 150.575 76.010 151.525 ;
        RECT 76.180 150.665 76.350 151.770 ;
        RECT 76.520 150.985 76.760 151.580 ;
        RECT 76.930 151.515 77.460 151.880 ;
        RECT 76.930 150.815 77.100 151.515 ;
        RECT 77.630 151.435 77.800 152.050 ;
        RECT 77.970 151.695 78.140 152.495 ;
        RECT 78.310 151.995 78.560 152.325 ;
        RECT 78.785 152.025 79.670 152.195 ;
        RECT 77.630 151.345 78.140 151.435 ;
        RECT 76.180 150.535 76.405 150.665 ;
        RECT 76.575 150.595 77.100 150.815 ;
        RECT 77.270 151.175 78.140 151.345 ;
        RECT 75.815 149.945 76.065 150.405 ;
        RECT 76.235 150.395 76.405 150.535 ;
        RECT 77.270 150.395 77.440 151.175 ;
        RECT 77.970 151.105 78.140 151.175 ;
        RECT 77.650 150.925 77.850 150.955 ;
        RECT 78.310 150.925 78.480 151.995 ;
        RECT 78.650 151.105 78.840 151.825 ;
        RECT 77.650 150.625 78.480 150.925 ;
        RECT 79.010 150.895 79.330 151.855 ;
        RECT 76.235 150.225 76.570 150.395 ;
        RECT 76.765 150.225 77.440 150.395 ;
        RECT 77.760 149.945 78.130 150.445 ;
        RECT 78.310 150.395 78.480 150.625 ;
        RECT 78.865 150.565 79.330 150.895 ;
        RECT 79.500 151.185 79.670 152.025 ;
        RECT 79.850 151.995 80.165 152.495 ;
        RECT 80.395 151.765 80.735 152.325 ;
        RECT 79.840 151.390 80.735 151.765 ;
        RECT 80.905 151.485 81.075 152.495 ;
        RECT 80.545 151.185 80.735 151.390 ;
        RECT 81.245 151.435 81.575 152.280 ;
        RECT 81.245 151.355 81.635 151.435 ;
        RECT 81.420 151.305 81.635 151.355 ;
        RECT 81.805 151.330 82.095 152.495 ;
        RECT 82.275 151.525 82.605 152.310 ;
        RECT 82.275 151.355 82.955 151.525 ;
        RECT 83.135 151.355 83.465 152.495 ;
        RECT 83.645 151.405 85.315 152.495 ;
        RECT 79.500 150.855 80.375 151.185 ;
        RECT 80.545 150.855 81.295 151.185 ;
        RECT 79.500 150.395 79.670 150.855 ;
        RECT 80.545 150.685 80.745 150.855 ;
        RECT 81.465 150.725 81.635 151.305 ;
        RECT 82.265 150.935 82.615 151.185 ;
        RECT 82.785 150.755 82.955 151.355 ;
        RECT 83.125 150.935 83.475 151.185 ;
        RECT 81.410 150.685 81.635 150.725 ;
        RECT 78.310 150.225 78.715 150.395 ;
        RECT 78.885 150.225 79.670 150.395 ;
        RECT 79.945 149.945 80.155 150.475 ;
        RECT 80.415 150.160 80.745 150.685 ;
        RECT 81.255 150.600 81.635 150.685 ;
        RECT 80.915 149.945 81.085 150.555 ;
        RECT 81.255 150.165 81.585 150.600 ;
        RECT 81.805 149.945 82.095 150.670 ;
        RECT 82.285 149.945 82.525 150.755 ;
        RECT 82.695 150.115 83.025 150.755 ;
        RECT 83.195 149.945 83.465 150.755 ;
        RECT 83.645 150.715 84.395 151.235 ;
        RECT 84.565 150.885 85.315 151.405 ;
        RECT 85.495 151.545 85.770 152.315 ;
        RECT 85.940 151.885 86.270 152.315 ;
        RECT 86.440 152.055 86.635 152.495 ;
        RECT 86.815 151.885 87.145 152.315 ;
        RECT 85.940 151.715 87.145 151.885 ;
        RECT 85.495 151.355 86.080 151.545 ;
        RECT 86.250 151.385 87.145 151.715 ;
        RECT 83.645 149.945 85.315 150.715 ;
        RECT 85.495 150.535 85.735 151.185 ;
        RECT 85.905 150.685 86.080 151.355 ;
        RECT 87.785 151.290 88.075 152.495 ;
        RECT 88.245 151.355 88.520 152.325 ;
        RECT 88.730 151.695 89.010 152.495 ;
        RECT 89.180 151.985 90.375 152.275 ;
        RECT 90.635 151.825 90.805 152.325 ;
        RECT 90.975 151.995 91.305 152.495 ;
        RECT 89.190 151.645 90.355 151.815 ;
        RECT 90.635 151.655 91.300 151.825 ;
        RECT 89.190 151.525 89.360 151.645 ;
        RECT 88.690 151.355 89.360 151.525 ;
        RECT 86.250 150.855 86.665 151.185 ;
        RECT 86.845 150.855 87.140 151.185 ;
        RECT 85.905 150.505 86.235 150.685 ;
        RECT 85.510 149.945 85.840 150.335 ;
        RECT 86.010 150.125 86.235 150.505 ;
        RECT 86.435 150.235 86.665 150.855 ;
        RECT 86.845 149.945 87.145 150.675 ;
        RECT 87.785 149.945 88.075 150.775 ;
        RECT 88.245 150.620 88.415 151.355 ;
        RECT 88.690 151.185 88.860 151.355 ;
        RECT 89.630 151.185 89.855 151.475 ;
        RECT 90.025 151.355 90.355 151.645 ;
        RECT 88.585 150.855 88.860 151.185 ;
        RECT 89.030 150.855 89.855 151.185 ;
        RECT 90.025 150.855 90.375 151.185 ;
        RECT 88.690 150.685 88.860 150.855 ;
        RECT 90.550 150.835 90.900 151.485 ;
        RECT 88.245 150.275 88.520 150.620 ;
        RECT 88.690 150.515 90.355 150.685 ;
        RECT 91.070 150.665 91.300 151.655 ;
        RECT 88.710 149.945 89.090 150.345 ;
        RECT 89.260 150.165 89.430 150.515 ;
        RECT 89.600 149.945 89.930 150.345 ;
        RECT 90.100 150.165 90.355 150.515 ;
        RECT 90.635 150.495 91.300 150.665 ;
        RECT 90.635 150.205 90.805 150.495 ;
        RECT 90.975 149.945 91.305 150.325 ;
        RECT 91.475 150.205 91.660 152.325 ;
        RECT 91.900 152.035 92.165 152.495 ;
        RECT 92.335 151.900 92.585 152.325 ;
        RECT 92.795 152.050 93.900 152.220 ;
        RECT 92.280 151.770 92.585 151.900 ;
        RECT 91.830 150.575 92.110 151.525 ;
        RECT 92.280 150.665 92.450 151.770 ;
        RECT 92.620 150.985 92.860 151.580 ;
        RECT 93.030 151.515 93.560 151.880 ;
        RECT 93.030 150.815 93.200 151.515 ;
        RECT 93.730 151.435 93.900 152.050 ;
        RECT 94.070 151.695 94.240 152.495 ;
        RECT 94.410 151.995 94.660 152.325 ;
        RECT 94.885 152.025 95.770 152.195 ;
        RECT 93.730 151.345 94.240 151.435 ;
        RECT 92.280 150.535 92.505 150.665 ;
        RECT 92.675 150.595 93.200 150.815 ;
        RECT 93.370 151.175 94.240 151.345 ;
        RECT 91.915 149.945 92.165 150.405 ;
        RECT 92.335 150.395 92.505 150.535 ;
        RECT 93.370 150.395 93.540 151.175 ;
        RECT 94.070 151.105 94.240 151.175 ;
        RECT 93.750 150.925 93.950 150.955 ;
        RECT 94.410 150.925 94.580 151.995 ;
        RECT 94.750 151.105 94.940 151.825 ;
        RECT 93.750 150.625 94.580 150.925 ;
        RECT 95.110 150.895 95.430 151.855 ;
        RECT 92.335 150.225 92.670 150.395 ;
        RECT 92.865 150.225 93.540 150.395 ;
        RECT 93.860 149.945 94.230 150.445 ;
        RECT 94.410 150.395 94.580 150.625 ;
        RECT 94.965 150.565 95.430 150.895 ;
        RECT 95.600 151.185 95.770 152.025 ;
        RECT 95.950 151.995 96.265 152.495 ;
        RECT 96.495 151.765 96.835 152.325 ;
        RECT 95.940 151.390 96.835 151.765 ;
        RECT 97.005 151.485 97.175 152.495 ;
        RECT 96.645 151.185 96.835 151.390 ;
        RECT 97.345 151.435 97.675 152.280 ;
        RECT 98.885 151.435 99.215 152.280 ;
        RECT 99.385 151.485 99.555 152.495 ;
        RECT 99.725 151.765 100.065 152.325 ;
        RECT 100.295 151.995 100.610 152.495 ;
        RECT 100.790 152.025 101.675 152.195 ;
        RECT 97.345 151.355 97.735 151.435 ;
        RECT 97.520 151.305 97.735 151.355 ;
        RECT 95.600 150.855 96.475 151.185 ;
        RECT 96.645 150.855 97.395 151.185 ;
        RECT 95.600 150.395 95.770 150.855 ;
        RECT 96.645 150.685 96.845 150.855 ;
        RECT 97.565 150.725 97.735 151.305 ;
        RECT 97.510 150.685 97.735 150.725 ;
        RECT 94.410 150.225 94.815 150.395 ;
        RECT 94.985 150.225 95.770 150.395 ;
        RECT 96.045 149.945 96.255 150.475 ;
        RECT 96.515 150.160 96.845 150.685 ;
        RECT 97.355 150.600 97.735 150.685 ;
        RECT 98.825 151.355 99.215 151.435 ;
        RECT 99.725 151.390 100.620 151.765 ;
        RECT 98.825 151.305 99.040 151.355 ;
        RECT 98.825 150.725 98.995 151.305 ;
        RECT 99.725 151.185 99.915 151.390 ;
        RECT 100.790 151.185 100.960 152.025 ;
        RECT 101.900 151.995 102.150 152.325 ;
        RECT 99.165 150.855 99.915 151.185 ;
        RECT 100.085 150.855 100.960 151.185 ;
        RECT 98.825 150.685 99.050 150.725 ;
        RECT 99.715 150.685 99.915 150.855 ;
        RECT 98.825 150.600 99.205 150.685 ;
        RECT 97.015 149.945 97.185 150.555 ;
        RECT 97.355 150.165 97.685 150.600 ;
        RECT 98.875 150.165 99.205 150.600 ;
        RECT 99.375 149.945 99.545 150.555 ;
        RECT 99.715 150.160 100.045 150.685 ;
        RECT 100.305 149.945 100.515 150.475 ;
        RECT 100.790 150.395 100.960 150.855 ;
        RECT 101.130 150.895 101.450 151.855 ;
        RECT 101.620 151.105 101.810 151.825 ;
        RECT 101.980 150.925 102.150 151.995 ;
        RECT 102.320 151.695 102.490 152.495 ;
        RECT 102.660 152.050 103.765 152.220 ;
        RECT 102.660 151.435 102.830 152.050 ;
        RECT 103.975 151.900 104.225 152.325 ;
        RECT 104.395 152.035 104.660 152.495 ;
        RECT 103.000 151.515 103.530 151.880 ;
        RECT 103.975 151.770 104.280 151.900 ;
        RECT 102.320 151.345 102.830 151.435 ;
        RECT 102.320 151.175 103.190 151.345 ;
        RECT 102.320 151.105 102.490 151.175 ;
        RECT 102.610 150.925 102.810 150.955 ;
        RECT 101.130 150.565 101.595 150.895 ;
        RECT 101.980 150.625 102.810 150.925 ;
        RECT 101.980 150.395 102.150 150.625 ;
        RECT 100.790 150.225 101.575 150.395 ;
        RECT 101.745 150.225 102.150 150.395 ;
        RECT 102.330 149.945 102.700 150.445 ;
        RECT 103.020 150.395 103.190 151.175 ;
        RECT 103.360 150.815 103.530 151.515 ;
        RECT 103.700 150.985 103.940 151.580 ;
        RECT 103.360 150.595 103.885 150.815 ;
        RECT 104.110 150.665 104.280 151.770 ;
        RECT 104.055 150.535 104.280 150.665 ;
        RECT 104.450 150.575 104.730 151.525 ;
        RECT 104.055 150.395 104.225 150.535 ;
        RECT 103.020 150.225 103.695 150.395 ;
        RECT 103.890 150.225 104.225 150.395 ;
        RECT 104.395 149.945 104.645 150.405 ;
        RECT 104.900 150.205 105.085 152.325 ;
        RECT 105.255 151.995 105.585 152.495 ;
        RECT 105.755 151.825 105.925 152.325 ;
        RECT 105.260 151.655 105.925 151.825 ;
        RECT 105.260 150.665 105.490 151.655 ;
        RECT 105.660 150.835 106.010 151.485 ;
        RECT 106.185 151.405 107.395 152.495 ;
        RECT 106.185 150.695 106.705 151.235 ;
        RECT 106.875 150.865 107.395 151.405 ;
        RECT 107.565 151.330 107.855 152.495 ;
        RECT 108.030 151.355 108.365 152.325 ;
        RECT 108.535 151.355 108.705 152.495 ;
        RECT 108.875 152.155 110.905 152.325 ;
        RECT 105.260 150.495 105.925 150.665 ;
        RECT 105.255 149.945 105.585 150.325 ;
        RECT 105.755 150.205 105.925 150.495 ;
        RECT 106.185 149.945 107.395 150.695 ;
        RECT 108.030 150.685 108.200 151.355 ;
        RECT 108.875 151.185 109.045 152.155 ;
        RECT 108.370 150.855 108.625 151.185 ;
        RECT 108.850 150.855 109.045 151.185 ;
        RECT 109.215 151.815 110.340 151.985 ;
        RECT 108.455 150.685 108.625 150.855 ;
        RECT 109.215 150.685 109.385 151.815 ;
        RECT 107.565 149.945 107.855 150.670 ;
        RECT 108.030 150.115 108.285 150.685 ;
        RECT 108.455 150.515 109.385 150.685 ;
        RECT 109.555 151.475 110.565 151.645 ;
        RECT 109.555 150.675 109.725 151.475 ;
        RECT 109.930 151.135 110.205 151.275 ;
        RECT 109.925 150.965 110.205 151.135 ;
        RECT 109.210 150.480 109.385 150.515 ;
        RECT 108.455 149.945 108.785 150.345 ;
        RECT 109.210 150.115 109.740 150.480 ;
        RECT 109.930 150.115 110.205 150.965 ;
        RECT 110.375 150.115 110.565 151.475 ;
        RECT 110.735 151.490 110.905 152.155 ;
        RECT 111.075 151.735 111.245 152.495 ;
        RECT 111.480 151.735 111.995 152.145 ;
        RECT 110.735 151.300 111.485 151.490 ;
        RECT 111.655 150.925 111.995 151.735 ;
        RECT 112.175 151.525 112.505 152.310 ;
        RECT 112.175 151.355 112.855 151.525 ;
        RECT 113.035 151.355 113.365 152.495 ;
        RECT 113.545 152.060 118.890 152.495 ;
        RECT 112.165 150.935 112.515 151.185 ;
        RECT 110.765 150.755 111.995 150.925 ;
        RECT 112.685 150.755 112.855 151.355 ;
        RECT 113.025 150.935 113.375 151.185 ;
        RECT 110.745 149.945 111.255 150.480 ;
        RECT 111.475 150.150 111.720 150.755 ;
        RECT 112.185 149.945 112.425 150.755 ;
        RECT 112.595 150.115 112.925 150.755 ;
        RECT 113.095 149.945 113.365 150.755 ;
        RECT 115.130 150.490 115.470 151.320 ;
        RECT 116.950 150.810 117.300 152.060 ;
        RECT 119.065 151.355 119.345 152.495 ;
        RECT 119.515 151.345 119.845 152.325 ;
        RECT 120.015 151.355 120.275 152.495 ;
        RECT 120.445 151.405 122.115 152.495 ;
        RECT 119.075 150.915 119.410 151.185 ;
        RECT 119.580 150.745 119.750 151.345 ;
        RECT 119.920 150.935 120.255 151.185 ;
        RECT 113.545 149.945 118.890 150.490 ;
        RECT 119.065 149.945 119.375 150.745 ;
        RECT 119.580 150.115 120.275 150.745 ;
        RECT 120.445 150.715 121.195 151.235 ;
        RECT 121.365 150.885 122.115 151.405 ;
        RECT 122.785 151.355 123.015 152.495 ;
        RECT 123.185 151.345 123.515 152.325 ;
        RECT 123.685 151.355 123.895 152.495 ;
        RECT 125.345 151.855 125.675 152.285 ;
        RECT 125.220 151.685 125.675 151.855 ;
        RECT 125.855 151.855 126.105 152.275 ;
        RECT 126.335 152.025 126.665 152.495 ;
        RECT 126.895 151.855 127.145 152.275 ;
        RECT 125.855 151.685 127.145 151.855 ;
        RECT 122.765 150.935 123.095 151.185 ;
        RECT 120.445 149.945 122.115 150.715 ;
        RECT 122.785 149.945 123.015 150.765 ;
        RECT 123.265 150.745 123.515 151.345 ;
        RECT 123.185 150.115 123.515 150.745 ;
        RECT 123.685 149.945 123.895 150.765 ;
        RECT 125.220 150.685 125.390 151.685 ;
        RECT 125.560 150.855 125.805 151.515 ;
        RECT 126.020 150.855 126.285 151.515 ;
        RECT 126.480 150.855 126.765 151.515 ;
        RECT 126.940 151.185 127.155 151.515 ;
        RECT 127.335 151.355 127.585 152.495 ;
        RECT 127.755 151.435 128.085 152.285 ;
        RECT 126.940 150.855 127.245 151.185 ;
        RECT 127.415 150.855 127.725 151.185 ;
        RECT 127.415 150.685 127.585 150.855 ;
        RECT 125.220 150.515 127.585 150.685 ;
        RECT 127.895 150.670 128.085 151.435 ;
        RECT 128.265 151.355 128.525 152.495 ;
        RECT 128.695 151.345 129.025 152.325 ;
        RECT 129.195 151.355 129.475 152.495 ;
        RECT 129.645 151.405 133.155 152.495 ;
        RECT 128.285 150.935 128.620 151.185 ;
        RECT 128.790 150.795 128.960 151.345 ;
        RECT 129.130 150.915 129.465 151.185 ;
        RECT 128.785 150.745 128.960 150.795 ;
        RECT 125.375 149.945 125.705 150.345 ;
        RECT 125.875 150.175 126.205 150.515 ;
        RECT 127.255 149.945 127.585 150.345 ;
        RECT 127.755 150.160 128.085 150.670 ;
        RECT 128.265 150.115 128.960 150.745 ;
        RECT 129.165 149.945 129.475 150.745 ;
        RECT 129.645 150.715 131.295 151.235 ;
        RECT 131.465 150.885 133.155 151.405 ;
        RECT 133.325 151.330 133.615 152.495 ;
        RECT 133.875 151.825 134.045 152.325 ;
        RECT 134.215 151.995 134.545 152.495 ;
        RECT 133.875 151.655 134.540 151.825 ;
        RECT 133.790 150.835 134.140 151.485 ;
        RECT 129.645 149.945 133.155 150.715 ;
        RECT 133.325 149.945 133.615 150.670 ;
        RECT 134.310 150.665 134.540 151.655 ;
        RECT 133.875 150.495 134.540 150.665 ;
        RECT 133.875 150.205 134.045 150.495 ;
        RECT 134.215 149.945 134.545 150.325 ;
        RECT 134.715 150.205 134.900 152.325 ;
        RECT 135.140 152.035 135.405 152.495 ;
        RECT 135.575 151.900 135.825 152.325 ;
        RECT 136.035 152.050 137.140 152.220 ;
        RECT 135.520 151.770 135.825 151.900 ;
        RECT 135.070 150.575 135.350 151.525 ;
        RECT 135.520 150.665 135.690 151.770 ;
        RECT 135.860 150.985 136.100 151.580 ;
        RECT 136.270 151.515 136.800 151.880 ;
        RECT 136.270 150.815 136.440 151.515 ;
        RECT 136.970 151.435 137.140 152.050 ;
        RECT 137.310 151.695 137.480 152.495 ;
        RECT 137.650 151.995 137.900 152.325 ;
        RECT 138.125 152.025 139.010 152.195 ;
        RECT 136.970 151.345 137.480 151.435 ;
        RECT 135.520 150.535 135.745 150.665 ;
        RECT 135.915 150.595 136.440 150.815 ;
        RECT 136.610 151.175 137.480 151.345 ;
        RECT 135.155 149.945 135.405 150.405 ;
        RECT 135.575 150.395 135.745 150.535 ;
        RECT 136.610 150.395 136.780 151.175 ;
        RECT 137.310 151.105 137.480 151.175 ;
        RECT 136.990 150.925 137.190 150.955 ;
        RECT 137.650 150.925 137.820 151.995 ;
        RECT 137.990 151.105 138.180 151.825 ;
        RECT 136.990 150.625 137.820 150.925 ;
        RECT 138.350 150.895 138.670 151.855 ;
        RECT 135.575 150.225 135.910 150.395 ;
        RECT 136.105 150.225 136.780 150.395 ;
        RECT 137.100 149.945 137.470 150.445 ;
        RECT 137.650 150.395 137.820 150.625 ;
        RECT 138.205 150.565 138.670 150.895 ;
        RECT 138.840 151.185 139.010 152.025 ;
        RECT 139.190 151.995 139.505 152.495 ;
        RECT 139.735 151.765 140.075 152.325 ;
        RECT 139.180 151.390 140.075 151.765 ;
        RECT 140.245 151.485 140.415 152.495 ;
        RECT 139.885 151.185 140.075 151.390 ;
        RECT 140.585 151.435 140.915 152.280 ;
        RECT 140.585 151.355 140.975 151.435 ;
        RECT 140.760 151.305 140.975 151.355 ;
        RECT 138.840 150.855 139.715 151.185 ;
        RECT 139.885 150.855 140.635 151.185 ;
        RECT 138.840 150.395 139.010 150.855 ;
        RECT 139.885 150.685 140.085 150.855 ;
        RECT 140.805 150.725 140.975 151.305 ;
        RECT 140.750 150.685 140.975 150.725 ;
        RECT 137.650 150.225 138.055 150.395 ;
        RECT 138.225 150.225 139.010 150.395 ;
        RECT 139.285 149.945 139.495 150.475 ;
        RECT 139.755 150.160 140.085 150.685 ;
        RECT 140.595 150.600 140.975 150.685 ;
        RECT 141.150 151.355 141.485 152.325 ;
        RECT 141.655 151.355 141.825 152.495 ;
        RECT 141.995 152.155 144.025 152.325 ;
        RECT 141.150 150.685 141.320 151.355 ;
        RECT 141.995 151.185 142.165 152.155 ;
        RECT 141.490 150.855 141.745 151.185 ;
        RECT 141.970 150.855 142.165 151.185 ;
        RECT 142.335 151.815 143.460 151.985 ;
        RECT 141.575 150.685 141.745 150.855 ;
        RECT 142.335 150.685 142.505 151.815 ;
        RECT 140.255 149.945 140.425 150.555 ;
        RECT 140.595 150.165 140.925 150.600 ;
        RECT 141.150 150.115 141.405 150.685 ;
        RECT 141.575 150.515 142.505 150.685 ;
        RECT 142.675 151.475 143.685 151.645 ;
        RECT 142.675 150.675 142.845 151.475 ;
        RECT 142.330 150.480 142.505 150.515 ;
        RECT 141.575 149.945 141.905 150.345 ;
        RECT 142.330 150.115 142.860 150.480 ;
        RECT 143.050 150.455 143.325 151.275 ;
        RECT 143.045 150.285 143.325 150.455 ;
        RECT 143.050 150.115 143.325 150.285 ;
        RECT 143.495 150.115 143.685 151.475 ;
        RECT 143.855 151.490 144.025 152.155 ;
        RECT 144.195 151.735 144.365 152.495 ;
        RECT 144.600 151.735 145.115 152.145 ;
        RECT 143.855 151.300 144.605 151.490 ;
        RECT 144.775 150.925 145.115 151.735 ;
        RECT 143.885 150.755 145.115 150.925 ;
        RECT 145.745 151.405 146.955 152.495 ;
        RECT 145.745 150.865 146.265 151.405 ;
        RECT 143.865 149.945 144.375 150.480 ;
        RECT 144.595 150.150 144.840 150.755 ;
        RECT 146.435 150.695 146.955 151.235 ;
        RECT 145.745 149.945 146.955 150.695 ;
        RECT 17.320 149.775 147.040 149.945 ;
        RECT 17.405 149.025 18.615 149.775 ;
        RECT 18.785 149.230 24.130 149.775 ;
        RECT 24.305 149.230 29.650 149.775 ;
        RECT 17.405 148.485 17.925 149.025 ;
        RECT 18.095 148.315 18.615 148.855 ;
        RECT 20.370 148.400 20.710 149.230 ;
        RECT 17.405 147.225 18.615 148.315 ;
        RECT 22.190 147.660 22.540 148.910 ;
        RECT 25.890 148.400 26.230 149.230 ;
        RECT 30.745 148.975 31.440 149.605 ;
        RECT 31.645 148.975 31.955 149.775 ;
        RECT 32.125 149.395 33.015 149.565 ;
        RECT 31.265 148.925 31.440 148.975 ;
        RECT 27.710 147.660 28.060 148.910 ;
        RECT 30.765 148.535 31.100 148.785 ;
        RECT 31.270 148.375 31.440 148.925 ;
        RECT 32.125 148.840 32.675 149.225 ;
        RECT 31.610 148.535 31.945 148.805 ;
        RECT 32.845 148.670 33.015 149.395 ;
        RECT 32.125 148.600 33.015 148.670 ;
        RECT 33.185 149.095 33.405 149.555 ;
        RECT 33.575 149.235 33.825 149.775 ;
        RECT 33.995 149.125 34.255 149.605 ;
        RECT 33.185 149.070 33.435 149.095 ;
        RECT 33.185 148.645 33.515 149.070 ;
        RECT 32.125 148.575 33.020 148.600 ;
        RECT 32.125 148.560 33.030 148.575 ;
        RECT 32.125 148.545 33.035 148.560 ;
        RECT 32.125 148.540 33.045 148.545 ;
        RECT 32.125 148.530 33.050 148.540 ;
        RECT 32.125 148.520 33.055 148.530 ;
        RECT 32.125 148.515 33.065 148.520 ;
        RECT 32.125 148.505 33.075 148.515 ;
        RECT 32.125 148.500 33.085 148.505 ;
        RECT 18.785 147.225 24.130 147.660 ;
        RECT 24.305 147.225 29.650 147.660 ;
        RECT 30.745 147.225 31.005 148.365 ;
        RECT 31.175 147.395 31.505 148.375 ;
        RECT 31.675 147.225 31.955 148.365 ;
        RECT 32.125 148.050 32.385 148.500 ;
        RECT 32.750 148.495 33.085 148.500 ;
        RECT 32.750 148.490 33.100 148.495 ;
        RECT 32.750 148.480 33.115 148.490 ;
        RECT 32.750 148.475 33.140 148.480 ;
        RECT 33.685 148.475 33.915 148.870 ;
        RECT 32.750 148.470 33.915 148.475 ;
        RECT 32.780 148.435 33.915 148.470 ;
        RECT 32.815 148.410 33.915 148.435 ;
        RECT 32.845 148.380 33.915 148.410 ;
        RECT 32.865 148.350 33.915 148.380 ;
        RECT 32.885 148.320 33.915 148.350 ;
        RECT 32.955 148.310 33.915 148.320 ;
        RECT 32.980 148.300 33.915 148.310 ;
        RECT 33.000 148.285 33.915 148.300 ;
        RECT 33.020 148.270 33.915 148.285 ;
        RECT 33.025 148.260 33.810 148.270 ;
        RECT 33.040 148.225 33.810 148.260 ;
        RECT 32.555 147.905 32.885 148.150 ;
        RECT 33.055 147.975 33.810 148.225 ;
        RECT 34.085 148.095 34.255 149.125 ;
        RECT 34.515 149.225 34.685 149.515 ;
        RECT 34.855 149.395 35.185 149.775 ;
        RECT 34.515 149.055 35.180 149.225 ;
        RECT 34.430 148.235 34.780 148.885 ;
        RECT 32.555 147.880 32.740 147.905 ;
        RECT 32.125 147.780 32.740 147.880 ;
        RECT 32.125 147.225 32.730 147.780 ;
        RECT 32.905 147.395 33.385 147.735 ;
        RECT 33.555 147.225 33.810 147.770 ;
        RECT 33.980 147.395 34.255 148.095 ;
        RECT 34.950 148.065 35.180 149.055 ;
        RECT 34.515 147.895 35.180 148.065 ;
        RECT 34.515 147.395 34.685 147.895 ;
        RECT 34.855 147.225 35.185 147.725 ;
        RECT 35.355 147.395 35.540 149.515 ;
        RECT 35.795 149.315 36.045 149.775 ;
        RECT 36.215 149.325 36.550 149.495 ;
        RECT 36.745 149.325 37.420 149.495 ;
        RECT 36.215 149.185 36.385 149.325 ;
        RECT 35.710 148.195 35.990 149.145 ;
        RECT 36.160 149.055 36.385 149.185 ;
        RECT 36.160 147.950 36.330 149.055 ;
        RECT 36.555 148.905 37.080 149.125 ;
        RECT 36.500 148.140 36.740 148.735 ;
        RECT 36.910 148.205 37.080 148.905 ;
        RECT 37.250 148.545 37.420 149.325 ;
        RECT 37.740 149.275 38.110 149.775 ;
        RECT 38.290 149.325 38.695 149.495 ;
        RECT 38.865 149.325 39.650 149.495 ;
        RECT 38.290 149.095 38.460 149.325 ;
        RECT 37.630 148.795 38.460 149.095 ;
        RECT 38.845 148.825 39.310 149.155 ;
        RECT 37.630 148.765 37.830 148.795 ;
        RECT 37.950 148.545 38.120 148.615 ;
        RECT 37.250 148.375 38.120 148.545 ;
        RECT 37.610 148.285 38.120 148.375 ;
        RECT 36.160 147.820 36.465 147.950 ;
        RECT 36.910 147.840 37.440 148.205 ;
        RECT 35.780 147.225 36.045 147.685 ;
        RECT 36.215 147.395 36.465 147.820 ;
        RECT 37.610 147.670 37.780 148.285 ;
        RECT 36.675 147.500 37.780 147.670 ;
        RECT 37.950 147.225 38.120 148.025 ;
        RECT 38.290 147.725 38.460 148.795 ;
        RECT 38.630 147.895 38.820 148.615 ;
        RECT 38.990 147.865 39.310 148.825 ;
        RECT 39.480 148.865 39.650 149.325 ;
        RECT 39.925 149.245 40.135 149.775 ;
        RECT 40.395 149.035 40.725 149.560 ;
        RECT 40.895 149.165 41.065 149.775 ;
        RECT 41.235 149.120 41.565 149.555 ;
        RECT 41.235 149.035 41.615 149.120 ;
        RECT 40.525 148.865 40.725 149.035 ;
        RECT 41.390 148.995 41.615 149.035 ;
        RECT 39.480 148.535 40.355 148.865 ;
        RECT 40.525 148.535 41.275 148.865 ;
        RECT 38.290 147.395 38.540 147.725 ;
        RECT 39.480 147.695 39.650 148.535 ;
        RECT 40.525 148.330 40.715 148.535 ;
        RECT 41.445 148.415 41.615 148.995 ;
        RECT 41.785 149.025 42.995 149.775 ;
        RECT 43.165 149.050 43.455 149.775 ;
        RECT 41.785 148.485 42.305 149.025 ;
        RECT 43.625 149.005 45.295 149.775 ;
        RECT 41.400 148.365 41.615 148.415 ;
        RECT 39.820 147.955 40.715 148.330 ;
        RECT 41.225 148.285 41.615 148.365 ;
        RECT 42.475 148.315 42.995 148.855 ;
        RECT 43.625 148.485 44.375 149.005 ;
        RECT 38.765 147.525 39.650 147.695 ;
        RECT 39.830 147.225 40.145 147.725 ;
        RECT 40.375 147.395 40.715 147.955 ;
        RECT 40.885 147.225 41.055 148.235 ;
        RECT 41.225 147.440 41.555 148.285 ;
        RECT 41.785 147.225 42.995 148.315 ;
        RECT 43.165 147.225 43.455 148.390 ;
        RECT 44.545 148.315 45.295 148.835 ;
        RECT 43.625 147.225 45.295 148.315 ;
        RECT 45.465 147.395 45.745 149.495 ;
        RECT 45.975 149.315 46.145 149.775 ;
        RECT 46.415 149.385 47.665 149.565 ;
        RECT 46.800 149.145 47.165 149.215 ;
        RECT 45.915 148.965 47.165 149.145 ;
        RECT 47.335 149.165 47.665 149.385 ;
        RECT 47.835 149.335 48.005 149.775 ;
        RECT 48.175 149.165 48.515 149.580 ;
        RECT 47.335 148.995 48.515 149.165 ;
        RECT 48.685 149.025 49.895 149.775 ;
        RECT 50.155 149.125 50.325 149.605 ;
        RECT 50.495 149.295 50.825 149.775 ;
        RECT 51.050 149.355 52.585 149.605 ;
        RECT 51.050 149.125 51.220 149.355 ;
        RECT 45.915 148.365 46.190 148.965 ;
        RECT 46.360 148.535 46.715 148.785 ;
        RECT 46.910 148.755 47.375 148.785 ;
        RECT 46.905 148.585 47.375 148.755 ;
        RECT 46.910 148.535 47.375 148.585 ;
        RECT 47.545 148.535 47.875 148.785 ;
        RECT 48.050 148.585 48.515 148.785 ;
        RECT 47.695 148.415 47.875 148.535 ;
        RECT 48.685 148.485 49.205 149.025 ;
        RECT 50.155 148.955 51.220 149.125 ;
        RECT 45.915 148.155 47.525 148.365 ;
        RECT 47.695 148.245 48.025 148.415 ;
        RECT 47.115 148.055 47.525 148.155 ;
        RECT 45.935 147.225 46.720 147.985 ;
        RECT 47.115 147.395 47.500 148.055 ;
        RECT 47.825 147.455 48.025 148.245 ;
        RECT 48.195 147.225 48.515 148.405 ;
        RECT 49.375 148.315 49.895 148.855 ;
        RECT 51.400 148.785 51.680 149.185 ;
        RECT 50.070 148.575 50.420 148.785 ;
        RECT 50.590 148.585 51.035 148.785 ;
        RECT 51.205 148.585 51.680 148.785 ;
        RECT 51.950 148.785 52.235 149.185 ;
        RECT 52.415 149.125 52.585 149.355 ;
        RECT 52.755 149.295 53.085 149.775 ;
        RECT 53.300 149.275 53.555 149.605 ;
        RECT 53.370 149.195 53.555 149.275 ;
        RECT 52.415 148.955 53.215 149.125 ;
        RECT 51.950 148.585 52.280 148.785 ;
        RECT 52.450 148.585 52.815 148.785 ;
        RECT 53.045 148.405 53.215 148.955 ;
        RECT 48.685 147.225 49.895 148.315 ;
        RECT 50.155 148.235 53.215 148.405 ;
        RECT 50.155 147.395 50.325 148.235 ;
        RECT 53.385 148.075 53.555 149.195 ;
        RECT 53.755 149.045 54.055 149.775 ;
        RECT 54.235 148.865 54.465 149.485 ;
        RECT 54.665 149.215 54.890 149.595 ;
        RECT 55.060 149.385 55.390 149.775 ;
        RECT 54.665 149.035 54.995 149.215 ;
        RECT 53.760 148.535 54.055 148.865 ;
        RECT 54.235 148.535 54.650 148.865 ;
        RECT 54.820 148.365 54.995 149.035 ;
        RECT 55.165 148.535 55.405 149.185 ;
        RECT 56.595 149.125 56.765 149.605 ;
        RECT 56.935 149.295 57.265 149.775 ;
        RECT 57.490 149.355 59.025 149.605 ;
        RECT 57.490 149.125 57.660 149.355 ;
        RECT 56.595 148.955 57.660 149.125 ;
        RECT 57.840 148.785 58.120 149.185 ;
        RECT 56.510 148.575 56.860 148.785 ;
        RECT 57.030 148.585 57.475 148.785 ;
        RECT 57.645 148.585 58.120 148.785 ;
        RECT 58.390 148.785 58.675 149.185 ;
        RECT 58.855 149.125 59.025 149.355 ;
        RECT 59.195 149.295 59.525 149.775 ;
        RECT 59.740 149.275 59.995 149.605 ;
        RECT 59.810 149.195 59.995 149.275 ;
        RECT 58.855 148.955 59.655 149.125 ;
        RECT 58.390 148.585 58.720 148.785 ;
        RECT 58.890 148.755 59.255 148.785 ;
        RECT 58.890 148.585 59.265 148.755 ;
        RECT 59.485 148.405 59.655 148.955 ;
        RECT 53.345 148.065 53.555 148.075 ;
        RECT 50.495 147.565 50.825 148.065 ;
        RECT 50.995 147.825 52.630 148.065 ;
        RECT 50.995 147.735 51.225 147.825 ;
        RECT 51.335 147.565 51.665 147.605 ;
        RECT 50.495 147.395 51.665 147.565 ;
        RECT 51.855 147.225 52.210 147.645 ;
        RECT 52.380 147.395 52.630 147.825 ;
        RECT 52.800 147.225 53.130 147.985 ;
        RECT 53.300 147.395 53.555 148.065 ;
        RECT 53.755 148.005 54.650 148.335 ;
        RECT 54.820 148.175 55.405 148.365 ;
        RECT 53.755 147.835 54.960 148.005 ;
        RECT 53.755 147.405 54.085 147.835 ;
        RECT 54.265 147.225 54.460 147.665 ;
        RECT 54.630 147.405 54.960 147.835 ;
        RECT 55.130 147.405 55.405 148.175 ;
        RECT 56.595 148.235 59.655 148.405 ;
        RECT 56.595 147.395 56.765 148.235 ;
        RECT 59.825 148.075 59.995 149.195 ;
        RECT 61.110 149.010 61.565 149.775 ;
        RECT 61.840 149.395 63.140 149.605 ;
        RECT 63.395 149.415 63.725 149.775 ;
        RECT 62.970 149.245 63.140 149.395 ;
        RECT 63.895 149.275 64.155 149.605 ;
        RECT 62.040 148.785 62.260 149.185 ;
        RECT 61.105 148.585 61.595 148.785 ;
        RECT 61.785 148.575 62.260 148.785 ;
        RECT 62.505 148.785 62.715 149.185 ;
        RECT 62.970 149.120 63.725 149.245 ;
        RECT 62.970 149.075 63.815 149.120 ;
        RECT 63.545 148.955 63.815 149.075 ;
        RECT 62.505 148.575 62.835 148.785 ;
        RECT 63.005 148.515 63.415 148.820 ;
        RECT 59.785 148.065 59.995 148.075 ;
        RECT 56.935 147.565 57.265 148.065 ;
        RECT 57.435 147.825 59.070 148.065 ;
        RECT 57.435 147.735 57.665 147.825 ;
        RECT 57.775 147.565 58.105 147.605 ;
        RECT 56.935 147.395 58.105 147.565 ;
        RECT 58.295 147.225 58.650 147.645 ;
        RECT 58.820 147.395 59.070 147.825 ;
        RECT 59.240 147.225 59.570 147.985 ;
        RECT 59.740 147.395 59.995 148.065 ;
        RECT 61.110 148.345 62.285 148.405 ;
        RECT 63.645 148.380 63.815 148.955 ;
        RECT 63.615 148.345 63.815 148.380 ;
        RECT 61.110 148.235 63.815 148.345 ;
        RECT 61.110 147.615 61.365 148.235 ;
        RECT 61.955 148.175 63.755 148.235 ;
        RECT 61.955 148.145 62.285 148.175 ;
        RECT 63.985 148.075 64.155 149.275 ;
        RECT 61.615 147.975 61.800 148.065 ;
        RECT 62.390 147.975 63.225 147.985 ;
        RECT 61.615 147.775 63.225 147.975 ;
        RECT 61.615 147.735 61.845 147.775 ;
        RECT 61.110 147.395 61.445 147.615 ;
        RECT 62.450 147.225 62.805 147.605 ;
        RECT 62.975 147.395 63.225 147.775 ;
        RECT 63.475 147.225 63.725 148.005 ;
        RECT 63.895 147.395 64.155 148.075 ;
        RECT 64.360 149.035 64.975 149.605 ;
        RECT 65.145 149.265 65.360 149.775 ;
        RECT 65.590 149.265 65.870 149.595 ;
        RECT 66.050 149.265 66.290 149.775 ;
        RECT 64.360 148.015 64.675 149.035 ;
        RECT 64.845 148.365 65.015 148.865 ;
        RECT 65.265 148.535 65.530 149.095 ;
        RECT 65.700 148.365 65.870 149.265 ;
        RECT 66.040 148.535 66.395 149.095 ;
        RECT 66.625 149.005 68.295 149.775 ;
        RECT 68.925 149.050 69.215 149.775 ;
        RECT 69.935 149.225 70.105 149.515 ;
        RECT 70.275 149.395 70.605 149.775 ;
        RECT 69.935 149.055 70.600 149.225 ;
        RECT 66.625 148.485 67.375 149.005 ;
        RECT 64.845 148.195 66.270 148.365 ;
        RECT 67.545 148.315 68.295 148.835 ;
        RECT 64.360 147.395 64.895 148.015 ;
        RECT 65.065 147.225 65.395 148.025 ;
        RECT 65.880 148.020 66.270 148.195 ;
        RECT 66.625 147.225 68.295 148.315 ;
        RECT 68.925 147.225 69.215 148.390 ;
        RECT 69.850 148.235 70.200 148.885 ;
        RECT 70.370 148.065 70.600 149.055 ;
        RECT 69.935 147.895 70.600 148.065 ;
        RECT 69.935 147.395 70.105 147.895 ;
        RECT 70.275 147.225 70.605 147.725 ;
        RECT 70.775 147.395 70.960 149.515 ;
        RECT 71.215 149.315 71.465 149.775 ;
        RECT 71.635 149.325 71.970 149.495 ;
        RECT 72.165 149.325 72.840 149.495 ;
        RECT 71.635 149.185 71.805 149.325 ;
        RECT 71.130 148.195 71.410 149.145 ;
        RECT 71.580 149.055 71.805 149.185 ;
        RECT 71.580 147.950 71.750 149.055 ;
        RECT 71.975 148.905 72.500 149.125 ;
        RECT 71.920 148.140 72.160 148.735 ;
        RECT 72.330 148.205 72.500 148.905 ;
        RECT 72.670 148.545 72.840 149.325 ;
        RECT 73.160 149.275 73.530 149.775 ;
        RECT 73.710 149.325 74.115 149.495 ;
        RECT 74.285 149.325 75.070 149.495 ;
        RECT 73.710 149.095 73.880 149.325 ;
        RECT 73.050 148.795 73.880 149.095 ;
        RECT 74.265 148.825 74.730 149.155 ;
        RECT 73.050 148.765 73.250 148.795 ;
        RECT 73.370 148.545 73.540 148.615 ;
        RECT 72.670 148.375 73.540 148.545 ;
        RECT 73.030 148.285 73.540 148.375 ;
        RECT 71.580 147.820 71.885 147.950 ;
        RECT 72.330 147.840 72.860 148.205 ;
        RECT 71.200 147.225 71.465 147.685 ;
        RECT 71.635 147.395 71.885 147.820 ;
        RECT 73.030 147.670 73.200 148.285 ;
        RECT 72.095 147.500 73.200 147.670 ;
        RECT 73.370 147.225 73.540 148.025 ;
        RECT 73.710 147.725 73.880 148.795 ;
        RECT 74.050 147.895 74.240 148.615 ;
        RECT 74.410 147.865 74.730 148.825 ;
        RECT 74.900 148.865 75.070 149.325 ;
        RECT 75.345 149.245 75.555 149.775 ;
        RECT 75.815 149.035 76.145 149.560 ;
        RECT 76.315 149.165 76.485 149.775 ;
        RECT 76.655 149.120 76.985 149.555 ;
        RECT 76.655 149.035 77.035 149.120 ;
        RECT 75.945 148.865 76.145 149.035 ;
        RECT 76.810 148.995 77.035 149.035 ;
        RECT 74.900 148.535 75.775 148.865 ;
        RECT 75.945 148.535 76.695 148.865 ;
        RECT 73.710 147.395 73.960 147.725 ;
        RECT 74.900 147.695 75.070 148.535 ;
        RECT 75.945 148.330 76.135 148.535 ;
        RECT 76.865 148.415 77.035 148.995 ;
        RECT 77.205 149.005 79.795 149.775 ;
        RECT 80.425 149.265 80.730 149.775 ;
        RECT 77.205 148.485 78.415 149.005 ;
        RECT 76.820 148.365 77.035 148.415 ;
        RECT 75.240 147.955 76.135 148.330 ;
        RECT 76.645 148.285 77.035 148.365 ;
        RECT 78.585 148.315 79.795 148.835 ;
        RECT 80.425 148.535 80.740 149.095 ;
        RECT 80.910 148.785 81.160 149.595 ;
        RECT 81.330 149.250 81.590 149.775 ;
        RECT 81.770 148.785 82.020 149.595 ;
        RECT 82.190 149.215 82.450 149.775 ;
        RECT 82.620 149.125 82.880 149.580 ;
        RECT 83.050 149.295 83.310 149.775 ;
        RECT 83.480 149.125 83.740 149.580 ;
        RECT 83.910 149.295 84.170 149.775 ;
        RECT 84.340 149.125 84.600 149.580 ;
        RECT 84.770 149.295 85.015 149.775 ;
        RECT 85.185 149.125 85.460 149.580 ;
        RECT 85.630 149.295 85.875 149.775 ;
        RECT 86.045 149.125 86.305 149.580 ;
        RECT 86.485 149.295 86.735 149.775 ;
        RECT 86.905 149.125 87.165 149.580 ;
        RECT 87.345 149.295 87.595 149.775 ;
        RECT 87.765 149.125 88.025 149.580 ;
        RECT 88.205 149.295 88.465 149.775 ;
        RECT 88.635 149.125 88.895 149.580 ;
        RECT 89.065 149.295 89.365 149.775 ;
        RECT 89.740 149.145 90.025 149.605 ;
        RECT 90.195 149.315 90.465 149.775 ;
        RECT 82.620 148.955 89.365 149.125 ;
        RECT 89.740 148.975 90.695 149.145 ;
        RECT 80.910 148.535 88.030 148.785 ;
        RECT 74.185 147.525 75.070 147.695 ;
        RECT 75.250 147.225 75.565 147.725 ;
        RECT 75.795 147.395 76.135 147.955 ;
        RECT 76.305 147.225 76.475 148.235 ;
        RECT 76.645 147.440 76.975 148.285 ;
        RECT 77.205 147.225 79.795 148.315 ;
        RECT 80.435 147.225 80.730 148.035 ;
        RECT 80.910 147.395 81.155 148.535 ;
        RECT 81.330 147.225 81.590 148.035 ;
        RECT 81.770 147.400 82.020 148.535 ;
        RECT 88.200 148.365 89.365 148.955 ;
        RECT 82.620 148.140 89.365 148.365 ;
        RECT 89.625 148.245 90.315 148.805 ;
        RECT 82.620 148.125 88.025 148.140 ;
        RECT 82.190 147.230 82.450 148.025 ;
        RECT 82.620 147.400 82.880 148.125 ;
        RECT 83.050 147.230 83.310 147.955 ;
        RECT 83.480 147.400 83.740 148.125 ;
        RECT 83.910 147.230 84.170 147.955 ;
        RECT 84.340 147.400 84.600 148.125 ;
        RECT 84.770 147.230 85.030 147.955 ;
        RECT 85.200 147.400 85.460 148.125 ;
        RECT 85.630 147.230 85.875 147.955 ;
        RECT 86.045 147.400 86.305 148.125 ;
        RECT 86.490 147.230 86.735 147.955 ;
        RECT 86.905 147.400 87.165 148.125 ;
        RECT 87.350 147.230 87.595 147.955 ;
        RECT 87.765 147.400 88.025 148.125 ;
        RECT 88.210 147.230 88.465 147.955 ;
        RECT 88.635 147.400 88.925 148.140 ;
        RECT 90.485 148.075 90.695 148.975 ;
        RECT 82.190 147.225 88.465 147.230 ;
        RECT 89.095 147.225 89.365 147.970 ;
        RECT 89.740 147.855 90.695 148.075 ;
        RECT 90.865 148.805 91.265 149.605 ;
        RECT 91.455 149.145 91.735 149.605 ;
        RECT 92.255 149.315 92.580 149.775 ;
        RECT 91.455 148.975 92.580 149.145 ;
        RECT 92.750 149.035 93.135 149.605 ;
        RECT 92.130 148.865 92.580 148.975 ;
        RECT 90.865 148.245 91.960 148.805 ;
        RECT 92.130 148.535 92.685 148.865 ;
        RECT 89.740 147.395 90.025 147.855 ;
        RECT 90.195 147.225 90.465 147.685 ;
        RECT 90.865 147.395 91.265 148.245 ;
        RECT 92.130 148.075 92.580 148.535 ;
        RECT 92.855 148.365 93.135 149.035 ;
        RECT 93.305 149.025 94.515 149.775 ;
        RECT 94.685 149.050 94.975 149.775 ;
        RECT 95.150 149.035 95.405 149.605 ;
        RECT 95.575 149.375 95.905 149.775 ;
        RECT 96.330 149.240 96.860 149.605 ;
        RECT 96.330 149.205 96.505 149.240 ;
        RECT 95.575 149.035 96.505 149.205 ;
        RECT 93.305 148.485 93.825 149.025 ;
        RECT 91.455 147.855 92.580 148.075 ;
        RECT 91.455 147.395 91.735 147.855 ;
        RECT 92.255 147.225 92.580 147.685 ;
        RECT 92.750 147.395 93.135 148.365 ;
        RECT 93.995 148.315 94.515 148.855 ;
        RECT 93.305 147.225 94.515 148.315 ;
        RECT 94.685 147.225 94.975 148.390 ;
        RECT 95.150 148.365 95.320 149.035 ;
        RECT 95.575 148.865 95.745 149.035 ;
        RECT 95.490 148.535 95.745 148.865 ;
        RECT 95.970 148.535 96.165 148.865 ;
        RECT 95.150 147.395 95.485 148.365 ;
        RECT 95.655 147.225 95.825 148.365 ;
        RECT 95.995 147.565 96.165 148.535 ;
        RECT 96.335 147.905 96.505 149.035 ;
        RECT 96.675 148.245 96.845 149.045 ;
        RECT 97.050 148.755 97.325 149.605 ;
        RECT 97.045 148.585 97.325 148.755 ;
        RECT 97.050 148.445 97.325 148.585 ;
        RECT 97.495 148.245 97.685 149.605 ;
        RECT 97.865 149.240 98.375 149.775 ;
        RECT 98.595 148.965 98.840 149.570 ;
        RECT 99.290 149.035 99.545 149.605 ;
        RECT 99.715 149.375 100.045 149.775 ;
        RECT 100.470 149.240 101.000 149.605 ;
        RECT 100.470 149.205 100.645 149.240 ;
        RECT 99.715 149.035 100.645 149.205 ;
        RECT 97.885 148.795 99.115 148.965 ;
        RECT 96.675 148.075 97.685 148.245 ;
        RECT 97.855 148.230 98.605 148.420 ;
        RECT 96.335 147.735 97.460 147.905 ;
        RECT 97.855 147.565 98.025 148.230 ;
        RECT 98.775 147.985 99.115 148.795 ;
        RECT 95.995 147.395 98.025 147.565 ;
        RECT 98.195 147.225 98.365 147.985 ;
        RECT 98.600 147.575 99.115 147.985 ;
        RECT 99.290 148.365 99.460 149.035 ;
        RECT 99.715 148.865 99.885 149.035 ;
        RECT 99.630 148.535 99.885 148.865 ;
        RECT 100.110 148.535 100.305 148.865 ;
        RECT 99.290 147.395 99.625 148.365 ;
        RECT 99.795 147.225 99.965 148.365 ;
        RECT 100.135 147.565 100.305 148.535 ;
        RECT 100.475 147.905 100.645 149.035 ;
        RECT 100.815 148.245 100.985 149.045 ;
        RECT 101.190 148.755 101.465 149.605 ;
        RECT 101.185 148.585 101.465 148.755 ;
        RECT 101.190 148.445 101.465 148.585 ;
        RECT 101.635 148.245 101.825 149.605 ;
        RECT 102.005 149.240 102.515 149.775 ;
        RECT 102.735 148.965 102.980 149.570 ;
        RECT 102.025 148.795 103.255 148.965 ;
        RECT 103.485 148.955 103.695 149.775 ;
        RECT 103.865 148.975 104.195 149.605 ;
        RECT 100.815 148.075 101.825 148.245 ;
        RECT 101.995 148.230 102.745 148.420 ;
        RECT 100.475 147.735 101.600 147.905 ;
        RECT 101.995 147.565 102.165 148.230 ;
        RECT 102.915 147.985 103.255 148.795 ;
        RECT 103.865 148.375 104.115 148.975 ;
        RECT 104.365 148.955 104.595 149.775 ;
        RECT 104.810 149.035 105.065 149.605 ;
        RECT 105.235 149.375 105.565 149.775 ;
        RECT 105.990 149.240 106.520 149.605 ;
        RECT 105.990 149.205 106.165 149.240 ;
        RECT 105.235 149.035 106.165 149.205 ;
        RECT 104.285 148.535 104.615 148.785 ;
        RECT 100.135 147.395 102.165 147.565 ;
        RECT 102.335 147.225 102.505 147.985 ;
        RECT 102.740 147.575 103.255 147.985 ;
        RECT 103.485 147.225 103.695 148.365 ;
        RECT 103.865 147.395 104.195 148.375 ;
        RECT 104.810 148.365 104.980 149.035 ;
        RECT 105.235 148.865 105.405 149.035 ;
        RECT 105.150 148.535 105.405 148.865 ;
        RECT 105.630 148.535 105.825 148.865 ;
        RECT 104.365 147.225 104.595 148.365 ;
        RECT 104.810 147.395 105.145 148.365 ;
        RECT 105.315 147.225 105.485 148.365 ;
        RECT 105.655 147.565 105.825 148.535 ;
        RECT 105.995 147.905 106.165 149.035 ;
        RECT 106.335 148.245 106.505 149.045 ;
        RECT 106.710 148.755 106.985 149.605 ;
        RECT 106.705 148.585 106.985 148.755 ;
        RECT 106.710 148.445 106.985 148.585 ;
        RECT 107.155 148.245 107.345 149.605 ;
        RECT 107.525 149.240 108.035 149.775 ;
        RECT 108.255 148.965 108.500 149.570 ;
        RECT 108.945 149.005 110.615 149.775 ;
        RECT 110.900 149.145 111.185 149.605 ;
        RECT 111.355 149.315 111.625 149.775 ;
        RECT 107.545 148.795 108.775 148.965 ;
        RECT 106.335 148.075 107.345 148.245 ;
        RECT 107.515 148.230 108.265 148.420 ;
        RECT 105.995 147.735 107.120 147.905 ;
        RECT 107.515 147.565 107.685 148.230 ;
        RECT 108.435 147.985 108.775 148.795 ;
        RECT 108.945 148.485 109.695 149.005 ;
        RECT 110.900 148.975 111.855 149.145 ;
        RECT 109.865 148.315 110.615 148.835 ;
        RECT 105.655 147.395 107.685 147.565 ;
        RECT 107.855 147.225 108.025 147.985 ;
        RECT 108.260 147.575 108.775 147.985 ;
        RECT 108.945 147.225 110.615 148.315 ;
        RECT 110.785 148.245 111.475 148.805 ;
        RECT 111.645 148.075 111.855 148.975 ;
        RECT 110.900 147.855 111.855 148.075 ;
        RECT 112.025 148.805 112.425 149.605 ;
        RECT 112.615 149.145 112.895 149.605 ;
        RECT 113.415 149.315 113.740 149.775 ;
        RECT 112.615 148.975 113.740 149.145 ;
        RECT 113.910 149.035 114.295 149.605 ;
        RECT 114.470 149.245 114.760 149.595 ;
        RECT 114.955 149.415 115.285 149.775 ;
        RECT 115.455 149.245 115.685 149.550 ;
        RECT 114.470 149.075 115.685 149.245 ;
        RECT 113.290 148.865 113.740 148.975 ;
        RECT 112.025 148.245 113.120 148.805 ;
        RECT 113.290 148.535 113.845 148.865 ;
        RECT 110.900 147.395 111.185 147.855 ;
        RECT 111.355 147.225 111.625 147.685 ;
        RECT 112.025 147.395 112.425 148.245 ;
        RECT 113.290 148.075 113.740 148.535 ;
        RECT 114.015 148.365 114.295 149.035 ;
        RECT 115.875 148.905 116.045 149.470 ;
        RECT 114.530 148.755 114.790 148.865 ;
        RECT 114.525 148.585 114.790 148.755 ;
        RECT 114.530 148.535 114.790 148.585 ;
        RECT 114.970 148.535 115.355 148.865 ;
        RECT 115.525 148.735 116.045 148.905 ;
        RECT 116.395 148.905 116.565 149.470 ;
        RECT 116.755 149.245 116.985 149.550 ;
        RECT 117.155 149.415 117.485 149.775 ;
        RECT 117.680 149.245 117.970 149.595 ;
        RECT 116.755 149.075 117.970 149.245 ;
        RECT 118.150 149.245 118.440 149.595 ;
        RECT 118.635 149.415 118.965 149.775 ;
        RECT 119.135 149.245 119.365 149.550 ;
        RECT 118.150 149.075 119.365 149.245 ;
        RECT 119.555 148.905 119.725 149.470 ;
        RECT 120.445 149.050 120.735 149.775 ;
        RECT 121.695 149.375 122.025 149.775 ;
        RECT 122.195 149.205 122.525 149.545 ;
        RECT 123.575 149.375 123.905 149.775 ;
        RECT 116.395 148.735 116.915 148.905 ;
        RECT 112.615 147.855 113.740 148.075 ;
        RECT 112.615 147.395 112.895 147.855 ;
        RECT 113.415 147.225 113.740 147.685 ;
        RECT 113.910 147.395 114.295 148.365 ;
        RECT 114.470 147.225 114.790 148.365 ;
        RECT 114.970 147.485 115.165 148.535 ;
        RECT 115.525 148.355 115.695 148.735 ;
        RECT 115.345 148.075 115.695 148.355 ;
        RECT 115.885 148.205 116.130 148.565 ;
        RECT 116.310 148.205 116.555 148.565 ;
        RECT 116.745 148.355 116.915 148.735 ;
        RECT 117.085 148.535 117.470 148.865 ;
        RECT 117.650 148.755 117.910 148.865 ;
        RECT 118.210 148.755 118.470 148.865 ;
        RECT 117.650 148.585 117.915 148.755 ;
        RECT 118.205 148.585 118.470 148.755 ;
        RECT 117.650 148.535 117.910 148.585 ;
        RECT 118.210 148.535 118.470 148.585 ;
        RECT 118.650 148.535 119.035 148.865 ;
        RECT 119.205 148.735 119.725 148.905 ;
        RECT 121.540 149.035 123.905 149.205 ;
        RECT 124.075 149.050 124.405 149.560 ;
        RECT 116.745 148.075 117.095 148.355 ;
        RECT 115.345 147.395 115.675 148.075 ;
        RECT 115.875 147.225 116.130 148.025 ;
        RECT 116.310 147.225 116.565 148.025 ;
        RECT 116.765 147.395 117.095 148.075 ;
        RECT 117.275 147.485 117.470 148.535 ;
        RECT 117.650 147.225 117.970 148.365 ;
        RECT 118.150 147.225 118.470 148.365 ;
        RECT 118.650 147.485 118.845 148.535 ;
        RECT 119.205 148.355 119.375 148.735 ;
        RECT 119.025 148.075 119.375 148.355 ;
        RECT 119.565 148.205 119.810 148.565 ;
        RECT 119.025 147.395 119.355 148.075 ;
        RECT 119.555 147.225 119.810 148.025 ;
        RECT 120.445 147.225 120.735 148.390 ;
        RECT 121.540 148.035 121.710 149.035 ;
        RECT 123.735 148.865 123.905 149.035 ;
        RECT 121.880 148.205 122.125 148.865 ;
        RECT 122.340 148.205 122.605 148.865 ;
        RECT 122.800 148.205 123.085 148.865 ;
        RECT 123.260 148.535 123.565 148.865 ;
        RECT 123.735 148.535 124.045 148.865 ;
        RECT 123.260 148.205 123.475 148.535 ;
        RECT 121.540 147.865 121.995 148.035 ;
        RECT 121.665 147.435 121.995 147.865 ;
        RECT 122.175 147.865 123.465 148.035 ;
        RECT 122.175 147.445 122.425 147.865 ;
        RECT 122.655 147.225 122.985 147.695 ;
        RECT 123.215 147.445 123.465 147.865 ;
        RECT 123.655 147.225 123.905 148.365 ;
        RECT 124.215 148.285 124.405 149.050 ;
        RECT 124.585 148.975 124.895 149.775 ;
        RECT 125.100 148.975 125.795 149.605 ;
        RECT 127.050 149.265 127.290 149.775 ;
        RECT 127.470 149.265 127.750 149.595 ;
        RECT 127.980 149.265 128.195 149.775 ;
        RECT 124.595 148.535 124.930 148.805 ;
        RECT 125.100 148.375 125.270 148.975 ;
        RECT 125.440 148.535 125.775 148.785 ;
        RECT 126.945 148.535 127.300 149.095 ;
        RECT 124.075 147.435 124.405 148.285 ;
        RECT 124.585 147.225 124.865 148.365 ;
        RECT 125.035 147.395 125.365 148.375 ;
        RECT 127.470 148.365 127.640 149.265 ;
        RECT 127.810 148.535 128.075 149.095 ;
        RECT 128.365 149.035 128.980 149.605 ;
        RECT 128.325 148.365 128.495 148.865 ;
        RECT 125.535 147.225 125.795 148.365 ;
        RECT 127.070 148.195 128.495 148.365 ;
        RECT 127.070 148.020 127.460 148.195 ;
        RECT 127.945 147.225 128.275 148.025 ;
        RECT 128.665 148.015 128.980 149.035 ;
        RECT 129.190 149.010 129.645 149.775 ;
        RECT 129.920 149.395 131.220 149.605 ;
        RECT 131.475 149.415 131.805 149.775 ;
        RECT 131.050 149.245 131.220 149.395 ;
        RECT 131.975 149.275 132.235 149.605 ;
        RECT 132.005 149.265 132.235 149.275 ;
        RECT 130.120 148.785 130.340 149.185 ;
        RECT 129.185 148.585 129.675 148.785 ;
        RECT 129.865 148.575 130.340 148.785 ;
        RECT 130.585 148.785 130.795 149.185 ;
        RECT 131.050 149.120 131.805 149.245 ;
        RECT 131.050 149.075 131.895 149.120 ;
        RECT 131.625 148.955 131.895 149.075 ;
        RECT 130.585 148.575 130.915 148.785 ;
        RECT 131.085 148.515 131.495 148.820 ;
        RECT 128.445 147.395 128.980 148.015 ;
        RECT 129.190 148.345 130.365 148.405 ;
        RECT 131.725 148.380 131.895 148.955 ;
        RECT 131.695 148.345 131.895 148.380 ;
        RECT 129.190 148.235 131.895 148.345 ;
        RECT 129.190 147.615 129.445 148.235 ;
        RECT 130.035 148.175 131.835 148.235 ;
        RECT 130.035 148.145 130.365 148.175 ;
        RECT 132.065 148.075 132.235 149.265 ;
        RECT 132.405 149.005 134.075 149.775 ;
        RECT 134.335 149.225 134.505 149.515 ;
        RECT 134.675 149.395 135.005 149.775 ;
        RECT 134.335 149.055 135.000 149.225 ;
        RECT 132.405 148.485 133.155 149.005 ;
        RECT 133.325 148.315 134.075 148.835 ;
        RECT 129.695 147.975 129.880 148.065 ;
        RECT 130.470 147.975 131.305 147.985 ;
        RECT 129.695 147.775 131.305 147.975 ;
        RECT 129.695 147.735 129.925 147.775 ;
        RECT 129.190 147.395 129.525 147.615 ;
        RECT 130.530 147.225 130.885 147.605 ;
        RECT 131.055 147.395 131.305 147.775 ;
        RECT 131.555 147.225 131.805 148.005 ;
        RECT 131.975 147.395 132.235 148.075 ;
        RECT 132.405 147.225 134.075 148.315 ;
        RECT 134.250 148.235 134.600 148.885 ;
        RECT 134.770 148.065 135.000 149.055 ;
        RECT 134.335 147.895 135.000 148.065 ;
        RECT 134.335 147.395 134.505 147.895 ;
        RECT 134.675 147.225 135.005 147.725 ;
        RECT 135.175 147.395 135.360 149.515 ;
        RECT 135.615 149.315 135.865 149.775 ;
        RECT 136.035 149.325 136.370 149.495 ;
        RECT 136.565 149.325 137.240 149.495 ;
        RECT 136.035 149.185 136.205 149.325 ;
        RECT 135.530 148.195 135.810 149.145 ;
        RECT 135.980 149.055 136.205 149.185 ;
        RECT 135.980 147.950 136.150 149.055 ;
        RECT 136.375 148.905 136.900 149.125 ;
        RECT 136.320 148.140 136.560 148.735 ;
        RECT 136.730 148.205 136.900 148.905 ;
        RECT 137.070 148.545 137.240 149.325 ;
        RECT 137.560 149.275 137.930 149.775 ;
        RECT 138.110 149.325 138.515 149.495 ;
        RECT 138.685 149.325 139.470 149.495 ;
        RECT 138.110 149.095 138.280 149.325 ;
        RECT 137.450 148.795 138.280 149.095 ;
        RECT 138.665 148.825 139.130 149.155 ;
        RECT 137.450 148.765 137.650 148.795 ;
        RECT 137.770 148.545 137.940 148.615 ;
        RECT 137.070 148.375 137.940 148.545 ;
        RECT 137.430 148.285 137.940 148.375 ;
        RECT 135.980 147.820 136.285 147.950 ;
        RECT 136.730 147.840 137.260 148.205 ;
        RECT 135.600 147.225 135.865 147.685 ;
        RECT 136.035 147.395 136.285 147.820 ;
        RECT 137.430 147.670 137.600 148.285 ;
        RECT 136.495 147.500 137.600 147.670 ;
        RECT 137.770 147.225 137.940 148.025 ;
        RECT 138.110 147.725 138.280 148.795 ;
        RECT 138.450 147.895 138.640 148.615 ;
        RECT 138.810 147.865 139.130 148.825 ;
        RECT 139.300 148.865 139.470 149.325 ;
        RECT 139.745 149.245 139.955 149.775 ;
        RECT 140.215 149.035 140.545 149.560 ;
        RECT 140.715 149.165 140.885 149.775 ;
        RECT 141.055 149.120 141.385 149.555 ;
        RECT 141.055 149.035 141.435 149.120 ;
        RECT 140.345 148.865 140.545 149.035 ;
        RECT 141.210 148.995 141.435 149.035 ;
        RECT 139.300 148.535 140.175 148.865 ;
        RECT 140.345 148.535 141.095 148.865 ;
        RECT 138.110 147.395 138.360 147.725 ;
        RECT 139.300 147.695 139.470 148.535 ;
        RECT 140.345 148.330 140.535 148.535 ;
        RECT 141.265 148.415 141.435 148.995 ;
        RECT 141.220 148.365 141.435 148.415 ;
        RECT 139.640 147.955 140.535 148.330 ;
        RECT 141.045 148.285 141.435 148.365 ;
        RECT 141.610 149.035 141.865 149.605 ;
        RECT 142.035 149.375 142.365 149.775 ;
        RECT 142.790 149.240 143.320 149.605 ;
        RECT 142.790 149.205 142.965 149.240 ;
        RECT 142.035 149.035 142.965 149.205 ;
        RECT 141.610 148.365 141.780 149.035 ;
        RECT 142.035 148.865 142.205 149.035 ;
        RECT 141.950 148.535 142.205 148.865 ;
        RECT 142.430 148.535 142.625 148.865 ;
        RECT 138.585 147.525 139.470 147.695 ;
        RECT 139.650 147.225 139.965 147.725 ;
        RECT 140.195 147.395 140.535 147.955 ;
        RECT 140.705 147.225 140.875 148.235 ;
        RECT 141.045 147.440 141.375 148.285 ;
        RECT 141.610 147.395 141.945 148.365 ;
        RECT 142.115 147.225 142.285 148.365 ;
        RECT 142.455 147.565 142.625 148.535 ;
        RECT 142.795 147.905 142.965 149.035 ;
        RECT 143.135 148.245 143.305 149.045 ;
        RECT 143.510 148.755 143.785 149.605 ;
        RECT 143.505 148.585 143.785 148.755 ;
        RECT 143.510 148.445 143.785 148.585 ;
        RECT 143.955 148.245 144.145 149.605 ;
        RECT 144.325 149.240 144.835 149.775 ;
        RECT 145.055 148.965 145.300 149.570 ;
        RECT 145.745 149.025 146.955 149.775 ;
        RECT 144.345 148.795 145.575 148.965 ;
        RECT 143.135 148.075 144.145 148.245 ;
        RECT 144.315 148.230 145.065 148.420 ;
        RECT 142.795 147.735 143.920 147.905 ;
        RECT 144.315 147.565 144.485 148.230 ;
        RECT 145.235 147.985 145.575 148.795 ;
        RECT 142.455 147.395 144.485 147.565 ;
        RECT 144.655 147.225 144.825 147.985 ;
        RECT 145.060 147.575 145.575 147.985 ;
        RECT 145.745 148.315 146.265 148.855 ;
        RECT 146.435 148.485 146.955 149.025 ;
        RECT 145.745 147.225 146.955 148.315 ;
        RECT 17.320 147.055 147.040 147.225 ;
        RECT 17.405 145.965 18.615 147.055 ;
        RECT 18.785 146.620 24.130 147.055 ;
        RECT 24.305 146.620 29.650 147.055 ;
        RECT 17.405 145.255 17.925 145.795 ;
        RECT 18.095 145.425 18.615 145.965 ;
        RECT 17.405 144.505 18.615 145.255 ;
        RECT 20.370 145.050 20.710 145.880 ;
        RECT 22.190 145.370 22.540 146.620 ;
        RECT 25.890 145.050 26.230 145.880 ;
        RECT 27.710 145.370 28.060 146.620 ;
        RECT 30.285 145.890 30.575 147.055 ;
        RECT 31.265 145.995 31.595 146.840 ;
        RECT 31.765 146.045 31.935 147.055 ;
        RECT 32.105 146.325 32.445 146.885 ;
        RECT 32.675 146.555 32.990 147.055 ;
        RECT 33.170 146.585 34.055 146.755 ;
        RECT 31.205 145.915 31.595 145.995 ;
        RECT 32.105 145.950 33.000 146.325 ;
        RECT 31.205 145.865 31.420 145.915 ;
        RECT 31.205 145.285 31.375 145.865 ;
        RECT 32.105 145.745 32.295 145.950 ;
        RECT 33.170 145.745 33.340 146.585 ;
        RECT 34.280 146.555 34.530 146.885 ;
        RECT 31.545 145.415 32.295 145.745 ;
        RECT 32.465 145.415 33.340 145.745 ;
        RECT 31.205 145.245 31.430 145.285 ;
        RECT 32.095 145.245 32.295 145.415 ;
        RECT 18.785 144.505 24.130 145.050 ;
        RECT 24.305 144.505 29.650 145.050 ;
        RECT 30.285 144.505 30.575 145.230 ;
        RECT 31.205 145.160 31.585 145.245 ;
        RECT 31.255 144.725 31.585 145.160 ;
        RECT 31.755 144.505 31.925 145.115 ;
        RECT 32.095 144.720 32.425 145.245 ;
        RECT 32.685 144.505 32.895 145.035 ;
        RECT 33.170 144.955 33.340 145.415 ;
        RECT 33.510 145.455 33.830 146.415 ;
        RECT 34.000 145.665 34.190 146.385 ;
        RECT 34.360 145.485 34.530 146.555 ;
        RECT 34.700 146.255 34.870 147.055 ;
        RECT 35.040 146.610 36.145 146.780 ;
        RECT 35.040 145.995 35.210 146.610 ;
        RECT 36.355 146.460 36.605 146.885 ;
        RECT 36.775 146.595 37.040 147.055 ;
        RECT 35.380 146.075 35.910 146.440 ;
        RECT 36.355 146.330 36.660 146.460 ;
        RECT 34.700 145.905 35.210 145.995 ;
        RECT 34.700 145.735 35.570 145.905 ;
        RECT 34.700 145.665 34.870 145.735 ;
        RECT 34.990 145.485 35.190 145.515 ;
        RECT 33.510 145.125 33.975 145.455 ;
        RECT 34.360 145.185 35.190 145.485 ;
        RECT 34.360 144.955 34.530 145.185 ;
        RECT 33.170 144.785 33.955 144.955 ;
        RECT 34.125 144.785 34.530 144.955 ;
        RECT 34.710 144.505 35.080 145.005 ;
        RECT 35.400 144.955 35.570 145.735 ;
        RECT 35.740 145.375 35.910 146.075 ;
        RECT 36.080 145.545 36.320 146.140 ;
        RECT 35.740 145.155 36.265 145.375 ;
        RECT 36.490 145.225 36.660 146.330 ;
        RECT 36.435 145.095 36.660 145.225 ;
        RECT 36.830 145.135 37.110 146.085 ;
        RECT 36.435 144.955 36.605 145.095 ;
        RECT 35.400 144.785 36.075 144.955 ;
        RECT 36.270 144.785 36.605 144.955 ;
        RECT 36.775 144.505 37.025 144.965 ;
        RECT 37.280 144.765 37.465 146.885 ;
        RECT 37.635 146.555 37.965 147.055 ;
        RECT 38.135 146.385 38.305 146.885 ;
        RECT 37.640 146.215 38.305 146.385 ;
        RECT 37.640 145.225 37.870 146.215 ;
        RECT 38.040 145.395 38.390 146.045 ;
        RECT 38.575 145.995 38.905 146.845 ;
        RECT 38.575 145.230 38.765 145.995 ;
        RECT 39.075 145.915 39.325 147.055 ;
        RECT 39.515 146.415 39.765 146.835 ;
        RECT 39.995 146.585 40.325 147.055 ;
        RECT 40.555 146.415 40.805 146.835 ;
        RECT 39.515 146.245 40.805 146.415 ;
        RECT 40.985 146.415 41.315 146.845 ;
        RECT 40.985 146.245 41.440 146.415 ;
        RECT 39.505 145.745 39.720 146.075 ;
        RECT 38.935 145.415 39.245 145.745 ;
        RECT 39.415 145.415 39.720 145.745 ;
        RECT 39.895 145.415 40.180 146.075 ;
        RECT 40.375 145.415 40.640 146.075 ;
        RECT 40.855 145.415 41.100 146.075 ;
        RECT 39.075 145.245 39.245 145.415 ;
        RECT 41.270 145.245 41.440 146.245 ;
        RECT 42.285 146.105 42.575 146.875 ;
        RECT 43.145 146.515 43.405 146.875 ;
        RECT 43.575 146.685 43.905 147.055 ;
        RECT 44.075 146.515 44.335 146.875 ;
        RECT 43.145 146.285 44.335 146.515 ;
        RECT 44.525 146.335 44.855 147.055 ;
        RECT 45.025 146.105 45.290 146.875 ;
        RECT 42.285 145.925 44.780 146.105 ;
        RECT 42.255 145.415 42.525 145.745 ;
        RECT 42.705 145.415 43.140 145.745 ;
        RECT 43.320 145.415 43.895 145.745 ;
        RECT 44.075 145.415 44.355 145.745 ;
        RECT 37.640 145.055 38.305 145.225 ;
        RECT 37.635 144.505 37.965 144.885 ;
        RECT 38.135 144.765 38.305 145.055 ;
        RECT 38.575 144.720 38.905 145.230 ;
        RECT 39.075 145.075 41.440 145.245 ;
        RECT 44.555 145.235 44.780 145.925 ;
        RECT 39.075 144.505 39.405 144.905 ;
        RECT 40.455 144.735 40.785 145.075 ;
        RECT 42.295 145.045 44.780 145.235 ;
        RECT 40.955 144.505 41.285 144.905 ;
        RECT 42.295 144.685 42.520 145.045 ;
        RECT 42.700 144.505 43.030 144.875 ;
        RECT 43.210 144.685 43.465 145.045 ;
        RECT 44.030 144.505 44.775 144.875 ;
        RECT 44.955 144.685 45.290 146.105 ;
        RECT 45.485 146.165 45.745 146.875 ;
        RECT 45.915 146.345 46.245 147.055 ;
        RECT 46.415 146.165 46.645 146.875 ;
        RECT 45.485 145.925 46.645 146.165 ;
        RECT 46.825 146.145 47.095 146.875 ;
        RECT 47.275 146.325 47.615 147.055 ;
        RECT 46.825 145.925 47.595 146.145 ;
        RECT 45.475 145.415 45.775 145.745 ;
        RECT 45.955 145.435 46.480 145.745 ;
        RECT 46.660 145.435 47.125 145.745 ;
        RECT 45.485 144.505 45.775 145.235 ;
        RECT 45.955 144.795 46.185 145.435 ;
        RECT 47.305 145.255 47.595 145.925 ;
        RECT 46.365 145.055 47.595 145.255 ;
        RECT 46.365 144.685 46.675 145.055 ;
        RECT 46.855 144.505 47.525 144.875 ;
        RECT 47.785 144.685 48.045 146.875 ;
        RECT 48.225 146.620 53.570 147.055 ;
        RECT 49.810 145.050 50.150 145.880 ;
        RECT 51.630 145.370 51.980 146.620 ;
        RECT 53.745 145.965 55.415 147.055 ;
        RECT 53.745 145.275 54.495 145.795 ;
        RECT 54.665 145.445 55.415 145.965 ;
        RECT 56.045 145.890 56.335 147.055 ;
        RECT 57.625 146.385 57.905 147.055 ;
        RECT 58.075 146.165 58.375 146.715 ;
        RECT 58.575 146.335 58.905 147.055 ;
        RECT 59.095 146.335 59.555 146.885 ;
        RECT 59.725 146.545 59.985 147.055 ;
        RECT 57.440 145.745 57.705 146.105 ;
        RECT 58.075 145.995 59.015 146.165 ;
        RECT 58.845 145.745 59.015 145.995 ;
        RECT 57.440 145.495 58.115 145.745 ;
        RECT 58.335 145.495 58.675 145.745 ;
        RECT 58.845 145.415 59.135 145.745 ;
        RECT 58.845 145.325 59.015 145.415 ;
        RECT 48.225 144.505 53.570 145.050 ;
        RECT 53.745 144.505 55.415 145.275 ;
        RECT 56.045 144.505 56.335 145.230 ;
        RECT 57.625 145.135 59.015 145.325 ;
        RECT 57.625 144.775 57.955 145.135 ;
        RECT 59.305 144.965 59.555 146.335 ;
        RECT 59.725 145.495 60.065 146.375 ;
        RECT 60.235 145.665 60.405 146.885 ;
        RECT 60.645 146.550 61.260 147.055 ;
        RECT 60.645 146.015 60.895 146.380 ;
        RECT 61.065 146.375 61.260 146.550 ;
        RECT 61.430 146.545 61.905 146.885 ;
        RECT 62.075 146.510 62.290 147.055 ;
        RECT 61.065 146.185 61.395 146.375 ;
        RECT 61.615 146.015 62.330 146.310 ;
        RECT 62.500 146.185 62.775 146.885 ;
        RECT 60.645 145.845 62.435 146.015 ;
        RECT 60.235 145.415 61.030 145.665 ;
        RECT 60.235 145.325 60.485 145.415 ;
        RECT 58.575 144.505 58.825 144.965 ;
        RECT 58.995 144.675 59.555 144.965 ;
        RECT 59.725 144.505 59.985 145.325 ;
        RECT 60.155 144.905 60.485 145.325 ;
        RECT 61.200 144.990 61.455 145.845 ;
        RECT 60.665 144.725 61.455 144.990 ;
        RECT 61.625 145.145 62.035 145.665 ;
        RECT 62.205 145.415 62.435 145.845 ;
        RECT 62.605 145.155 62.775 146.185 ;
        RECT 61.625 144.725 61.825 145.145 ;
        RECT 62.015 144.505 62.345 144.965 ;
        RECT 62.515 144.675 62.775 145.155 ;
        RECT 62.980 146.265 63.515 146.885 ;
        RECT 62.980 145.245 63.295 146.265 ;
        RECT 63.685 146.255 64.015 147.055 ;
        RECT 65.245 146.620 70.590 147.055 ;
        RECT 70.765 146.620 76.110 147.055 ;
        RECT 64.500 146.085 64.890 146.260 ;
        RECT 63.465 145.915 64.890 146.085 ;
        RECT 63.465 145.415 63.635 145.915 ;
        RECT 62.980 144.675 63.595 145.245 ;
        RECT 63.885 145.185 64.150 145.745 ;
        RECT 64.320 145.015 64.490 145.915 ;
        RECT 64.660 145.185 65.015 145.745 ;
        RECT 66.830 145.050 67.170 145.880 ;
        RECT 68.650 145.370 69.000 146.620 ;
        RECT 72.350 145.050 72.690 145.880 ;
        RECT 74.170 145.370 74.520 146.620 ;
        RECT 76.780 146.265 77.315 146.885 ;
        RECT 76.780 145.245 77.095 146.265 ;
        RECT 77.485 146.255 77.815 147.055 ;
        RECT 78.300 146.085 78.690 146.260 ;
        RECT 77.265 145.915 78.690 146.085 ;
        RECT 79.105 145.915 79.315 147.055 ;
        RECT 77.265 145.415 77.435 145.915 ;
        RECT 63.765 144.505 63.980 145.015 ;
        RECT 64.210 144.685 64.490 145.015 ;
        RECT 64.670 144.505 64.910 145.015 ;
        RECT 65.245 144.505 70.590 145.050 ;
        RECT 70.765 144.505 76.110 145.050 ;
        RECT 76.780 144.675 77.395 145.245 ;
        RECT 77.685 145.185 77.950 145.745 ;
        RECT 78.120 145.015 78.290 145.915 ;
        RECT 79.485 145.905 79.815 146.885 ;
        RECT 79.985 145.915 80.215 147.055 ;
        RECT 80.425 145.965 81.635 147.055 ;
        RECT 78.460 145.185 78.815 145.745 ;
        RECT 77.565 144.505 77.780 145.015 ;
        RECT 78.010 144.685 78.290 145.015 ;
        RECT 78.470 144.505 78.710 145.015 ;
        RECT 79.105 144.505 79.315 145.325 ;
        RECT 79.485 145.305 79.735 145.905 ;
        RECT 79.905 145.495 80.235 145.745 ;
        RECT 79.485 144.675 79.815 145.305 ;
        RECT 79.985 144.505 80.215 145.325 ;
        RECT 80.425 145.255 80.945 145.795 ;
        RECT 81.115 145.425 81.635 145.965 ;
        RECT 81.805 145.890 82.095 147.055 ;
        RECT 82.265 145.965 85.775 147.055 ;
        RECT 85.945 145.965 87.155 147.055 ;
        RECT 87.385 145.995 87.715 146.840 ;
        RECT 87.885 146.045 88.055 147.055 ;
        RECT 88.225 146.325 88.565 146.885 ;
        RECT 88.795 146.555 89.110 147.055 ;
        RECT 89.290 146.585 90.175 146.755 ;
        RECT 82.265 145.275 83.915 145.795 ;
        RECT 84.085 145.445 85.775 145.965 ;
        RECT 80.425 144.505 81.635 145.255 ;
        RECT 81.805 144.505 82.095 145.230 ;
        RECT 82.265 144.505 85.775 145.275 ;
        RECT 85.945 145.255 86.465 145.795 ;
        RECT 86.635 145.425 87.155 145.965 ;
        RECT 87.325 145.915 87.715 145.995 ;
        RECT 88.225 145.950 89.120 146.325 ;
        RECT 87.325 145.865 87.540 145.915 ;
        RECT 87.325 145.285 87.495 145.865 ;
        RECT 88.225 145.745 88.415 145.950 ;
        RECT 89.290 145.745 89.460 146.585 ;
        RECT 90.400 146.555 90.650 146.885 ;
        RECT 87.665 145.415 88.415 145.745 ;
        RECT 88.585 145.415 89.460 145.745 ;
        RECT 85.945 144.505 87.155 145.255 ;
        RECT 87.325 145.245 87.550 145.285 ;
        RECT 88.215 145.245 88.415 145.415 ;
        RECT 87.325 145.160 87.705 145.245 ;
        RECT 87.375 144.725 87.705 145.160 ;
        RECT 87.875 144.505 88.045 145.115 ;
        RECT 88.215 144.720 88.545 145.245 ;
        RECT 88.805 144.505 89.015 145.035 ;
        RECT 89.290 144.955 89.460 145.415 ;
        RECT 89.630 145.455 89.950 146.415 ;
        RECT 90.120 145.665 90.310 146.385 ;
        RECT 90.480 145.485 90.650 146.555 ;
        RECT 90.820 146.255 90.990 147.055 ;
        RECT 91.160 146.610 92.265 146.780 ;
        RECT 91.160 145.995 91.330 146.610 ;
        RECT 92.475 146.460 92.725 146.885 ;
        RECT 92.895 146.595 93.160 147.055 ;
        RECT 91.500 146.075 92.030 146.440 ;
        RECT 92.475 146.330 92.780 146.460 ;
        RECT 90.820 145.905 91.330 145.995 ;
        RECT 90.820 145.735 91.690 145.905 ;
        RECT 90.820 145.665 90.990 145.735 ;
        RECT 91.110 145.485 91.310 145.515 ;
        RECT 89.630 145.125 90.095 145.455 ;
        RECT 90.480 145.185 91.310 145.485 ;
        RECT 90.480 144.955 90.650 145.185 ;
        RECT 89.290 144.785 90.075 144.955 ;
        RECT 90.245 144.785 90.650 144.955 ;
        RECT 90.830 144.505 91.200 145.005 ;
        RECT 91.520 144.955 91.690 145.735 ;
        RECT 91.860 145.375 92.030 146.075 ;
        RECT 92.200 145.545 92.440 146.140 ;
        RECT 91.860 145.155 92.385 145.375 ;
        RECT 92.610 145.225 92.780 146.330 ;
        RECT 92.555 145.095 92.780 145.225 ;
        RECT 92.950 145.135 93.230 146.085 ;
        RECT 92.555 144.955 92.725 145.095 ;
        RECT 91.520 144.785 92.195 144.955 ;
        RECT 92.390 144.785 92.725 144.955 ;
        RECT 92.895 144.505 93.145 144.965 ;
        RECT 93.400 144.765 93.585 146.885 ;
        RECT 93.755 146.555 94.085 147.055 ;
        RECT 94.255 146.385 94.425 146.885 ;
        RECT 93.760 146.215 94.425 146.385 ;
        RECT 94.775 146.385 94.945 146.885 ;
        RECT 95.115 146.555 95.445 147.055 ;
        RECT 94.775 146.215 95.440 146.385 ;
        RECT 93.760 145.225 93.990 146.215 ;
        RECT 94.160 145.395 94.510 146.045 ;
        RECT 94.690 145.395 95.040 146.045 ;
        RECT 95.210 145.225 95.440 146.215 ;
        RECT 93.760 145.055 94.425 145.225 ;
        RECT 93.755 144.505 94.085 144.885 ;
        RECT 94.255 144.765 94.425 145.055 ;
        RECT 94.775 145.055 95.440 145.225 ;
        RECT 94.775 144.765 94.945 145.055 ;
        RECT 95.115 144.505 95.445 144.885 ;
        RECT 95.615 144.765 95.800 146.885 ;
        RECT 96.040 146.595 96.305 147.055 ;
        RECT 96.475 146.460 96.725 146.885 ;
        RECT 96.935 146.610 98.040 146.780 ;
        RECT 96.420 146.330 96.725 146.460 ;
        RECT 95.970 145.135 96.250 146.085 ;
        RECT 96.420 145.225 96.590 146.330 ;
        RECT 96.760 145.545 97.000 146.140 ;
        RECT 97.170 146.075 97.700 146.440 ;
        RECT 97.170 145.375 97.340 146.075 ;
        RECT 97.870 145.995 98.040 146.610 ;
        RECT 98.210 146.255 98.380 147.055 ;
        RECT 98.550 146.555 98.800 146.885 ;
        RECT 99.025 146.585 99.910 146.755 ;
        RECT 97.870 145.905 98.380 145.995 ;
        RECT 96.420 145.095 96.645 145.225 ;
        RECT 96.815 145.155 97.340 145.375 ;
        RECT 97.510 145.735 98.380 145.905 ;
        RECT 96.055 144.505 96.305 144.965 ;
        RECT 96.475 144.955 96.645 145.095 ;
        RECT 97.510 144.955 97.680 145.735 ;
        RECT 98.210 145.665 98.380 145.735 ;
        RECT 97.890 145.485 98.090 145.515 ;
        RECT 98.550 145.485 98.720 146.555 ;
        RECT 98.890 145.665 99.080 146.385 ;
        RECT 97.890 145.185 98.720 145.485 ;
        RECT 99.250 145.455 99.570 146.415 ;
        RECT 96.475 144.785 96.810 144.955 ;
        RECT 97.005 144.785 97.680 144.955 ;
        RECT 98.000 144.505 98.370 145.005 ;
        RECT 98.550 144.955 98.720 145.185 ;
        RECT 99.105 145.125 99.570 145.455 ;
        RECT 99.740 145.745 99.910 146.585 ;
        RECT 100.090 146.555 100.405 147.055 ;
        RECT 100.635 146.325 100.975 146.885 ;
        RECT 100.080 145.950 100.975 146.325 ;
        RECT 101.145 146.045 101.315 147.055 ;
        RECT 100.785 145.745 100.975 145.950 ;
        RECT 101.485 145.995 101.815 146.840 ;
        RECT 103.080 146.425 103.365 146.885 ;
        RECT 103.535 146.595 103.805 147.055 ;
        RECT 103.080 146.205 104.035 146.425 ;
        RECT 101.485 145.915 101.875 145.995 ;
        RECT 101.660 145.865 101.875 145.915 ;
        RECT 99.740 145.415 100.615 145.745 ;
        RECT 100.785 145.415 101.535 145.745 ;
        RECT 99.740 144.955 99.910 145.415 ;
        RECT 100.785 145.245 100.985 145.415 ;
        RECT 101.705 145.285 101.875 145.865 ;
        RECT 102.965 145.475 103.655 146.035 ;
        RECT 103.825 145.305 104.035 146.205 ;
        RECT 101.650 145.245 101.875 145.285 ;
        RECT 98.550 144.785 98.955 144.955 ;
        RECT 99.125 144.785 99.910 144.955 ;
        RECT 100.185 144.505 100.395 145.035 ;
        RECT 100.655 144.720 100.985 145.245 ;
        RECT 101.495 145.160 101.875 145.245 ;
        RECT 101.155 144.505 101.325 145.115 ;
        RECT 101.495 144.725 101.825 145.160 ;
        RECT 103.080 145.135 104.035 145.305 ;
        RECT 104.205 146.035 104.605 146.885 ;
        RECT 104.795 146.425 105.075 146.885 ;
        RECT 105.595 146.595 105.920 147.055 ;
        RECT 104.795 146.205 105.920 146.425 ;
        RECT 104.205 145.475 105.300 146.035 ;
        RECT 105.470 145.745 105.920 146.205 ;
        RECT 106.090 145.915 106.475 146.885 ;
        RECT 103.080 144.675 103.365 145.135 ;
        RECT 103.535 144.505 103.805 144.965 ;
        RECT 104.205 144.675 104.605 145.475 ;
        RECT 105.470 145.415 106.025 145.745 ;
        RECT 105.470 145.305 105.920 145.415 ;
        RECT 104.795 145.135 105.920 145.305 ;
        RECT 106.195 145.245 106.475 145.915 ;
        RECT 107.565 145.890 107.855 147.055 ;
        RECT 108.085 145.995 108.415 146.840 ;
        RECT 108.585 146.045 108.755 147.055 ;
        RECT 108.925 146.325 109.265 146.885 ;
        RECT 109.495 146.555 109.810 147.055 ;
        RECT 109.990 146.585 110.875 146.755 ;
        RECT 108.025 145.915 108.415 145.995 ;
        RECT 108.925 145.950 109.820 146.325 ;
        RECT 104.795 144.675 105.075 145.135 ;
        RECT 105.595 144.505 105.920 144.965 ;
        RECT 106.090 144.675 106.475 145.245 ;
        RECT 108.025 145.865 108.240 145.915 ;
        RECT 108.025 145.285 108.195 145.865 ;
        RECT 108.925 145.745 109.115 145.950 ;
        RECT 109.990 145.745 110.160 146.585 ;
        RECT 111.100 146.555 111.350 146.885 ;
        RECT 108.365 145.415 109.115 145.745 ;
        RECT 109.285 145.415 110.160 145.745 ;
        RECT 108.025 145.245 108.250 145.285 ;
        RECT 108.915 145.245 109.115 145.415 ;
        RECT 107.565 144.505 107.855 145.230 ;
        RECT 108.025 145.160 108.405 145.245 ;
        RECT 108.075 144.725 108.405 145.160 ;
        RECT 108.575 144.505 108.745 145.115 ;
        RECT 108.915 144.720 109.245 145.245 ;
        RECT 109.505 144.505 109.715 145.035 ;
        RECT 109.990 144.955 110.160 145.415 ;
        RECT 110.330 145.455 110.650 146.415 ;
        RECT 110.820 145.665 111.010 146.385 ;
        RECT 111.180 145.485 111.350 146.555 ;
        RECT 111.520 146.255 111.690 147.055 ;
        RECT 111.860 146.610 112.965 146.780 ;
        RECT 111.860 145.995 112.030 146.610 ;
        RECT 113.175 146.460 113.425 146.885 ;
        RECT 113.595 146.595 113.860 147.055 ;
        RECT 112.200 146.075 112.730 146.440 ;
        RECT 113.175 146.330 113.480 146.460 ;
        RECT 111.520 145.905 112.030 145.995 ;
        RECT 111.520 145.735 112.390 145.905 ;
        RECT 111.520 145.665 111.690 145.735 ;
        RECT 111.810 145.485 112.010 145.515 ;
        RECT 110.330 145.125 110.795 145.455 ;
        RECT 111.180 145.185 112.010 145.485 ;
        RECT 111.180 144.955 111.350 145.185 ;
        RECT 109.990 144.785 110.775 144.955 ;
        RECT 110.945 144.785 111.350 144.955 ;
        RECT 111.530 144.505 111.900 145.005 ;
        RECT 112.220 144.955 112.390 145.735 ;
        RECT 112.560 145.375 112.730 146.075 ;
        RECT 112.900 145.545 113.140 146.140 ;
        RECT 112.560 145.155 113.085 145.375 ;
        RECT 113.310 145.225 113.480 146.330 ;
        RECT 113.255 145.095 113.480 145.225 ;
        RECT 113.650 145.135 113.930 146.085 ;
        RECT 113.255 144.955 113.425 145.095 ;
        RECT 112.220 144.785 112.895 144.955 ;
        RECT 113.090 144.785 113.425 144.955 ;
        RECT 113.595 144.505 113.845 144.965 ;
        RECT 114.100 144.765 114.285 146.885 ;
        RECT 114.455 146.555 114.785 147.055 ;
        RECT 114.955 146.385 115.125 146.885 ;
        RECT 114.460 146.215 115.125 146.385 ;
        RECT 114.460 145.225 114.690 146.215 ;
        RECT 114.860 145.395 115.210 146.045 ;
        RECT 115.390 145.915 115.725 146.885 ;
        RECT 115.895 145.915 116.065 147.055 ;
        RECT 116.235 146.715 118.265 146.885 ;
        RECT 115.390 145.245 115.560 145.915 ;
        RECT 116.235 145.745 116.405 146.715 ;
        RECT 115.730 145.415 115.985 145.745 ;
        RECT 116.210 145.415 116.405 145.745 ;
        RECT 116.575 146.375 117.700 146.545 ;
        RECT 115.815 145.245 115.985 145.415 ;
        RECT 116.575 145.245 116.745 146.375 ;
        RECT 114.460 145.055 115.125 145.225 ;
        RECT 114.455 144.505 114.785 144.885 ;
        RECT 114.955 144.765 115.125 145.055 ;
        RECT 115.390 144.675 115.645 145.245 ;
        RECT 115.815 145.075 116.745 145.245 ;
        RECT 116.915 146.035 117.925 146.205 ;
        RECT 116.915 145.235 117.085 146.035 ;
        RECT 116.570 145.040 116.745 145.075 ;
        RECT 115.815 144.505 116.145 144.905 ;
        RECT 116.570 144.675 117.100 145.040 ;
        RECT 117.290 145.015 117.565 145.835 ;
        RECT 117.285 144.845 117.565 145.015 ;
        RECT 117.290 144.675 117.565 144.845 ;
        RECT 117.735 144.675 117.925 146.035 ;
        RECT 118.095 146.050 118.265 146.715 ;
        RECT 118.435 146.295 118.605 147.055 ;
        RECT 118.840 146.295 119.355 146.705 ;
        RECT 118.095 145.860 118.845 146.050 ;
        RECT 119.015 145.485 119.355 146.295 ;
        RECT 119.640 146.425 119.925 146.885 ;
        RECT 120.095 146.595 120.365 147.055 ;
        RECT 119.640 146.205 120.595 146.425 ;
        RECT 118.125 145.315 119.355 145.485 ;
        RECT 119.525 145.475 120.215 146.035 ;
        RECT 118.105 144.505 118.615 145.040 ;
        RECT 118.835 144.710 119.080 145.315 ;
        RECT 120.385 145.305 120.595 146.205 ;
        RECT 119.640 145.135 120.595 145.305 ;
        RECT 120.765 146.035 121.165 146.885 ;
        RECT 121.355 146.425 121.635 146.885 ;
        RECT 122.155 146.595 122.480 147.055 ;
        RECT 121.355 146.205 122.480 146.425 ;
        RECT 120.765 145.475 121.860 146.035 ;
        RECT 122.030 145.745 122.480 146.205 ;
        RECT 122.650 145.915 123.035 146.885 ;
        RECT 123.210 146.255 123.465 147.055 ;
        RECT 123.665 146.205 123.995 146.885 ;
        RECT 119.640 144.675 119.925 145.135 ;
        RECT 120.095 144.505 120.365 144.965 ;
        RECT 120.765 144.675 121.165 145.475 ;
        RECT 122.030 145.415 122.585 145.745 ;
        RECT 122.030 145.305 122.480 145.415 ;
        RECT 121.355 145.135 122.480 145.305 ;
        RECT 122.755 145.245 123.035 145.915 ;
        RECT 123.210 145.715 123.455 146.075 ;
        RECT 123.645 145.925 123.995 146.205 ;
        RECT 123.645 145.545 123.815 145.925 ;
        RECT 124.175 145.745 124.370 146.795 ;
        RECT 124.550 145.915 124.870 147.055 ;
        RECT 125.050 145.915 125.385 146.885 ;
        RECT 125.555 145.915 125.725 147.055 ;
        RECT 125.895 146.715 127.925 146.885 ;
        RECT 121.355 144.675 121.635 145.135 ;
        RECT 122.155 144.505 122.480 144.965 ;
        RECT 122.650 144.675 123.035 145.245 ;
        RECT 123.295 145.375 123.815 145.545 ;
        RECT 123.985 145.415 124.370 145.745 ;
        RECT 124.550 145.695 124.810 145.745 ;
        RECT 124.550 145.525 124.815 145.695 ;
        RECT 124.550 145.415 124.810 145.525 ;
        RECT 123.295 144.810 123.465 145.375 ;
        RECT 125.050 145.245 125.220 145.915 ;
        RECT 125.895 145.745 126.065 146.715 ;
        RECT 125.390 145.415 125.645 145.745 ;
        RECT 125.870 145.415 126.065 145.745 ;
        RECT 126.235 146.375 127.360 146.545 ;
        RECT 125.475 145.245 125.645 145.415 ;
        RECT 126.235 145.245 126.405 146.375 ;
        RECT 123.655 145.035 124.870 145.205 ;
        RECT 123.655 144.730 123.885 145.035 ;
        RECT 124.055 144.505 124.385 144.865 ;
        RECT 124.580 144.685 124.870 145.035 ;
        RECT 125.050 144.675 125.305 145.245 ;
        RECT 125.475 145.075 126.405 145.245 ;
        RECT 126.575 146.035 127.585 146.205 ;
        RECT 126.575 145.235 126.745 146.035 ;
        RECT 126.230 145.040 126.405 145.075 ;
        RECT 125.475 144.505 125.805 144.905 ;
        RECT 126.230 144.675 126.760 145.040 ;
        RECT 126.950 145.015 127.225 145.835 ;
        RECT 126.945 144.845 127.225 145.015 ;
        RECT 126.950 144.675 127.225 144.845 ;
        RECT 127.395 144.675 127.585 146.035 ;
        RECT 127.755 146.050 127.925 146.715 ;
        RECT 128.095 146.295 128.265 147.055 ;
        RECT 128.500 146.295 129.015 146.705 ;
        RECT 127.755 145.860 128.505 146.050 ;
        RECT 128.675 145.485 129.015 146.295 ;
        RECT 127.785 145.315 129.015 145.485 ;
        RECT 129.185 145.915 129.570 146.885 ;
        RECT 129.740 146.595 130.065 147.055 ;
        RECT 130.585 146.425 130.865 146.885 ;
        RECT 129.740 146.205 130.865 146.425 ;
        RECT 127.765 144.505 128.275 145.040 ;
        RECT 128.495 144.710 128.740 145.315 ;
        RECT 129.185 145.245 129.465 145.915 ;
        RECT 129.740 145.745 130.190 146.205 ;
        RECT 131.055 146.035 131.455 146.885 ;
        RECT 131.855 146.595 132.125 147.055 ;
        RECT 132.295 146.425 132.580 146.885 ;
        RECT 129.635 145.415 130.190 145.745 ;
        RECT 130.360 145.475 131.455 146.035 ;
        RECT 129.740 145.305 130.190 145.415 ;
        RECT 129.185 144.675 129.570 145.245 ;
        RECT 129.740 145.135 130.865 145.305 ;
        RECT 129.740 144.505 130.065 144.965 ;
        RECT 130.585 144.675 130.865 145.135 ;
        RECT 131.055 144.675 131.455 145.475 ;
        RECT 131.625 146.205 132.580 146.425 ;
        RECT 131.625 145.305 131.835 146.205 ;
        RECT 132.005 145.475 132.695 146.035 ;
        RECT 133.325 145.890 133.615 147.055 ;
        RECT 134.335 146.385 134.505 146.885 ;
        RECT 134.675 146.555 135.005 147.055 ;
        RECT 134.335 146.215 135.000 146.385 ;
        RECT 134.250 145.395 134.600 146.045 ;
        RECT 131.625 145.135 132.580 145.305 ;
        RECT 131.855 144.505 132.125 144.965 ;
        RECT 132.295 144.675 132.580 145.135 ;
        RECT 133.325 144.505 133.615 145.230 ;
        RECT 134.770 145.225 135.000 146.215 ;
        RECT 134.335 145.055 135.000 145.225 ;
        RECT 134.335 144.765 134.505 145.055 ;
        RECT 134.675 144.505 135.005 144.885 ;
        RECT 135.175 144.765 135.360 146.885 ;
        RECT 135.600 146.595 135.865 147.055 ;
        RECT 136.035 146.460 136.285 146.885 ;
        RECT 136.495 146.610 137.600 146.780 ;
        RECT 135.980 146.330 136.285 146.460 ;
        RECT 135.530 145.135 135.810 146.085 ;
        RECT 135.980 145.225 136.150 146.330 ;
        RECT 136.320 145.545 136.560 146.140 ;
        RECT 136.730 146.075 137.260 146.440 ;
        RECT 136.730 145.375 136.900 146.075 ;
        RECT 137.430 145.995 137.600 146.610 ;
        RECT 137.770 146.255 137.940 147.055 ;
        RECT 138.110 146.555 138.360 146.885 ;
        RECT 138.585 146.585 139.470 146.755 ;
        RECT 137.430 145.905 137.940 145.995 ;
        RECT 135.980 145.095 136.205 145.225 ;
        RECT 136.375 145.155 136.900 145.375 ;
        RECT 137.070 145.735 137.940 145.905 ;
        RECT 135.615 144.505 135.865 144.965 ;
        RECT 136.035 144.955 136.205 145.095 ;
        RECT 137.070 144.955 137.240 145.735 ;
        RECT 137.770 145.665 137.940 145.735 ;
        RECT 137.450 145.485 137.650 145.515 ;
        RECT 138.110 145.485 138.280 146.555 ;
        RECT 138.450 145.665 138.640 146.385 ;
        RECT 137.450 145.185 138.280 145.485 ;
        RECT 138.810 145.455 139.130 146.415 ;
        RECT 136.035 144.785 136.370 144.955 ;
        RECT 136.565 144.785 137.240 144.955 ;
        RECT 137.560 144.505 137.930 145.005 ;
        RECT 138.110 144.955 138.280 145.185 ;
        RECT 138.665 145.125 139.130 145.455 ;
        RECT 139.300 145.745 139.470 146.585 ;
        RECT 139.650 146.555 139.965 147.055 ;
        RECT 140.195 146.325 140.535 146.885 ;
        RECT 139.640 145.950 140.535 146.325 ;
        RECT 140.705 146.045 140.875 147.055 ;
        RECT 140.345 145.745 140.535 145.950 ;
        RECT 141.045 145.995 141.375 146.840 ;
        RECT 142.180 146.425 142.465 146.885 ;
        RECT 142.635 146.595 142.905 147.055 ;
        RECT 142.180 146.205 143.135 146.425 ;
        RECT 141.045 145.915 141.435 145.995 ;
        RECT 141.220 145.865 141.435 145.915 ;
        RECT 139.300 145.415 140.175 145.745 ;
        RECT 140.345 145.415 141.095 145.745 ;
        RECT 139.300 144.955 139.470 145.415 ;
        RECT 140.345 145.245 140.545 145.415 ;
        RECT 141.265 145.285 141.435 145.865 ;
        RECT 142.065 145.475 142.755 146.035 ;
        RECT 142.925 145.305 143.135 146.205 ;
        RECT 141.210 145.245 141.435 145.285 ;
        RECT 138.110 144.785 138.515 144.955 ;
        RECT 138.685 144.785 139.470 144.955 ;
        RECT 139.745 144.505 139.955 145.035 ;
        RECT 140.215 144.720 140.545 145.245 ;
        RECT 141.055 145.160 141.435 145.245 ;
        RECT 140.715 144.505 140.885 145.115 ;
        RECT 141.055 144.725 141.385 145.160 ;
        RECT 142.180 145.135 143.135 145.305 ;
        RECT 143.305 146.035 143.705 146.885 ;
        RECT 143.895 146.425 144.175 146.885 ;
        RECT 144.695 146.595 145.020 147.055 ;
        RECT 143.895 146.205 145.020 146.425 ;
        RECT 143.305 145.475 144.400 146.035 ;
        RECT 144.570 145.745 145.020 146.205 ;
        RECT 145.190 145.915 145.575 146.885 ;
        RECT 142.180 144.675 142.465 145.135 ;
        RECT 142.635 144.505 142.905 144.965 ;
        RECT 143.305 144.675 143.705 145.475 ;
        RECT 144.570 145.415 145.125 145.745 ;
        RECT 144.570 145.305 145.020 145.415 ;
        RECT 143.895 145.135 145.020 145.305 ;
        RECT 145.295 145.245 145.575 145.915 ;
        RECT 145.745 145.965 146.955 147.055 ;
        RECT 145.745 145.425 146.265 145.965 ;
        RECT 146.435 145.255 146.955 145.795 ;
        RECT 143.895 144.675 144.175 145.135 ;
        RECT 144.695 144.505 145.020 144.965 ;
        RECT 145.190 144.675 145.575 145.245 ;
        RECT 145.745 144.505 146.955 145.255 ;
        RECT 17.320 144.335 147.040 144.505 ;
        RECT 17.405 143.585 18.615 144.335 ;
        RECT 18.785 143.790 24.130 144.335 ;
        RECT 24.305 143.790 29.650 144.335 ;
        RECT 17.405 143.045 17.925 143.585 ;
        RECT 18.095 142.875 18.615 143.415 ;
        RECT 20.370 142.960 20.710 143.790 ;
        RECT 17.405 141.785 18.615 142.875 ;
        RECT 22.190 142.220 22.540 143.470 ;
        RECT 25.890 142.960 26.230 143.790 ;
        RECT 29.825 143.565 31.495 144.335 ;
        RECT 32.130 143.830 32.465 144.335 ;
        RECT 32.635 143.765 32.875 144.140 ;
        RECT 33.155 144.005 33.325 144.150 ;
        RECT 33.155 143.810 33.530 144.005 ;
        RECT 33.890 143.840 34.285 144.335 ;
        RECT 27.710 142.220 28.060 143.470 ;
        RECT 29.825 143.045 30.575 143.565 ;
        RECT 30.745 142.875 31.495 143.395 ;
        RECT 18.785 141.785 24.130 142.220 ;
        RECT 24.305 141.785 29.650 142.220 ;
        RECT 29.825 141.785 31.495 142.875 ;
        RECT 32.185 142.805 32.485 143.655 ;
        RECT 32.655 143.615 32.875 143.765 ;
        RECT 32.655 143.285 33.190 143.615 ;
        RECT 33.360 143.475 33.530 143.810 ;
        RECT 34.455 143.645 34.695 144.165 ;
        RECT 32.655 142.635 32.890 143.285 ;
        RECT 33.360 143.115 34.345 143.475 ;
        RECT 32.215 142.405 32.890 142.635 ;
        RECT 33.060 143.095 34.345 143.115 ;
        RECT 33.060 142.945 33.920 143.095 ;
        RECT 32.215 141.975 32.385 142.405 ;
        RECT 32.555 141.785 32.885 142.235 ;
        RECT 33.060 142.000 33.345 142.945 ;
        RECT 34.520 142.840 34.695 143.645 ;
        RECT 35.825 143.605 36.115 144.335 ;
        RECT 35.815 143.095 36.115 143.425 ;
        RECT 36.295 143.405 36.525 144.045 ;
        RECT 36.705 143.785 37.015 144.155 ;
        RECT 37.195 143.965 37.865 144.335 ;
        RECT 36.705 143.585 37.935 143.785 ;
        RECT 36.295 143.095 36.820 143.405 ;
        RECT 37.000 143.095 37.465 143.405 ;
        RECT 37.645 142.915 37.935 143.585 ;
        RECT 33.520 142.465 34.215 142.775 ;
        RECT 33.525 141.785 34.210 142.255 ;
        RECT 34.390 142.055 34.695 142.840 ;
        RECT 35.825 142.675 36.985 142.915 ;
        RECT 35.825 141.965 36.085 142.675 ;
        RECT 36.255 141.785 36.585 142.495 ;
        RECT 36.755 141.965 36.985 142.675 ;
        RECT 37.165 142.695 37.935 142.915 ;
        RECT 37.165 141.965 37.435 142.695 ;
        RECT 37.615 141.785 37.955 142.515 ;
        RECT 38.125 141.965 38.385 144.155 ;
        RECT 38.565 143.615 38.905 144.125 ;
        RECT 38.565 142.215 38.825 143.615 ;
        RECT 39.075 143.535 39.345 144.335 ;
        RECT 39.000 143.095 39.330 143.345 ;
        RECT 39.525 143.095 39.805 144.065 ;
        RECT 39.985 143.095 40.285 144.065 ;
        RECT 40.465 143.095 40.815 144.060 ;
        RECT 41.035 143.835 41.530 144.165 ;
        RECT 39.015 142.925 39.330 143.095 ;
        RECT 41.035 142.925 41.205 143.835 ;
        RECT 39.015 142.755 41.205 142.925 ;
        RECT 38.565 141.955 38.905 142.215 ;
        RECT 39.075 141.785 39.405 142.585 ;
        RECT 39.870 141.955 40.120 142.755 ;
        RECT 40.305 141.785 40.635 142.505 ;
        RECT 40.855 141.955 41.105 142.755 ;
        RECT 41.375 142.345 41.615 143.655 ;
        RECT 41.785 143.585 42.995 144.335 ;
        RECT 43.165 143.610 43.455 144.335 ;
        RECT 43.625 143.790 48.970 144.335 ;
        RECT 49.145 143.790 54.490 144.335 ;
        RECT 41.785 143.045 42.305 143.585 ;
        RECT 42.475 142.875 42.995 143.415 ;
        RECT 45.210 142.960 45.550 143.790 ;
        RECT 41.275 141.785 41.610 142.165 ;
        RECT 41.785 141.785 42.995 142.875 ;
        RECT 43.165 141.785 43.455 142.950 ;
        RECT 47.030 142.220 47.380 143.470 ;
        RECT 50.730 142.960 51.070 143.790 ;
        RECT 54.665 143.535 55.360 144.165 ;
        RECT 55.565 143.535 55.875 144.335 ;
        RECT 52.550 142.220 52.900 143.470 ;
        RECT 54.685 143.095 55.020 143.345 ;
        RECT 55.190 142.935 55.360 143.535 ;
        RECT 56.505 143.515 56.765 144.335 ;
        RECT 56.935 143.515 57.265 143.935 ;
        RECT 57.445 143.850 58.235 144.115 ;
        RECT 57.015 143.425 57.265 143.515 ;
        RECT 55.530 143.095 55.865 143.365 ;
        RECT 43.625 141.785 48.970 142.220 ;
        RECT 49.145 141.785 54.490 142.220 ;
        RECT 54.665 141.785 54.925 142.925 ;
        RECT 55.095 141.955 55.425 142.935 ;
        RECT 55.595 141.785 55.875 142.925 ;
        RECT 56.505 142.465 56.845 143.345 ;
        RECT 57.015 143.175 57.810 143.425 ;
        RECT 56.505 141.785 56.765 142.295 ;
        RECT 57.015 141.955 57.185 143.175 ;
        RECT 57.980 142.995 58.235 143.850 ;
        RECT 58.405 143.695 58.605 144.115 ;
        RECT 58.795 143.875 59.125 144.335 ;
        RECT 58.405 143.175 58.815 143.695 ;
        RECT 59.295 143.685 59.555 144.165 ;
        RECT 58.985 142.995 59.215 143.425 ;
        RECT 57.425 142.825 59.215 142.995 ;
        RECT 57.425 142.460 57.675 142.825 ;
        RECT 57.845 142.465 58.175 142.655 ;
        RECT 58.395 142.530 59.110 142.825 ;
        RECT 59.385 142.655 59.555 143.685 ;
        RECT 60.275 143.785 60.445 144.075 ;
        RECT 60.615 143.955 60.945 144.335 ;
        RECT 60.275 143.615 60.940 143.785 ;
        RECT 60.190 142.795 60.540 143.445 ;
        RECT 57.845 142.290 58.040 142.465 ;
        RECT 57.425 141.785 58.040 142.290 ;
        RECT 58.210 141.955 58.685 142.295 ;
        RECT 58.855 141.785 59.070 142.330 ;
        RECT 59.280 141.955 59.555 142.655 ;
        RECT 60.710 142.625 60.940 143.615 ;
        RECT 60.275 142.455 60.940 142.625 ;
        RECT 60.275 141.955 60.445 142.455 ;
        RECT 60.615 141.785 60.945 142.285 ;
        RECT 61.115 141.955 61.300 144.075 ;
        RECT 61.555 143.875 61.805 144.335 ;
        RECT 61.975 143.885 62.310 144.055 ;
        RECT 62.505 143.885 63.180 144.055 ;
        RECT 61.975 143.745 62.145 143.885 ;
        RECT 61.470 142.755 61.750 143.705 ;
        RECT 61.920 143.615 62.145 143.745 ;
        RECT 61.920 142.510 62.090 143.615 ;
        RECT 62.315 143.465 62.840 143.685 ;
        RECT 62.260 142.700 62.500 143.295 ;
        RECT 62.670 142.765 62.840 143.465 ;
        RECT 63.010 143.105 63.180 143.885 ;
        RECT 63.500 143.835 63.870 144.335 ;
        RECT 64.050 143.885 64.455 144.055 ;
        RECT 64.625 143.885 65.410 144.055 ;
        RECT 64.050 143.655 64.220 143.885 ;
        RECT 63.390 143.355 64.220 143.655 ;
        RECT 64.605 143.385 65.070 143.715 ;
        RECT 63.390 143.325 63.590 143.355 ;
        RECT 63.710 143.105 63.880 143.175 ;
        RECT 63.010 142.935 63.880 143.105 ;
        RECT 63.370 142.845 63.880 142.935 ;
        RECT 61.920 142.380 62.225 142.510 ;
        RECT 62.670 142.400 63.200 142.765 ;
        RECT 61.540 141.785 61.805 142.245 ;
        RECT 61.975 141.955 62.225 142.380 ;
        RECT 63.370 142.230 63.540 142.845 ;
        RECT 62.435 142.060 63.540 142.230 ;
        RECT 63.710 141.785 63.880 142.585 ;
        RECT 64.050 142.285 64.220 143.355 ;
        RECT 64.390 142.455 64.580 143.175 ;
        RECT 64.750 142.425 65.070 143.385 ;
        RECT 65.240 143.425 65.410 143.885 ;
        RECT 65.685 143.805 65.895 144.335 ;
        RECT 66.155 143.595 66.485 144.120 ;
        RECT 66.655 143.725 66.825 144.335 ;
        RECT 66.995 143.680 67.325 144.115 ;
        RECT 66.995 143.595 67.375 143.680 ;
        RECT 66.285 143.425 66.485 143.595 ;
        RECT 67.150 143.555 67.375 143.595 ;
        RECT 65.240 143.095 66.115 143.425 ;
        RECT 66.285 143.095 67.035 143.425 ;
        RECT 64.050 141.955 64.300 142.285 ;
        RECT 65.240 142.255 65.410 143.095 ;
        RECT 66.285 142.890 66.475 143.095 ;
        RECT 67.205 142.975 67.375 143.555 ;
        RECT 67.545 143.585 68.755 144.335 ;
        RECT 68.925 143.610 69.215 144.335 ;
        RECT 67.545 143.045 68.065 143.585 ;
        RECT 69.385 143.565 71.975 144.335 ;
        RECT 67.160 142.925 67.375 142.975 ;
        RECT 65.580 142.515 66.475 142.890 ;
        RECT 66.985 142.845 67.375 142.925 ;
        RECT 68.235 142.875 68.755 143.415 ;
        RECT 69.385 143.045 70.595 143.565 ;
        RECT 72.145 143.535 72.455 144.335 ;
        RECT 72.660 143.535 73.355 144.165 ;
        RECT 64.525 142.085 65.410 142.255 ;
        RECT 65.590 141.785 65.905 142.285 ;
        RECT 66.135 141.955 66.475 142.515 ;
        RECT 66.645 141.785 66.815 142.795 ;
        RECT 66.985 142.000 67.315 142.845 ;
        RECT 67.545 141.785 68.755 142.875 ;
        RECT 68.925 141.785 69.215 142.950 ;
        RECT 70.765 142.875 71.975 143.395 ;
        RECT 72.155 143.095 72.490 143.365 ;
        RECT 72.660 142.975 72.830 143.535 ;
        RECT 73.525 143.390 73.865 144.165 ;
        RECT 74.035 143.875 74.205 144.335 ;
        RECT 74.445 143.900 74.805 144.165 ;
        RECT 74.445 143.895 74.800 143.900 ;
        RECT 74.445 143.885 74.795 143.895 ;
        RECT 74.445 143.880 74.790 143.885 ;
        RECT 74.445 143.870 74.785 143.880 ;
        RECT 75.435 143.875 75.605 144.335 ;
        RECT 74.445 143.865 74.780 143.870 ;
        RECT 74.445 143.855 74.770 143.865 ;
        RECT 74.445 143.845 74.760 143.855 ;
        RECT 74.445 143.705 74.745 143.845 ;
        RECT 74.035 143.515 74.745 143.705 ;
        RECT 74.935 143.705 75.265 143.785 ;
        RECT 75.775 143.705 76.115 144.165 ;
        RECT 74.935 143.515 76.115 143.705 ;
        RECT 76.750 143.595 77.005 144.165 ;
        RECT 77.175 143.935 77.505 144.335 ;
        RECT 77.930 143.800 78.460 144.165 ;
        RECT 78.650 143.995 78.925 144.165 ;
        RECT 78.645 143.825 78.925 143.995 ;
        RECT 77.930 143.765 78.105 143.800 ;
        RECT 77.175 143.595 78.105 143.765 ;
        RECT 73.000 143.095 73.335 143.345 ;
        RECT 72.660 142.935 72.835 142.975 ;
        RECT 69.385 141.785 71.975 142.875 ;
        RECT 72.145 141.785 72.425 142.925 ;
        RECT 72.595 141.955 72.925 142.935 ;
        RECT 73.095 141.785 73.355 142.925 ;
        RECT 73.525 141.955 73.805 143.390 ;
        RECT 74.035 142.945 74.320 143.515 ;
        RECT 74.505 143.115 74.975 143.345 ;
        RECT 75.145 143.325 75.475 143.345 ;
        RECT 75.145 143.145 75.595 143.325 ;
        RECT 75.785 143.145 76.115 143.345 ;
        RECT 74.035 142.730 75.185 142.945 ;
        RECT 73.975 141.785 74.685 142.560 ;
        RECT 74.855 141.955 75.185 142.730 ;
        RECT 75.380 142.030 75.595 143.145 ;
        RECT 75.885 142.805 76.115 143.145 ;
        RECT 76.750 142.925 76.920 143.595 ;
        RECT 77.175 143.425 77.345 143.595 ;
        RECT 77.090 143.095 77.345 143.425 ;
        RECT 77.570 143.095 77.765 143.425 ;
        RECT 75.775 141.785 76.105 142.505 ;
        RECT 76.750 141.955 77.085 142.925 ;
        RECT 77.255 141.785 77.425 142.925 ;
        RECT 77.595 142.125 77.765 143.095 ;
        RECT 77.935 142.465 78.105 143.595 ;
        RECT 78.275 142.805 78.445 143.605 ;
        RECT 78.650 143.005 78.925 143.825 ;
        RECT 79.095 142.805 79.285 144.165 ;
        RECT 79.465 143.800 79.975 144.335 ;
        RECT 80.195 143.525 80.440 144.130 ;
        RECT 81.515 143.820 81.685 144.335 ;
        RECT 81.855 143.680 82.185 144.115 ;
        RECT 82.355 143.725 82.525 144.335 ;
        RECT 81.805 143.595 82.185 143.680 ;
        RECT 82.695 143.595 83.025 144.120 ;
        RECT 83.285 143.805 83.495 144.335 ;
        RECT 83.770 143.885 84.555 144.055 ;
        RECT 84.725 143.885 85.130 144.055 ;
        RECT 81.805 143.555 82.030 143.595 ;
        RECT 79.485 143.355 80.715 143.525 ;
        RECT 78.275 142.635 79.285 142.805 ;
        RECT 79.455 142.790 80.205 142.980 ;
        RECT 77.935 142.295 79.060 142.465 ;
        RECT 79.455 142.125 79.625 142.790 ;
        RECT 80.375 142.545 80.715 143.355 ;
        RECT 81.805 142.975 81.975 143.555 ;
        RECT 82.695 143.425 82.895 143.595 ;
        RECT 83.770 143.425 83.940 143.885 ;
        RECT 82.145 143.095 82.895 143.425 ;
        RECT 83.065 143.095 83.940 143.425 ;
        RECT 81.805 142.925 82.020 142.975 ;
        RECT 81.805 142.845 82.195 142.925 ;
        RECT 77.595 141.955 79.625 142.125 ;
        RECT 79.795 141.785 79.965 142.545 ;
        RECT 80.200 142.135 80.715 142.545 ;
        RECT 81.525 141.785 81.695 142.700 ;
        RECT 81.865 142.000 82.195 142.845 ;
        RECT 82.705 142.890 82.895 143.095 ;
        RECT 82.365 141.785 82.535 142.795 ;
        RECT 82.705 142.515 83.600 142.890 ;
        RECT 82.705 141.955 83.045 142.515 ;
        RECT 83.275 141.785 83.590 142.285 ;
        RECT 83.770 142.255 83.940 143.095 ;
        RECT 84.110 143.385 84.575 143.715 ;
        RECT 84.960 143.655 85.130 143.885 ;
        RECT 85.310 143.835 85.680 144.335 ;
        RECT 86.000 143.885 86.675 144.055 ;
        RECT 86.870 143.885 87.205 144.055 ;
        RECT 84.110 142.425 84.430 143.385 ;
        RECT 84.960 143.355 85.790 143.655 ;
        RECT 84.600 142.455 84.790 143.175 ;
        RECT 84.960 142.285 85.130 143.355 ;
        RECT 85.590 143.325 85.790 143.355 ;
        RECT 85.300 143.105 85.470 143.175 ;
        RECT 86.000 143.105 86.170 143.885 ;
        RECT 87.035 143.745 87.205 143.885 ;
        RECT 87.375 143.875 87.625 144.335 ;
        RECT 85.300 142.935 86.170 143.105 ;
        RECT 86.340 143.465 86.865 143.685 ;
        RECT 87.035 143.615 87.260 143.745 ;
        RECT 85.300 142.845 85.810 142.935 ;
        RECT 83.770 142.085 84.655 142.255 ;
        RECT 84.880 141.955 85.130 142.285 ;
        RECT 85.300 141.785 85.470 142.585 ;
        RECT 85.640 142.230 85.810 142.845 ;
        RECT 86.340 142.765 86.510 143.465 ;
        RECT 85.980 142.400 86.510 142.765 ;
        RECT 86.680 142.700 86.920 143.295 ;
        RECT 87.090 142.510 87.260 143.615 ;
        RECT 87.430 142.755 87.710 143.705 ;
        RECT 86.955 142.380 87.260 142.510 ;
        RECT 85.640 142.060 86.745 142.230 ;
        RECT 86.955 141.955 87.205 142.380 ;
        RECT 87.375 141.785 87.640 142.245 ;
        RECT 87.880 141.955 88.065 144.075 ;
        RECT 88.235 143.955 88.565 144.335 ;
        RECT 88.735 143.785 88.905 144.075 ;
        RECT 88.240 143.615 88.905 143.785 ;
        RECT 88.240 142.625 88.470 143.615 ;
        RECT 89.165 143.565 91.755 144.335 ;
        RECT 88.640 142.795 88.990 143.445 ;
        RECT 89.165 143.045 90.375 143.565 ;
        RECT 90.545 142.875 91.755 143.395 ;
        RECT 88.240 142.455 88.905 142.625 ;
        RECT 88.235 141.785 88.565 142.285 ;
        RECT 88.735 141.955 88.905 142.455 ;
        RECT 89.165 141.785 91.755 142.875 ;
        RECT 91.925 143.390 92.265 144.165 ;
        RECT 92.435 143.875 92.605 144.335 ;
        RECT 92.845 143.900 93.205 144.165 ;
        RECT 92.845 143.895 93.200 143.900 ;
        RECT 92.845 143.885 93.195 143.895 ;
        RECT 92.845 143.880 93.190 143.885 ;
        RECT 92.845 143.870 93.185 143.880 ;
        RECT 93.835 143.875 94.005 144.335 ;
        RECT 92.845 143.865 93.180 143.870 ;
        RECT 92.845 143.855 93.170 143.865 ;
        RECT 92.845 143.845 93.160 143.855 ;
        RECT 92.845 143.705 93.145 143.845 ;
        RECT 92.435 143.515 93.145 143.705 ;
        RECT 93.335 143.705 93.665 143.785 ;
        RECT 94.175 143.705 94.515 144.165 ;
        RECT 93.335 143.515 94.515 143.705 ;
        RECT 94.685 143.610 94.975 144.335 ;
        RECT 95.145 143.595 95.530 144.165 ;
        RECT 95.700 143.875 96.025 144.335 ;
        RECT 96.545 143.705 96.825 144.165 ;
        RECT 91.925 141.955 92.205 143.390 ;
        RECT 92.435 142.945 92.720 143.515 ;
        RECT 92.905 143.115 93.375 143.345 ;
        RECT 93.545 143.325 93.875 143.345 ;
        RECT 93.545 143.145 93.995 143.325 ;
        RECT 94.185 143.145 94.515 143.345 ;
        RECT 92.435 142.730 93.585 142.945 ;
        RECT 92.375 141.785 93.085 142.560 ;
        RECT 93.255 141.955 93.585 142.730 ;
        RECT 93.780 142.030 93.995 143.145 ;
        RECT 94.285 142.805 94.515 143.145 ;
        RECT 94.175 141.785 94.505 142.505 ;
        RECT 94.685 141.785 94.975 142.950 ;
        RECT 95.145 142.925 95.425 143.595 ;
        RECT 95.700 143.535 96.825 143.705 ;
        RECT 95.700 143.425 96.150 143.535 ;
        RECT 95.595 143.095 96.150 143.425 ;
        RECT 97.015 143.365 97.415 144.165 ;
        RECT 97.815 143.875 98.085 144.335 ;
        RECT 98.255 143.705 98.540 144.165 ;
        RECT 95.145 141.955 95.530 142.925 ;
        RECT 95.700 142.635 96.150 143.095 ;
        RECT 96.320 142.805 97.415 143.365 ;
        RECT 95.700 142.415 96.825 142.635 ;
        RECT 95.700 141.785 96.025 142.245 ;
        RECT 96.545 141.955 96.825 142.415 ;
        RECT 97.015 141.955 97.415 142.805 ;
        RECT 97.585 143.535 98.540 143.705 ;
        RECT 98.825 143.585 100.035 144.335 ;
        RECT 100.320 143.705 100.605 144.165 ;
        RECT 100.775 143.875 101.045 144.335 ;
        RECT 97.585 142.635 97.795 143.535 ;
        RECT 97.965 142.805 98.655 143.365 ;
        RECT 98.825 143.045 99.345 143.585 ;
        RECT 100.320 143.535 101.275 143.705 ;
        RECT 99.515 142.875 100.035 143.415 ;
        RECT 97.585 142.415 98.540 142.635 ;
        RECT 97.815 141.785 98.085 142.245 ;
        RECT 98.255 141.955 98.540 142.415 ;
        RECT 98.825 141.785 100.035 142.875 ;
        RECT 100.205 142.805 100.895 143.365 ;
        RECT 101.065 142.635 101.275 143.535 ;
        RECT 100.320 142.415 101.275 142.635 ;
        RECT 101.445 143.365 101.845 144.165 ;
        RECT 102.035 143.705 102.315 144.165 ;
        RECT 102.835 143.875 103.160 144.335 ;
        RECT 102.035 143.535 103.160 143.705 ;
        RECT 103.330 143.595 103.715 144.165 ;
        RECT 102.710 143.425 103.160 143.535 ;
        RECT 101.445 142.805 102.540 143.365 ;
        RECT 102.710 143.095 103.265 143.425 ;
        RECT 100.320 141.955 100.605 142.415 ;
        RECT 100.775 141.785 101.045 142.245 ;
        RECT 101.445 141.955 101.845 142.805 ;
        RECT 102.710 142.635 103.160 143.095 ;
        RECT 103.435 142.925 103.715 143.595 ;
        RECT 102.035 142.415 103.160 142.635 ;
        RECT 102.035 141.955 102.315 142.415 ;
        RECT 102.835 141.785 103.160 142.245 ;
        RECT 103.330 141.955 103.715 142.925 ;
        RECT 103.885 143.390 104.225 144.165 ;
        RECT 104.395 143.875 104.565 144.335 ;
        RECT 104.805 143.900 105.165 144.165 ;
        RECT 104.805 143.895 105.160 143.900 ;
        RECT 104.805 143.885 105.155 143.895 ;
        RECT 104.805 143.880 105.150 143.885 ;
        RECT 104.805 143.870 105.145 143.880 ;
        RECT 105.795 143.875 105.965 144.335 ;
        RECT 104.805 143.865 105.140 143.870 ;
        RECT 104.805 143.855 105.130 143.865 ;
        RECT 104.805 143.845 105.120 143.855 ;
        RECT 104.805 143.705 105.105 143.845 ;
        RECT 104.395 143.515 105.105 143.705 ;
        RECT 105.295 143.705 105.625 143.785 ;
        RECT 106.135 143.705 106.475 144.165 ;
        RECT 106.645 143.790 111.990 144.335 ;
        RECT 105.295 143.515 106.475 143.705 ;
        RECT 103.885 141.955 104.165 143.390 ;
        RECT 104.395 142.945 104.680 143.515 ;
        RECT 104.865 143.115 105.335 143.345 ;
        RECT 105.505 143.325 105.835 143.345 ;
        RECT 105.505 143.145 105.955 143.325 ;
        RECT 106.145 143.145 106.475 143.345 ;
        RECT 104.395 142.730 105.545 142.945 ;
        RECT 104.335 141.785 105.045 142.560 ;
        RECT 105.215 141.955 105.545 142.730 ;
        RECT 105.740 142.030 105.955 143.145 ;
        RECT 106.245 142.805 106.475 143.145 ;
        RECT 108.230 142.960 108.570 143.790 ;
        RECT 112.255 143.785 112.425 144.075 ;
        RECT 112.595 143.955 112.925 144.335 ;
        RECT 112.255 143.615 112.920 143.785 ;
        RECT 106.135 141.785 106.465 142.505 ;
        RECT 110.050 142.220 110.400 143.470 ;
        RECT 112.170 142.795 112.520 143.445 ;
        RECT 112.690 142.625 112.920 143.615 ;
        RECT 112.255 142.455 112.920 142.625 ;
        RECT 106.645 141.785 111.990 142.220 ;
        RECT 112.255 141.955 112.425 142.455 ;
        RECT 112.595 141.785 112.925 142.285 ;
        RECT 113.095 141.955 113.280 144.075 ;
        RECT 113.535 143.875 113.785 144.335 ;
        RECT 113.955 143.885 114.290 144.055 ;
        RECT 114.485 143.885 115.160 144.055 ;
        RECT 113.955 143.745 114.125 143.885 ;
        RECT 113.450 142.755 113.730 143.705 ;
        RECT 113.900 143.615 114.125 143.745 ;
        RECT 113.900 142.510 114.070 143.615 ;
        RECT 114.295 143.465 114.820 143.685 ;
        RECT 114.240 142.700 114.480 143.295 ;
        RECT 114.650 142.765 114.820 143.465 ;
        RECT 114.990 143.105 115.160 143.885 ;
        RECT 115.480 143.835 115.850 144.335 ;
        RECT 116.030 143.885 116.435 144.055 ;
        RECT 116.605 143.885 117.390 144.055 ;
        RECT 116.030 143.655 116.200 143.885 ;
        RECT 115.370 143.355 116.200 143.655 ;
        RECT 116.585 143.385 117.050 143.715 ;
        RECT 115.370 143.325 115.570 143.355 ;
        RECT 115.690 143.105 115.860 143.175 ;
        RECT 114.990 142.935 115.860 143.105 ;
        RECT 115.350 142.845 115.860 142.935 ;
        RECT 113.900 142.380 114.205 142.510 ;
        RECT 114.650 142.400 115.180 142.765 ;
        RECT 113.520 141.785 113.785 142.245 ;
        RECT 113.955 141.955 114.205 142.380 ;
        RECT 115.350 142.230 115.520 142.845 ;
        RECT 114.415 142.060 115.520 142.230 ;
        RECT 115.690 141.785 115.860 142.585 ;
        RECT 116.030 142.285 116.200 143.355 ;
        RECT 116.370 142.455 116.560 143.175 ;
        RECT 116.730 142.425 117.050 143.385 ;
        RECT 117.220 143.425 117.390 143.885 ;
        RECT 117.665 143.805 117.875 144.335 ;
        RECT 118.135 143.595 118.465 144.120 ;
        RECT 118.635 143.725 118.805 144.335 ;
        RECT 118.975 143.680 119.305 144.115 ;
        RECT 118.975 143.595 119.355 143.680 ;
        RECT 120.445 143.610 120.735 144.335 ;
        RECT 118.265 143.425 118.465 143.595 ;
        RECT 119.130 143.555 119.355 143.595 ;
        RECT 120.910 143.570 121.365 144.335 ;
        RECT 121.640 143.955 122.940 144.165 ;
        RECT 123.195 143.975 123.525 144.335 ;
        RECT 122.770 143.805 122.940 143.955 ;
        RECT 123.695 143.835 123.955 144.165 ;
        RECT 123.725 143.825 123.955 143.835 ;
        RECT 117.220 143.095 118.095 143.425 ;
        RECT 118.265 143.095 119.015 143.425 ;
        RECT 116.030 141.955 116.280 142.285 ;
        RECT 117.220 142.255 117.390 143.095 ;
        RECT 118.265 142.890 118.455 143.095 ;
        RECT 119.185 142.975 119.355 143.555 ;
        RECT 121.840 143.345 122.060 143.745 ;
        RECT 120.905 143.145 121.395 143.345 ;
        RECT 121.585 143.135 122.060 143.345 ;
        RECT 122.305 143.345 122.515 143.745 ;
        RECT 122.770 143.680 123.525 143.805 ;
        RECT 122.770 143.635 123.615 143.680 ;
        RECT 123.345 143.515 123.615 143.635 ;
        RECT 122.305 143.135 122.635 143.345 ;
        RECT 122.805 143.075 123.215 143.380 ;
        RECT 119.140 142.925 119.355 142.975 ;
        RECT 117.560 142.515 118.455 142.890 ;
        RECT 118.965 142.845 119.355 142.925 ;
        RECT 116.505 142.085 117.390 142.255 ;
        RECT 117.570 141.785 117.885 142.285 ;
        RECT 118.115 141.955 118.455 142.515 ;
        RECT 118.625 141.785 118.795 142.795 ;
        RECT 118.965 142.000 119.295 142.845 ;
        RECT 120.445 141.785 120.735 142.950 ;
        RECT 120.910 142.905 122.085 142.965 ;
        RECT 123.445 142.940 123.615 143.515 ;
        RECT 123.415 142.905 123.615 142.940 ;
        RECT 120.910 142.795 123.615 142.905 ;
        RECT 120.910 142.175 121.165 142.795 ;
        RECT 121.755 142.735 123.555 142.795 ;
        RECT 121.755 142.705 122.085 142.735 ;
        RECT 123.785 142.635 123.955 143.825 ;
        RECT 124.215 143.785 124.385 144.075 ;
        RECT 124.555 143.955 124.885 144.335 ;
        RECT 124.215 143.615 124.880 143.785 ;
        RECT 124.130 142.795 124.480 143.445 ;
        RECT 121.415 142.535 121.600 142.625 ;
        RECT 122.190 142.535 123.025 142.545 ;
        RECT 121.415 142.335 123.025 142.535 ;
        RECT 121.415 142.295 121.645 142.335 ;
        RECT 120.910 141.955 121.245 142.175 ;
        RECT 122.250 141.785 122.605 142.165 ;
        RECT 122.775 141.955 123.025 142.335 ;
        RECT 123.275 141.785 123.525 142.565 ;
        RECT 123.695 141.955 123.955 142.635 ;
        RECT 124.650 142.625 124.880 143.615 ;
        RECT 124.215 142.455 124.880 142.625 ;
        RECT 124.215 141.955 124.385 142.455 ;
        RECT 124.555 141.785 124.885 142.285 ;
        RECT 125.055 141.955 125.240 144.075 ;
        RECT 125.495 143.875 125.745 144.335 ;
        RECT 125.915 143.885 126.250 144.055 ;
        RECT 126.445 143.885 127.120 144.055 ;
        RECT 125.915 143.745 126.085 143.885 ;
        RECT 125.410 142.755 125.690 143.705 ;
        RECT 125.860 143.615 126.085 143.745 ;
        RECT 125.860 142.510 126.030 143.615 ;
        RECT 126.255 143.465 126.780 143.685 ;
        RECT 126.200 142.700 126.440 143.295 ;
        RECT 126.610 142.765 126.780 143.465 ;
        RECT 126.950 143.105 127.120 143.885 ;
        RECT 127.440 143.835 127.810 144.335 ;
        RECT 127.990 143.885 128.395 144.055 ;
        RECT 128.565 143.885 129.350 144.055 ;
        RECT 127.990 143.655 128.160 143.885 ;
        RECT 127.330 143.355 128.160 143.655 ;
        RECT 128.545 143.385 129.010 143.715 ;
        RECT 127.330 143.325 127.530 143.355 ;
        RECT 127.650 143.105 127.820 143.175 ;
        RECT 126.950 142.935 127.820 143.105 ;
        RECT 127.310 142.845 127.820 142.935 ;
        RECT 125.860 142.380 126.165 142.510 ;
        RECT 126.610 142.400 127.140 142.765 ;
        RECT 125.480 141.785 125.745 142.245 ;
        RECT 125.915 141.955 126.165 142.380 ;
        RECT 127.310 142.230 127.480 142.845 ;
        RECT 126.375 142.060 127.480 142.230 ;
        RECT 127.650 141.785 127.820 142.585 ;
        RECT 127.990 142.285 128.160 143.355 ;
        RECT 128.330 142.455 128.520 143.175 ;
        RECT 128.690 142.425 129.010 143.385 ;
        RECT 129.180 143.425 129.350 143.885 ;
        RECT 129.625 143.805 129.835 144.335 ;
        RECT 130.095 143.595 130.425 144.120 ;
        RECT 130.595 143.725 130.765 144.335 ;
        RECT 130.935 143.680 131.265 144.115 ;
        RECT 131.485 143.790 136.830 144.335 ;
        RECT 130.935 143.595 131.315 143.680 ;
        RECT 130.225 143.425 130.425 143.595 ;
        RECT 131.090 143.555 131.315 143.595 ;
        RECT 129.180 143.095 130.055 143.425 ;
        RECT 130.225 143.095 130.975 143.425 ;
        RECT 127.990 141.955 128.240 142.285 ;
        RECT 129.180 142.255 129.350 143.095 ;
        RECT 130.225 142.890 130.415 143.095 ;
        RECT 131.145 142.975 131.315 143.555 ;
        RECT 131.100 142.925 131.315 142.975 ;
        RECT 133.070 142.960 133.410 143.790 ;
        RECT 137.555 143.785 137.725 144.165 ;
        RECT 137.905 143.955 138.235 144.335 ;
        RECT 137.555 143.615 138.220 143.785 ;
        RECT 138.415 143.660 138.675 144.165 ;
        RECT 129.520 142.515 130.415 142.890 ;
        RECT 130.925 142.845 131.315 142.925 ;
        RECT 128.465 142.085 129.350 142.255 ;
        RECT 129.530 141.785 129.845 142.285 ;
        RECT 130.075 141.955 130.415 142.515 ;
        RECT 130.585 141.785 130.755 142.795 ;
        RECT 130.925 142.000 131.255 142.845 ;
        RECT 134.890 142.220 135.240 143.470 ;
        RECT 137.485 143.065 137.815 143.435 ;
        RECT 138.050 143.360 138.220 143.615 ;
        RECT 138.050 143.030 138.335 143.360 ;
        RECT 138.050 142.885 138.220 143.030 ;
        RECT 137.555 142.715 138.220 142.885 ;
        RECT 138.505 142.860 138.675 143.660 ;
        RECT 131.485 141.785 136.830 142.220 ;
        RECT 137.555 141.955 137.725 142.715 ;
        RECT 137.905 141.785 138.235 142.545 ;
        RECT 138.405 141.955 138.675 142.860 ;
        RECT 138.845 143.660 139.105 144.165 ;
        RECT 139.285 143.955 139.615 144.335 ;
        RECT 139.795 143.785 139.965 144.165 ;
        RECT 138.845 142.860 139.015 143.660 ;
        RECT 139.300 143.615 139.965 143.785 ;
        RECT 140.315 143.785 140.485 144.165 ;
        RECT 140.700 143.955 141.030 144.335 ;
        RECT 140.315 143.615 141.030 143.785 ;
        RECT 139.300 143.360 139.470 143.615 ;
        RECT 139.185 143.030 139.470 143.360 ;
        RECT 139.705 143.065 140.035 143.435 ;
        RECT 140.225 143.065 140.580 143.435 ;
        RECT 140.860 143.425 141.030 143.615 ;
        RECT 141.200 143.590 141.455 144.165 ;
        RECT 140.860 143.095 141.115 143.425 ;
        RECT 139.300 142.885 139.470 143.030 ;
        RECT 140.860 142.885 141.030 143.095 ;
        RECT 138.845 141.955 139.115 142.860 ;
        RECT 139.300 142.715 139.965 142.885 ;
        RECT 139.285 141.785 139.615 142.545 ;
        RECT 139.795 141.955 139.965 142.715 ;
        RECT 140.315 142.715 141.030 142.885 ;
        RECT 141.285 142.860 141.455 143.590 ;
        RECT 141.630 143.495 141.890 144.335 ;
        RECT 142.180 143.705 142.465 144.165 ;
        RECT 142.635 143.875 142.905 144.335 ;
        RECT 142.180 143.535 143.135 143.705 ;
        RECT 140.315 141.955 140.485 142.715 ;
        RECT 140.700 141.785 141.030 142.545 ;
        RECT 141.200 141.955 141.455 142.860 ;
        RECT 141.630 141.785 141.890 142.935 ;
        RECT 142.065 142.805 142.755 143.365 ;
        RECT 142.925 142.635 143.135 143.535 ;
        RECT 142.180 142.415 143.135 142.635 ;
        RECT 143.305 143.365 143.705 144.165 ;
        RECT 143.895 143.705 144.175 144.165 ;
        RECT 144.695 143.875 145.020 144.335 ;
        RECT 143.895 143.535 145.020 143.705 ;
        RECT 145.190 143.595 145.575 144.165 ;
        RECT 144.570 143.425 145.020 143.535 ;
        RECT 143.305 142.805 144.400 143.365 ;
        RECT 144.570 143.095 145.125 143.425 ;
        RECT 142.180 141.955 142.465 142.415 ;
        RECT 142.635 141.785 142.905 142.245 ;
        RECT 143.305 141.955 143.705 142.805 ;
        RECT 144.570 142.635 145.020 143.095 ;
        RECT 145.295 142.925 145.575 143.595 ;
        RECT 145.745 143.585 146.955 144.335 ;
        RECT 143.895 142.415 145.020 142.635 ;
        RECT 143.895 141.955 144.175 142.415 ;
        RECT 144.695 141.785 145.020 142.245 ;
        RECT 145.190 141.955 145.575 142.925 ;
        RECT 145.745 142.875 146.265 143.415 ;
        RECT 146.435 143.045 146.955 143.585 ;
        RECT 145.745 141.785 146.955 142.875 ;
        RECT 17.320 141.615 147.040 141.785 ;
        RECT 17.405 140.525 18.615 141.615 ;
        RECT 18.785 141.180 24.130 141.615 ;
        RECT 24.305 141.180 29.650 141.615 ;
        RECT 17.405 139.815 17.925 140.355 ;
        RECT 18.095 139.985 18.615 140.525 ;
        RECT 17.405 139.065 18.615 139.815 ;
        RECT 20.370 139.610 20.710 140.440 ;
        RECT 22.190 139.930 22.540 141.180 ;
        RECT 25.890 139.610 26.230 140.440 ;
        RECT 27.710 139.930 28.060 141.180 ;
        RECT 30.285 140.450 30.575 141.615 ;
        RECT 30.745 140.525 32.415 141.615 ;
        RECT 32.585 141.105 32.845 141.615 ;
        RECT 30.745 139.835 31.495 140.355 ;
        RECT 31.665 140.005 32.415 140.525 ;
        RECT 32.585 140.055 32.925 140.935 ;
        RECT 33.095 140.225 33.265 141.445 ;
        RECT 33.505 141.110 34.120 141.615 ;
        RECT 33.505 140.575 33.755 140.940 ;
        RECT 33.925 140.935 34.120 141.110 ;
        RECT 34.290 141.105 34.765 141.445 ;
        RECT 34.935 141.070 35.150 141.615 ;
        RECT 33.925 140.745 34.255 140.935 ;
        RECT 34.475 140.575 35.190 140.870 ;
        RECT 35.360 140.745 35.635 141.445 ;
        RECT 35.895 140.945 36.065 141.445 ;
        RECT 36.235 141.115 36.565 141.615 ;
        RECT 35.895 140.775 36.560 140.945 ;
        RECT 33.505 140.405 35.295 140.575 ;
        RECT 33.095 139.975 33.890 140.225 ;
        RECT 33.095 139.885 33.345 139.975 ;
        RECT 18.785 139.065 24.130 139.610 ;
        RECT 24.305 139.065 29.650 139.610 ;
        RECT 30.285 139.065 30.575 139.790 ;
        RECT 30.745 139.065 32.415 139.835 ;
        RECT 32.585 139.065 32.845 139.885 ;
        RECT 33.015 139.465 33.345 139.885 ;
        RECT 34.060 139.550 34.315 140.405 ;
        RECT 33.525 139.285 34.315 139.550 ;
        RECT 34.485 139.705 34.895 140.225 ;
        RECT 35.065 139.975 35.295 140.405 ;
        RECT 35.465 139.715 35.635 140.745 ;
        RECT 35.810 139.955 36.160 140.605 ;
        RECT 36.330 139.785 36.560 140.775 ;
        RECT 34.485 139.285 34.685 139.705 ;
        RECT 34.875 139.065 35.205 139.525 ;
        RECT 35.375 139.235 35.635 139.715 ;
        RECT 35.895 139.615 36.560 139.785 ;
        RECT 35.895 139.325 36.065 139.615 ;
        RECT 36.235 139.065 36.565 139.445 ;
        RECT 36.735 139.325 36.920 141.445 ;
        RECT 37.160 141.155 37.425 141.615 ;
        RECT 37.595 141.020 37.845 141.445 ;
        RECT 38.055 141.170 39.160 141.340 ;
        RECT 37.540 140.890 37.845 141.020 ;
        RECT 37.090 139.695 37.370 140.645 ;
        RECT 37.540 139.785 37.710 140.890 ;
        RECT 37.880 140.105 38.120 140.700 ;
        RECT 38.290 140.635 38.820 141.000 ;
        RECT 38.290 139.935 38.460 140.635 ;
        RECT 38.990 140.555 39.160 141.170 ;
        RECT 39.330 140.815 39.500 141.615 ;
        RECT 39.670 141.115 39.920 141.445 ;
        RECT 40.145 141.145 41.030 141.315 ;
        RECT 38.990 140.465 39.500 140.555 ;
        RECT 37.540 139.655 37.765 139.785 ;
        RECT 37.935 139.715 38.460 139.935 ;
        RECT 38.630 140.295 39.500 140.465 ;
        RECT 37.175 139.065 37.425 139.525 ;
        RECT 37.595 139.515 37.765 139.655 ;
        RECT 38.630 139.515 38.800 140.295 ;
        RECT 39.330 140.225 39.500 140.295 ;
        RECT 39.010 140.045 39.210 140.075 ;
        RECT 39.670 140.045 39.840 141.115 ;
        RECT 40.010 140.225 40.200 140.945 ;
        RECT 39.010 139.745 39.840 140.045 ;
        RECT 40.370 140.015 40.690 140.975 ;
        RECT 37.595 139.345 37.930 139.515 ;
        RECT 38.125 139.345 38.800 139.515 ;
        RECT 39.120 139.065 39.490 139.565 ;
        RECT 39.670 139.515 39.840 139.745 ;
        RECT 40.225 139.685 40.690 140.015 ;
        RECT 40.860 140.305 41.030 141.145 ;
        RECT 41.210 141.115 41.525 141.615 ;
        RECT 41.755 140.885 42.095 141.445 ;
        RECT 41.200 140.510 42.095 140.885 ;
        RECT 42.265 140.605 42.435 141.615 ;
        RECT 41.905 140.305 42.095 140.510 ;
        RECT 42.605 140.555 42.935 141.400 ;
        RECT 42.605 140.475 42.995 140.555 ;
        RECT 43.165 140.525 44.375 141.615 ;
        RECT 44.795 140.885 45.090 141.615 ;
        RECT 45.260 140.715 45.520 141.440 ;
        RECT 45.690 140.885 45.950 141.615 ;
        RECT 46.120 140.715 46.380 141.440 ;
        RECT 46.550 140.885 46.810 141.615 ;
        RECT 46.980 140.715 47.240 141.440 ;
        RECT 47.410 140.885 47.670 141.615 ;
        RECT 47.840 140.715 48.100 141.440 ;
        RECT 42.780 140.425 42.995 140.475 ;
        RECT 40.860 139.975 41.735 140.305 ;
        RECT 41.905 139.975 42.655 140.305 ;
        RECT 40.860 139.515 41.030 139.975 ;
        RECT 41.905 139.805 42.105 139.975 ;
        RECT 42.825 139.845 42.995 140.425 ;
        RECT 42.770 139.805 42.995 139.845 ;
        RECT 39.670 139.345 40.075 139.515 ;
        RECT 40.245 139.345 41.030 139.515 ;
        RECT 41.305 139.065 41.515 139.595 ;
        RECT 41.775 139.280 42.105 139.805 ;
        RECT 42.615 139.720 42.995 139.805 ;
        RECT 43.165 139.815 43.685 140.355 ;
        RECT 43.855 139.985 44.375 140.525 ;
        RECT 44.790 140.475 48.100 140.715 ;
        RECT 48.270 140.505 48.530 141.615 ;
        RECT 44.790 139.885 45.760 140.475 ;
        RECT 48.700 140.305 48.950 141.440 ;
        RECT 49.130 140.505 49.425 141.615 ;
        RECT 49.605 140.525 52.195 141.615 ;
        RECT 45.930 140.055 48.950 140.305 ;
        RECT 42.275 139.065 42.445 139.675 ;
        RECT 42.615 139.285 42.945 139.720 ;
        RECT 43.165 139.065 44.375 139.815 ;
        RECT 44.790 139.715 48.100 139.885 ;
        RECT 44.790 139.065 45.090 139.545 ;
        RECT 45.260 139.260 45.520 139.715 ;
        RECT 45.690 139.065 45.950 139.545 ;
        RECT 46.120 139.260 46.380 139.715 ;
        RECT 46.550 139.065 46.810 139.545 ;
        RECT 46.980 139.260 47.240 139.715 ;
        RECT 47.410 139.065 47.670 139.545 ;
        RECT 47.840 139.260 48.100 139.715 ;
        RECT 48.270 139.065 48.530 139.590 ;
        RECT 48.700 139.245 48.950 140.055 ;
        RECT 49.120 139.695 49.435 140.305 ;
        RECT 49.605 139.835 50.815 140.355 ;
        RECT 50.985 140.005 52.195 140.525 ;
        RECT 52.835 140.555 53.165 141.405 ;
        RECT 49.130 139.065 49.375 139.525 ;
        RECT 49.605 139.065 52.195 139.835 ;
        RECT 52.835 139.790 53.025 140.555 ;
        RECT 53.335 140.475 53.585 141.615 ;
        RECT 53.775 140.975 54.025 141.395 ;
        RECT 54.255 141.145 54.585 141.615 ;
        RECT 54.815 140.975 55.065 141.395 ;
        RECT 53.775 140.805 55.065 140.975 ;
        RECT 55.245 140.975 55.575 141.405 ;
        RECT 55.245 140.805 55.700 140.975 ;
        RECT 53.765 140.305 53.980 140.635 ;
        RECT 53.195 139.975 53.505 140.305 ;
        RECT 53.675 139.975 53.980 140.305 ;
        RECT 54.155 139.975 54.440 140.635 ;
        RECT 54.635 139.975 54.900 140.635 ;
        RECT 55.115 139.975 55.360 140.635 ;
        RECT 53.335 139.805 53.505 139.975 ;
        RECT 55.530 139.805 55.700 140.805 ;
        RECT 56.045 140.450 56.335 141.615 ;
        RECT 56.505 140.525 57.715 141.615 ;
        RECT 52.835 139.280 53.165 139.790 ;
        RECT 53.335 139.635 55.700 139.805 ;
        RECT 56.505 139.815 57.025 140.355 ;
        RECT 57.195 139.985 57.715 140.525 ;
        RECT 57.895 140.505 58.190 141.615 ;
        RECT 58.370 140.305 58.620 141.440 ;
        RECT 58.790 140.505 59.050 141.615 ;
        RECT 59.220 140.715 59.480 141.440 ;
        RECT 59.650 140.885 59.910 141.615 ;
        RECT 60.080 140.715 60.340 141.440 ;
        RECT 60.510 140.885 60.770 141.615 ;
        RECT 60.940 140.715 61.200 141.440 ;
        RECT 61.370 140.885 61.630 141.615 ;
        RECT 61.800 140.715 62.060 141.440 ;
        RECT 62.230 140.885 62.525 141.615 ;
        RECT 63.000 140.815 63.300 141.615 ;
        RECT 59.220 140.475 62.530 140.715 ;
        RECT 63.470 140.645 63.800 141.445 ;
        RECT 63.970 140.815 64.140 141.615 ;
        RECT 64.310 140.645 64.640 141.445 ;
        RECT 64.810 140.815 64.980 141.615 ;
        RECT 65.150 140.645 65.480 141.445 ;
        RECT 65.650 140.815 65.820 141.615 ;
        RECT 65.990 140.645 66.320 141.445 ;
        RECT 66.490 140.815 66.745 141.615 ;
        RECT 67.085 140.745 67.360 141.445 ;
        RECT 67.530 141.070 67.785 141.615 ;
        RECT 67.955 141.105 68.435 141.445 ;
        RECT 68.610 141.060 69.215 141.615 ;
        RECT 68.600 140.960 69.215 141.060 ;
        RECT 68.600 140.935 68.785 140.960 ;
        RECT 53.335 139.065 53.665 139.465 ;
        RECT 54.715 139.295 55.045 139.635 ;
        RECT 55.215 139.065 55.545 139.465 ;
        RECT 56.045 139.065 56.335 139.790 ;
        RECT 56.505 139.065 57.715 139.815 ;
        RECT 57.885 139.695 58.200 140.305 ;
        RECT 58.370 140.055 61.390 140.305 ;
        RECT 57.945 139.065 58.190 139.525 ;
        RECT 58.370 139.245 58.620 140.055 ;
        RECT 61.560 139.885 62.530 140.475 ;
        RECT 59.220 139.715 62.530 139.885 ;
        RECT 62.945 140.475 66.915 140.645 ;
        RECT 62.945 139.885 63.265 140.475 ;
        RECT 63.465 140.055 66.320 140.305 ;
        RECT 66.570 139.885 66.915 140.475 ;
        RECT 58.790 139.065 59.050 139.590 ;
        RECT 59.220 139.260 59.480 139.715 ;
        RECT 59.650 139.065 59.910 139.545 ;
        RECT 60.080 139.260 60.340 139.715 ;
        RECT 60.510 139.065 60.770 139.545 ;
        RECT 60.940 139.260 61.200 139.715 ;
        RECT 61.370 139.065 61.630 139.545 ;
        RECT 61.800 139.260 62.060 139.715 ;
        RECT 62.945 139.695 66.915 139.885 ;
        RECT 67.085 139.715 67.255 140.745 ;
        RECT 67.530 140.615 68.285 140.865 ;
        RECT 68.455 140.690 68.785 140.935 ;
        RECT 67.530 140.580 68.300 140.615 ;
        RECT 67.530 140.570 68.315 140.580 ;
        RECT 67.425 140.555 68.320 140.570 ;
        RECT 67.425 140.540 68.340 140.555 ;
        RECT 67.425 140.530 68.360 140.540 ;
        RECT 67.425 140.520 68.385 140.530 ;
        RECT 67.425 140.490 68.455 140.520 ;
        RECT 67.425 140.460 68.475 140.490 ;
        RECT 67.425 140.430 68.495 140.460 ;
        RECT 67.425 140.405 68.525 140.430 ;
        RECT 67.425 140.370 68.560 140.405 ;
        RECT 67.425 140.365 68.590 140.370 ;
        RECT 67.425 139.970 67.655 140.365 ;
        RECT 68.200 140.360 68.590 140.365 ;
        RECT 68.225 140.350 68.590 140.360 ;
        RECT 68.240 140.345 68.590 140.350 ;
        RECT 68.255 140.340 68.590 140.345 ;
        RECT 68.955 140.340 69.215 140.790 ;
        RECT 69.390 140.475 69.710 141.615 ;
        RECT 68.255 140.335 69.215 140.340 ;
        RECT 68.265 140.325 69.215 140.335 ;
        RECT 68.275 140.320 69.215 140.325 ;
        RECT 68.285 140.310 69.215 140.320 ;
        RECT 68.290 140.300 69.215 140.310 ;
        RECT 69.890 140.305 70.085 141.355 ;
        RECT 70.265 140.765 70.595 141.445 ;
        RECT 70.795 140.815 71.050 141.615 ;
        RECT 71.315 140.945 71.485 141.445 ;
        RECT 71.655 141.115 71.985 141.615 ;
        RECT 71.315 140.775 71.980 140.945 ;
        RECT 70.265 140.485 70.615 140.765 ;
        RECT 68.295 140.295 69.215 140.300 ;
        RECT 68.305 140.280 69.215 140.295 ;
        RECT 68.310 140.265 69.215 140.280 ;
        RECT 68.320 140.240 69.215 140.265 ;
        RECT 69.450 140.255 69.710 140.305 ;
        RECT 67.825 139.770 68.155 140.195 ;
        RECT 62.230 139.065 62.530 139.545 ;
        RECT 62.995 139.065 63.300 139.525 ;
        RECT 63.470 139.235 63.800 139.695 ;
        RECT 63.970 139.065 64.140 139.525 ;
        RECT 64.310 139.235 64.640 139.695 ;
        RECT 64.810 139.065 64.980 139.525 ;
        RECT 65.150 139.235 65.480 139.695 ;
        RECT 65.650 139.065 65.820 139.525 ;
        RECT 65.990 139.235 66.320 139.695 ;
        RECT 66.490 139.065 66.745 139.525 ;
        RECT 67.085 139.235 67.345 139.715 ;
        RECT 67.515 139.065 67.765 139.605 ;
        RECT 67.935 139.285 68.155 139.770 ;
        RECT 68.325 140.170 69.215 140.240 ;
        RECT 68.325 139.445 68.495 140.170 ;
        RECT 69.445 140.085 69.710 140.255 ;
        RECT 68.665 139.615 69.215 140.000 ;
        RECT 69.450 139.975 69.710 140.085 ;
        RECT 69.890 139.975 70.275 140.305 ;
        RECT 70.445 140.105 70.615 140.485 ;
        RECT 70.805 140.275 71.050 140.635 ;
        RECT 70.445 139.935 70.965 140.105 ;
        RECT 71.230 139.955 71.580 140.605 ;
        RECT 70.795 139.915 70.965 139.935 ;
        RECT 69.390 139.595 70.605 139.765 ;
        RECT 68.325 139.275 69.215 139.445 ;
        RECT 69.390 139.245 69.680 139.595 ;
        RECT 69.875 139.065 70.205 139.425 ;
        RECT 70.375 139.290 70.605 139.595 ;
        RECT 70.795 139.745 70.995 139.915 ;
        RECT 71.750 139.785 71.980 140.775 ;
        RECT 70.795 139.370 70.965 139.745 ;
        RECT 71.315 139.615 71.980 139.785 ;
        RECT 71.315 139.325 71.485 139.615 ;
        RECT 71.655 139.065 71.985 139.445 ;
        RECT 72.155 139.325 72.340 141.445 ;
        RECT 72.580 141.155 72.845 141.615 ;
        RECT 73.015 141.020 73.265 141.445 ;
        RECT 73.475 141.170 74.580 141.340 ;
        RECT 72.960 140.890 73.265 141.020 ;
        RECT 72.510 139.695 72.790 140.645 ;
        RECT 72.960 139.785 73.130 140.890 ;
        RECT 73.300 140.105 73.540 140.700 ;
        RECT 73.710 140.635 74.240 141.000 ;
        RECT 73.710 139.935 73.880 140.635 ;
        RECT 74.410 140.555 74.580 141.170 ;
        RECT 74.750 140.815 74.920 141.615 ;
        RECT 75.090 141.115 75.340 141.445 ;
        RECT 75.565 141.145 76.450 141.315 ;
        RECT 74.410 140.465 74.920 140.555 ;
        RECT 72.960 139.655 73.185 139.785 ;
        RECT 73.355 139.715 73.880 139.935 ;
        RECT 74.050 140.295 74.920 140.465 ;
        RECT 72.595 139.065 72.845 139.525 ;
        RECT 73.015 139.515 73.185 139.655 ;
        RECT 74.050 139.515 74.220 140.295 ;
        RECT 74.750 140.225 74.920 140.295 ;
        RECT 74.430 140.045 74.630 140.075 ;
        RECT 75.090 140.045 75.260 141.115 ;
        RECT 75.430 140.225 75.620 140.945 ;
        RECT 74.430 139.745 75.260 140.045 ;
        RECT 75.790 140.015 76.110 140.975 ;
        RECT 73.015 139.345 73.350 139.515 ;
        RECT 73.545 139.345 74.220 139.515 ;
        RECT 74.540 139.065 74.910 139.565 ;
        RECT 75.090 139.515 75.260 139.745 ;
        RECT 75.645 139.685 76.110 140.015 ;
        RECT 76.280 140.305 76.450 141.145 ;
        RECT 76.630 141.115 76.945 141.615 ;
        RECT 77.175 140.885 77.515 141.445 ;
        RECT 76.620 140.510 77.515 140.885 ;
        RECT 77.685 140.605 77.855 141.615 ;
        RECT 77.325 140.305 77.515 140.510 ;
        RECT 78.025 140.555 78.355 141.400 ;
        RECT 78.590 141.235 78.925 141.615 ;
        RECT 78.025 140.475 78.415 140.555 ;
        RECT 78.200 140.425 78.415 140.475 ;
        RECT 76.280 139.975 77.155 140.305 ;
        RECT 77.325 139.975 78.075 140.305 ;
        RECT 76.280 139.515 76.450 139.975 ;
        RECT 77.325 139.805 77.525 139.975 ;
        RECT 78.245 139.845 78.415 140.425 ;
        RECT 78.190 139.805 78.415 139.845 ;
        RECT 75.090 139.345 75.495 139.515 ;
        RECT 75.665 139.345 76.450 139.515 ;
        RECT 76.725 139.065 76.935 139.595 ;
        RECT 77.195 139.280 77.525 139.805 ;
        RECT 78.035 139.720 78.415 139.805 ;
        RECT 78.585 139.745 78.825 141.055 ;
        RECT 79.095 140.645 79.345 141.445 ;
        RECT 79.565 140.895 79.895 141.615 ;
        RECT 80.080 140.645 80.330 141.445 ;
        RECT 80.795 140.815 81.125 141.615 ;
        RECT 81.295 141.185 81.635 141.445 ;
        RECT 78.995 140.475 81.185 140.645 ;
        RECT 77.695 139.065 77.865 139.675 ;
        RECT 78.035 139.285 78.365 139.720 ;
        RECT 78.995 139.565 79.165 140.475 ;
        RECT 80.870 140.305 81.185 140.475 ;
        RECT 78.670 139.235 79.165 139.565 ;
        RECT 79.385 139.340 79.735 140.305 ;
        RECT 79.915 139.335 80.215 140.305 ;
        RECT 80.395 139.335 80.675 140.305 ;
        RECT 80.870 140.055 81.200 140.305 ;
        RECT 80.855 139.065 81.125 139.865 ;
        RECT 81.375 139.785 81.635 141.185 ;
        RECT 81.805 140.450 82.095 141.615 ;
        RECT 82.265 140.855 82.780 141.265 ;
        RECT 83.015 140.855 83.185 141.615 ;
        RECT 83.355 141.275 85.385 141.445 ;
        RECT 82.265 140.045 82.605 140.855 ;
        RECT 83.355 140.610 83.525 141.275 ;
        RECT 83.920 140.935 85.045 141.105 ;
        RECT 82.775 140.420 83.525 140.610 ;
        RECT 83.695 140.595 84.705 140.765 ;
        RECT 82.265 139.875 83.495 140.045 ;
        RECT 81.295 139.275 81.635 139.785 ;
        RECT 81.805 139.065 82.095 139.790 ;
        RECT 82.540 139.270 82.785 139.875 ;
        RECT 83.005 139.065 83.515 139.600 ;
        RECT 83.695 139.235 83.885 140.595 ;
        RECT 84.055 139.915 84.330 140.395 ;
        RECT 84.055 139.745 84.335 139.915 ;
        RECT 84.535 139.795 84.705 140.595 ;
        RECT 84.875 139.805 85.045 140.935 ;
        RECT 85.215 140.305 85.385 141.275 ;
        RECT 85.555 140.475 85.725 141.615 ;
        RECT 85.895 140.475 86.230 141.445 ;
        RECT 86.425 140.725 86.685 141.435 ;
        RECT 86.855 140.905 87.185 141.615 ;
        RECT 87.355 140.725 87.585 141.435 ;
        RECT 86.425 140.485 87.585 140.725 ;
        RECT 87.765 140.705 88.035 141.435 ;
        RECT 88.215 140.885 88.555 141.615 ;
        RECT 87.765 140.485 88.535 140.705 ;
        RECT 85.215 139.975 85.410 140.305 ;
        RECT 85.635 139.975 85.890 140.305 ;
        RECT 85.635 139.805 85.805 139.975 ;
        RECT 86.060 139.805 86.230 140.475 ;
        RECT 86.415 139.975 86.715 140.305 ;
        RECT 86.895 139.995 87.420 140.305 ;
        RECT 87.600 139.995 88.065 140.305 ;
        RECT 84.055 139.235 84.330 139.745 ;
        RECT 84.875 139.635 85.805 139.805 ;
        RECT 84.875 139.600 85.050 139.635 ;
        RECT 84.520 139.235 85.050 139.600 ;
        RECT 85.475 139.065 85.805 139.465 ;
        RECT 85.975 139.235 86.230 139.805 ;
        RECT 86.425 139.065 86.715 139.795 ;
        RECT 86.895 139.355 87.125 139.995 ;
        RECT 88.245 139.815 88.535 140.485 ;
        RECT 87.305 139.615 88.535 139.815 ;
        RECT 87.305 139.245 87.615 139.615 ;
        RECT 87.795 139.065 88.465 139.435 ;
        RECT 88.725 139.245 88.985 141.435 ;
        RECT 89.165 140.525 90.375 141.615 ;
        RECT 90.635 140.945 90.805 141.445 ;
        RECT 90.975 141.115 91.305 141.615 ;
        RECT 90.635 140.775 91.300 140.945 ;
        RECT 89.165 139.815 89.685 140.355 ;
        RECT 89.855 139.985 90.375 140.525 ;
        RECT 90.550 139.955 90.900 140.605 ;
        RECT 89.165 139.065 90.375 139.815 ;
        RECT 91.070 139.785 91.300 140.775 ;
        RECT 90.635 139.615 91.300 139.785 ;
        RECT 90.635 139.325 90.805 139.615 ;
        RECT 90.975 139.065 91.305 139.445 ;
        RECT 91.475 139.325 91.660 141.445 ;
        RECT 91.900 141.155 92.165 141.615 ;
        RECT 92.335 141.020 92.585 141.445 ;
        RECT 92.795 141.170 93.900 141.340 ;
        RECT 92.280 140.890 92.585 141.020 ;
        RECT 91.830 139.695 92.110 140.645 ;
        RECT 92.280 139.785 92.450 140.890 ;
        RECT 92.620 140.105 92.860 140.700 ;
        RECT 93.030 140.635 93.560 141.000 ;
        RECT 93.030 139.935 93.200 140.635 ;
        RECT 93.730 140.555 93.900 141.170 ;
        RECT 94.070 140.815 94.240 141.615 ;
        RECT 94.410 141.115 94.660 141.445 ;
        RECT 94.885 141.145 95.770 141.315 ;
        RECT 93.730 140.465 94.240 140.555 ;
        RECT 92.280 139.655 92.505 139.785 ;
        RECT 92.675 139.715 93.200 139.935 ;
        RECT 93.370 140.295 94.240 140.465 ;
        RECT 91.915 139.065 92.165 139.525 ;
        RECT 92.335 139.515 92.505 139.655 ;
        RECT 93.370 139.515 93.540 140.295 ;
        RECT 94.070 140.225 94.240 140.295 ;
        RECT 93.750 140.045 93.950 140.075 ;
        RECT 94.410 140.045 94.580 141.115 ;
        RECT 94.750 140.225 94.940 140.945 ;
        RECT 93.750 139.745 94.580 140.045 ;
        RECT 95.110 140.015 95.430 140.975 ;
        RECT 92.335 139.345 92.670 139.515 ;
        RECT 92.865 139.345 93.540 139.515 ;
        RECT 93.860 139.065 94.230 139.565 ;
        RECT 94.410 139.515 94.580 139.745 ;
        RECT 94.965 139.685 95.430 140.015 ;
        RECT 95.600 140.305 95.770 141.145 ;
        RECT 95.950 141.115 96.265 141.615 ;
        RECT 96.495 140.885 96.835 141.445 ;
        RECT 95.940 140.510 96.835 140.885 ;
        RECT 97.005 140.605 97.175 141.615 ;
        RECT 96.645 140.305 96.835 140.510 ;
        RECT 97.345 140.555 97.675 141.400 ;
        RECT 97.905 140.645 98.215 141.445 ;
        RECT 98.385 140.815 98.695 141.615 ;
        RECT 98.865 140.985 99.125 141.445 ;
        RECT 99.295 141.155 99.550 141.615 ;
        RECT 99.725 140.985 99.985 141.445 ;
        RECT 98.865 140.815 99.985 140.985 ;
        RECT 97.345 140.475 97.735 140.555 ;
        RECT 97.520 140.425 97.735 140.475 ;
        RECT 95.600 139.975 96.475 140.305 ;
        RECT 96.645 139.975 97.395 140.305 ;
        RECT 95.600 139.515 95.770 139.975 ;
        RECT 96.645 139.805 96.845 139.975 ;
        RECT 97.565 139.845 97.735 140.425 ;
        RECT 97.510 139.805 97.735 139.845 ;
        RECT 94.410 139.345 94.815 139.515 ;
        RECT 94.985 139.345 95.770 139.515 ;
        RECT 96.045 139.065 96.255 139.595 ;
        RECT 96.515 139.280 96.845 139.805 ;
        RECT 97.355 139.720 97.735 139.805 ;
        RECT 97.905 140.475 98.935 140.645 ;
        RECT 97.015 139.065 97.185 139.675 ;
        RECT 97.355 139.285 97.685 139.720 ;
        RECT 97.905 139.565 98.075 140.475 ;
        RECT 98.245 139.735 98.595 140.305 ;
        RECT 98.765 140.225 98.935 140.475 ;
        RECT 99.725 140.565 99.985 140.815 ;
        RECT 100.155 140.745 100.440 141.615 ;
        RECT 99.725 140.395 100.480 140.565 ;
        RECT 98.765 140.055 99.905 140.225 ;
        RECT 100.075 139.885 100.480 140.395 ;
        RECT 98.830 139.715 100.480 139.885 ;
        RECT 101.605 140.560 101.910 141.345 ;
        RECT 102.090 141.145 102.775 141.615 ;
        RECT 102.085 140.625 102.780 140.935 ;
        RECT 101.605 139.755 101.780 140.560 ;
        RECT 102.955 140.455 103.240 141.400 ;
        RECT 103.415 141.165 103.745 141.615 ;
        RECT 103.915 140.995 104.085 141.425 ;
        RECT 102.380 140.305 103.240 140.455 ;
        RECT 101.955 140.285 103.240 140.305 ;
        RECT 103.410 140.765 104.085 140.995 ;
        RECT 104.435 140.995 104.605 141.425 ;
        RECT 104.775 141.165 105.105 141.615 ;
        RECT 104.435 140.765 105.110 140.995 ;
        RECT 101.955 139.925 102.940 140.285 ;
        RECT 103.410 140.115 103.645 140.765 ;
        RECT 97.905 139.235 98.205 139.565 ;
        RECT 98.375 139.065 98.650 139.545 ;
        RECT 98.830 139.325 99.125 139.715 ;
        RECT 99.295 139.065 99.550 139.545 ;
        RECT 99.725 139.325 99.985 139.715 ;
        RECT 100.155 139.065 100.435 139.545 ;
        RECT 101.605 139.235 101.845 139.755 ;
        RECT 102.770 139.590 102.940 139.925 ;
        RECT 103.110 139.785 103.645 140.115 ;
        RECT 103.425 139.635 103.645 139.785 ;
        RECT 103.815 139.745 104.115 140.595 ;
        RECT 104.405 139.745 104.705 140.595 ;
        RECT 104.875 140.115 105.110 140.765 ;
        RECT 105.280 140.455 105.565 141.400 ;
        RECT 105.745 141.145 106.430 141.615 ;
        RECT 105.740 140.625 106.435 140.935 ;
        RECT 106.610 140.560 106.915 141.345 ;
        RECT 105.280 140.305 106.140 140.455 ;
        RECT 105.280 140.285 106.565 140.305 ;
        RECT 104.875 139.785 105.410 140.115 ;
        RECT 105.580 139.925 106.565 140.285 ;
        RECT 104.875 139.635 105.095 139.785 ;
        RECT 102.015 139.065 102.410 139.560 ;
        RECT 102.770 139.395 103.145 139.590 ;
        RECT 102.975 139.250 103.145 139.395 ;
        RECT 103.425 139.260 103.665 139.635 ;
        RECT 103.835 139.065 104.170 139.570 ;
        RECT 104.350 139.065 104.685 139.570 ;
        RECT 104.855 139.260 105.095 139.635 ;
        RECT 105.580 139.590 105.750 139.925 ;
        RECT 106.740 139.755 106.915 140.560 ;
        RECT 107.565 140.450 107.855 141.615 ;
        RECT 108.025 141.180 113.370 141.615 ;
        RECT 113.545 141.180 118.890 141.615 ;
        RECT 105.375 139.395 105.750 139.590 ;
        RECT 105.375 139.250 105.545 139.395 ;
        RECT 106.110 139.065 106.505 139.560 ;
        RECT 106.675 139.235 106.915 139.755 ;
        RECT 107.565 139.065 107.855 139.790 ;
        RECT 109.610 139.610 109.950 140.440 ;
        RECT 111.430 139.930 111.780 141.180 ;
        RECT 115.130 139.610 115.470 140.440 ;
        RECT 116.950 139.930 117.300 141.180 ;
        RECT 119.065 140.525 120.275 141.615 ;
        RECT 119.065 139.815 119.585 140.355 ;
        RECT 119.755 139.985 120.275 140.525 ;
        RECT 120.450 141.225 120.785 141.445 ;
        RECT 121.790 141.235 122.145 141.615 ;
        RECT 120.450 140.605 120.705 141.225 ;
        RECT 120.955 141.065 121.185 141.105 ;
        RECT 122.315 141.065 122.565 141.445 ;
        RECT 120.955 140.865 122.565 141.065 ;
        RECT 120.955 140.775 121.140 140.865 ;
        RECT 121.730 140.855 122.565 140.865 ;
        RECT 122.815 140.835 123.065 141.615 ;
        RECT 123.235 140.765 123.495 141.445 ;
        RECT 121.295 140.665 121.625 140.695 ;
        RECT 121.295 140.605 123.095 140.665 ;
        RECT 120.450 140.495 123.155 140.605 ;
        RECT 120.450 140.435 121.625 140.495 ;
        RECT 122.955 140.460 123.155 140.495 ;
        RECT 120.445 140.055 120.935 140.255 ;
        RECT 121.125 140.055 121.600 140.265 ;
        RECT 108.025 139.065 113.370 139.610 ;
        RECT 113.545 139.065 118.890 139.610 ;
        RECT 119.065 139.065 120.275 139.815 ;
        RECT 120.450 139.065 120.905 139.830 ;
        RECT 121.380 139.655 121.600 140.055 ;
        RECT 121.845 140.055 122.175 140.265 ;
        RECT 121.845 139.655 122.055 140.055 ;
        RECT 122.345 140.020 122.755 140.325 ;
        RECT 122.985 139.885 123.155 140.460 ;
        RECT 122.885 139.765 123.155 139.885 ;
        RECT 122.310 139.720 123.155 139.765 ;
        RECT 122.310 139.595 123.065 139.720 ;
        RECT 122.310 139.445 122.480 139.595 ;
        RECT 123.325 139.565 123.495 140.765 ;
        RECT 123.665 140.475 123.945 141.615 ;
        RECT 124.115 140.465 124.445 141.445 ;
        RECT 124.615 140.475 124.875 141.615 ;
        RECT 125.045 140.525 128.555 141.615 ;
        RECT 128.725 140.525 129.935 141.615 ;
        RECT 123.675 140.035 124.010 140.305 ;
        RECT 124.180 139.865 124.350 140.465 ;
        RECT 124.520 140.055 124.855 140.305 ;
        RECT 121.180 139.235 122.480 139.445 ;
        RECT 122.735 139.065 123.065 139.425 ;
        RECT 123.235 139.235 123.495 139.565 ;
        RECT 123.665 139.065 123.975 139.865 ;
        RECT 124.180 139.235 124.875 139.865 ;
        RECT 125.045 139.835 126.695 140.355 ;
        RECT 126.865 140.005 128.555 140.525 ;
        RECT 125.045 139.065 128.555 139.835 ;
        RECT 128.725 139.815 129.245 140.355 ;
        RECT 129.415 139.985 129.935 140.525 ;
        RECT 130.110 141.225 130.445 141.445 ;
        RECT 131.450 141.235 131.805 141.615 ;
        RECT 130.110 140.605 130.365 141.225 ;
        RECT 130.615 141.065 130.845 141.105 ;
        RECT 131.975 141.065 132.225 141.445 ;
        RECT 130.615 140.865 132.225 141.065 ;
        RECT 130.615 140.775 130.800 140.865 ;
        RECT 131.390 140.855 132.225 140.865 ;
        RECT 132.475 140.835 132.725 141.615 ;
        RECT 132.895 140.765 133.155 141.445 ;
        RECT 130.955 140.665 131.285 140.695 ;
        RECT 130.955 140.605 132.755 140.665 ;
        RECT 130.110 140.495 132.815 140.605 ;
        RECT 130.110 140.435 131.285 140.495 ;
        RECT 132.615 140.460 132.815 140.495 ;
        RECT 130.105 140.055 130.595 140.255 ;
        RECT 130.785 140.055 131.260 140.265 ;
        RECT 128.725 139.065 129.935 139.815 ;
        RECT 130.110 139.065 130.565 139.830 ;
        RECT 131.040 139.655 131.260 140.055 ;
        RECT 131.505 140.055 131.835 140.265 ;
        RECT 131.505 139.655 131.715 140.055 ;
        RECT 132.005 140.020 132.415 140.325 ;
        RECT 132.645 139.885 132.815 140.460 ;
        RECT 132.545 139.765 132.815 139.885 ;
        RECT 131.970 139.720 132.815 139.765 ;
        RECT 131.970 139.595 132.725 139.720 ;
        RECT 131.970 139.445 132.140 139.595 ;
        RECT 132.985 139.575 133.155 140.765 ;
        RECT 133.325 140.450 133.615 141.615 ;
        RECT 134.710 140.475 135.045 141.445 ;
        RECT 135.215 140.475 135.385 141.615 ;
        RECT 135.555 141.275 137.585 141.445 ;
        RECT 134.710 139.805 134.880 140.475 ;
        RECT 135.555 140.305 135.725 141.275 ;
        RECT 135.050 139.975 135.305 140.305 ;
        RECT 135.530 139.975 135.725 140.305 ;
        RECT 135.895 140.935 137.020 141.105 ;
        RECT 135.135 139.805 135.305 139.975 ;
        RECT 135.895 139.805 136.065 140.935 ;
        RECT 132.925 139.565 133.155 139.575 ;
        RECT 130.840 139.235 132.140 139.445 ;
        RECT 132.395 139.065 132.725 139.425 ;
        RECT 132.895 139.235 133.155 139.565 ;
        RECT 133.325 139.065 133.615 139.790 ;
        RECT 134.710 139.235 134.965 139.805 ;
        RECT 135.135 139.635 136.065 139.805 ;
        RECT 136.235 140.595 137.245 140.765 ;
        RECT 136.235 139.795 136.405 140.595 ;
        RECT 136.610 139.915 136.885 140.395 ;
        RECT 136.605 139.745 136.885 139.915 ;
        RECT 135.890 139.600 136.065 139.635 ;
        RECT 135.135 139.065 135.465 139.465 ;
        RECT 135.890 139.235 136.420 139.600 ;
        RECT 136.610 139.235 136.885 139.745 ;
        RECT 137.055 139.235 137.245 140.595 ;
        RECT 137.415 140.610 137.585 141.275 ;
        RECT 137.755 140.855 137.925 141.615 ;
        RECT 138.160 140.855 138.675 141.265 ;
        RECT 137.415 140.420 138.165 140.610 ;
        RECT 138.335 140.045 138.675 140.855 ;
        RECT 137.445 139.875 138.675 140.045 ;
        RECT 138.845 140.475 139.230 141.445 ;
        RECT 139.400 141.155 139.725 141.615 ;
        RECT 140.245 140.985 140.525 141.445 ;
        RECT 139.400 140.765 140.525 140.985 ;
        RECT 137.425 139.065 137.935 139.600 ;
        RECT 138.155 139.270 138.400 139.875 ;
        RECT 138.845 139.805 139.125 140.475 ;
        RECT 139.400 140.305 139.850 140.765 ;
        RECT 140.715 140.595 141.115 141.445 ;
        RECT 141.515 141.155 141.785 141.615 ;
        RECT 141.955 140.985 142.240 141.445 ;
        RECT 139.295 139.975 139.850 140.305 ;
        RECT 140.020 140.035 141.115 140.595 ;
        RECT 139.400 139.865 139.850 139.975 ;
        RECT 138.845 139.235 139.230 139.805 ;
        RECT 139.400 139.695 140.525 139.865 ;
        RECT 139.400 139.065 139.725 139.525 ;
        RECT 140.245 139.235 140.525 139.695 ;
        RECT 140.715 139.235 141.115 140.035 ;
        RECT 141.285 140.765 142.240 140.985 ;
        RECT 141.285 139.865 141.495 140.765 ;
        RECT 141.665 140.035 142.355 140.595 ;
        RECT 142.525 140.540 142.795 141.445 ;
        RECT 142.965 140.855 143.295 141.615 ;
        RECT 143.475 140.685 143.645 141.445 ;
        RECT 141.285 139.695 142.240 139.865 ;
        RECT 141.515 139.065 141.785 139.525 ;
        RECT 141.955 139.235 142.240 139.695 ;
        RECT 142.525 139.740 142.695 140.540 ;
        RECT 142.980 140.515 143.645 140.685 ;
        RECT 143.995 140.685 144.165 141.445 ;
        RECT 144.380 140.855 144.710 141.615 ;
        RECT 143.995 140.515 144.710 140.685 ;
        RECT 144.880 140.540 145.135 141.445 ;
        RECT 142.980 140.370 143.150 140.515 ;
        RECT 142.865 140.040 143.150 140.370 ;
        RECT 142.980 139.785 143.150 140.040 ;
        RECT 143.385 139.965 143.715 140.335 ;
        RECT 143.905 139.965 144.260 140.335 ;
        RECT 144.540 140.305 144.710 140.515 ;
        RECT 144.540 139.975 144.795 140.305 ;
        RECT 144.540 139.785 144.710 139.975 ;
        RECT 144.965 139.810 145.135 140.540 ;
        RECT 145.310 140.465 145.570 141.615 ;
        RECT 145.745 140.525 146.955 141.615 ;
        RECT 145.745 139.985 146.265 140.525 ;
        RECT 142.525 139.235 142.785 139.740 ;
        RECT 142.980 139.615 143.645 139.785 ;
        RECT 142.965 139.065 143.295 139.445 ;
        RECT 143.475 139.235 143.645 139.615 ;
        RECT 143.995 139.615 144.710 139.785 ;
        RECT 143.995 139.235 144.165 139.615 ;
        RECT 144.380 139.065 144.710 139.445 ;
        RECT 144.880 139.235 145.135 139.810 ;
        RECT 145.310 139.065 145.570 139.905 ;
        RECT 146.435 139.815 146.955 140.355 ;
        RECT 145.745 139.065 146.955 139.815 ;
        RECT 17.320 138.895 147.040 139.065 ;
        RECT 17.405 138.145 18.615 138.895 ;
        RECT 17.405 137.605 17.925 138.145 ;
        RECT 18.790 138.055 19.050 138.895 ;
        RECT 19.225 138.150 19.480 138.725 ;
        RECT 19.650 138.515 19.980 138.895 ;
        RECT 20.195 138.345 20.365 138.725 ;
        RECT 20.625 138.350 25.970 138.895 ;
        RECT 19.650 138.175 20.365 138.345 ;
        RECT 18.095 137.435 18.615 137.975 ;
        RECT 17.405 136.345 18.615 137.435 ;
        RECT 18.790 136.345 19.050 137.495 ;
        RECT 19.225 137.420 19.395 138.150 ;
        RECT 19.650 137.985 19.820 138.175 ;
        RECT 19.565 137.655 19.820 137.985 ;
        RECT 19.650 137.445 19.820 137.655 ;
        RECT 20.100 137.625 20.455 137.995 ;
        RECT 22.210 137.520 22.550 138.350 ;
        RECT 26.145 138.125 28.735 138.895 ;
        RECT 29.415 138.240 29.745 138.675 ;
        RECT 29.915 138.285 30.085 138.895 ;
        RECT 29.365 138.155 29.745 138.240 ;
        RECT 30.255 138.155 30.585 138.680 ;
        RECT 30.845 138.365 31.055 138.895 ;
        RECT 31.330 138.445 32.115 138.615 ;
        RECT 32.285 138.445 32.690 138.615 ;
        RECT 19.225 136.515 19.480 137.420 ;
        RECT 19.650 137.275 20.365 137.445 ;
        RECT 19.650 136.345 19.980 137.105 ;
        RECT 20.195 136.515 20.365 137.275 ;
        RECT 24.030 136.780 24.380 138.030 ;
        RECT 26.145 137.605 27.355 138.125 ;
        RECT 29.365 138.115 29.590 138.155 ;
        RECT 27.525 137.435 28.735 137.955 ;
        RECT 20.625 136.345 25.970 136.780 ;
        RECT 26.145 136.345 28.735 137.435 ;
        RECT 29.365 137.535 29.535 138.115 ;
        RECT 30.255 137.985 30.455 138.155 ;
        RECT 31.330 137.985 31.500 138.445 ;
        RECT 29.705 137.655 30.455 137.985 ;
        RECT 30.625 137.655 31.500 137.985 ;
        RECT 29.365 137.485 29.580 137.535 ;
        RECT 29.365 137.405 29.755 137.485 ;
        RECT 29.425 136.560 29.755 137.405 ;
        RECT 30.265 137.450 30.455 137.655 ;
        RECT 29.925 136.345 30.095 137.355 ;
        RECT 30.265 137.075 31.160 137.450 ;
        RECT 30.265 136.515 30.605 137.075 ;
        RECT 30.835 136.345 31.150 136.845 ;
        RECT 31.330 136.815 31.500 137.655 ;
        RECT 31.670 137.945 32.135 138.275 ;
        RECT 32.520 138.215 32.690 138.445 ;
        RECT 32.870 138.395 33.240 138.895 ;
        RECT 33.560 138.445 34.235 138.615 ;
        RECT 34.430 138.445 34.765 138.615 ;
        RECT 31.670 136.985 31.990 137.945 ;
        RECT 32.520 137.915 33.350 138.215 ;
        RECT 32.160 137.015 32.350 137.735 ;
        RECT 32.520 136.845 32.690 137.915 ;
        RECT 33.150 137.885 33.350 137.915 ;
        RECT 32.860 137.665 33.030 137.735 ;
        RECT 33.560 137.665 33.730 138.445 ;
        RECT 34.595 138.305 34.765 138.445 ;
        RECT 34.935 138.435 35.185 138.895 ;
        RECT 32.860 137.495 33.730 137.665 ;
        RECT 33.900 138.025 34.425 138.245 ;
        RECT 34.595 138.175 34.820 138.305 ;
        RECT 32.860 137.405 33.370 137.495 ;
        RECT 31.330 136.645 32.215 136.815 ;
        RECT 32.440 136.515 32.690 136.845 ;
        RECT 32.860 136.345 33.030 137.145 ;
        RECT 33.200 136.790 33.370 137.405 ;
        RECT 33.900 137.325 34.070 138.025 ;
        RECT 33.540 136.960 34.070 137.325 ;
        RECT 34.240 137.260 34.480 137.855 ;
        RECT 34.650 137.070 34.820 138.175 ;
        RECT 34.990 137.315 35.270 138.265 ;
        RECT 34.515 136.940 34.820 137.070 ;
        RECT 33.200 136.620 34.305 136.790 ;
        RECT 34.515 136.515 34.765 136.940 ;
        RECT 34.935 136.345 35.200 136.805 ;
        RECT 35.440 136.515 35.625 138.635 ;
        RECT 35.795 138.515 36.125 138.895 ;
        RECT 36.295 138.345 36.465 138.635 ;
        RECT 35.800 138.175 36.465 138.345 ;
        RECT 35.800 137.185 36.030 138.175 ;
        RECT 36.725 138.145 37.935 138.895 ;
        RECT 38.140 138.155 38.755 138.725 ;
        RECT 38.925 138.385 39.140 138.895 ;
        RECT 39.370 138.385 39.650 138.715 ;
        RECT 39.830 138.385 40.070 138.895 ;
        RECT 36.200 137.355 36.550 138.005 ;
        RECT 36.725 137.605 37.245 138.145 ;
        RECT 37.415 137.435 37.935 137.975 ;
        RECT 35.800 137.015 36.465 137.185 ;
        RECT 35.795 136.345 36.125 136.845 ;
        RECT 36.295 136.515 36.465 137.015 ;
        RECT 36.725 136.345 37.935 137.435 ;
        RECT 38.140 137.135 38.455 138.155 ;
        RECT 38.625 137.485 38.795 137.985 ;
        RECT 39.045 137.655 39.310 138.215 ;
        RECT 39.480 137.485 39.650 138.385 ;
        RECT 39.820 137.655 40.175 138.215 ;
        RECT 38.625 137.315 40.050 137.485 ;
        RECT 38.140 136.515 38.675 137.135 ;
        RECT 38.845 136.345 39.175 137.145 ;
        RECT 39.660 137.140 40.050 137.315 ;
        RECT 40.415 136.525 40.675 138.715 ;
        RECT 40.935 138.525 41.605 138.895 ;
        RECT 41.785 138.345 42.095 138.715 ;
        RECT 40.865 138.145 42.095 138.345 ;
        RECT 40.865 137.475 41.155 138.145 ;
        RECT 42.275 137.965 42.505 138.605 ;
        RECT 42.685 138.165 42.975 138.895 ;
        RECT 43.165 138.170 43.455 138.895 ;
        RECT 44.715 138.435 44.970 138.895 ;
        RECT 45.140 138.265 45.470 138.725 ;
        RECT 45.640 138.435 45.810 138.895 ;
        RECT 45.980 138.265 46.310 138.725 ;
        RECT 46.480 138.435 46.650 138.895 ;
        RECT 46.820 138.265 47.150 138.725 ;
        RECT 47.320 138.435 47.490 138.895 ;
        RECT 47.660 138.265 47.990 138.725 ;
        RECT 48.160 138.435 48.465 138.895 ;
        RECT 49.345 138.265 49.675 138.625 ;
        RECT 50.295 138.435 50.545 138.895 ;
        RECT 50.715 138.435 51.275 138.725 ;
        RECT 44.545 138.075 48.515 138.265 ;
        RECT 49.345 138.075 50.735 138.265 ;
        RECT 41.335 137.655 41.800 137.965 ;
        RECT 41.980 137.655 42.505 137.965 ;
        RECT 42.685 137.655 42.985 137.985 ;
        RECT 40.865 137.255 41.635 137.475 ;
        RECT 40.845 136.345 41.185 137.075 ;
        RECT 41.365 136.525 41.635 137.255 ;
        RECT 41.815 137.235 42.975 137.475 ;
        RECT 41.815 136.525 42.045 137.235 ;
        RECT 42.215 136.345 42.545 137.055 ;
        RECT 42.715 136.525 42.975 137.235 ;
        RECT 43.165 136.345 43.455 137.510 ;
        RECT 44.545 137.485 44.890 138.075 ;
        RECT 45.140 137.655 47.995 137.905 ;
        RECT 48.195 137.485 48.515 138.075 ;
        RECT 50.565 137.985 50.735 138.075 ;
        RECT 44.545 137.315 48.515 137.485 ;
        RECT 49.160 137.655 49.835 137.905 ;
        RECT 50.055 137.655 50.395 137.905 ;
        RECT 50.565 137.655 50.855 137.985 ;
        RECT 44.715 136.345 44.970 137.145 ;
        RECT 45.140 136.515 45.470 137.315 ;
        RECT 45.640 136.345 45.810 137.145 ;
        RECT 45.980 136.515 46.310 137.315 ;
        RECT 46.480 136.345 46.650 137.145 ;
        RECT 46.820 136.515 47.150 137.315 ;
        RECT 47.320 136.345 47.490 137.145 ;
        RECT 47.660 136.515 47.990 137.315 ;
        RECT 49.160 137.295 49.425 137.655 ;
        RECT 50.565 137.405 50.735 137.655 ;
        RECT 49.795 137.235 50.735 137.405 ;
        RECT 48.160 136.345 48.460 137.145 ;
        RECT 49.345 136.345 49.625 137.015 ;
        RECT 49.795 136.685 50.095 137.235 ;
        RECT 51.025 137.065 51.275 138.435 ;
        RECT 51.445 138.075 51.705 138.895 ;
        RECT 51.875 138.075 52.205 138.495 ;
        RECT 52.385 138.410 53.175 138.675 ;
        RECT 51.955 137.985 52.205 138.075 ;
        RECT 50.295 136.345 50.625 137.065 ;
        RECT 50.815 136.515 51.275 137.065 ;
        RECT 51.445 137.025 51.785 137.905 ;
        RECT 51.955 137.735 52.750 137.985 ;
        RECT 51.445 136.345 51.705 136.855 ;
        RECT 51.955 136.515 52.125 137.735 ;
        RECT 52.920 137.555 53.175 138.410 ;
        RECT 53.345 138.255 53.545 138.675 ;
        RECT 53.735 138.435 54.065 138.895 ;
        RECT 53.345 137.735 53.755 138.255 ;
        RECT 54.235 138.245 54.495 138.725 ;
        RECT 53.925 137.555 54.155 137.985 ;
        RECT 52.365 137.385 54.155 137.555 ;
        RECT 52.365 137.020 52.615 137.385 ;
        RECT 52.785 137.025 53.115 137.215 ;
        RECT 53.335 137.090 54.050 137.385 ;
        RECT 54.325 137.215 54.495 138.245 ;
        RECT 55.635 138.240 55.965 138.675 ;
        RECT 56.135 138.285 56.305 138.895 ;
        RECT 55.585 138.155 55.965 138.240 ;
        RECT 56.475 138.155 56.805 138.680 ;
        RECT 57.065 138.365 57.275 138.895 ;
        RECT 57.550 138.445 58.335 138.615 ;
        RECT 58.505 138.445 58.910 138.615 ;
        RECT 55.585 138.115 55.810 138.155 ;
        RECT 55.585 137.535 55.755 138.115 ;
        RECT 56.475 137.985 56.675 138.155 ;
        RECT 57.550 137.985 57.720 138.445 ;
        RECT 55.925 137.655 56.675 137.985 ;
        RECT 56.845 137.655 57.720 137.985 ;
        RECT 55.585 137.485 55.800 137.535 ;
        RECT 55.585 137.405 55.975 137.485 ;
        RECT 52.785 136.850 52.980 137.025 ;
        RECT 52.365 136.345 52.980 136.850 ;
        RECT 53.150 136.515 53.625 136.855 ;
        RECT 53.795 136.345 54.010 136.890 ;
        RECT 54.220 136.515 54.495 137.215 ;
        RECT 55.645 136.560 55.975 137.405 ;
        RECT 56.485 137.450 56.675 137.655 ;
        RECT 56.145 136.345 56.315 137.355 ;
        RECT 56.485 137.075 57.380 137.450 ;
        RECT 56.485 136.515 56.825 137.075 ;
        RECT 57.055 136.345 57.370 136.845 ;
        RECT 57.550 136.815 57.720 137.655 ;
        RECT 57.890 137.945 58.355 138.275 ;
        RECT 58.740 138.215 58.910 138.445 ;
        RECT 59.090 138.395 59.460 138.895 ;
        RECT 59.780 138.445 60.455 138.615 ;
        RECT 60.650 138.445 60.985 138.615 ;
        RECT 57.890 136.985 58.210 137.945 ;
        RECT 58.740 137.915 59.570 138.215 ;
        RECT 58.380 137.015 58.570 137.735 ;
        RECT 58.740 136.845 58.910 137.915 ;
        RECT 59.370 137.885 59.570 137.915 ;
        RECT 59.080 137.665 59.250 137.735 ;
        RECT 59.780 137.665 59.950 138.445 ;
        RECT 60.815 138.305 60.985 138.445 ;
        RECT 61.155 138.435 61.405 138.895 ;
        RECT 59.080 137.495 59.950 137.665 ;
        RECT 60.120 138.025 60.645 138.245 ;
        RECT 60.815 138.175 61.040 138.305 ;
        RECT 59.080 137.405 59.590 137.495 ;
        RECT 57.550 136.645 58.435 136.815 ;
        RECT 58.660 136.515 58.910 136.845 ;
        RECT 59.080 136.345 59.250 137.145 ;
        RECT 59.420 136.790 59.590 137.405 ;
        RECT 60.120 137.325 60.290 138.025 ;
        RECT 59.760 136.960 60.290 137.325 ;
        RECT 60.460 137.260 60.700 137.855 ;
        RECT 60.870 137.070 61.040 138.175 ;
        RECT 61.210 137.315 61.490 138.265 ;
        RECT 60.735 136.940 61.040 137.070 ;
        RECT 59.420 136.620 60.525 136.790 ;
        RECT 60.735 136.515 60.985 136.940 ;
        RECT 61.155 136.345 61.420 136.805 ;
        RECT 61.660 136.515 61.845 138.635 ;
        RECT 62.015 138.515 62.345 138.895 ;
        RECT 62.515 138.345 62.685 138.635 ;
        RECT 62.020 138.175 62.685 138.345 ;
        RECT 62.020 137.185 62.250 138.175 ;
        RECT 62.980 138.155 63.595 138.725 ;
        RECT 63.765 138.385 63.980 138.895 ;
        RECT 64.210 138.385 64.490 138.715 ;
        RECT 64.670 138.385 64.910 138.895 ;
        RECT 62.420 137.355 62.770 138.005 ;
        RECT 62.020 137.015 62.685 137.185 ;
        RECT 62.015 136.345 62.345 136.845 ;
        RECT 62.515 136.515 62.685 137.015 ;
        RECT 62.980 137.135 63.295 138.155 ;
        RECT 63.465 137.485 63.635 137.985 ;
        RECT 63.885 137.655 64.150 138.215 ;
        RECT 64.320 137.485 64.490 138.385 ;
        RECT 64.660 137.655 65.015 138.215 ;
        RECT 65.245 138.125 68.755 138.895 ;
        RECT 68.925 138.170 69.215 138.895 ;
        RECT 70.395 138.345 70.565 138.635 ;
        RECT 70.735 138.515 71.065 138.895 ;
        RECT 70.395 138.175 71.060 138.345 ;
        RECT 65.245 137.605 66.895 138.125 ;
        RECT 63.465 137.315 64.890 137.485 ;
        RECT 67.065 137.435 68.755 137.955 ;
        RECT 62.980 136.515 63.515 137.135 ;
        RECT 63.685 136.345 64.015 137.145 ;
        RECT 64.500 137.140 64.890 137.315 ;
        RECT 65.245 136.345 68.755 137.435 ;
        RECT 68.925 136.345 69.215 137.510 ;
        RECT 70.310 137.355 70.660 138.005 ;
        RECT 70.830 137.185 71.060 138.175 ;
        RECT 70.395 137.015 71.060 137.185 ;
        RECT 70.395 136.515 70.565 137.015 ;
        RECT 70.735 136.345 71.065 136.845 ;
        RECT 71.235 136.515 71.420 138.635 ;
        RECT 71.675 138.435 71.925 138.895 ;
        RECT 72.095 138.445 72.430 138.615 ;
        RECT 72.625 138.445 73.300 138.615 ;
        RECT 72.095 138.305 72.265 138.445 ;
        RECT 71.590 137.315 71.870 138.265 ;
        RECT 72.040 138.175 72.265 138.305 ;
        RECT 72.040 137.070 72.210 138.175 ;
        RECT 72.435 138.025 72.960 138.245 ;
        RECT 72.380 137.260 72.620 137.855 ;
        RECT 72.790 137.325 72.960 138.025 ;
        RECT 73.130 137.665 73.300 138.445 ;
        RECT 73.620 138.395 73.990 138.895 ;
        RECT 74.170 138.445 74.575 138.615 ;
        RECT 74.745 138.445 75.530 138.615 ;
        RECT 74.170 138.215 74.340 138.445 ;
        RECT 73.510 137.915 74.340 138.215 ;
        RECT 74.725 137.945 75.190 138.275 ;
        RECT 73.510 137.885 73.710 137.915 ;
        RECT 73.830 137.665 74.000 137.735 ;
        RECT 73.130 137.495 74.000 137.665 ;
        RECT 73.490 137.405 74.000 137.495 ;
        RECT 72.040 136.940 72.345 137.070 ;
        RECT 72.790 136.960 73.320 137.325 ;
        RECT 71.660 136.345 71.925 136.805 ;
        RECT 72.095 136.515 72.345 136.940 ;
        RECT 73.490 136.790 73.660 137.405 ;
        RECT 72.555 136.620 73.660 136.790 ;
        RECT 73.830 136.345 74.000 137.145 ;
        RECT 74.170 136.845 74.340 137.915 ;
        RECT 74.510 137.015 74.700 137.735 ;
        RECT 74.870 136.985 75.190 137.945 ;
        RECT 75.360 137.985 75.530 138.445 ;
        RECT 75.805 138.365 76.015 138.895 ;
        RECT 76.275 138.155 76.605 138.680 ;
        RECT 76.775 138.285 76.945 138.895 ;
        RECT 77.115 138.240 77.445 138.675 ;
        RECT 78.700 138.265 78.985 138.725 ;
        RECT 79.155 138.435 79.425 138.895 ;
        RECT 77.115 138.155 77.495 138.240 ;
        RECT 76.405 137.985 76.605 138.155 ;
        RECT 77.270 138.115 77.495 138.155 ;
        RECT 75.360 137.655 76.235 137.985 ;
        RECT 76.405 137.655 77.155 137.985 ;
        RECT 74.170 136.515 74.420 136.845 ;
        RECT 75.360 136.815 75.530 137.655 ;
        RECT 76.405 137.450 76.595 137.655 ;
        RECT 77.325 137.535 77.495 138.115 ;
        RECT 78.700 138.095 79.655 138.265 ;
        RECT 77.280 137.485 77.495 137.535 ;
        RECT 75.700 137.075 76.595 137.450 ;
        RECT 77.105 137.405 77.495 137.485 ;
        RECT 74.645 136.645 75.530 136.815 ;
        RECT 75.710 136.345 76.025 136.845 ;
        RECT 76.255 136.515 76.595 137.075 ;
        RECT 76.765 136.345 76.935 137.355 ;
        RECT 77.105 136.560 77.435 137.405 ;
        RECT 78.585 137.365 79.275 137.925 ;
        RECT 79.445 137.195 79.655 138.095 ;
        RECT 78.700 136.975 79.655 137.195 ;
        RECT 79.825 137.925 80.225 138.725 ;
        RECT 80.415 138.265 80.695 138.725 ;
        RECT 81.215 138.435 81.540 138.895 ;
        RECT 80.415 138.095 81.540 138.265 ;
        RECT 81.710 138.155 82.095 138.725 ;
        RECT 81.090 137.985 81.540 138.095 ;
        RECT 79.825 137.365 80.920 137.925 ;
        RECT 81.090 137.655 81.645 137.985 ;
        RECT 78.700 136.515 78.985 136.975 ;
        RECT 79.155 136.345 79.425 136.805 ;
        RECT 79.825 136.515 80.225 137.365 ;
        RECT 81.090 137.195 81.540 137.655 ;
        RECT 81.815 137.485 82.095 138.155 ;
        RECT 82.380 138.265 82.665 138.725 ;
        RECT 82.835 138.435 83.105 138.895 ;
        RECT 82.380 138.095 83.335 138.265 ;
        RECT 80.415 136.975 81.540 137.195 ;
        RECT 80.415 136.515 80.695 136.975 ;
        RECT 81.215 136.345 81.540 136.805 ;
        RECT 81.710 136.515 82.095 137.485 ;
        RECT 82.265 137.365 82.955 137.925 ;
        RECT 83.125 137.195 83.335 138.095 ;
        RECT 82.380 136.975 83.335 137.195 ;
        RECT 83.505 137.925 83.905 138.725 ;
        RECT 84.095 138.265 84.375 138.725 ;
        RECT 84.895 138.435 85.220 138.895 ;
        RECT 84.095 138.095 85.220 138.265 ;
        RECT 85.390 138.155 85.775 138.725 ;
        RECT 85.965 138.325 86.220 138.675 ;
        RECT 86.390 138.495 86.720 138.895 ;
        RECT 86.890 138.325 87.060 138.675 ;
        RECT 87.230 138.495 87.610 138.895 ;
        RECT 85.965 138.155 87.630 138.325 ;
        RECT 87.800 138.220 88.075 138.565 ;
        RECT 84.770 137.985 85.220 138.095 ;
        RECT 83.505 137.365 84.600 137.925 ;
        RECT 84.770 137.655 85.325 137.985 ;
        RECT 82.380 136.515 82.665 136.975 ;
        RECT 82.835 136.345 83.105 136.805 ;
        RECT 83.505 136.515 83.905 137.365 ;
        RECT 84.770 137.195 85.220 137.655 ;
        RECT 85.495 137.485 85.775 138.155 ;
        RECT 87.460 137.985 87.630 138.155 ;
        RECT 85.945 137.655 86.295 137.985 ;
        RECT 86.465 137.655 87.290 137.985 ;
        RECT 87.460 137.655 87.735 137.985 ;
        RECT 84.095 136.975 85.220 137.195 ;
        RECT 84.095 136.515 84.375 136.975 ;
        RECT 84.895 136.345 85.220 136.805 ;
        RECT 85.390 136.515 85.775 137.485 ;
        RECT 85.965 137.195 86.295 137.485 ;
        RECT 86.465 137.365 86.690 137.655 ;
        RECT 87.460 137.485 87.630 137.655 ;
        RECT 87.905 137.485 88.075 138.220 ;
        RECT 88.245 138.065 88.535 138.895 ;
        RECT 88.705 138.350 94.050 138.895 ;
        RECT 86.960 137.315 87.630 137.485 ;
        RECT 86.960 137.195 87.130 137.315 ;
        RECT 85.965 137.025 87.130 137.195 ;
        RECT 85.945 136.565 87.140 136.855 ;
        RECT 87.310 136.345 87.590 137.145 ;
        RECT 87.800 136.515 88.075 137.485 ;
        RECT 88.245 136.345 88.535 137.550 ;
        RECT 90.290 137.520 90.630 138.350 ;
        RECT 94.685 138.170 94.975 138.895 ;
        RECT 95.145 138.125 97.735 138.895 ;
        RECT 97.955 138.355 98.180 138.715 ;
        RECT 98.360 138.525 98.690 138.895 ;
        RECT 98.870 138.355 99.125 138.715 ;
        RECT 99.690 138.525 100.435 138.895 ;
        RECT 97.955 138.165 100.440 138.355 ;
        RECT 92.110 136.780 92.460 138.030 ;
        RECT 95.145 137.605 96.355 138.125 ;
        RECT 88.705 136.345 94.050 136.780 ;
        RECT 94.685 136.345 94.975 137.510 ;
        RECT 96.525 137.435 97.735 137.955 ;
        RECT 97.915 137.655 98.185 137.985 ;
        RECT 98.365 137.655 98.800 137.985 ;
        RECT 98.980 137.655 99.555 137.985 ;
        RECT 99.735 137.655 100.015 137.985 ;
        RECT 100.215 137.475 100.440 138.165 ;
        RECT 95.145 136.345 97.735 137.435 ;
        RECT 97.945 137.295 100.440 137.475 ;
        RECT 100.615 137.295 100.950 138.715 ;
        RECT 102.135 138.345 102.305 138.635 ;
        RECT 102.475 138.515 102.805 138.895 ;
        RECT 102.135 138.175 102.800 138.345 ;
        RECT 102.050 137.355 102.400 138.005 ;
        RECT 97.945 136.525 98.235 137.295 ;
        RECT 98.805 136.885 99.995 137.115 ;
        RECT 98.805 136.525 99.065 136.885 ;
        RECT 99.235 136.345 99.565 136.715 ;
        RECT 99.735 136.525 99.995 136.885 ;
        RECT 100.185 136.345 100.515 137.065 ;
        RECT 100.685 136.525 100.950 137.295 ;
        RECT 102.570 137.185 102.800 138.175 ;
        RECT 102.135 137.015 102.800 137.185 ;
        RECT 102.135 136.515 102.305 137.015 ;
        RECT 102.475 136.345 102.805 136.845 ;
        RECT 102.975 136.515 103.160 138.635 ;
        RECT 103.415 138.435 103.665 138.895 ;
        RECT 103.835 138.445 104.170 138.615 ;
        RECT 104.365 138.445 105.040 138.615 ;
        RECT 103.835 138.305 104.005 138.445 ;
        RECT 103.330 137.315 103.610 138.265 ;
        RECT 103.780 138.175 104.005 138.305 ;
        RECT 103.780 137.070 103.950 138.175 ;
        RECT 104.175 138.025 104.700 138.245 ;
        RECT 104.120 137.260 104.360 137.855 ;
        RECT 104.530 137.325 104.700 138.025 ;
        RECT 104.870 137.665 105.040 138.445 ;
        RECT 105.360 138.395 105.730 138.895 ;
        RECT 105.910 138.445 106.315 138.615 ;
        RECT 106.485 138.445 107.270 138.615 ;
        RECT 105.910 138.215 106.080 138.445 ;
        RECT 105.250 137.915 106.080 138.215 ;
        RECT 106.465 137.945 106.930 138.275 ;
        RECT 105.250 137.885 105.450 137.915 ;
        RECT 105.570 137.665 105.740 137.735 ;
        RECT 104.870 137.495 105.740 137.665 ;
        RECT 105.230 137.405 105.740 137.495 ;
        RECT 103.780 136.940 104.085 137.070 ;
        RECT 104.530 136.960 105.060 137.325 ;
        RECT 103.400 136.345 103.665 136.805 ;
        RECT 103.835 136.515 104.085 136.940 ;
        RECT 105.230 136.790 105.400 137.405 ;
        RECT 104.295 136.620 105.400 136.790 ;
        RECT 105.570 136.345 105.740 137.145 ;
        RECT 105.910 136.845 106.080 137.915 ;
        RECT 106.250 137.015 106.440 137.735 ;
        RECT 106.610 136.985 106.930 137.945 ;
        RECT 107.100 137.985 107.270 138.445 ;
        RECT 107.545 138.365 107.755 138.895 ;
        RECT 108.015 138.155 108.345 138.680 ;
        RECT 108.515 138.285 108.685 138.895 ;
        RECT 108.855 138.240 109.185 138.675 ;
        RECT 109.495 138.345 109.665 138.635 ;
        RECT 109.835 138.515 110.165 138.895 ;
        RECT 108.855 138.155 109.235 138.240 ;
        RECT 109.495 138.175 110.160 138.345 ;
        RECT 108.145 137.985 108.345 138.155 ;
        RECT 109.010 138.115 109.235 138.155 ;
        RECT 107.100 137.655 107.975 137.985 ;
        RECT 108.145 137.655 108.895 137.985 ;
        RECT 105.910 136.515 106.160 136.845 ;
        RECT 107.100 136.815 107.270 137.655 ;
        RECT 108.145 137.450 108.335 137.655 ;
        RECT 109.065 137.535 109.235 138.115 ;
        RECT 109.020 137.485 109.235 137.535 ;
        RECT 107.440 137.075 108.335 137.450 ;
        RECT 108.845 137.405 109.235 137.485 ;
        RECT 106.385 136.645 107.270 136.815 ;
        RECT 107.450 136.345 107.765 136.845 ;
        RECT 107.995 136.515 108.335 137.075 ;
        RECT 108.505 136.345 108.675 137.355 ;
        RECT 108.845 136.560 109.175 137.405 ;
        RECT 109.410 137.355 109.760 138.005 ;
        RECT 109.930 137.185 110.160 138.175 ;
        RECT 109.495 137.015 110.160 137.185 ;
        RECT 109.495 136.515 109.665 137.015 ;
        RECT 109.835 136.345 110.165 136.845 ;
        RECT 110.335 136.515 110.520 138.635 ;
        RECT 110.775 138.435 111.025 138.895 ;
        RECT 111.195 138.445 111.530 138.615 ;
        RECT 111.725 138.445 112.400 138.615 ;
        RECT 111.195 138.305 111.365 138.445 ;
        RECT 110.690 137.315 110.970 138.265 ;
        RECT 111.140 138.175 111.365 138.305 ;
        RECT 111.140 137.070 111.310 138.175 ;
        RECT 111.535 138.025 112.060 138.245 ;
        RECT 111.480 137.260 111.720 137.855 ;
        RECT 111.890 137.325 112.060 138.025 ;
        RECT 112.230 137.665 112.400 138.445 ;
        RECT 112.720 138.395 113.090 138.895 ;
        RECT 113.270 138.445 113.675 138.615 ;
        RECT 113.845 138.445 114.630 138.615 ;
        RECT 113.270 138.215 113.440 138.445 ;
        RECT 112.610 137.915 113.440 138.215 ;
        RECT 113.825 137.945 114.290 138.275 ;
        RECT 112.610 137.885 112.810 137.915 ;
        RECT 112.930 137.665 113.100 137.735 ;
        RECT 112.230 137.495 113.100 137.665 ;
        RECT 112.590 137.405 113.100 137.495 ;
        RECT 111.140 136.940 111.445 137.070 ;
        RECT 111.890 136.960 112.420 137.325 ;
        RECT 110.760 136.345 111.025 136.805 ;
        RECT 111.195 136.515 111.445 136.940 ;
        RECT 112.590 136.790 112.760 137.405 ;
        RECT 111.655 136.620 112.760 136.790 ;
        RECT 112.930 136.345 113.100 137.145 ;
        RECT 113.270 136.845 113.440 137.915 ;
        RECT 113.610 137.015 113.800 137.735 ;
        RECT 113.970 136.985 114.290 137.945 ;
        RECT 114.460 137.985 114.630 138.445 ;
        RECT 114.905 138.365 115.115 138.895 ;
        RECT 115.375 138.155 115.705 138.680 ;
        RECT 115.875 138.285 116.045 138.895 ;
        RECT 116.215 138.240 116.545 138.675 ;
        RECT 116.215 138.155 116.595 138.240 ;
        RECT 115.505 137.985 115.705 138.155 ;
        RECT 116.370 138.115 116.595 138.155 ;
        RECT 114.460 137.655 115.335 137.985 ;
        RECT 115.505 137.655 116.255 137.985 ;
        RECT 113.270 136.515 113.520 136.845 ;
        RECT 114.460 136.815 114.630 137.655 ;
        RECT 115.505 137.450 115.695 137.655 ;
        RECT 116.425 137.535 116.595 138.115 ;
        RECT 116.765 138.125 120.275 138.895 ;
        RECT 120.445 138.170 120.735 138.895 ;
        RECT 120.905 138.155 121.290 138.725 ;
        RECT 121.460 138.435 121.785 138.895 ;
        RECT 122.305 138.265 122.585 138.725 ;
        RECT 116.765 137.605 118.415 138.125 ;
        RECT 116.380 137.485 116.595 137.535 ;
        RECT 114.800 137.075 115.695 137.450 ;
        RECT 116.205 137.405 116.595 137.485 ;
        RECT 118.585 137.435 120.275 137.955 ;
        RECT 113.745 136.645 114.630 136.815 ;
        RECT 114.810 136.345 115.125 136.845 ;
        RECT 115.355 136.515 115.695 137.075 ;
        RECT 115.865 136.345 116.035 137.355 ;
        RECT 116.205 136.560 116.535 137.405 ;
        RECT 116.765 136.345 120.275 137.435 ;
        RECT 120.445 136.345 120.735 137.510 ;
        RECT 120.905 137.485 121.185 138.155 ;
        RECT 121.460 138.095 122.585 138.265 ;
        RECT 121.460 137.985 121.910 138.095 ;
        RECT 121.355 137.655 121.910 137.985 ;
        RECT 122.775 137.925 123.175 138.725 ;
        RECT 123.575 138.435 123.845 138.895 ;
        RECT 124.015 138.265 124.300 138.725 ;
        RECT 120.905 136.515 121.290 137.485 ;
        RECT 121.460 137.195 121.910 137.655 ;
        RECT 122.080 137.365 123.175 137.925 ;
        RECT 121.460 136.975 122.585 137.195 ;
        RECT 121.460 136.345 121.785 136.805 ;
        RECT 122.305 136.515 122.585 136.975 ;
        RECT 122.775 136.515 123.175 137.365 ;
        RECT 123.345 138.095 124.300 138.265 ;
        RECT 124.585 138.125 128.095 138.895 ;
        RECT 128.265 138.145 129.475 138.895 ;
        RECT 123.345 137.195 123.555 138.095 ;
        RECT 123.725 137.365 124.415 137.925 ;
        RECT 124.585 137.605 126.235 138.125 ;
        RECT 126.405 137.435 128.095 137.955 ;
        RECT 128.265 137.605 128.785 138.145 ;
        RECT 129.650 138.130 130.105 138.895 ;
        RECT 130.380 138.515 131.680 138.725 ;
        RECT 131.935 138.535 132.265 138.895 ;
        RECT 131.510 138.365 131.680 138.515 ;
        RECT 132.435 138.395 132.695 138.725 ;
        RECT 128.955 137.435 129.475 137.975 ;
        RECT 130.580 137.905 130.800 138.305 ;
        RECT 129.645 137.705 130.135 137.905 ;
        RECT 130.325 137.695 130.800 137.905 ;
        RECT 131.045 137.905 131.255 138.305 ;
        RECT 131.510 138.240 132.265 138.365 ;
        RECT 131.510 138.195 132.355 138.240 ;
        RECT 132.085 138.075 132.355 138.195 ;
        RECT 131.045 137.695 131.375 137.905 ;
        RECT 131.545 137.635 131.955 137.940 ;
        RECT 123.345 136.975 124.300 137.195 ;
        RECT 123.575 136.345 123.845 136.805 ;
        RECT 124.015 136.515 124.300 136.975 ;
        RECT 124.585 136.345 128.095 137.435 ;
        RECT 128.265 136.345 129.475 137.435 ;
        RECT 129.650 137.465 130.825 137.525 ;
        RECT 132.185 137.500 132.355 138.075 ;
        RECT 132.155 137.465 132.355 137.500 ;
        RECT 129.650 137.355 132.355 137.465 ;
        RECT 129.650 136.735 129.905 137.355 ;
        RECT 130.495 137.295 132.295 137.355 ;
        RECT 130.495 137.265 130.825 137.295 ;
        RECT 132.525 137.195 132.695 138.395 ;
        RECT 133.415 138.345 133.585 138.635 ;
        RECT 133.755 138.515 134.085 138.895 ;
        RECT 133.415 138.175 134.080 138.345 ;
        RECT 133.330 137.355 133.680 138.005 ;
        RECT 130.155 137.095 130.340 137.185 ;
        RECT 130.930 137.095 131.765 137.105 ;
        RECT 130.155 136.895 131.765 137.095 ;
        RECT 130.155 136.855 130.385 136.895 ;
        RECT 129.650 136.515 129.985 136.735 ;
        RECT 130.990 136.345 131.345 136.725 ;
        RECT 131.515 136.515 131.765 136.895 ;
        RECT 132.015 136.345 132.265 137.125 ;
        RECT 132.435 136.515 132.695 137.195 ;
        RECT 133.850 137.185 134.080 138.175 ;
        RECT 133.415 137.015 134.080 137.185 ;
        RECT 133.415 136.515 133.585 137.015 ;
        RECT 133.755 136.345 134.085 136.845 ;
        RECT 134.255 136.515 134.440 138.635 ;
        RECT 134.695 138.435 134.945 138.895 ;
        RECT 135.115 138.445 135.450 138.615 ;
        RECT 135.645 138.445 136.320 138.615 ;
        RECT 135.115 138.305 135.285 138.445 ;
        RECT 134.610 137.315 134.890 138.265 ;
        RECT 135.060 138.175 135.285 138.305 ;
        RECT 135.060 137.070 135.230 138.175 ;
        RECT 135.455 138.025 135.980 138.245 ;
        RECT 135.400 137.260 135.640 137.855 ;
        RECT 135.810 137.325 135.980 138.025 ;
        RECT 136.150 137.665 136.320 138.445 ;
        RECT 136.640 138.395 137.010 138.895 ;
        RECT 137.190 138.445 137.595 138.615 ;
        RECT 137.765 138.445 138.550 138.615 ;
        RECT 137.190 138.215 137.360 138.445 ;
        RECT 136.530 137.915 137.360 138.215 ;
        RECT 137.745 137.945 138.210 138.275 ;
        RECT 136.530 137.885 136.730 137.915 ;
        RECT 136.850 137.665 137.020 137.735 ;
        RECT 136.150 137.495 137.020 137.665 ;
        RECT 136.510 137.405 137.020 137.495 ;
        RECT 135.060 136.940 135.365 137.070 ;
        RECT 135.810 136.960 136.340 137.325 ;
        RECT 134.680 136.345 134.945 136.805 ;
        RECT 135.115 136.515 135.365 136.940 ;
        RECT 136.510 136.790 136.680 137.405 ;
        RECT 135.575 136.620 136.680 136.790 ;
        RECT 136.850 136.345 137.020 137.145 ;
        RECT 137.190 136.845 137.360 137.915 ;
        RECT 137.530 137.015 137.720 137.735 ;
        RECT 137.890 136.985 138.210 137.945 ;
        RECT 138.380 137.985 138.550 138.445 ;
        RECT 138.825 138.365 139.035 138.895 ;
        RECT 139.295 138.155 139.625 138.680 ;
        RECT 139.795 138.285 139.965 138.895 ;
        RECT 140.135 138.240 140.465 138.675 ;
        RECT 140.775 138.345 140.945 138.725 ;
        RECT 141.125 138.515 141.455 138.895 ;
        RECT 140.135 138.155 140.515 138.240 ;
        RECT 140.775 138.175 141.440 138.345 ;
        RECT 141.635 138.220 141.895 138.725 ;
        RECT 139.425 137.985 139.625 138.155 ;
        RECT 140.290 138.115 140.515 138.155 ;
        RECT 138.380 137.655 139.255 137.985 ;
        RECT 139.425 137.655 140.175 137.985 ;
        RECT 137.190 136.515 137.440 136.845 ;
        RECT 138.380 136.815 138.550 137.655 ;
        RECT 139.425 137.450 139.615 137.655 ;
        RECT 140.345 137.535 140.515 138.115 ;
        RECT 140.705 137.625 141.035 137.995 ;
        RECT 141.270 137.920 141.440 138.175 ;
        RECT 140.300 137.485 140.515 137.535 ;
        RECT 138.720 137.075 139.615 137.450 ;
        RECT 140.125 137.405 140.515 137.485 ;
        RECT 141.270 137.590 141.555 137.920 ;
        RECT 141.270 137.445 141.440 137.590 ;
        RECT 137.665 136.645 138.550 136.815 ;
        RECT 138.730 136.345 139.045 136.845 ;
        RECT 139.275 136.515 139.615 137.075 ;
        RECT 139.785 136.345 139.955 137.355 ;
        RECT 140.125 136.560 140.455 137.405 ;
        RECT 140.775 137.275 141.440 137.445 ;
        RECT 141.725 137.420 141.895 138.220 ;
        RECT 142.155 138.345 142.325 138.725 ;
        RECT 142.540 138.515 142.870 138.895 ;
        RECT 142.155 138.175 142.870 138.345 ;
        RECT 142.065 137.625 142.420 137.995 ;
        RECT 142.700 137.985 142.870 138.175 ;
        RECT 143.040 138.150 143.295 138.725 ;
        RECT 142.700 137.655 142.955 137.985 ;
        RECT 142.700 137.445 142.870 137.655 ;
        RECT 140.775 136.515 140.945 137.275 ;
        RECT 141.125 136.345 141.455 137.105 ;
        RECT 141.625 136.515 141.895 137.420 ;
        RECT 142.155 137.275 142.870 137.445 ;
        RECT 143.125 137.420 143.295 138.150 ;
        RECT 143.470 138.055 143.730 138.895 ;
        RECT 143.995 138.345 144.165 138.725 ;
        RECT 144.380 138.515 144.710 138.895 ;
        RECT 143.995 138.175 144.710 138.345 ;
        RECT 143.905 137.625 144.260 137.995 ;
        RECT 144.540 137.985 144.710 138.175 ;
        RECT 144.880 138.150 145.135 138.725 ;
        RECT 144.540 137.655 144.795 137.985 ;
        RECT 142.155 136.515 142.325 137.275 ;
        RECT 142.540 136.345 142.870 137.105 ;
        RECT 143.040 136.515 143.295 137.420 ;
        RECT 143.470 136.345 143.730 137.495 ;
        RECT 144.540 137.445 144.710 137.655 ;
        RECT 143.995 137.275 144.710 137.445 ;
        RECT 144.965 137.420 145.135 138.150 ;
        RECT 145.310 138.055 145.570 138.895 ;
        RECT 145.745 138.145 146.955 138.895 ;
        RECT 143.995 136.515 144.165 137.275 ;
        RECT 144.380 136.345 144.710 137.105 ;
        RECT 144.880 136.515 145.135 137.420 ;
        RECT 145.310 136.345 145.570 137.495 ;
        RECT 145.745 137.435 146.265 137.975 ;
        RECT 146.435 137.605 146.955 138.145 ;
        RECT 145.745 136.345 146.955 137.435 ;
        RECT 17.320 136.175 147.040 136.345 ;
        RECT 17.405 135.085 18.615 136.175 ;
        RECT 17.405 134.375 17.925 134.915 ;
        RECT 18.095 134.545 18.615 135.085 ;
        RECT 18.790 135.025 19.050 136.175 ;
        RECT 19.225 135.100 19.480 136.005 ;
        RECT 19.650 135.415 19.980 136.175 ;
        RECT 20.195 135.245 20.365 136.005 ;
        RECT 20.625 135.740 25.970 136.175 ;
        RECT 17.405 133.625 18.615 134.375 ;
        RECT 18.790 133.625 19.050 134.465 ;
        RECT 19.225 134.370 19.395 135.100 ;
        RECT 19.650 135.075 20.365 135.245 ;
        RECT 19.650 134.865 19.820 135.075 ;
        RECT 19.565 134.535 19.820 134.865 ;
        RECT 19.225 133.795 19.480 134.370 ;
        RECT 19.650 134.345 19.820 134.535 ;
        RECT 20.100 134.525 20.455 134.895 ;
        RECT 19.650 134.175 20.365 134.345 ;
        RECT 19.650 133.625 19.980 134.005 ;
        RECT 20.195 133.795 20.365 134.175 ;
        RECT 22.210 134.170 22.550 135.000 ;
        RECT 24.030 134.490 24.380 135.740 ;
        RECT 26.145 135.085 29.655 136.175 ;
        RECT 26.145 134.395 27.795 134.915 ;
        RECT 27.965 134.565 29.655 135.085 ;
        RECT 30.285 135.010 30.575 136.175 ;
        RECT 30.745 135.085 34.255 136.175 ;
        RECT 35.345 135.620 35.950 136.175 ;
        RECT 36.125 135.665 36.605 136.005 ;
        RECT 36.775 135.630 37.030 136.175 ;
        RECT 35.345 135.520 35.960 135.620 ;
        RECT 35.775 135.495 35.960 135.520 ;
        RECT 30.745 134.395 32.395 134.915 ;
        RECT 32.565 134.565 34.255 135.085 ;
        RECT 35.345 134.900 35.605 135.350 ;
        RECT 35.775 135.250 36.105 135.495 ;
        RECT 36.275 135.175 37.030 135.425 ;
        RECT 37.200 135.305 37.475 136.005 ;
        RECT 37.645 135.665 37.905 136.175 ;
        RECT 36.260 135.140 37.030 135.175 ;
        RECT 36.245 135.130 37.030 135.140 ;
        RECT 36.240 135.115 37.135 135.130 ;
        RECT 36.220 135.100 37.135 135.115 ;
        RECT 36.200 135.090 37.135 135.100 ;
        RECT 36.175 135.080 37.135 135.090 ;
        RECT 36.105 135.050 37.135 135.080 ;
        RECT 36.085 135.020 37.135 135.050 ;
        RECT 36.065 134.990 37.135 135.020 ;
        RECT 36.035 134.965 37.135 134.990 ;
        RECT 36.000 134.930 37.135 134.965 ;
        RECT 35.970 134.925 37.135 134.930 ;
        RECT 35.970 134.920 36.360 134.925 ;
        RECT 35.970 134.910 36.335 134.920 ;
        RECT 35.970 134.905 36.320 134.910 ;
        RECT 35.970 134.900 36.305 134.905 ;
        RECT 35.345 134.895 36.305 134.900 ;
        RECT 35.345 134.885 36.295 134.895 ;
        RECT 35.345 134.880 36.285 134.885 ;
        RECT 35.345 134.870 36.275 134.880 ;
        RECT 35.345 134.860 36.270 134.870 ;
        RECT 35.345 134.855 36.265 134.860 ;
        RECT 35.345 134.840 36.255 134.855 ;
        RECT 35.345 134.825 36.250 134.840 ;
        RECT 35.345 134.800 36.240 134.825 ;
        RECT 35.345 134.730 36.235 134.800 ;
        RECT 20.625 133.625 25.970 134.170 ;
        RECT 26.145 133.625 29.655 134.395 ;
        RECT 30.285 133.625 30.575 134.350 ;
        RECT 30.745 133.625 34.255 134.395 ;
        RECT 35.345 134.175 35.895 134.560 ;
        RECT 36.065 134.005 36.235 134.730 ;
        RECT 35.345 133.835 36.235 134.005 ;
        RECT 36.405 134.330 36.735 134.755 ;
        RECT 36.905 134.530 37.135 134.925 ;
        RECT 36.405 133.845 36.625 134.330 ;
        RECT 37.305 134.275 37.475 135.305 ;
        RECT 37.645 134.615 37.985 135.495 ;
        RECT 38.155 134.785 38.325 136.005 ;
        RECT 38.565 135.670 39.180 136.175 ;
        RECT 38.565 135.135 38.815 135.500 ;
        RECT 38.985 135.495 39.180 135.670 ;
        RECT 39.350 135.665 39.825 136.005 ;
        RECT 39.995 135.630 40.210 136.175 ;
        RECT 38.985 135.305 39.315 135.495 ;
        RECT 39.535 135.135 40.250 135.430 ;
        RECT 40.420 135.305 40.695 136.005 ;
        RECT 40.955 135.505 41.125 136.005 ;
        RECT 41.295 135.675 41.625 136.175 ;
        RECT 40.955 135.335 41.620 135.505 ;
        RECT 38.565 134.965 40.355 135.135 ;
        RECT 38.155 134.535 38.950 134.785 ;
        RECT 38.155 134.445 38.405 134.535 ;
        RECT 36.795 133.625 37.045 134.165 ;
        RECT 37.215 133.795 37.475 134.275 ;
        RECT 37.645 133.625 37.905 134.445 ;
        RECT 38.075 134.025 38.405 134.445 ;
        RECT 39.120 134.110 39.375 134.965 ;
        RECT 38.585 133.845 39.375 134.110 ;
        RECT 39.545 134.265 39.955 134.785 ;
        RECT 40.125 134.535 40.355 134.965 ;
        RECT 40.525 134.275 40.695 135.305 ;
        RECT 40.870 134.515 41.220 135.165 ;
        RECT 41.390 134.345 41.620 135.335 ;
        RECT 39.545 133.845 39.745 134.265 ;
        RECT 39.935 133.625 40.265 134.085 ;
        RECT 40.435 133.795 40.695 134.275 ;
        RECT 40.955 134.175 41.620 134.345 ;
        RECT 40.955 133.885 41.125 134.175 ;
        RECT 41.295 133.625 41.625 134.005 ;
        RECT 41.795 133.885 41.980 136.005 ;
        RECT 42.220 135.715 42.485 136.175 ;
        RECT 42.655 135.580 42.905 136.005 ;
        RECT 43.115 135.730 44.220 135.900 ;
        RECT 42.600 135.450 42.905 135.580 ;
        RECT 42.150 134.255 42.430 135.205 ;
        RECT 42.600 134.345 42.770 135.450 ;
        RECT 42.940 134.665 43.180 135.260 ;
        RECT 43.350 135.195 43.880 135.560 ;
        RECT 43.350 134.495 43.520 135.195 ;
        RECT 44.050 135.115 44.220 135.730 ;
        RECT 44.390 135.375 44.560 136.175 ;
        RECT 44.730 135.675 44.980 136.005 ;
        RECT 45.205 135.705 46.090 135.875 ;
        RECT 44.050 135.025 44.560 135.115 ;
        RECT 42.600 134.215 42.825 134.345 ;
        RECT 42.995 134.275 43.520 134.495 ;
        RECT 43.690 134.855 44.560 135.025 ;
        RECT 42.235 133.625 42.485 134.085 ;
        RECT 42.655 134.075 42.825 134.215 ;
        RECT 43.690 134.075 43.860 134.855 ;
        RECT 44.390 134.785 44.560 134.855 ;
        RECT 44.070 134.605 44.270 134.635 ;
        RECT 44.730 134.605 44.900 135.675 ;
        RECT 45.070 134.785 45.260 135.505 ;
        RECT 44.070 134.305 44.900 134.605 ;
        RECT 45.430 134.575 45.750 135.535 ;
        RECT 42.655 133.905 42.990 134.075 ;
        RECT 43.185 133.905 43.860 134.075 ;
        RECT 44.180 133.625 44.550 134.125 ;
        RECT 44.730 134.075 44.900 134.305 ;
        RECT 45.285 134.245 45.750 134.575 ;
        RECT 45.920 134.865 46.090 135.705 ;
        RECT 46.270 135.675 46.585 136.175 ;
        RECT 46.815 135.445 47.155 136.005 ;
        RECT 46.260 135.070 47.155 135.445 ;
        RECT 47.325 135.165 47.495 136.175 ;
        RECT 46.965 134.865 47.155 135.070 ;
        RECT 47.665 135.115 47.995 135.960 ;
        RECT 48.225 135.620 48.830 136.175 ;
        RECT 49.005 135.665 49.485 136.005 ;
        RECT 49.655 135.630 49.910 136.175 ;
        RECT 48.225 135.520 48.840 135.620 ;
        RECT 48.655 135.495 48.840 135.520 ;
        RECT 47.665 135.035 48.055 135.115 ;
        RECT 47.840 134.985 48.055 135.035 ;
        RECT 45.920 134.535 46.795 134.865 ;
        RECT 46.965 134.535 47.715 134.865 ;
        RECT 45.920 134.075 46.090 134.535 ;
        RECT 46.965 134.365 47.165 134.535 ;
        RECT 47.885 134.405 48.055 134.985 ;
        RECT 48.225 134.900 48.485 135.350 ;
        RECT 48.655 135.250 48.985 135.495 ;
        RECT 49.155 135.175 49.910 135.425 ;
        RECT 50.080 135.305 50.355 136.005 ;
        RECT 49.140 135.140 49.910 135.175 ;
        RECT 49.125 135.130 49.910 135.140 ;
        RECT 49.120 135.115 50.015 135.130 ;
        RECT 49.100 135.100 50.015 135.115 ;
        RECT 49.080 135.090 50.015 135.100 ;
        RECT 49.055 135.080 50.015 135.090 ;
        RECT 48.985 135.050 50.015 135.080 ;
        RECT 48.965 135.020 50.015 135.050 ;
        RECT 48.945 134.990 50.015 135.020 ;
        RECT 48.915 134.965 50.015 134.990 ;
        RECT 48.880 134.930 50.015 134.965 ;
        RECT 48.850 134.925 50.015 134.930 ;
        RECT 48.850 134.920 49.240 134.925 ;
        RECT 48.850 134.910 49.215 134.920 ;
        RECT 48.850 134.905 49.200 134.910 ;
        RECT 48.850 134.900 49.185 134.905 ;
        RECT 48.225 134.895 49.185 134.900 ;
        RECT 48.225 134.885 49.175 134.895 ;
        RECT 48.225 134.880 49.165 134.885 ;
        RECT 48.225 134.870 49.155 134.880 ;
        RECT 48.225 134.860 49.150 134.870 ;
        RECT 48.225 134.855 49.145 134.860 ;
        RECT 48.225 134.840 49.135 134.855 ;
        RECT 48.225 134.825 49.130 134.840 ;
        RECT 48.225 134.800 49.120 134.825 ;
        RECT 48.225 134.730 49.115 134.800 ;
        RECT 47.830 134.365 48.055 134.405 ;
        RECT 44.730 133.905 45.135 134.075 ;
        RECT 45.305 133.905 46.090 134.075 ;
        RECT 46.365 133.625 46.575 134.155 ;
        RECT 46.835 133.840 47.165 134.365 ;
        RECT 47.675 134.280 48.055 134.365 ;
        RECT 47.335 133.625 47.505 134.235 ;
        RECT 47.675 133.845 48.005 134.280 ;
        RECT 48.225 134.175 48.775 134.560 ;
        RECT 48.945 134.005 49.115 134.730 ;
        RECT 48.225 133.835 49.115 134.005 ;
        RECT 49.285 134.330 49.615 134.755 ;
        RECT 49.785 134.530 50.015 134.925 ;
        RECT 49.285 133.845 49.505 134.330 ;
        RECT 50.185 134.275 50.355 135.305 ;
        RECT 51.630 135.205 52.020 135.380 ;
        RECT 52.505 135.375 52.835 136.175 ;
        RECT 53.005 135.385 53.540 136.005 ;
        RECT 53.745 135.620 54.350 136.175 ;
        RECT 54.525 135.665 55.005 136.005 ;
        RECT 55.175 135.630 55.430 136.175 ;
        RECT 53.745 135.520 54.360 135.620 ;
        RECT 51.630 135.035 53.055 135.205 ;
        RECT 51.505 134.305 51.860 134.865 ;
        RECT 49.675 133.625 49.925 134.165 ;
        RECT 50.095 133.795 50.355 134.275 ;
        RECT 52.030 134.135 52.200 135.035 ;
        RECT 52.370 134.305 52.635 134.865 ;
        RECT 52.885 134.535 53.055 135.035 ;
        RECT 53.225 134.365 53.540 135.385 ;
        RECT 54.175 135.495 54.360 135.520 ;
        RECT 53.745 134.900 54.005 135.350 ;
        RECT 54.175 135.250 54.505 135.495 ;
        RECT 54.675 135.175 55.430 135.425 ;
        RECT 55.600 135.305 55.875 136.005 ;
        RECT 54.660 135.140 55.430 135.175 ;
        RECT 54.645 135.130 55.430 135.140 ;
        RECT 54.640 135.115 55.535 135.130 ;
        RECT 54.620 135.100 55.535 135.115 ;
        RECT 54.600 135.090 55.535 135.100 ;
        RECT 54.575 135.080 55.535 135.090 ;
        RECT 54.505 135.050 55.535 135.080 ;
        RECT 54.485 135.020 55.535 135.050 ;
        RECT 54.465 134.990 55.535 135.020 ;
        RECT 54.435 134.965 55.535 134.990 ;
        RECT 54.400 134.930 55.535 134.965 ;
        RECT 54.370 134.925 55.535 134.930 ;
        RECT 54.370 134.920 54.760 134.925 ;
        RECT 54.370 134.910 54.735 134.920 ;
        RECT 54.370 134.905 54.720 134.910 ;
        RECT 54.370 134.900 54.705 134.905 ;
        RECT 53.745 134.895 54.705 134.900 ;
        RECT 53.745 134.885 54.695 134.895 ;
        RECT 53.745 134.880 54.685 134.885 ;
        RECT 53.745 134.870 54.675 134.880 ;
        RECT 53.745 134.860 54.670 134.870 ;
        RECT 53.745 134.855 54.665 134.860 ;
        RECT 53.745 134.840 54.655 134.855 ;
        RECT 53.745 134.825 54.650 134.840 ;
        RECT 53.745 134.800 54.640 134.825 ;
        RECT 53.745 134.730 54.635 134.800 ;
        RECT 51.610 133.625 51.850 134.135 ;
        RECT 52.030 133.805 52.310 134.135 ;
        RECT 52.540 133.625 52.755 134.135 ;
        RECT 52.925 133.795 53.540 134.365 ;
        RECT 53.745 134.175 54.295 134.560 ;
        RECT 54.465 134.005 54.635 134.730 ;
        RECT 53.745 133.835 54.635 134.005 ;
        RECT 54.805 134.330 55.135 134.755 ;
        RECT 55.305 134.530 55.535 134.925 ;
        RECT 54.805 133.845 55.025 134.330 ;
        RECT 55.705 134.275 55.875 135.305 ;
        RECT 56.045 135.010 56.335 136.175 ;
        RECT 56.595 135.505 56.765 136.005 ;
        RECT 56.935 135.675 57.265 136.175 ;
        RECT 56.595 135.335 57.260 135.505 ;
        RECT 56.510 134.515 56.860 135.165 ;
        RECT 55.195 133.625 55.445 134.165 ;
        RECT 55.615 133.795 55.875 134.275 ;
        RECT 56.045 133.625 56.335 134.350 ;
        RECT 57.030 134.345 57.260 135.335 ;
        RECT 56.595 134.175 57.260 134.345 ;
        RECT 56.595 133.885 56.765 134.175 ;
        RECT 56.935 133.625 57.265 134.005 ;
        RECT 57.435 133.885 57.620 136.005 ;
        RECT 57.860 135.715 58.125 136.175 ;
        RECT 58.295 135.580 58.545 136.005 ;
        RECT 58.755 135.730 59.860 135.900 ;
        RECT 58.240 135.450 58.545 135.580 ;
        RECT 57.790 134.255 58.070 135.205 ;
        RECT 58.240 134.345 58.410 135.450 ;
        RECT 58.580 134.665 58.820 135.260 ;
        RECT 58.990 135.195 59.520 135.560 ;
        RECT 58.990 134.495 59.160 135.195 ;
        RECT 59.690 135.115 59.860 135.730 ;
        RECT 60.030 135.375 60.200 136.175 ;
        RECT 60.370 135.675 60.620 136.005 ;
        RECT 60.845 135.705 61.730 135.875 ;
        RECT 59.690 135.025 60.200 135.115 ;
        RECT 58.240 134.215 58.465 134.345 ;
        RECT 58.635 134.275 59.160 134.495 ;
        RECT 59.330 134.855 60.200 135.025 ;
        RECT 57.875 133.625 58.125 134.085 ;
        RECT 58.295 134.075 58.465 134.215 ;
        RECT 59.330 134.075 59.500 134.855 ;
        RECT 60.030 134.785 60.200 134.855 ;
        RECT 59.710 134.605 59.910 134.635 ;
        RECT 60.370 134.605 60.540 135.675 ;
        RECT 60.710 134.785 60.900 135.505 ;
        RECT 59.710 134.305 60.540 134.605 ;
        RECT 61.070 134.575 61.390 135.535 ;
        RECT 58.295 133.905 58.630 134.075 ;
        RECT 58.825 133.905 59.500 134.075 ;
        RECT 59.820 133.625 60.190 134.125 ;
        RECT 60.370 134.075 60.540 134.305 ;
        RECT 60.925 134.245 61.390 134.575 ;
        RECT 61.560 134.865 61.730 135.705 ;
        RECT 61.910 135.675 62.225 136.175 ;
        RECT 62.455 135.445 62.795 136.005 ;
        RECT 61.900 135.070 62.795 135.445 ;
        RECT 62.965 135.165 63.135 136.175 ;
        RECT 62.605 134.865 62.795 135.070 ;
        RECT 63.305 135.115 63.635 135.960 ;
        RECT 63.865 135.740 69.210 136.175 ;
        RECT 63.305 135.035 63.695 135.115 ;
        RECT 63.480 134.985 63.695 135.035 ;
        RECT 61.560 134.535 62.435 134.865 ;
        RECT 62.605 134.535 63.355 134.865 ;
        RECT 61.560 134.075 61.730 134.535 ;
        RECT 62.605 134.365 62.805 134.535 ;
        RECT 63.525 134.405 63.695 134.985 ;
        RECT 63.470 134.365 63.695 134.405 ;
        RECT 60.370 133.905 60.775 134.075 ;
        RECT 60.945 133.905 61.730 134.075 ;
        RECT 62.005 133.625 62.215 134.155 ;
        RECT 62.475 133.840 62.805 134.365 ;
        RECT 63.315 134.280 63.695 134.365 ;
        RECT 62.975 133.625 63.145 134.235 ;
        RECT 63.315 133.845 63.645 134.280 ;
        RECT 65.450 134.170 65.790 135.000 ;
        RECT 67.270 134.490 67.620 135.740 ;
        RECT 69.385 135.085 71.975 136.175 ;
        RECT 72.235 135.505 72.405 136.005 ;
        RECT 72.575 135.675 72.905 136.175 ;
        RECT 72.235 135.335 72.900 135.505 ;
        RECT 69.385 134.395 70.595 134.915 ;
        RECT 70.765 134.565 71.975 135.085 ;
        RECT 72.150 134.515 72.500 135.165 ;
        RECT 63.865 133.625 69.210 134.170 ;
        RECT 69.385 133.625 71.975 134.395 ;
        RECT 72.670 134.345 72.900 135.335 ;
        RECT 72.235 134.175 72.900 134.345 ;
        RECT 72.235 133.885 72.405 134.175 ;
        RECT 72.575 133.625 72.905 134.005 ;
        RECT 73.075 133.885 73.260 136.005 ;
        RECT 73.500 135.715 73.765 136.175 ;
        RECT 73.935 135.580 74.185 136.005 ;
        RECT 74.395 135.730 75.500 135.900 ;
        RECT 73.880 135.450 74.185 135.580 ;
        RECT 73.430 134.255 73.710 135.205 ;
        RECT 73.880 134.345 74.050 135.450 ;
        RECT 74.220 134.665 74.460 135.260 ;
        RECT 74.630 135.195 75.160 135.560 ;
        RECT 74.630 134.495 74.800 135.195 ;
        RECT 75.330 135.115 75.500 135.730 ;
        RECT 75.670 135.375 75.840 136.175 ;
        RECT 76.010 135.675 76.260 136.005 ;
        RECT 76.485 135.705 77.370 135.875 ;
        RECT 75.330 135.025 75.840 135.115 ;
        RECT 73.880 134.215 74.105 134.345 ;
        RECT 74.275 134.275 74.800 134.495 ;
        RECT 74.970 134.855 75.840 135.025 ;
        RECT 73.515 133.625 73.765 134.085 ;
        RECT 73.935 134.075 74.105 134.215 ;
        RECT 74.970 134.075 75.140 134.855 ;
        RECT 75.670 134.785 75.840 134.855 ;
        RECT 75.350 134.605 75.550 134.635 ;
        RECT 76.010 134.605 76.180 135.675 ;
        RECT 76.350 134.785 76.540 135.505 ;
        RECT 75.350 134.305 76.180 134.605 ;
        RECT 76.710 134.575 77.030 135.535 ;
        RECT 73.935 133.905 74.270 134.075 ;
        RECT 74.465 133.905 75.140 134.075 ;
        RECT 75.460 133.625 75.830 134.125 ;
        RECT 76.010 134.075 76.180 134.305 ;
        RECT 76.565 134.245 77.030 134.575 ;
        RECT 77.200 134.865 77.370 135.705 ;
        RECT 77.550 135.675 77.865 136.175 ;
        RECT 78.095 135.445 78.435 136.005 ;
        RECT 77.540 135.070 78.435 135.445 ;
        RECT 78.605 135.165 78.775 136.175 ;
        RECT 78.245 134.865 78.435 135.070 ;
        RECT 78.945 135.115 79.275 135.960 ;
        RECT 78.945 135.035 79.335 135.115 ;
        RECT 79.510 135.035 79.830 136.175 ;
        RECT 79.120 134.985 79.335 135.035 ;
        RECT 77.200 134.535 78.075 134.865 ;
        RECT 78.245 134.535 78.995 134.865 ;
        RECT 77.200 134.075 77.370 134.535 ;
        RECT 78.245 134.365 78.445 134.535 ;
        RECT 79.165 134.405 79.335 134.985 ;
        RECT 80.010 134.865 80.205 135.915 ;
        RECT 80.385 135.325 80.715 136.005 ;
        RECT 80.915 135.375 81.170 136.175 ;
        RECT 80.385 135.045 80.735 135.325 ;
        RECT 79.570 134.815 79.830 134.865 ;
        RECT 79.565 134.645 79.830 134.815 ;
        RECT 79.570 134.535 79.830 134.645 ;
        RECT 80.010 134.535 80.395 134.865 ;
        RECT 80.565 134.665 80.735 135.045 ;
        RECT 80.925 134.835 81.170 135.195 ;
        RECT 81.805 135.010 82.095 136.175 ;
        RECT 82.265 135.035 82.650 136.005 ;
        RECT 82.820 135.715 83.145 136.175 ;
        RECT 83.665 135.545 83.945 136.005 ;
        RECT 82.820 135.325 83.945 135.545 ;
        RECT 80.565 134.495 81.085 134.665 ;
        RECT 79.110 134.365 79.335 134.405 ;
        RECT 76.010 133.905 76.415 134.075 ;
        RECT 76.585 133.905 77.370 134.075 ;
        RECT 77.645 133.625 77.855 134.155 ;
        RECT 78.115 133.840 78.445 134.365 ;
        RECT 78.955 134.280 79.335 134.365 ;
        RECT 78.615 133.625 78.785 134.235 ;
        RECT 78.955 133.845 79.285 134.280 ;
        RECT 79.510 134.155 80.725 134.325 ;
        RECT 79.510 133.805 79.800 134.155 ;
        RECT 79.995 133.625 80.325 133.985 ;
        RECT 80.495 133.850 80.725 134.155 ;
        RECT 80.915 133.930 81.085 134.495 ;
        RECT 82.265 134.365 82.545 135.035 ;
        RECT 82.820 134.865 83.270 135.325 ;
        RECT 84.135 135.155 84.535 136.005 ;
        RECT 84.935 135.715 85.205 136.175 ;
        RECT 85.375 135.545 85.660 136.005 ;
        RECT 82.715 134.535 83.270 134.865 ;
        RECT 83.440 134.595 84.535 135.155 ;
        RECT 82.820 134.425 83.270 134.535 ;
        RECT 81.805 133.625 82.095 134.350 ;
        RECT 82.265 133.795 82.650 134.365 ;
        RECT 82.820 134.255 83.945 134.425 ;
        RECT 82.820 133.625 83.145 134.085 ;
        RECT 83.665 133.795 83.945 134.255 ;
        RECT 84.135 133.795 84.535 134.595 ;
        RECT 84.705 135.325 85.660 135.545 ;
        RECT 84.705 134.425 84.915 135.325 ;
        RECT 85.085 134.595 85.775 135.155 ;
        RECT 85.945 135.035 86.225 136.175 ;
        RECT 86.395 135.025 86.725 136.005 ;
        RECT 86.895 135.035 87.155 136.175 ;
        RECT 88.335 135.505 88.505 136.005 ;
        RECT 88.675 135.675 89.005 136.175 ;
        RECT 88.335 135.335 89.000 135.505 ;
        RECT 85.955 134.595 86.290 134.865 ;
        RECT 86.460 134.475 86.630 135.025 ;
        RECT 86.800 134.615 87.135 134.865 ;
        RECT 88.250 134.515 88.600 135.165 ;
        RECT 86.460 134.425 86.635 134.475 ;
        RECT 84.705 134.255 85.660 134.425 ;
        RECT 84.935 133.625 85.205 134.085 ;
        RECT 85.375 133.795 85.660 134.255 ;
        RECT 85.945 133.625 86.255 134.425 ;
        RECT 86.460 133.795 87.155 134.425 ;
        RECT 88.770 134.345 89.000 135.335 ;
        RECT 88.335 134.175 89.000 134.345 ;
        RECT 88.335 133.885 88.505 134.175 ;
        RECT 88.675 133.625 89.005 134.005 ;
        RECT 89.175 133.885 89.360 136.005 ;
        RECT 89.600 135.715 89.865 136.175 ;
        RECT 90.035 135.580 90.285 136.005 ;
        RECT 90.495 135.730 91.600 135.900 ;
        RECT 89.980 135.450 90.285 135.580 ;
        RECT 89.530 134.255 89.810 135.205 ;
        RECT 89.980 134.345 90.150 135.450 ;
        RECT 90.320 134.665 90.560 135.260 ;
        RECT 90.730 135.195 91.260 135.560 ;
        RECT 90.730 134.495 90.900 135.195 ;
        RECT 91.430 135.115 91.600 135.730 ;
        RECT 91.770 135.375 91.940 136.175 ;
        RECT 92.110 135.675 92.360 136.005 ;
        RECT 92.585 135.705 93.470 135.875 ;
        RECT 91.430 135.025 91.940 135.115 ;
        RECT 89.980 134.215 90.205 134.345 ;
        RECT 90.375 134.275 90.900 134.495 ;
        RECT 91.070 134.855 91.940 135.025 ;
        RECT 89.615 133.625 89.865 134.085 ;
        RECT 90.035 134.075 90.205 134.215 ;
        RECT 91.070 134.075 91.240 134.855 ;
        RECT 91.770 134.785 91.940 134.855 ;
        RECT 91.450 134.605 91.650 134.635 ;
        RECT 92.110 134.605 92.280 135.675 ;
        RECT 92.450 134.785 92.640 135.505 ;
        RECT 91.450 134.305 92.280 134.605 ;
        RECT 92.810 134.575 93.130 135.535 ;
        RECT 90.035 133.905 90.370 134.075 ;
        RECT 90.565 133.905 91.240 134.075 ;
        RECT 91.560 133.625 91.930 134.125 ;
        RECT 92.110 134.075 92.280 134.305 ;
        RECT 92.665 134.245 93.130 134.575 ;
        RECT 93.300 134.865 93.470 135.705 ;
        RECT 93.650 135.675 93.965 136.175 ;
        RECT 94.195 135.445 94.535 136.005 ;
        RECT 93.640 135.070 94.535 135.445 ;
        RECT 94.705 135.165 94.875 136.175 ;
        RECT 94.345 134.865 94.535 135.070 ;
        RECT 95.045 135.115 95.375 135.960 ;
        RECT 95.045 135.035 95.435 135.115 ;
        RECT 95.605 135.085 96.815 136.175 ;
        RECT 95.220 134.985 95.435 135.035 ;
        RECT 93.300 134.535 94.175 134.865 ;
        RECT 94.345 134.535 95.095 134.865 ;
        RECT 93.300 134.075 93.470 134.535 ;
        RECT 94.345 134.365 94.545 134.535 ;
        RECT 95.265 134.405 95.435 134.985 ;
        RECT 95.210 134.365 95.435 134.405 ;
        RECT 92.110 133.905 92.515 134.075 ;
        RECT 92.685 133.905 93.470 134.075 ;
        RECT 93.745 133.625 93.955 134.155 ;
        RECT 94.215 133.840 94.545 134.365 ;
        RECT 95.055 134.280 95.435 134.365 ;
        RECT 95.605 134.375 96.125 134.915 ;
        RECT 96.295 134.545 96.815 135.085 ;
        RECT 96.990 135.225 97.255 135.995 ;
        RECT 97.425 135.455 97.755 136.175 ;
        RECT 97.945 135.635 98.205 135.995 ;
        RECT 98.375 135.805 98.705 136.175 ;
        RECT 98.875 135.635 99.135 135.995 ;
        RECT 97.945 135.405 99.135 135.635 ;
        RECT 99.705 135.225 99.995 135.995 ;
        RECT 94.715 133.625 94.885 134.235 ;
        RECT 95.055 133.845 95.385 134.280 ;
        RECT 95.605 133.625 96.815 134.375 ;
        RECT 96.990 133.805 97.325 135.225 ;
        RECT 97.500 135.045 99.995 135.225 ;
        RECT 100.205 135.085 102.795 136.175 ;
        RECT 97.500 134.355 97.725 135.045 ;
        RECT 97.925 134.535 98.205 134.865 ;
        RECT 98.385 134.535 98.960 134.865 ;
        RECT 99.140 134.535 99.575 134.865 ;
        RECT 99.755 134.535 100.025 134.865 ;
        RECT 100.205 134.395 101.415 134.915 ;
        RECT 101.585 134.565 102.795 135.085 ;
        RECT 103.430 135.035 103.765 136.005 ;
        RECT 103.935 135.035 104.105 136.175 ;
        RECT 104.275 135.835 106.305 136.005 ;
        RECT 97.500 134.165 99.985 134.355 ;
        RECT 97.505 133.625 98.250 133.995 ;
        RECT 98.815 133.805 99.070 134.165 ;
        RECT 99.250 133.625 99.580 133.995 ;
        RECT 99.760 133.805 99.985 134.165 ;
        RECT 100.205 133.625 102.795 134.395 ;
        RECT 103.430 134.365 103.600 135.035 ;
        RECT 104.275 134.865 104.445 135.835 ;
        RECT 103.770 134.535 104.025 134.865 ;
        RECT 104.250 134.535 104.445 134.865 ;
        RECT 104.615 135.495 105.740 135.665 ;
        RECT 103.855 134.365 104.025 134.535 ;
        RECT 104.615 134.365 104.785 135.495 ;
        RECT 103.430 133.795 103.685 134.365 ;
        RECT 103.855 134.195 104.785 134.365 ;
        RECT 104.955 135.155 105.965 135.325 ;
        RECT 104.955 134.355 105.125 135.155 ;
        RECT 105.330 134.815 105.605 134.955 ;
        RECT 105.325 134.645 105.605 134.815 ;
        RECT 104.610 134.160 104.785 134.195 ;
        RECT 103.855 133.625 104.185 134.025 ;
        RECT 104.610 133.795 105.140 134.160 ;
        RECT 105.330 133.795 105.605 134.645 ;
        RECT 105.775 133.795 105.965 135.155 ;
        RECT 106.135 135.170 106.305 135.835 ;
        RECT 106.475 135.415 106.645 136.175 ;
        RECT 106.880 135.415 107.395 135.825 ;
        RECT 106.135 134.980 106.885 135.170 ;
        RECT 107.055 134.605 107.395 135.415 ;
        RECT 107.565 135.010 107.855 136.175 ;
        RECT 108.030 135.035 108.365 136.005 ;
        RECT 108.535 135.035 108.705 136.175 ;
        RECT 108.875 135.835 110.905 136.005 ;
        RECT 106.165 134.435 107.395 134.605 ;
        RECT 106.145 133.625 106.655 134.160 ;
        RECT 106.875 133.830 107.120 134.435 ;
        RECT 108.030 134.365 108.200 135.035 ;
        RECT 108.875 134.865 109.045 135.835 ;
        RECT 108.370 134.535 108.625 134.865 ;
        RECT 108.850 134.535 109.045 134.865 ;
        RECT 109.215 135.495 110.340 135.665 ;
        RECT 108.455 134.365 108.625 134.535 ;
        RECT 109.215 134.365 109.385 135.495 ;
        RECT 107.565 133.625 107.855 134.350 ;
        RECT 108.030 133.795 108.285 134.365 ;
        RECT 108.455 134.195 109.385 134.365 ;
        RECT 109.555 135.155 110.565 135.325 ;
        RECT 109.555 134.355 109.725 135.155 ;
        RECT 109.210 134.160 109.385 134.195 ;
        RECT 108.455 133.625 108.785 134.025 ;
        RECT 109.210 133.795 109.740 134.160 ;
        RECT 109.930 134.135 110.205 134.955 ;
        RECT 109.925 133.965 110.205 134.135 ;
        RECT 109.930 133.795 110.205 133.965 ;
        RECT 110.375 133.795 110.565 135.155 ;
        RECT 110.735 135.170 110.905 135.835 ;
        RECT 111.075 135.415 111.245 136.175 ;
        RECT 111.480 135.415 111.995 135.825 ;
        RECT 112.165 135.740 117.510 136.175 ;
        RECT 110.735 134.980 111.485 135.170 ;
        RECT 111.655 134.605 111.995 135.415 ;
        RECT 110.765 134.435 111.995 134.605 ;
        RECT 110.745 133.625 111.255 134.160 ;
        RECT 111.475 133.830 111.720 134.435 ;
        RECT 113.750 134.170 114.090 135.000 ;
        RECT 115.570 134.490 115.920 135.740 ;
        RECT 118.665 135.115 118.995 135.960 ;
        RECT 119.165 135.165 119.335 136.175 ;
        RECT 119.505 135.445 119.845 136.005 ;
        RECT 120.075 135.675 120.390 136.175 ;
        RECT 120.570 135.705 121.455 135.875 ;
        RECT 118.605 135.035 118.995 135.115 ;
        RECT 119.505 135.070 120.400 135.445 ;
        RECT 118.605 134.985 118.820 135.035 ;
        RECT 118.605 134.405 118.775 134.985 ;
        RECT 119.505 134.865 119.695 135.070 ;
        RECT 120.570 134.865 120.740 135.705 ;
        RECT 121.680 135.675 121.930 136.005 ;
        RECT 118.945 134.535 119.695 134.865 ;
        RECT 119.865 134.535 120.740 134.865 ;
        RECT 118.605 134.365 118.830 134.405 ;
        RECT 119.495 134.365 119.695 134.535 ;
        RECT 118.605 134.280 118.985 134.365 ;
        RECT 112.165 133.625 117.510 134.170 ;
        RECT 118.655 133.845 118.985 134.280 ;
        RECT 119.155 133.625 119.325 134.235 ;
        RECT 119.495 133.840 119.825 134.365 ;
        RECT 120.085 133.625 120.295 134.155 ;
        RECT 120.570 134.075 120.740 134.535 ;
        RECT 120.910 134.575 121.230 135.535 ;
        RECT 121.400 134.785 121.590 135.505 ;
        RECT 121.760 134.605 121.930 135.675 ;
        RECT 122.100 135.375 122.270 136.175 ;
        RECT 122.440 135.730 123.545 135.900 ;
        RECT 122.440 135.115 122.610 135.730 ;
        RECT 123.755 135.580 124.005 136.005 ;
        RECT 124.175 135.715 124.440 136.175 ;
        RECT 122.780 135.195 123.310 135.560 ;
        RECT 123.755 135.450 124.060 135.580 ;
        RECT 122.100 135.025 122.610 135.115 ;
        RECT 122.100 134.855 122.970 135.025 ;
        RECT 122.100 134.785 122.270 134.855 ;
        RECT 122.390 134.605 122.590 134.635 ;
        RECT 120.910 134.245 121.375 134.575 ;
        RECT 121.760 134.305 122.590 134.605 ;
        RECT 121.760 134.075 121.930 134.305 ;
        RECT 120.570 133.905 121.355 134.075 ;
        RECT 121.525 133.905 121.930 134.075 ;
        RECT 122.110 133.625 122.480 134.125 ;
        RECT 122.800 134.075 122.970 134.855 ;
        RECT 123.140 134.495 123.310 135.195 ;
        RECT 123.480 134.665 123.720 135.260 ;
        RECT 123.140 134.275 123.665 134.495 ;
        RECT 123.890 134.345 124.060 135.450 ;
        RECT 123.835 134.215 124.060 134.345 ;
        RECT 124.230 134.255 124.510 135.205 ;
        RECT 123.835 134.075 124.005 134.215 ;
        RECT 122.800 133.905 123.475 134.075 ;
        RECT 123.670 133.905 124.005 134.075 ;
        RECT 124.175 133.625 124.425 134.085 ;
        RECT 124.680 133.885 124.865 136.005 ;
        RECT 125.035 135.675 125.365 136.175 ;
        RECT 125.535 135.505 125.705 136.005 ;
        RECT 125.040 135.335 125.705 135.505 ;
        RECT 126.080 135.545 126.365 136.005 ;
        RECT 126.535 135.715 126.805 136.175 ;
        RECT 125.040 134.345 125.270 135.335 ;
        RECT 126.080 135.325 127.035 135.545 ;
        RECT 125.440 134.515 125.790 135.165 ;
        RECT 125.965 134.595 126.655 135.155 ;
        RECT 126.825 134.425 127.035 135.325 ;
        RECT 125.040 134.175 125.705 134.345 ;
        RECT 125.035 133.625 125.365 134.005 ;
        RECT 125.535 133.885 125.705 134.175 ;
        RECT 126.080 134.255 127.035 134.425 ;
        RECT 127.205 135.155 127.605 136.005 ;
        RECT 127.795 135.545 128.075 136.005 ;
        RECT 128.595 135.715 128.920 136.175 ;
        RECT 127.795 135.325 128.920 135.545 ;
        RECT 127.205 134.595 128.300 135.155 ;
        RECT 128.470 134.865 128.920 135.325 ;
        RECT 129.090 135.035 129.475 136.005 ;
        RECT 129.645 135.085 133.155 136.175 ;
        RECT 126.080 133.795 126.365 134.255 ;
        RECT 126.535 133.625 126.805 134.085 ;
        RECT 127.205 133.795 127.605 134.595 ;
        RECT 128.470 134.535 129.025 134.865 ;
        RECT 128.470 134.425 128.920 134.535 ;
        RECT 127.795 134.255 128.920 134.425 ;
        RECT 129.195 134.365 129.475 135.035 ;
        RECT 127.795 133.795 128.075 134.255 ;
        RECT 128.595 133.625 128.920 134.085 ;
        RECT 129.090 133.795 129.475 134.365 ;
        RECT 129.645 134.395 131.295 134.915 ;
        RECT 131.465 134.565 133.155 135.085 ;
        RECT 133.325 135.010 133.615 136.175 ;
        RECT 133.875 135.505 134.045 136.005 ;
        RECT 134.215 135.675 134.545 136.175 ;
        RECT 133.875 135.335 134.540 135.505 ;
        RECT 133.790 134.515 134.140 135.165 ;
        RECT 129.645 133.625 133.155 134.395 ;
        RECT 133.325 133.625 133.615 134.350 ;
        RECT 134.310 134.345 134.540 135.335 ;
        RECT 133.875 134.175 134.540 134.345 ;
        RECT 133.875 133.885 134.045 134.175 ;
        RECT 134.215 133.625 134.545 134.005 ;
        RECT 134.715 133.885 134.900 136.005 ;
        RECT 135.140 135.715 135.405 136.175 ;
        RECT 135.575 135.580 135.825 136.005 ;
        RECT 136.035 135.730 137.140 135.900 ;
        RECT 135.520 135.450 135.825 135.580 ;
        RECT 135.070 134.255 135.350 135.205 ;
        RECT 135.520 134.345 135.690 135.450 ;
        RECT 135.860 134.665 136.100 135.260 ;
        RECT 136.270 135.195 136.800 135.560 ;
        RECT 136.270 134.495 136.440 135.195 ;
        RECT 136.970 135.115 137.140 135.730 ;
        RECT 137.310 135.375 137.480 136.175 ;
        RECT 137.650 135.675 137.900 136.005 ;
        RECT 138.125 135.705 139.010 135.875 ;
        RECT 136.970 135.025 137.480 135.115 ;
        RECT 135.520 134.215 135.745 134.345 ;
        RECT 135.915 134.275 136.440 134.495 ;
        RECT 136.610 134.855 137.480 135.025 ;
        RECT 135.155 133.625 135.405 134.085 ;
        RECT 135.575 134.075 135.745 134.215 ;
        RECT 136.610 134.075 136.780 134.855 ;
        RECT 137.310 134.785 137.480 134.855 ;
        RECT 136.990 134.605 137.190 134.635 ;
        RECT 137.650 134.605 137.820 135.675 ;
        RECT 137.990 134.785 138.180 135.505 ;
        RECT 136.990 134.305 137.820 134.605 ;
        RECT 138.350 134.575 138.670 135.535 ;
        RECT 135.575 133.905 135.910 134.075 ;
        RECT 136.105 133.905 136.780 134.075 ;
        RECT 137.100 133.625 137.470 134.125 ;
        RECT 137.650 134.075 137.820 134.305 ;
        RECT 138.205 134.245 138.670 134.575 ;
        RECT 138.840 134.865 139.010 135.705 ;
        RECT 139.190 135.675 139.505 136.175 ;
        RECT 139.735 135.445 140.075 136.005 ;
        RECT 139.180 135.070 140.075 135.445 ;
        RECT 140.245 135.165 140.415 136.175 ;
        RECT 139.885 134.865 140.075 135.070 ;
        RECT 140.585 135.115 140.915 135.960 ;
        RECT 140.585 135.035 140.975 135.115 ;
        RECT 140.760 134.985 140.975 135.035 ;
        RECT 138.840 134.535 139.715 134.865 ;
        RECT 139.885 134.535 140.635 134.865 ;
        RECT 138.840 134.075 139.010 134.535 ;
        RECT 139.885 134.365 140.085 134.535 ;
        RECT 140.805 134.405 140.975 134.985 ;
        RECT 140.750 134.365 140.975 134.405 ;
        RECT 137.650 133.905 138.055 134.075 ;
        RECT 138.225 133.905 139.010 134.075 ;
        RECT 139.285 133.625 139.495 134.155 ;
        RECT 139.755 133.840 140.085 134.365 ;
        RECT 140.595 134.280 140.975 134.365 ;
        RECT 141.145 135.035 141.530 136.005 ;
        RECT 141.700 135.715 142.025 136.175 ;
        RECT 142.545 135.545 142.825 136.005 ;
        RECT 141.700 135.325 142.825 135.545 ;
        RECT 141.145 134.365 141.425 135.035 ;
        RECT 141.700 134.865 142.150 135.325 ;
        RECT 143.015 135.155 143.415 136.005 ;
        RECT 143.815 135.715 144.085 136.175 ;
        RECT 144.255 135.545 144.540 136.005 ;
        RECT 141.595 134.535 142.150 134.865 ;
        RECT 142.320 134.595 143.415 135.155 ;
        RECT 141.700 134.425 142.150 134.535 ;
        RECT 140.255 133.625 140.425 134.235 ;
        RECT 140.595 133.845 140.925 134.280 ;
        RECT 141.145 133.795 141.530 134.365 ;
        RECT 141.700 134.255 142.825 134.425 ;
        RECT 141.700 133.625 142.025 134.085 ;
        RECT 142.545 133.795 142.825 134.255 ;
        RECT 143.015 133.795 143.415 134.595 ;
        RECT 143.585 135.325 144.540 135.545 ;
        RECT 143.585 134.425 143.795 135.325 ;
        RECT 143.965 134.595 144.655 135.155 ;
        RECT 145.745 135.085 146.955 136.175 ;
        RECT 145.745 134.545 146.265 135.085 ;
        RECT 143.585 134.255 144.540 134.425 ;
        RECT 146.435 134.375 146.955 134.915 ;
        RECT 143.815 133.625 144.085 134.085 ;
        RECT 144.255 133.795 144.540 134.255 ;
        RECT 145.745 133.625 146.955 134.375 ;
        RECT 17.320 133.455 147.040 133.625 ;
        RECT 17.405 132.705 18.615 133.455 ;
        RECT 19.335 132.905 19.505 133.195 ;
        RECT 19.675 133.075 20.005 133.455 ;
        RECT 19.335 132.735 20.000 132.905 ;
        RECT 17.405 132.165 17.925 132.705 ;
        RECT 18.095 131.995 18.615 132.535 ;
        RECT 17.405 130.905 18.615 131.995 ;
        RECT 19.250 131.915 19.600 132.565 ;
        RECT 19.770 131.745 20.000 132.735 ;
        RECT 19.335 131.575 20.000 131.745 ;
        RECT 19.335 131.075 19.505 131.575 ;
        RECT 19.675 130.905 20.005 131.405 ;
        RECT 20.175 131.075 20.360 133.195 ;
        RECT 20.615 132.995 20.865 133.455 ;
        RECT 21.035 133.005 21.370 133.175 ;
        RECT 21.565 133.005 22.240 133.175 ;
        RECT 21.035 132.865 21.205 133.005 ;
        RECT 20.530 131.875 20.810 132.825 ;
        RECT 20.980 132.735 21.205 132.865 ;
        RECT 20.980 131.630 21.150 132.735 ;
        RECT 21.375 132.585 21.900 132.805 ;
        RECT 21.320 131.820 21.560 132.415 ;
        RECT 21.730 131.885 21.900 132.585 ;
        RECT 22.070 132.225 22.240 133.005 ;
        RECT 22.560 132.955 22.930 133.455 ;
        RECT 23.110 133.005 23.515 133.175 ;
        RECT 23.685 133.005 24.470 133.175 ;
        RECT 23.110 132.775 23.280 133.005 ;
        RECT 22.450 132.475 23.280 132.775 ;
        RECT 23.665 132.505 24.130 132.835 ;
        RECT 22.450 132.445 22.650 132.475 ;
        RECT 22.770 132.225 22.940 132.295 ;
        RECT 22.070 132.055 22.940 132.225 ;
        RECT 22.430 131.965 22.940 132.055 ;
        RECT 20.980 131.500 21.285 131.630 ;
        RECT 21.730 131.520 22.260 131.885 ;
        RECT 20.600 130.905 20.865 131.365 ;
        RECT 21.035 131.075 21.285 131.500 ;
        RECT 22.430 131.350 22.600 131.965 ;
        RECT 21.495 131.180 22.600 131.350 ;
        RECT 22.770 130.905 22.940 131.705 ;
        RECT 23.110 131.405 23.280 132.475 ;
        RECT 23.450 131.575 23.640 132.295 ;
        RECT 23.810 131.545 24.130 132.505 ;
        RECT 24.300 132.545 24.470 133.005 ;
        RECT 24.745 132.925 24.955 133.455 ;
        RECT 25.215 132.715 25.545 133.240 ;
        RECT 25.715 132.845 25.885 133.455 ;
        RECT 26.055 132.800 26.385 133.235 ;
        RECT 27.690 132.945 27.930 133.455 ;
        RECT 28.110 132.945 28.390 133.275 ;
        RECT 28.620 132.945 28.835 133.455 ;
        RECT 26.055 132.715 26.435 132.800 ;
        RECT 25.345 132.545 25.545 132.715 ;
        RECT 26.210 132.675 26.435 132.715 ;
        RECT 24.300 132.215 25.175 132.545 ;
        RECT 25.345 132.215 26.095 132.545 ;
        RECT 23.110 131.075 23.360 131.405 ;
        RECT 24.300 131.375 24.470 132.215 ;
        RECT 25.345 132.010 25.535 132.215 ;
        RECT 26.265 132.095 26.435 132.675 ;
        RECT 27.585 132.215 27.940 132.775 ;
        RECT 26.220 132.045 26.435 132.095 ;
        RECT 28.110 132.045 28.280 132.945 ;
        RECT 28.450 132.215 28.715 132.775 ;
        RECT 29.005 132.715 29.620 133.285 ;
        RECT 29.825 132.910 35.170 133.455 ;
        RECT 28.965 132.045 29.135 132.545 ;
        RECT 24.640 131.635 25.535 132.010 ;
        RECT 26.045 131.965 26.435 132.045 ;
        RECT 23.585 131.205 24.470 131.375 ;
        RECT 24.650 130.905 24.965 131.405 ;
        RECT 25.195 131.075 25.535 131.635 ;
        RECT 25.705 130.905 25.875 131.915 ;
        RECT 26.045 131.120 26.375 131.965 ;
        RECT 27.710 131.875 29.135 132.045 ;
        RECT 27.710 131.700 28.100 131.875 ;
        RECT 28.585 130.905 28.915 131.705 ;
        RECT 29.305 131.695 29.620 132.715 ;
        RECT 31.410 132.080 31.750 132.910 ;
        RECT 35.895 132.905 36.065 133.195 ;
        RECT 36.235 133.075 36.565 133.455 ;
        RECT 35.895 132.735 36.560 132.905 ;
        RECT 29.085 131.075 29.620 131.695 ;
        RECT 33.230 131.340 33.580 132.590 ;
        RECT 35.810 131.915 36.160 132.565 ;
        RECT 36.330 131.745 36.560 132.735 ;
        RECT 35.895 131.575 36.560 131.745 ;
        RECT 29.825 130.905 35.170 131.340 ;
        RECT 35.895 131.075 36.065 131.575 ;
        RECT 36.235 130.905 36.565 131.405 ;
        RECT 36.735 131.075 36.920 133.195 ;
        RECT 37.175 132.995 37.425 133.455 ;
        RECT 37.595 133.005 37.930 133.175 ;
        RECT 38.125 133.005 38.800 133.175 ;
        RECT 37.595 132.865 37.765 133.005 ;
        RECT 37.090 131.875 37.370 132.825 ;
        RECT 37.540 132.735 37.765 132.865 ;
        RECT 37.540 131.630 37.710 132.735 ;
        RECT 37.935 132.585 38.460 132.805 ;
        RECT 37.880 131.820 38.120 132.415 ;
        RECT 38.290 131.885 38.460 132.585 ;
        RECT 38.630 132.225 38.800 133.005 ;
        RECT 39.120 132.955 39.490 133.455 ;
        RECT 39.670 133.005 40.075 133.175 ;
        RECT 40.245 133.005 41.030 133.175 ;
        RECT 39.670 132.775 39.840 133.005 ;
        RECT 39.010 132.475 39.840 132.775 ;
        RECT 40.225 132.505 40.690 132.835 ;
        RECT 39.010 132.445 39.210 132.475 ;
        RECT 39.330 132.225 39.500 132.295 ;
        RECT 38.630 132.055 39.500 132.225 ;
        RECT 38.990 131.965 39.500 132.055 ;
        RECT 37.540 131.500 37.845 131.630 ;
        RECT 38.290 131.520 38.820 131.885 ;
        RECT 37.160 130.905 37.425 131.365 ;
        RECT 37.595 131.075 37.845 131.500 ;
        RECT 38.990 131.350 39.160 131.965 ;
        RECT 38.055 131.180 39.160 131.350 ;
        RECT 39.330 130.905 39.500 131.705 ;
        RECT 39.670 131.405 39.840 132.475 ;
        RECT 40.010 131.575 40.200 132.295 ;
        RECT 40.370 131.545 40.690 132.505 ;
        RECT 40.860 132.545 41.030 133.005 ;
        RECT 41.305 132.925 41.515 133.455 ;
        RECT 41.775 132.715 42.105 133.240 ;
        RECT 42.275 132.845 42.445 133.455 ;
        RECT 42.615 132.800 42.945 133.235 ;
        RECT 42.615 132.715 42.995 132.800 ;
        RECT 43.165 132.730 43.455 133.455 ;
        RECT 41.905 132.545 42.105 132.715 ;
        RECT 42.770 132.675 42.995 132.715 ;
        RECT 40.860 132.215 41.735 132.545 ;
        RECT 41.905 132.215 42.655 132.545 ;
        RECT 39.670 131.075 39.920 131.405 ;
        RECT 40.860 131.375 41.030 132.215 ;
        RECT 41.905 132.010 42.095 132.215 ;
        RECT 42.825 132.095 42.995 132.675 ;
        RECT 43.625 132.655 44.320 133.285 ;
        RECT 44.525 132.655 44.835 133.455 ;
        RECT 45.005 132.910 50.350 133.455 ;
        RECT 43.645 132.215 43.980 132.465 ;
        RECT 42.780 132.045 42.995 132.095 ;
        RECT 41.200 131.635 42.095 132.010 ;
        RECT 42.605 131.965 42.995 132.045 ;
        RECT 40.145 131.205 41.030 131.375 ;
        RECT 41.210 130.905 41.525 131.405 ;
        RECT 41.755 131.075 42.095 131.635 ;
        RECT 42.265 130.905 42.435 131.915 ;
        RECT 42.605 131.120 42.935 131.965 ;
        RECT 43.165 130.905 43.455 132.070 ;
        RECT 44.150 132.055 44.320 132.655 ;
        RECT 44.490 132.215 44.825 132.485 ;
        RECT 46.590 132.080 46.930 132.910 ;
        RECT 51.495 132.800 51.825 133.235 ;
        RECT 51.995 132.845 52.165 133.455 ;
        RECT 51.445 132.715 51.825 132.800 ;
        RECT 52.335 132.715 52.665 133.240 ;
        RECT 52.925 132.925 53.135 133.455 ;
        RECT 53.410 133.005 54.195 133.175 ;
        RECT 54.365 133.005 54.770 133.175 ;
        RECT 51.445 132.675 51.670 132.715 ;
        RECT 43.625 130.905 43.885 132.045 ;
        RECT 44.055 131.075 44.385 132.055 ;
        RECT 44.555 130.905 44.835 132.045 ;
        RECT 48.410 131.340 48.760 132.590 ;
        RECT 51.445 132.095 51.615 132.675 ;
        RECT 52.335 132.545 52.535 132.715 ;
        RECT 53.410 132.545 53.580 133.005 ;
        RECT 51.785 132.215 52.535 132.545 ;
        RECT 52.705 132.215 53.580 132.545 ;
        RECT 51.445 132.045 51.660 132.095 ;
        RECT 51.445 131.965 51.835 132.045 ;
        RECT 45.005 130.905 50.350 131.340 ;
        RECT 51.505 131.120 51.835 131.965 ;
        RECT 52.345 132.010 52.535 132.215 ;
        RECT 52.005 130.905 52.175 131.915 ;
        RECT 52.345 131.635 53.240 132.010 ;
        RECT 52.345 131.075 52.685 131.635 ;
        RECT 52.915 130.905 53.230 131.405 ;
        RECT 53.410 131.375 53.580 132.215 ;
        RECT 53.750 132.505 54.215 132.835 ;
        RECT 54.600 132.775 54.770 133.005 ;
        RECT 54.950 132.955 55.320 133.455 ;
        RECT 55.640 133.005 56.315 133.175 ;
        RECT 56.510 133.005 56.845 133.175 ;
        RECT 53.750 131.545 54.070 132.505 ;
        RECT 54.600 132.475 55.430 132.775 ;
        RECT 54.240 131.575 54.430 132.295 ;
        RECT 54.600 131.405 54.770 132.475 ;
        RECT 55.230 132.445 55.430 132.475 ;
        RECT 54.940 132.225 55.110 132.295 ;
        RECT 55.640 132.225 55.810 133.005 ;
        RECT 56.675 132.865 56.845 133.005 ;
        RECT 57.015 132.995 57.265 133.455 ;
        RECT 54.940 132.055 55.810 132.225 ;
        RECT 55.980 132.585 56.505 132.805 ;
        RECT 56.675 132.735 56.900 132.865 ;
        RECT 54.940 131.965 55.450 132.055 ;
        RECT 53.410 131.205 54.295 131.375 ;
        RECT 54.520 131.075 54.770 131.405 ;
        RECT 54.940 130.905 55.110 131.705 ;
        RECT 55.280 131.350 55.450 131.965 ;
        RECT 55.980 131.885 56.150 132.585 ;
        RECT 55.620 131.520 56.150 131.885 ;
        RECT 56.320 131.820 56.560 132.415 ;
        RECT 56.730 131.630 56.900 132.735 ;
        RECT 57.070 131.875 57.350 132.825 ;
        RECT 56.595 131.500 56.900 131.630 ;
        RECT 55.280 131.180 56.385 131.350 ;
        RECT 56.595 131.075 56.845 131.500 ;
        RECT 57.015 130.905 57.280 131.365 ;
        RECT 57.520 131.075 57.705 133.195 ;
        RECT 57.875 133.075 58.205 133.455 ;
        RECT 58.375 132.905 58.545 133.195 ;
        RECT 58.805 132.910 64.150 133.455 ;
        RECT 57.880 132.735 58.545 132.905 ;
        RECT 57.880 131.745 58.110 132.735 ;
        RECT 58.280 131.915 58.630 132.565 ;
        RECT 60.390 132.080 60.730 132.910 ;
        RECT 64.325 132.705 65.535 133.455 ;
        RECT 65.750 132.995 66.015 133.455 ;
        RECT 66.385 132.815 66.555 133.285 ;
        RECT 66.805 132.995 66.975 133.455 ;
        RECT 67.225 132.815 67.395 133.285 ;
        RECT 67.645 132.995 67.815 133.455 ;
        RECT 68.065 132.815 68.235 133.285 ;
        RECT 68.405 132.990 68.655 133.455 ;
        RECT 57.880 131.575 58.545 131.745 ;
        RECT 57.875 130.905 58.205 131.405 ;
        RECT 58.375 131.075 58.545 131.575 ;
        RECT 62.210 131.340 62.560 132.590 ;
        RECT 64.325 132.165 64.845 132.705 ;
        RECT 66.385 132.635 68.755 132.815 ;
        RECT 68.925 132.730 69.215 133.455 ;
        RECT 69.445 132.995 69.690 133.455 ;
        RECT 65.015 131.995 65.535 132.535 ;
        RECT 65.725 132.215 68.235 132.465 ;
        RECT 68.405 132.045 68.755 132.635 ;
        RECT 69.385 132.215 69.700 132.825 ;
        RECT 69.870 132.465 70.120 133.275 ;
        RECT 70.290 132.930 70.550 133.455 ;
        RECT 70.720 132.805 70.980 133.260 ;
        RECT 71.150 132.975 71.410 133.455 ;
        RECT 71.580 132.805 71.840 133.260 ;
        RECT 72.010 132.975 72.270 133.455 ;
        RECT 72.440 132.805 72.700 133.260 ;
        RECT 72.870 132.975 73.130 133.455 ;
        RECT 73.300 132.805 73.560 133.260 ;
        RECT 73.730 132.975 74.030 133.455 ;
        RECT 70.720 132.635 74.030 132.805 ;
        RECT 69.870 132.215 72.890 132.465 ;
        RECT 58.805 130.905 64.150 131.340 ;
        RECT 64.325 130.905 65.535 131.995 ;
        RECT 65.750 130.905 66.045 132.045 ;
        RECT 66.305 131.875 68.755 132.045 ;
        RECT 66.305 131.075 66.635 131.875 ;
        RECT 66.805 130.905 66.975 131.705 ;
        RECT 67.145 131.075 67.475 131.875 ;
        RECT 67.985 131.855 68.755 131.875 ;
        RECT 67.645 130.905 67.815 131.705 ;
        RECT 67.985 131.075 68.315 131.855 ;
        RECT 68.485 130.905 68.655 131.365 ;
        RECT 68.925 130.905 69.215 132.070 ;
        RECT 69.395 130.905 69.690 132.015 ;
        RECT 69.870 131.080 70.120 132.215 ;
        RECT 73.060 132.045 74.030 132.635 ;
        RECT 74.445 132.685 77.035 133.455 ;
        RECT 77.210 132.965 77.465 133.455 ;
        RECT 77.635 132.945 78.865 133.285 ;
        RECT 74.445 132.165 75.655 132.685 ;
        RECT 70.290 130.905 70.550 132.015 ;
        RECT 70.720 131.805 74.030 132.045 ;
        RECT 75.825 131.995 77.035 132.515 ;
        RECT 77.230 132.215 77.450 132.795 ;
        RECT 77.635 132.045 77.815 132.945 ;
        RECT 77.985 132.215 78.360 132.775 ;
        RECT 78.535 132.715 78.865 132.945 ;
        RECT 79.045 132.910 84.390 133.455 ;
        RECT 78.565 132.215 78.875 132.545 ;
        RECT 80.630 132.080 80.970 132.910 ;
        RECT 85.065 132.635 85.295 133.455 ;
        RECT 85.465 132.655 85.795 133.285 ;
        RECT 70.720 131.080 70.980 131.805 ;
        RECT 71.150 130.905 71.410 131.635 ;
        RECT 71.580 131.080 71.840 131.805 ;
        RECT 72.010 130.905 72.270 131.635 ;
        RECT 72.440 131.080 72.700 131.805 ;
        RECT 72.870 130.905 73.130 131.635 ;
        RECT 73.300 131.080 73.560 131.805 ;
        RECT 73.730 130.905 74.025 131.635 ;
        RECT 74.445 130.905 77.035 131.995 ;
        RECT 77.210 130.905 77.465 132.045 ;
        RECT 77.635 131.875 78.865 132.045 ;
        RECT 77.635 131.075 77.965 131.875 ;
        RECT 78.135 130.905 78.365 131.705 ;
        RECT 78.535 131.075 78.865 131.875 ;
        RECT 82.450 131.340 82.800 132.590 ;
        RECT 85.045 132.215 85.375 132.465 ;
        RECT 85.545 132.055 85.795 132.655 ;
        RECT 85.965 132.635 86.175 133.455 ;
        RECT 86.405 133.075 87.295 133.245 ;
        RECT 86.405 132.520 86.955 132.905 ;
        RECT 87.125 132.350 87.295 133.075 ;
        RECT 79.045 130.905 84.390 131.340 ;
        RECT 85.065 130.905 85.295 132.045 ;
        RECT 85.465 131.075 85.795 132.055 ;
        RECT 86.405 132.280 87.295 132.350 ;
        RECT 87.465 132.750 87.685 133.235 ;
        RECT 87.855 132.915 88.105 133.455 ;
        RECT 88.275 132.805 88.535 133.285 ;
        RECT 87.465 132.325 87.795 132.750 ;
        RECT 86.405 132.255 87.300 132.280 ;
        RECT 86.405 132.240 87.310 132.255 ;
        RECT 86.405 132.225 87.315 132.240 ;
        RECT 86.405 132.220 87.325 132.225 ;
        RECT 86.405 132.210 87.330 132.220 ;
        RECT 86.405 132.200 87.335 132.210 ;
        RECT 86.405 132.195 87.345 132.200 ;
        RECT 86.405 132.185 87.355 132.195 ;
        RECT 86.405 132.180 87.365 132.185 ;
        RECT 85.965 130.905 86.175 132.045 ;
        RECT 86.405 131.730 86.665 132.180 ;
        RECT 87.030 132.175 87.365 132.180 ;
        RECT 87.030 132.170 87.380 132.175 ;
        RECT 87.030 132.160 87.395 132.170 ;
        RECT 87.030 132.155 87.420 132.160 ;
        RECT 87.965 132.155 88.195 132.550 ;
        RECT 87.030 132.150 88.195 132.155 ;
        RECT 87.060 132.115 88.195 132.150 ;
        RECT 87.095 132.090 88.195 132.115 ;
        RECT 87.125 132.060 88.195 132.090 ;
        RECT 87.145 132.030 88.195 132.060 ;
        RECT 87.165 132.000 88.195 132.030 ;
        RECT 87.235 131.990 88.195 132.000 ;
        RECT 87.260 131.980 88.195 131.990 ;
        RECT 87.280 131.965 88.195 131.980 ;
        RECT 87.300 131.950 88.195 131.965 ;
        RECT 87.305 131.940 88.090 131.950 ;
        RECT 87.320 131.905 88.090 131.940 ;
        RECT 86.835 131.585 87.165 131.830 ;
        RECT 87.335 131.655 88.090 131.905 ;
        RECT 88.365 131.775 88.535 132.805 ;
        RECT 86.835 131.560 87.020 131.585 ;
        RECT 86.405 131.460 87.020 131.560 ;
        RECT 86.405 130.905 87.010 131.460 ;
        RECT 87.185 131.075 87.665 131.415 ;
        RECT 87.835 130.905 88.090 131.450 ;
        RECT 88.260 131.075 88.535 131.775 ;
        RECT 89.170 132.715 89.425 133.285 ;
        RECT 89.595 133.055 89.925 133.455 ;
        RECT 90.350 132.920 90.880 133.285 ;
        RECT 91.070 133.115 91.345 133.285 ;
        RECT 91.065 132.945 91.345 133.115 ;
        RECT 90.350 132.885 90.525 132.920 ;
        RECT 89.595 132.715 90.525 132.885 ;
        RECT 89.170 132.045 89.340 132.715 ;
        RECT 89.595 132.545 89.765 132.715 ;
        RECT 89.510 132.215 89.765 132.545 ;
        RECT 89.990 132.215 90.185 132.545 ;
        RECT 89.170 131.075 89.505 132.045 ;
        RECT 89.675 130.905 89.845 132.045 ;
        RECT 90.015 131.245 90.185 132.215 ;
        RECT 90.355 131.585 90.525 132.715 ;
        RECT 90.695 131.925 90.865 132.725 ;
        RECT 91.070 132.125 91.345 132.945 ;
        RECT 91.515 131.925 91.705 133.285 ;
        RECT 91.885 132.920 92.395 133.455 ;
        RECT 92.615 132.645 92.860 133.250 ;
        RECT 93.305 132.705 94.515 133.455 ;
        RECT 94.685 132.730 94.975 133.455 ;
        RECT 95.145 132.910 100.490 133.455 ;
        RECT 91.905 132.475 93.135 132.645 ;
        RECT 90.695 131.755 91.705 131.925 ;
        RECT 91.875 131.910 92.625 132.100 ;
        RECT 90.355 131.415 91.480 131.585 ;
        RECT 91.875 131.245 92.045 131.910 ;
        RECT 92.795 131.665 93.135 132.475 ;
        RECT 93.305 132.165 93.825 132.705 ;
        RECT 93.995 131.995 94.515 132.535 ;
        RECT 96.730 132.080 97.070 132.910 ;
        RECT 100.665 132.685 102.335 133.455 ;
        RECT 102.620 132.825 102.905 133.285 ;
        RECT 103.075 132.995 103.345 133.455 ;
        RECT 90.015 131.075 92.045 131.245 ;
        RECT 92.215 130.905 92.385 131.665 ;
        RECT 92.620 131.255 93.135 131.665 ;
        RECT 93.305 130.905 94.515 131.995 ;
        RECT 94.685 130.905 94.975 132.070 ;
        RECT 98.550 131.340 98.900 132.590 ;
        RECT 100.665 132.165 101.415 132.685 ;
        RECT 102.620 132.655 103.575 132.825 ;
        RECT 101.585 131.995 102.335 132.515 ;
        RECT 95.145 130.905 100.490 131.340 ;
        RECT 100.665 130.905 102.335 131.995 ;
        RECT 102.505 131.925 103.195 132.485 ;
        RECT 103.365 131.755 103.575 132.655 ;
        RECT 102.620 131.535 103.575 131.755 ;
        RECT 103.745 132.485 104.145 133.285 ;
        RECT 104.335 132.825 104.615 133.285 ;
        RECT 105.135 132.995 105.460 133.455 ;
        RECT 104.335 132.655 105.460 132.825 ;
        RECT 105.630 132.715 106.015 133.285 ;
        RECT 105.010 132.545 105.460 132.655 ;
        RECT 103.745 131.925 104.840 132.485 ;
        RECT 105.010 132.215 105.565 132.545 ;
        RECT 102.620 131.075 102.905 131.535 ;
        RECT 103.075 130.905 103.345 131.365 ;
        RECT 103.745 131.075 104.145 131.925 ;
        RECT 105.010 131.755 105.460 132.215 ;
        RECT 105.735 132.045 106.015 132.715 ;
        RECT 106.185 132.685 107.855 133.455 ;
        RECT 106.185 132.165 106.935 132.685 ;
        RECT 104.335 131.535 105.460 131.755 ;
        RECT 104.335 131.075 104.615 131.535 ;
        RECT 105.135 130.905 105.460 131.365 ;
        RECT 105.630 131.075 106.015 132.045 ;
        RECT 107.105 131.995 107.855 132.515 ;
        RECT 106.185 130.905 107.855 131.995 ;
        RECT 108.025 132.510 108.365 133.285 ;
        RECT 108.535 132.995 108.705 133.455 ;
        RECT 108.945 133.020 109.305 133.285 ;
        RECT 108.945 133.015 109.300 133.020 ;
        RECT 108.945 133.005 109.295 133.015 ;
        RECT 108.945 133.000 109.290 133.005 ;
        RECT 108.945 132.990 109.285 133.000 ;
        RECT 109.935 132.995 110.105 133.455 ;
        RECT 108.945 132.985 109.280 132.990 ;
        RECT 108.945 132.975 109.270 132.985 ;
        RECT 108.945 132.965 109.260 132.975 ;
        RECT 108.945 132.825 109.245 132.965 ;
        RECT 108.535 132.635 109.245 132.825 ;
        RECT 109.435 132.825 109.765 132.905 ;
        RECT 110.275 132.825 110.615 133.285 ;
        RECT 110.845 132.975 111.125 133.455 ;
        RECT 109.435 132.635 110.615 132.825 ;
        RECT 111.295 132.805 111.555 133.195 ;
        RECT 111.730 132.975 111.985 133.455 ;
        RECT 112.155 132.805 112.450 133.195 ;
        RECT 112.630 132.975 112.905 133.455 ;
        RECT 113.075 132.955 113.375 133.285 ;
        RECT 110.800 132.635 112.450 132.805 ;
        RECT 108.025 131.075 108.305 132.510 ;
        RECT 108.535 132.065 108.820 132.635 ;
        RECT 109.005 132.235 109.475 132.465 ;
        RECT 109.645 132.445 109.975 132.465 ;
        RECT 109.645 132.265 110.095 132.445 ;
        RECT 110.285 132.265 110.615 132.465 ;
        RECT 108.535 131.850 109.685 132.065 ;
        RECT 108.475 130.905 109.185 131.680 ;
        RECT 109.355 131.075 109.685 131.850 ;
        RECT 109.880 131.150 110.095 132.265 ;
        RECT 110.385 131.925 110.615 132.265 ;
        RECT 110.800 132.125 111.205 132.635 ;
        RECT 111.375 132.295 112.515 132.465 ;
        RECT 110.800 131.955 111.555 132.125 ;
        RECT 110.275 130.905 110.605 131.625 ;
        RECT 110.840 130.905 111.125 131.775 ;
        RECT 111.295 131.705 111.555 131.955 ;
        RECT 112.345 132.045 112.515 132.295 ;
        RECT 112.685 132.215 113.035 132.785 ;
        RECT 113.205 132.045 113.375 132.955 ;
        RECT 113.545 132.685 117.055 133.455 ;
        RECT 117.685 132.825 118.025 133.285 ;
        RECT 118.195 132.995 118.365 133.455 ;
        RECT 118.995 133.020 119.355 133.285 ;
        RECT 119.000 133.015 119.355 133.020 ;
        RECT 119.005 133.005 119.355 133.015 ;
        RECT 119.010 133.000 119.355 133.005 ;
        RECT 119.015 132.990 119.355 133.000 ;
        RECT 119.595 132.995 119.765 133.455 ;
        RECT 119.020 132.985 119.355 132.990 ;
        RECT 119.030 132.975 119.355 132.985 ;
        RECT 119.040 132.965 119.355 132.975 ;
        RECT 118.535 132.825 118.865 132.905 ;
        RECT 113.545 132.165 115.195 132.685 ;
        RECT 117.685 132.635 118.865 132.825 ;
        RECT 119.055 132.825 119.355 132.965 ;
        RECT 119.055 132.635 119.765 132.825 ;
        RECT 112.345 131.875 113.375 132.045 ;
        RECT 115.365 131.995 117.055 132.515 ;
        RECT 111.295 131.535 112.415 131.705 ;
        RECT 111.295 131.075 111.555 131.535 ;
        RECT 111.730 130.905 111.985 131.365 ;
        RECT 112.155 131.075 112.415 131.535 ;
        RECT 112.585 130.905 112.895 131.705 ;
        RECT 113.065 131.075 113.375 131.875 ;
        RECT 113.545 130.905 117.055 131.995 ;
        RECT 117.685 132.265 118.015 132.465 ;
        RECT 118.325 132.445 118.655 132.465 ;
        RECT 118.205 132.265 118.655 132.445 ;
        RECT 117.685 131.925 117.915 132.265 ;
        RECT 117.695 130.905 118.025 131.625 ;
        RECT 118.205 131.150 118.420 132.265 ;
        RECT 118.825 132.235 119.295 132.465 ;
        RECT 119.480 132.065 119.765 132.635 ;
        RECT 119.935 132.510 120.275 133.285 ;
        RECT 120.445 132.730 120.735 133.455 ;
        RECT 120.955 132.800 121.285 133.235 ;
        RECT 121.455 132.845 121.625 133.455 ;
        RECT 118.615 131.850 119.765 132.065 ;
        RECT 118.615 131.075 118.945 131.850 ;
        RECT 119.115 130.905 119.825 131.680 ;
        RECT 119.995 131.075 120.275 132.510 ;
        RECT 120.905 132.715 121.285 132.800 ;
        RECT 121.795 132.715 122.125 133.240 ;
        RECT 122.385 132.925 122.595 133.455 ;
        RECT 122.870 133.005 123.655 133.175 ;
        RECT 123.825 133.005 124.230 133.175 ;
        RECT 120.905 132.675 121.130 132.715 ;
        RECT 120.905 132.095 121.075 132.675 ;
        RECT 121.795 132.545 121.995 132.715 ;
        RECT 122.870 132.545 123.040 133.005 ;
        RECT 121.245 132.215 121.995 132.545 ;
        RECT 122.165 132.215 123.040 132.545 ;
        RECT 120.445 130.905 120.735 132.070 ;
        RECT 120.905 132.045 121.120 132.095 ;
        RECT 120.905 131.965 121.295 132.045 ;
        RECT 120.965 131.120 121.295 131.965 ;
        RECT 121.805 132.010 121.995 132.215 ;
        RECT 121.465 130.905 121.635 131.915 ;
        RECT 121.805 131.635 122.700 132.010 ;
        RECT 121.805 131.075 122.145 131.635 ;
        RECT 122.375 130.905 122.690 131.405 ;
        RECT 122.870 131.375 123.040 132.215 ;
        RECT 123.210 132.505 123.675 132.835 ;
        RECT 124.060 132.775 124.230 133.005 ;
        RECT 124.410 132.955 124.780 133.455 ;
        RECT 125.100 133.005 125.775 133.175 ;
        RECT 125.970 133.005 126.305 133.175 ;
        RECT 123.210 131.545 123.530 132.505 ;
        RECT 124.060 132.475 124.890 132.775 ;
        RECT 123.700 131.575 123.890 132.295 ;
        RECT 124.060 131.405 124.230 132.475 ;
        RECT 124.690 132.445 124.890 132.475 ;
        RECT 124.400 132.225 124.570 132.295 ;
        RECT 125.100 132.225 125.270 133.005 ;
        RECT 126.135 132.865 126.305 133.005 ;
        RECT 126.475 132.995 126.725 133.455 ;
        RECT 124.400 132.055 125.270 132.225 ;
        RECT 125.440 132.585 125.965 132.805 ;
        RECT 126.135 132.735 126.360 132.865 ;
        RECT 124.400 131.965 124.910 132.055 ;
        RECT 122.870 131.205 123.755 131.375 ;
        RECT 123.980 131.075 124.230 131.405 ;
        RECT 124.400 130.905 124.570 131.705 ;
        RECT 124.740 131.350 124.910 131.965 ;
        RECT 125.440 131.885 125.610 132.585 ;
        RECT 125.080 131.520 125.610 131.885 ;
        RECT 125.780 131.820 126.020 132.415 ;
        RECT 126.190 131.630 126.360 132.735 ;
        RECT 126.530 131.875 126.810 132.825 ;
        RECT 126.055 131.500 126.360 131.630 ;
        RECT 124.740 131.180 125.845 131.350 ;
        RECT 126.055 131.075 126.305 131.500 ;
        RECT 126.475 130.905 126.740 131.365 ;
        RECT 126.980 131.075 127.165 133.195 ;
        RECT 127.335 133.075 127.665 133.455 ;
        RECT 127.835 132.905 128.005 133.195 ;
        RECT 127.340 132.735 128.005 132.905 ;
        RECT 127.340 131.745 127.570 132.735 ;
        RECT 127.740 131.915 128.090 132.565 ;
        RECT 128.265 132.510 128.605 133.285 ;
        RECT 128.775 132.995 128.945 133.455 ;
        RECT 129.185 133.020 129.545 133.285 ;
        RECT 129.185 133.015 129.540 133.020 ;
        RECT 129.185 133.005 129.535 133.015 ;
        RECT 129.185 133.000 129.530 133.005 ;
        RECT 129.185 132.990 129.525 133.000 ;
        RECT 130.175 132.995 130.345 133.455 ;
        RECT 129.185 132.985 129.520 132.990 ;
        RECT 129.185 132.975 129.510 132.985 ;
        RECT 129.185 132.965 129.500 132.975 ;
        RECT 129.185 132.825 129.485 132.965 ;
        RECT 128.775 132.635 129.485 132.825 ;
        RECT 129.675 132.825 130.005 132.905 ;
        RECT 130.515 132.825 130.855 133.285 ;
        RECT 129.675 132.635 130.855 132.825 ;
        RECT 131.025 132.685 133.615 133.455 ;
        RECT 133.790 132.715 134.045 133.285 ;
        RECT 134.215 133.055 134.545 133.455 ;
        RECT 134.970 132.920 135.500 133.285 ;
        RECT 135.690 133.115 135.965 133.285 ;
        RECT 135.685 132.945 135.965 133.115 ;
        RECT 134.970 132.885 135.145 132.920 ;
        RECT 134.215 132.715 135.145 132.885 ;
        RECT 127.340 131.575 128.005 131.745 ;
        RECT 127.335 130.905 127.665 131.405 ;
        RECT 127.835 131.075 128.005 131.575 ;
        RECT 128.265 131.075 128.545 132.510 ;
        RECT 128.775 132.065 129.060 132.635 ;
        RECT 129.245 132.235 129.715 132.465 ;
        RECT 129.885 132.445 130.215 132.465 ;
        RECT 129.885 132.265 130.335 132.445 ;
        RECT 130.525 132.265 130.855 132.465 ;
        RECT 128.775 131.850 129.925 132.065 ;
        RECT 128.715 130.905 129.425 131.680 ;
        RECT 129.595 131.075 129.925 131.850 ;
        RECT 130.120 131.150 130.335 132.265 ;
        RECT 130.625 131.925 130.855 132.265 ;
        RECT 131.025 132.165 132.235 132.685 ;
        RECT 132.405 131.995 133.615 132.515 ;
        RECT 130.515 130.905 130.845 131.625 ;
        RECT 131.025 130.905 133.615 131.995 ;
        RECT 133.790 132.045 133.960 132.715 ;
        RECT 134.215 132.545 134.385 132.715 ;
        RECT 134.130 132.215 134.385 132.545 ;
        RECT 134.610 132.215 134.805 132.545 ;
        RECT 133.790 131.075 134.125 132.045 ;
        RECT 134.295 130.905 134.465 132.045 ;
        RECT 134.635 131.245 134.805 132.215 ;
        RECT 134.975 131.585 135.145 132.715 ;
        RECT 135.315 131.925 135.485 132.725 ;
        RECT 135.690 132.125 135.965 132.945 ;
        RECT 136.135 131.925 136.325 133.285 ;
        RECT 136.505 132.920 137.015 133.455 ;
        RECT 137.235 132.645 137.480 133.250 ;
        RECT 137.930 132.715 138.185 133.285 ;
        RECT 138.355 133.055 138.685 133.455 ;
        RECT 139.110 132.920 139.640 133.285 ;
        RECT 139.110 132.885 139.285 132.920 ;
        RECT 138.355 132.715 139.285 132.885 ;
        RECT 139.830 132.775 140.105 133.285 ;
        RECT 136.525 132.475 137.755 132.645 ;
        RECT 135.315 131.755 136.325 131.925 ;
        RECT 136.495 131.910 137.245 132.100 ;
        RECT 134.975 131.415 136.100 131.585 ;
        RECT 136.495 131.245 136.665 131.910 ;
        RECT 137.415 131.665 137.755 132.475 ;
        RECT 134.635 131.075 136.665 131.245 ;
        RECT 136.835 130.905 137.005 131.665 ;
        RECT 137.240 131.255 137.755 131.665 ;
        RECT 137.930 132.045 138.100 132.715 ;
        RECT 138.355 132.545 138.525 132.715 ;
        RECT 138.270 132.215 138.525 132.545 ;
        RECT 138.750 132.215 138.945 132.545 ;
        RECT 137.930 131.075 138.265 132.045 ;
        RECT 138.435 130.905 138.605 132.045 ;
        RECT 138.775 131.245 138.945 132.215 ;
        RECT 139.115 131.585 139.285 132.715 ;
        RECT 139.455 131.925 139.625 132.725 ;
        RECT 139.825 132.605 140.105 132.775 ;
        RECT 139.830 132.125 140.105 132.605 ;
        RECT 140.275 131.925 140.465 133.285 ;
        RECT 140.645 132.920 141.155 133.455 ;
        RECT 141.375 132.645 141.620 133.250 ;
        RECT 142.155 132.905 142.325 133.285 ;
        RECT 142.505 133.075 142.835 133.455 ;
        RECT 142.155 132.735 142.820 132.905 ;
        RECT 143.015 132.780 143.275 133.285 ;
        RECT 140.665 132.475 141.895 132.645 ;
        RECT 139.455 131.755 140.465 131.925 ;
        RECT 140.635 131.910 141.385 132.100 ;
        RECT 139.115 131.415 140.240 131.585 ;
        RECT 140.635 131.245 140.805 131.910 ;
        RECT 141.555 131.665 141.895 132.475 ;
        RECT 142.085 132.185 142.415 132.555 ;
        RECT 142.650 132.480 142.820 132.735 ;
        RECT 142.650 132.150 142.935 132.480 ;
        RECT 142.650 132.005 142.820 132.150 ;
        RECT 138.775 131.075 140.805 131.245 ;
        RECT 140.975 130.905 141.145 131.665 ;
        RECT 141.380 131.255 141.895 131.665 ;
        RECT 142.155 131.835 142.820 132.005 ;
        RECT 143.105 131.980 143.275 132.780 ;
        RECT 143.995 132.905 144.165 133.285 ;
        RECT 144.380 133.075 144.710 133.455 ;
        RECT 143.995 132.735 144.710 132.905 ;
        RECT 143.905 132.185 144.260 132.555 ;
        RECT 144.540 132.545 144.710 132.735 ;
        RECT 144.880 132.710 145.135 133.285 ;
        RECT 144.540 132.215 144.795 132.545 ;
        RECT 144.540 132.005 144.710 132.215 ;
        RECT 142.155 131.075 142.325 131.835 ;
        RECT 142.505 130.905 142.835 131.665 ;
        RECT 143.005 131.075 143.275 131.980 ;
        RECT 143.995 131.835 144.710 132.005 ;
        RECT 144.965 131.980 145.135 132.710 ;
        RECT 145.310 132.615 145.570 133.455 ;
        RECT 145.745 132.705 146.955 133.455 ;
        RECT 143.995 131.075 144.165 131.835 ;
        RECT 144.380 130.905 144.710 131.665 ;
        RECT 144.880 131.075 145.135 131.980 ;
        RECT 145.310 130.905 145.570 132.055 ;
        RECT 145.745 131.995 146.265 132.535 ;
        RECT 146.435 132.165 146.955 132.705 ;
        RECT 145.745 130.905 146.955 131.995 ;
        RECT 17.320 130.735 147.040 130.905 ;
        RECT 17.405 129.645 18.615 130.735 ;
        RECT 17.405 128.935 17.925 129.475 ;
        RECT 18.095 129.105 18.615 129.645 ;
        RECT 18.790 129.595 19.125 130.565 ;
        RECT 19.295 129.595 19.465 130.735 ;
        RECT 19.635 130.395 21.665 130.565 ;
        RECT 17.405 128.185 18.615 128.935 ;
        RECT 18.790 128.925 18.960 129.595 ;
        RECT 19.635 129.425 19.805 130.395 ;
        RECT 19.130 129.095 19.385 129.425 ;
        RECT 19.610 129.095 19.805 129.425 ;
        RECT 19.975 130.055 21.100 130.225 ;
        RECT 19.215 128.925 19.385 129.095 ;
        RECT 19.975 128.925 20.145 130.055 ;
        RECT 18.790 128.355 19.045 128.925 ;
        RECT 19.215 128.755 20.145 128.925 ;
        RECT 20.315 129.715 21.325 129.885 ;
        RECT 20.315 128.915 20.485 129.715 ;
        RECT 20.690 129.375 20.965 129.515 ;
        RECT 20.685 129.205 20.965 129.375 ;
        RECT 19.970 128.720 20.145 128.755 ;
        RECT 19.215 128.185 19.545 128.585 ;
        RECT 19.970 128.355 20.500 128.720 ;
        RECT 20.690 128.355 20.965 129.205 ;
        RECT 21.135 128.355 21.325 129.715 ;
        RECT 21.495 129.730 21.665 130.395 ;
        RECT 21.835 129.975 22.005 130.735 ;
        RECT 22.240 129.975 22.755 130.385 ;
        RECT 21.495 129.540 22.245 129.730 ;
        RECT 22.415 129.165 22.755 129.975 ;
        RECT 22.985 129.675 23.315 130.520 ;
        RECT 23.485 129.725 23.655 130.735 ;
        RECT 23.825 130.005 24.165 130.565 ;
        RECT 24.395 130.235 24.710 130.735 ;
        RECT 24.890 130.265 25.775 130.435 ;
        RECT 21.525 128.995 22.755 129.165 ;
        RECT 22.925 129.595 23.315 129.675 ;
        RECT 23.825 129.630 24.720 130.005 ;
        RECT 22.925 129.545 23.140 129.595 ;
        RECT 21.505 128.185 22.015 128.720 ;
        RECT 22.235 128.390 22.480 128.995 ;
        RECT 22.925 128.965 23.095 129.545 ;
        RECT 23.825 129.425 24.015 129.630 ;
        RECT 24.890 129.425 25.060 130.265 ;
        RECT 26.000 130.235 26.250 130.565 ;
        RECT 23.265 129.095 24.015 129.425 ;
        RECT 24.185 129.095 25.060 129.425 ;
        RECT 22.925 128.925 23.150 128.965 ;
        RECT 23.815 128.925 24.015 129.095 ;
        RECT 22.925 128.840 23.305 128.925 ;
        RECT 22.975 128.405 23.305 128.840 ;
        RECT 23.475 128.185 23.645 128.795 ;
        RECT 23.815 128.400 24.145 128.925 ;
        RECT 24.405 128.185 24.615 128.715 ;
        RECT 24.890 128.635 25.060 129.095 ;
        RECT 25.230 129.135 25.550 130.095 ;
        RECT 25.720 129.345 25.910 130.065 ;
        RECT 26.080 129.165 26.250 130.235 ;
        RECT 26.420 129.935 26.590 130.735 ;
        RECT 26.760 130.290 27.865 130.460 ;
        RECT 26.760 129.675 26.930 130.290 ;
        RECT 28.075 130.140 28.325 130.565 ;
        RECT 28.495 130.275 28.760 130.735 ;
        RECT 27.100 129.755 27.630 130.120 ;
        RECT 28.075 130.010 28.380 130.140 ;
        RECT 26.420 129.585 26.930 129.675 ;
        RECT 26.420 129.415 27.290 129.585 ;
        RECT 26.420 129.345 26.590 129.415 ;
        RECT 26.710 129.165 26.910 129.195 ;
        RECT 25.230 128.805 25.695 129.135 ;
        RECT 26.080 128.865 26.910 129.165 ;
        RECT 26.080 128.635 26.250 128.865 ;
        RECT 24.890 128.465 25.675 128.635 ;
        RECT 25.845 128.465 26.250 128.635 ;
        RECT 26.430 128.185 26.800 128.685 ;
        RECT 27.120 128.635 27.290 129.415 ;
        RECT 27.460 129.055 27.630 129.755 ;
        RECT 27.800 129.225 28.040 129.820 ;
        RECT 27.460 128.835 27.985 129.055 ;
        RECT 28.210 128.905 28.380 130.010 ;
        RECT 28.155 128.775 28.380 128.905 ;
        RECT 28.550 128.815 28.830 129.765 ;
        RECT 28.155 128.635 28.325 128.775 ;
        RECT 27.120 128.465 27.795 128.635 ;
        RECT 27.990 128.465 28.325 128.635 ;
        RECT 28.495 128.185 28.745 128.645 ;
        RECT 29.000 128.445 29.185 130.565 ;
        RECT 29.355 130.235 29.685 130.735 ;
        RECT 29.855 130.065 30.025 130.565 ;
        RECT 29.360 129.895 30.025 130.065 ;
        RECT 29.360 128.905 29.590 129.895 ;
        RECT 29.760 129.075 30.110 129.725 ;
        RECT 30.285 129.570 30.575 130.735 ;
        RECT 30.745 129.935 31.185 130.565 ;
        RECT 30.745 128.925 31.055 129.935 ;
        RECT 31.360 129.885 31.675 130.735 ;
        RECT 31.845 130.395 33.275 130.565 ;
        RECT 31.845 129.715 32.015 130.395 ;
        RECT 31.225 129.545 32.015 129.715 ;
        RECT 31.225 129.095 31.395 129.545 ;
        RECT 32.185 129.425 32.385 130.225 ;
        RECT 31.565 129.095 31.955 129.375 ;
        RECT 32.140 129.095 32.385 129.425 ;
        RECT 32.585 129.095 32.835 130.225 ;
        RECT 33.025 129.765 33.275 130.395 ;
        RECT 33.455 129.935 33.785 130.735 ;
        RECT 33.965 130.300 39.310 130.735 ;
        RECT 39.485 130.300 44.830 130.735 ;
        RECT 45.005 130.300 50.350 130.735 ;
        RECT 50.525 130.300 55.870 130.735 ;
        RECT 33.025 129.595 33.795 129.765 ;
        RECT 33.050 129.095 33.455 129.425 ;
        RECT 33.625 128.925 33.795 129.595 ;
        RECT 29.360 128.735 30.025 128.905 ;
        RECT 29.355 128.185 29.685 128.565 ;
        RECT 29.855 128.445 30.025 128.735 ;
        RECT 30.285 128.185 30.575 128.910 ;
        RECT 30.745 128.365 31.185 128.925 ;
        RECT 31.355 128.185 31.805 128.925 ;
        RECT 31.975 128.755 33.135 128.925 ;
        RECT 31.975 128.355 32.145 128.755 ;
        RECT 32.315 128.185 32.735 128.585 ;
        RECT 32.905 128.355 33.135 128.755 ;
        RECT 33.305 128.355 33.795 128.925 ;
        RECT 35.550 128.730 35.890 129.560 ;
        RECT 37.370 129.050 37.720 130.300 ;
        RECT 41.070 128.730 41.410 129.560 ;
        RECT 42.890 129.050 43.240 130.300 ;
        RECT 46.590 128.730 46.930 129.560 ;
        RECT 48.410 129.050 48.760 130.300 ;
        RECT 52.110 128.730 52.450 129.560 ;
        RECT 53.930 129.050 54.280 130.300 ;
        RECT 56.045 129.570 56.335 130.735 ;
        RECT 56.505 130.300 61.850 130.735 ;
        RECT 62.025 130.300 67.370 130.735 ;
        RECT 33.965 128.185 39.310 128.730 ;
        RECT 39.485 128.185 44.830 128.730 ;
        RECT 45.005 128.185 50.350 128.730 ;
        RECT 50.525 128.185 55.870 128.730 ;
        RECT 56.045 128.185 56.335 128.910 ;
        RECT 58.090 128.730 58.430 129.560 ;
        RECT 59.910 129.050 60.260 130.300 ;
        RECT 63.610 128.730 63.950 129.560 ;
        RECT 65.430 129.050 65.780 130.300 ;
        RECT 67.545 129.645 68.755 130.735 ;
        RECT 67.545 128.935 68.065 129.475 ;
        RECT 68.235 129.105 68.755 129.645 ;
        RECT 68.925 129.885 69.305 130.565 ;
        RECT 69.895 129.885 70.065 130.735 ;
        RECT 70.235 130.055 70.565 130.565 ;
        RECT 70.735 130.225 70.905 130.735 ;
        RECT 71.075 130.055 71.475 130.565 ;
        RECT 70.235 129.885 71.475 130.055 ;
        RECT 56.505 128.185 61.850 128.730 ;
        RECT 62.025 128.185 67.370 128.730 ;
        RECT 67.545 128.185 68.755 128.935 ;
        RECT 68.925 128.925 69.095 129.885 ;
        RECT 69.265 129.545 70.570 129.715 ;
        RECT 71.655 129.635 71.975 130.565 ;
        RECT 69.265 129.095 69.510 129.545 ;
        RECT 69.680 129.175 70.230 129.375 ;
        RECT 70.400 129.345 70.570 129.545 ;
        RECT 71.345 129.465 71.975 129.635 ;
        RECT 72.145 129.865 72.420 130.565 ;
        RECT 72.630 130.190 72.845 130.735 ;
        RECT 73.015 130.225 73.490 130.565 ;
        RECT 73.660 130.230 74.275 130.735 ;
        RECT 73.660 130.055 73.855 130.230 ;
        RECT 70.400 129.175 70.775 129.345 ;
        RECT 70.945 128.925 71.175 129.425 ;
        RECT 68.925 128.755 71.175 128.925 ;
        RECT 68.975 128.185 69.305 128.575 ;
        RECT 69.475 128.435 69.645 128.755 ;
        RECT 71.345 128.585 71.515 129.465 ;
        RECT 69.815 128.185 70.145 128.575 ;
        RECT 70.560 128.415 71.515 128.585 ;
        RECT 71.685 128.185 71.975 129.020 ;
        RECT 72.145 128.835 72.315 129.865 ;
        RECT 72.590 129.695 73.305 129.990 ;
        RECT 73.525 129.865 73.855 130.055 ;
        RECT 74.025 129.695 74.275 130.060 ;
        RECT 72.485 129.525 74.275 129.695 ;
        RECT 72.485 129.095 72.715 129.525 ;
        RECT 72.145 128.355 72.405 128.835 ;
        RECT 72.885 128.825 73.295 129.345 ;
        RECT 72.575 128.185 72.905 128.645 ;
        RECT 73.095 128.405 73.295 128.825 ;
        RECT 73.465 128.670 73.720 129.525 ;
        RECT 74.515 129.345 74.685 130.565 ;
        RECT 74.935 130.225 75.195 130.735 ;
        RECT 75.365 130.300 80.710 130.735 ;
        RECT 73.890 129.095 74.685 129.345 ;
        RECT 74.855 129.175 75.195 130.055 ;
        RECT 74.435 129.005 74.685 129.095 ;
        RECT 73.465 128.405 74.255 128.670 ;
        RECT 74.435 128.585 74.765 129.005 ;
        RECT 74.935 128.185 75.195 129.005 ;
        RECT 76.950 128.730 77.290 129.560 ;
        RECT 78.770 129.050 79.120 130.300 ;
        RECT 81.805 129.570 82.095 130.735 ;
        RECT 82.725 130.225 83.915 130.515 ;
        RECT 82.745 129.885 83.915 130.055 ;
        RECT 84.085 129.935 84.365 130.735 ;
        RECT 82.745 129.595 83.070 129.885 ;
        RECT 83.745 129.765 83.915 129.885 ;
        RECT 83.240 129.425 83.435 129.715 ;
        RECT 83.745 129.595 84.405 129.765 ;
        RECT 84.575 129.595 84.850 130.565 ;
        RECT 85.025 129.595 85.285 130.735 ;
        RECT 85.525 130.225 87.140 130.555 ;
        RECT 84.235 129.425 84.405 129.595 ;
        RECT 82.725 129.095 83.070 129.425 ;
        RECT 83.240 129.095 84.065 129.425 ;
        RECT 84.235 129.095 84.510 129.425 ;
        RECT 84.235 128.925 84.405 129.095 ;
        RECT 75.365 128.185 80.710 128.730 ;
        RECT 81.805 128.185 82.095 128.910 ;
        RECT 82.740 128.755 84.405 128.925 ;
        RECT 84.680 128.860 84.850 129.595 ;
        RECT 85.535 129.425 85.705 129.985 ;
        RECT 85.965 129.885 87.140 130.055 ;
        RECT 87.310 129.935 87.590 130.735 ;
        RECT 85.965 129.595 86.295 129.885 ;
        RECT 86.970 129.765 87.140 129.885 ;
        RECT 86.465 129.425 86.710 129.715 ;
        RECT 86.970 129.595 87.630 129.765 ;
        RECT 87.800 129.595 88.075 130.565 ;
        RECT 87.460 129.425 87.630 129.595 ;
        RECT 85.030 129.175 85.365 129.425 ;
        RECT 85.535 129.095 86.250 129.425 ;
        RECT 86.465 129.095 87.290 129.425 ;
        RECT 87.460 129.095 87.735 129.425 ;
        RECT 85.535 129.005 85.785 129.095 ;
        RECT 82.740 128.405 82.995 128.755 ;
        RECT 83.165 128.185 83.495 128.585 ;
        RECT 83.665 128.405 83.835 128.755 ;
        RECT 84.005 128.185 84.385 128.585 ;
        RECT 84.575 128.515 84.850 128.860 ;
        RECT 85.025 128.185 85.285 129.005 ;
        RECT 85.455 128.585 85.785 129.005 ;
        RECT 87.460 128.925 87.630 129.095 ;
        RECT 85.965 128.755 87.630 128.925 ;
        RECT 87.905 128.860 88.075 129.595 ;
        RECT 85.965 128.355 86.225 128.755 ;
        RECT 86.395 128.185 86.725 128.585 ;
        RECT 86.895 128.405 87.065 128.755 ;
        RECT 87.235 128.185 87.610 128.585 ;
        RECT 87.800 128.515 88.075 128.860 ;
        RECT 88.250 129.595 88.585 130.565 ;
        RECT 88.755 129.595 88.925 130.735 ;
        RECT 89.095 130.395 91.125 130.565 ;
        RECT 88.250 128.925 88.420 129.595 ;
        RECT 89.095 129.425 89.265 130.395 ;
        RECT 88.590 129.095 88.845 129.425 ;
        RECT 89.070 129.095 89.265 129.425 ;
        RECT 89.435 130.055 90.560 130.225 ;
        RECT 88.675 128.925 88.845 129.095 ;
        RECT 89.435 128.925 89.605 130.055 ;
        RECT 88.250 128.355 88.505 128.925 ;
        RECT 88.675 128.755 89.605 128.925 ;
        RECT 89.775 129.715 90.785 129.885 ;
        RECT 89.775 128.915 89.945 129.715 ;
        RECT 90.150 129.375 90.425 129.515 ;
        RECT 90.145 129.205 90.425 129.375 ;
        RECT 89.430 128.720 89.605 128.755 ;
        RECT 88.675 128.185 89.005 128.585 ;
        RECT 89.430 128.355 89.960 128.720 ;
        RECT 90.150 128.355 90.425 129.205 ;
        RECT 90.595 128.355 90.785 129.715 ;
        RECT 90.955 129.730 91.125 130.395 ;
        RECT 91.295 129.975 91.465 130.735 ;
        RECT 91.700 129.975 92.215 130.385 ;
        RECT 90.955 129.540 91.705 129.730 ;
        RECT 91.875 129.165 92.215 129.975 ;
        RECT 90.985 128.995 92.215 129.165 ;
        RECT 92.390 129.595 92.725 130.565 ;
        RECT 92.895 129.595 93.065 130.735 ;
        RECT 93.235 130.395 95.265 130.565 ;
        RECT 90.965 128.185 91.475 128.720 ;
        RECT 91.695 128.390 91.940 128.995 ;
        RECT 92.390 128.925 92.560 129.595 ;
        RECT 93.235 129.425 93.405 130.395 ;
        RECT 92.730 129.095 92.985 129.425 ;
        RECT 93.210 129.095 93.405 129.425 ;
        RECT 93.575 130.055 94.700 130.225 ;
        RECT 92.815 128.925 92.985 129.095 ;
        RECT 93.575 128.925 93.745 130.055 ;
        RECT 92.390 128.355 92.645 128.925 ;
        RECT 92.815 128.755 93.745 128.925 ;
        RECT 93.915 129.715 94.925 129.885 ;
        RECT 93.915 128.915 94.085 129.715 ;
        RECT 94.290 129.035 94.565 129.515 ;
        RECT 94.285 128.865 94.565 129.035 ;
        RECT 93.570 128.720 93.745 128.755 ;
        RECT 92.815 128.185 93.145 128.585 ;
        RECT 93.570 128.355 94.100 128.720 ;
        RECT 94.290 128.355 94.565 128.865 ;
        RECT 94.735 128.355 94.925 129.715 ;
        RECT 95.095 129.730 95.265 130.395 ;
        RECT 95.435 129.975 95.605 130.735 ;
        RECT 95.840 129.975 96.355 130.385 ;
        RECT 95.095 129.540 95.845 129.730 ;
        RECT 96.015 129.165 96.355 129.975 ;
        RECT 96.525 129.645 100.035 130.735 ;
        RECT 95.125 128.995 96.355 129.165 ;
        RECT 95.105 128.185 95.615 128.720 ;
        RECT 95.835 128.390 96.080 128.995 ;
        RECT 96.525 128.955 98.175 129.475 ;
        RECT 98.345 129.125 100.035 129.645 ;
        RECT 100.670 129.595 100.925 130.735 ;
        RECT 101.095 129.765 101.425 130.565 ;
        RECT 101.595 129.935 101.765 130.735 ;
        RECT 101.935 129.765 102.265 130.565 ;
        RECT 102.435 129.935 102.605 130.735 ;
        RECT 102.775 129.765 103.105 130.565 ;
        RECT 103.275 129.935 103.445 130.735 ;
        RECT 103.615 129.765 103.945 130.565 ;
        RECT 104.115 129.935 104.365 130.735 ;
        RECT 101.095 129.595 103.945 129.765 ;
        RECT 100.690 129.175 102.310 129.425 ;
        RECT 102.490 129.175 103.025 129.595 ;
        RECT 103.195 129.175 104.635 129.425 ;
        RECT 96.525 128.185 100.035 128.955 ;
        RECT 100.670 128.815 102.605 129.005 ;
        RECT 100.670 128.355 101.005 128.815 ;
        RECT 101.175 128.185 101.345 128.645 ;
        RECT 101.515 128.355 101.845 128.815 ;
        RECT 102.015 128.185 102.185 128.645 ;
        RECT 102.355 128.565 102.605 128.815 ;
        RECT 102.775 128.905 103.025 129.175 ;
        RECT 104.805 129.130 105.085 130.565 ;
        RECT 105.255 129.960 105.965 130.735 ;
        RECT 106.135 129.790 106.465 130.565 ;
        RECT 105.315 129.575 106.465 129.790 ;
        RECT 102.775 128.735 103.945 128.905 ;
        RECT 104.115 128.565 104.365 128.985 ;
        RECT 102.355 128.355 104.365 128.565 ;
        RECT 104.805 128.355 105.145 129.130 ;
        RECT 105.315 129.005 105.600 129.575 ;
        RECT 105.785 129.175 106.255 129.405 ;
        RECT 106.660 129.375 106.875 130.490 ;
        RECT 107.055 130.015 107.385 130.735 ;
        RECT 107.165 129.375 107.395 129.715 ;
        RECT 107.565 129.570 107.855 130.735 ;
        RECT 108.025 129.645 109.695 130.735 ;
        RECT 106.425 129.195 106.875 129.375 ;
        RECT 106.425 129.175 106.755 129.195 ;
        RECT 107.065 129.175 107.395 129.375 ;
        RECT 105.315 128.815 106.025 129.005 ;
        RECT 105.725 128.675 106.025 128.815 ;
        RECT 106.215 128.815 107.395 129.005 ;
        RECT 108.025 128.955 108.775 129.475 ;
        RECT 108.945 129.125 109.695 129.645 ;
        RECT 110.325 129.595 110.710 130.565 ;
        RECT 110.880 130.275 111.205 130.735 ;
        RECT 111.725 130.105 112.005 130.565 ;
        RECT 110.880 129.885 112.005 130.105 ;
        RECT 106.215 128.735 106.545 128.815 ;
        RECT 105.725 128.665 106.040 128.675 ;
        RECT 105.725 128.655 106.050 128.665 ;
        RECT 105.725 128.650 106.060 128.655 ;
        RECT 105.315 128.185 105.485 128.645 ;
        RECT 105.725 128.640 106.065 128.650 ;
        RECT 105.725 128.635 106.070 128.640 ;
        RECT 105.725 128.625 106.075 128.635 ;
        RECT 105.725 128.620 106.080 128.625 ;
        RECT 105.725 128.355 106.085 128.620 ;
        RECT 106.715 128.185 106.885 128.645 ;
        RECT 107.055 128.355 107.395 128.815 ;
        RECT 107.565 128.185 107.855 128.910 ;
        RECT 108.025 128.185 109.695 128.955 ;
        RECT 110.325 128.925 110.605 129.595 ;
        RECT 110.880 129.425 111.330 129.885 ;
        RECT 112.195 129.715 112.595 130.565 ;
        RECT 112.995 130.275 113.265 130.735 ;
        RECT 113.435 130.105 113.720 130.565 ;
        RECT 110.775 129.095 111.330 129.425 ;
        RECT 111.500 129.155 112.595 129.715 ;
        RECT 110.880 128.985 111.330 129.095 ;
        RECT 110.325 128.355 110.710 128.925 ;
        RECT 110.880 128.815 112.005 128.985 ;
        RECT 110.880 128.185 111.205 128.645 ;
        RECT 111.725 128.355 112.005 128.815 ;
        RECT 112.195 128.355 112.595 129.155 ;
        RECT 112.765 129.885 113.720 130.105 ;
        RECT 114.095 130.065 114.265 130.565 ;
        RECT 114.435 130.235 114.765 130.735 ;
        RECT 114.095 129.895 114.760 130.065 ;
        RECT 112.765 128.985 112.975 129.885 ;
        RECT 113.145 129.155 113.835 129.715 ;
        RECT 114.010 129.075 114.360 129.725 ;
        RECT 112.765 128.815 113.720 128.985 ;
        RECT 114.530 128.905 114.760 129.895 ;
        RECT 112.995 128.185 113.265 128.645 ;
        RECT 113.435 128.355 113.720 128.815 ;
        RECT 114.095 128.735 114.760 128.905 ;
        RECT 114.095 128.445 114.265 128.735 ;
        RECT 114.435 128.185 114.765 128.565 ;
        RECT 114.935 128.445 115.120 130.565 ;
        RECT 115.360 130.275 115.625 130.735 ;
        RECT 115.795 130.140 116.045 130.565 ;
        RECT 116.255 130.290 117.360 130.460 ;
        RECT 115.740 130.010 116.045 130.140 ;
        RECT 115.290 128.815 115.570 129.765 ;
        RECT 115.740 128.905 115.910 130.010 ;
        RECT 116.080 129.225 116.320 129.820 ;
        RECT 116.490 129.755 117.020 130.120 ;
        RECT 116.490 129.055 116.660 129.755 ;
        RECT 117.190 129.675 117.360 130.290 ;
        RECT 117.530 129.935 117.700 130.735 ;
        RECT 117.870 130.235 118.120 130.565 ;
        RECT 118.345 130.265 119.230 130.435 ;
        RECT 117.190 129.585 117.700 129.675 ;
        RECT 115.740 128.775 115.965 128.905 ;
        RECT 116.135 128.835 116.660 129.055 ;
        RECT 116.830 129.415 117.700 129.585 ;
        RECT 115.375 128.185 115.625 128.645 ;
        RECT 115.795 128.635 115.965 128.775 ;
        RECT 116.830 128.635 117.000 129.415 ;
        RECT 117.530 129.345 117.700 129.415 ;
        RECT 117.210 129.165 117.410 129.195 ;
        RECT 117.870 129.165 118.040 130.235 ;
        RECT 118.210 129.345 118.400 130.065 ;
        RECT 117.210 128.865 118.040 129.165 ;
        RECT 118.570 129.135 118.890 130.095 ;
        RECT 115.795 128.465 116.130 128.635 ;
        RECT 116.325 128.465 117.000 128.635 ;
        RECT 117.320 128.185 117.690 128.685 ;
        RECT 117.870 128.635 118.040 128.865 ;
        RECT 118.425 128.805 118.890 129.135 ;
        RECT 119.060 129.425 119.230 130.265 ;
        RECT 119.410 130.235 119.725 130.735 ;
        RECT 119.955 130.005 120.295 130.565 ;
        RECT 119.400 129.630 120.295 130.005 ;
        RECT 120.465 129.725 120.635 130.735 ;
        RECT 120.105 129.425 120.295 129.630 ;
        RECT 120.805 129.675 121.135 130.520 ;
        RECT 121.455 130.065 121.625 130.565 ;
        RECT 121.795 130.235 122.125 130.735 ;
        RECT 121.455 129.895 122.120 130.065 ;
        RECT 120.805 129.595 121.195 129.675 ;
        RECT 120.980 129.545 121.195 129.595 ;
        RECT 119.060 129.095 119.935 129.425 ;
        RECT 120.105 129.095 120.855 129.425 ;
        RECT 119.060 128.635 119.230 129.095 ;
        RECT 120.105 128.925 120.305 129.095 ;
        RECT 121.025 128.965 121.195 129.545 ;
        RECT 121.370 129.075 121.720 129.725 ;
        RECT 120.970 128.925 121.195 128.965 ;
        RECT 117.870 128.465 118.275 128.635 ;
        RECT 118.445 128.465 119.230 128.635 ;
        RECT 119.505 128.185 119.715 128.715 ;
        RECT 119.975 128.400 120.305 128.925 ;
        RECT 120.815 128.840 121.195 128.925 ;
        RECT 121.890 128.905 122.120 129.895 ;
        RECT 120.475 128.185 120.645 128.795 ;
        RECT 120.815 128.405 121.145 128.840 ;
        RECT 121.455 128.735 122.120 128.905 ;
        RECT 121.455 128.445 121.625 128.735 ;
        RECT 121.795 128.185 122.125 128.565 ;
        RECT 122.295 128.445 122.480 130.565 ;
        RECT 122.720 130.275 122.985 130.735 ;
        RECT 123.155 130.140 123.405 130.565 ;
        RECT 123.615 130.290 124.720 130.460 ;
        RECT 123.100 130.010 123.405 130.140 ;
        RECT 122.650 128.815 122.930 129.765 ;
        RECT 123.100 128.905 123.270 130.010 ;
        RECT 123.440 129.225 123.680 129.820 ;
        RECT 123.850 129.755 124.380 130.120 ;
        RECT 123.850 129.055 124.020 129.755 ;
        RECT 124.550 129.675 124.720 130.290 ;
        RECT 124.890 129.935 125.060 130.735 ;
        RECT 125.230 130.235 125.480 130.565 ;
        RECT 125.705 130.265 126.590 130.435 ;
        RECT 124.550 129.585 125.060 129.675 ;
        RECT 123.100 128.775 123.325 128.905 ;
        RECT 123.495 128.835 124.020 129.055 ;
        RECT 124.190 129.415 125.060 129.585 ;
        RECT 122.735 128.185 122.985 128.645 ;
        RECT 123.155 128.635 123.325 128.775 ;
        RECT 124.190 128.635 124.360 129.415 ;
        RECT 124.890 129.345 125.060 129.415 ;
        RECT 124.570 129.165 124.770 129.195 ;
        RECT 125.230 129.165 125.400 130.235 ;
        RECT 125.570 129.345 125.760 130.065 ;
        RECT 124.570 128.865 125.400 129.165 ;
        RECT 125.930 129.135 126.250 130.095 ;
        RECT 123.155 128.465 123.490 128.635 ;
        RECT 123.685 128.465 124.360 128.635 ;
        RECT 124.680 128.185 125.050 128.685 ;
        RECT 125.230 128.635 125.400 128.865 ;
        RECT 125.785 128.805 126.250 129.135 ;
        RECT 126.420 129.425 126.590 130.265 ;
        RECT 126.770 130.235 127.085 130.735 ;
        RECT 127.315 130.005 127.655 130.565 ;
        RECT 126.760 129.630 127.655 130.005 ;
        RECT 127.825 129.725 127.995 130.735 ;
        RECT 127.465 129.425 127.655 129.630 ;
        RECT 128.165 129.675 128.495 130.520 ;
        RECT 128.165 129.595 128.555 129.675 ;
        RECT 128.725 129.645 130.395 130.735 ;
        RECT 130.655 130.115 130.825 130.545 ;
        RECT 130.995 130.285 131.325 130.735 ;
        RECT 130.655 129.885 131.330 130.115 ;
        RECT 128.340 129.545 128.555 129.595 ;
        RECT 126.420 129.095 127.295 129.425 ;
        RECT 127.465 129.095 128.215 129.425 ;
        RECT 126.420 128.635 126.590 129.095 ;
        RECT 127.465 128.925 127.665 129.095 ;
        RECT 128.385 128.965 128.555 129.545 ;
        RECT 128.330 128.925 128.555 128.965 ;
        RECT 125.230 128.465 125.635 128.635 ;
        RECT 125.805 128.465 126.590 128.635 ;
        RECT 126.865 128.185 127.075 128.715 ;
        RECT 127.335 128.400 127.665 128.925 ;
        RECT 128.175 128.840 128.555 128.925 ;
        RECT 128.725 128.955 129.475 129.475 ;
        RECT 129.645 129.125 130.395 129.645 ;
        RECT 127.835 128.185 128.005 128.795 ;
        RECT 128.175 128.405 128.505 128.840 ;
        RECT 128.725 128.185 130.395 128.955 ;
        RECT 130.625 128.865 130.925 129.715 ;
        RECT 131.095 129.235 131.330 129.885 ;
        RECT 131.500 129.575 131.785 130.520 ;
        RECT 131.965 130.265 132.650 130.735 ;
        RECT 131.960 129.745 132.655 130.055 ;
        RECT 132.830 129.680 133.135 130.465 ;
        RECT 131.500 129.425 132.360 129.575 ;
        RECT 131.500 129.405 132.785 129.425 ;
        RECT 131.095 128.905 131.630 129.235 ;
        RECT 131.800 129.045 132.785 129.405 ;
        RECT 131.095 128.755 131.315 128.905 ;
        RECT 130.570 128.185 130.905 128.690 ;
        RECT 131.075 128.380 131.315 128.755 ;
        RECT 131.800 128.710 131.970 129.045 ;
        RECT 132.960 128.875 133.135 129.680 ;
        RECT 133.325 129.570 133.615 130.735 ;
        RECT 133.790 129.785 134.055 130.555 ;
        RECT 134.225 130.015 134.555 130.735 ;
        RECT 134.745 130.195 135.005 130.555 ;
        RECT 135.175 130.365 135.505 130.735 ;
        RECT 135.675 130.195 135.935 130.555 ;
        RECT 134.745 129.965 135.935 130.195 ;
        RECT 136.505 129.785 136.795 130.555 ;
        RECT 137.555 130.065 137.725 130.565 ;
        RECT 137.895 130.235 138.225 130.735 ;
        RECT 137.555 129.895 138.220 130.065 ;
        RECT 131.595 128.515 131.970 128.710 ;
        RECT 131.595 128.370 131.765 128.515 ;
        RECT 132.330 128.185 132.725 128.680 ;
        RECT 132.895 128.355 133.135 128.875 ;
        RECT 133.325 128.185 133.615 128.910 ;
        RECT 133.790 128.365 134.125 129.785 ;
        RECT 134.300 129.605 136.795 129.785 ;
        RECT 134.300 128.915 134.525 129.605 ;
        RECT 134.725 129.095 135.005 129.425 ;
        RECT 135.185 129.095 135.760 129.425 ;
        RECT 135.940 129.095 136.375 129.425 ;
        RECT 136.555 129.095 136.825 129.425 ;
        RECT 137.470 129.075 137.820 129.725 ;
        RECT 134.300 128.725 136.785 128.915 ;
        RECT 137.990 128.905 138.220 129.895 ;
        RECT 134.305 128.185 135.050 128.555 ;
        RECT 135.615 128.365 135.870 128.725 ;
        RECT 136.050 128.185 136.380 128.555 ;
        RECT 136.560 128.365 136.785 128.725 ;
        RECT 137.555 128.735 138.220 128.905 ;
        RECT 137.555 128.445 137.725 128.735 ;
        RECT 137.895 128.185 138.225 128.565 ;
        RECT 138.395 128.445 138.580 130.565 ;
        RECT 138.820 130.275 139.085 130.735 ;
        RECT 139.255 130.140 139.505 130.565 ;
        RECT 139.715 130.290 140.820 130.460 ;
        RECT 139.200 130.010 139.505 130.140 ;
        RECT 138.750 128.815 139.030 129.765 ;
        RECT 139.200 128.905 139.370 130.010 ;
        RECT 139.540 129.225 139.780 129.820 ;
        RECT 139.950 129.755 140.480 130.120 ;
        RECT 139.950 129.055 140.120 129.755 ;
        RECT 140.650 129.675 140.820 130.290 ;
        RECT 140.990 129.935 141.160 130.735 ;
        RECT 141.330 130.235 141.580 130.565 ;
        RECT 141.805 130.265 142.690 130.435 ;
        RECT 140.650 129.585 141.160 129.675 ;
        RECT 139.200 128.775 139.425 128.905 ;
        RECT 139.595 128.835 140.120 129.055 ;
        RECT 140.290 129.415 141.160 129.585 ;
        RECT 138.835 128.185 139.085 128.645 ;
        RECT 139.255 128.635 139.425 128.775 ;
        RECT 140.290 128.635 140.460 129.415 ;
        RECT 140.990 129.345 141.160 129.415 ;
        RECT 140.670 129.165 140.870 129.195 ;
        RECT 141.330 129.165 141.500 130.235 ;
        RECT 141.670 129.345 141.860 130.065 ;
        RECT 140.670 128.865 141.500 129.165 ;
        RECT 142.030 129.135 142.350 130.095 ;
        RECT 139.255 128.465 139.590 128.635 ;
        RECT 139.785 128.465 140.460 128.635 ;
        RECT 140.780 128.185 141.150 128.685 ;
        RECT 141.330 128.635 141.500 128.865 ;
        RECT 141.885 128.805 142.350 129.135 ;
        RECT 142.520 129.425 142.690 130.265 ;
        RECT 142.870 130.235 143.185 130.735 ;
        RECT 143.415 130.005 143.755 130.565 ;
        RECT 142.860 129.630 143.755 130.005 ;
        RECT 143.925 129.725 144.095 130.735 ;
        RECT 143.565 129.425 143.755 129.630 ;
        RECT 144.265 129.675 144.595 130.520 ;
        RECT 144.265 129.595 144.655 129.675 ;
        RECT 144.440 129.545 144.655 129.595 ;
        RECT 142.520 129.095 143.395 129.425 ;
        RECT 143.565 129.095 144.315 129.425 ;
        RECT 142.520 128.635 142.690 129.095 ;
        RECT 143.565 128.925 143.765 129.095 ;
        RECT 144.485 128.965 144.655 129.545 ;
        RECT 145.745 129.645 146.955 130.735 ;
        RECT 145.745 129.105 146.265 129.645 ;
        RECT 144.430 128.925 144.655 128.965 ;
        RECT 146.435 128.935 146.955 129.475 ;
        RECT 141.330 128.465 141.735 128.635 ;
        RECT 141.905 128.465 142.690 128.635 ;
        RECT 142.965 128.185 143.175 128.715 ;
        RECT 143.435 128.400 143.765 128.925 ;
        RECT 144.275 128.840 144.655 128.925 ;
        RECT 143.935 128.185 144.105 128.795 ;
        RECT 144.275 128.405 144.605 128.840 ;
        RECT 145.745 128.185 146.955 128.935 ;
        RECT 17.320 128.015 147.040 128.185 ;
        RECT 17.405 127.265 18.615 128.015 ;
        RECT 17.405 126.725 17.925 127.265 ;
        RECT 18.790 127.175 19.050 128.015 ;
        RECT 19.225 127.270 19.480 127.845 ;
        RECT 19.650 127.635 19.980 128.015 ;
        RECT 20.195 127.465 20.365 127.845 ;
        RECT 19.650 127.295 20.365 127.465 ;
        RECT 20.715 127.465 20.885 127.845 ;
        RECT 21.065 127.635 21.395 128.015 ;
        RECT 20.715 127.295 21.380 127.465 ;
        RECT 21.575 127.340 21.835 127.845 ;
        RECT 18.095 126.555 18.615 127.095 ;
        RECT 17.405 125.465 18.615 126.555 ;
        RECT 18.790 125.465 19.050 126.615 ;
        RECT 19.225 126.540 19.395 127.270 ;
        RECT 19.650 127.105 19.820 127.295 ;
        RECT 19.565 126.775 19.820 127.105 ;
        RECT 19.650 126.565 19.820 126.775 ;
        RECT 20.100 126.745 20.455 127.115 ;
        RECT 20.645 126.745 20.985 127.115 ;
        RECT 21.210 127.040 21.380 127.295 ;
        RECT 21.210 126.710 21.485 127.040 ;
        RECT 21.210 126.565 21.380 126.710 ;
        RECT 19.225 125.635 19.480 126.540 ;
        RECT 19.650 126.395 20.365 126.565 ;
        RECT 19.650 125.465 19.980 126.225 ;
        RECT 20.195 125.635 20.365 126.395 ;
        RECT 20.705 126.395 21.380 126.565 ;
        RECT 21.655 126.540 21.835 127.340 ;
        RECT 22.005 127.245 24.595 128.015 ;
        RECT 24.855 127.465 25.025 127.755 ;
        RECT 25.195 127.635 25.525 128.015 ;
        RECT 24.855 127.295 25.520 127.465 ;
        RECT 22.005 126.725 23.215 127.245 ;
        RECT 23.385 126.555 24.595 127.075 ;
        RECT 20.705 125.635 20.885 126.395 ;
        RECT 21.065 125.465 21.395 126.225 ;
        RECT 21.565 125.635 21.835 126.540 ;
        RECT 22.005 125.465 24.595 126.555 ;
        RECT 24.770 126.475 25.120 127.125 ;
        RECT 25.290 126.305 25.520 127.295 ;
        RECT 24.855 126.135 25.520 126.305 ;
        RECT 24.855 125.635 25.025 126.135 ;
        RECT 25.195 125.465 25.525 125.965 ;
        RECT 25.695 125.635 25.880 127.755 ;
        RECT 26.135 127.555 26.385 128.015 ;
        RECT 26.555 127.565 26.890 127.735 ;
        RECT 27.085 127.565 27.760 127.735 ;
        RECT 26.555 127.425 26.725 127.565 ;
        RECT 26.050 126.435 26.330 127.385 ;
        RECT 26.500 127.295 26.725 127.425 ;
        RECT 26.500 126.190 26.670 127.295 ;
        RECT 26.895 127.145 27.420 127.365 ;
        RECT 26.840 126.380 27.080 126.975 ;
        RECT 27.250 126.445 27.420 127.145 ;
        RECT 27.590 126.785 27.760 127.565 ;
        RECT 28.080 127.515 28.450 128.015 ;
        RECT 28.630 127.565 29.035 127.735 ;
        RECT 29.205 127.565 29.990 127.735 ;
        RECT 28.630 127.335 28.800 127.565 ;
        RECT 27.970 127.035 28.800 127.335 ;
        RECT 29.185 127.065 29.650 127.395 ;
        RECT 27.970 127.005 28.170 127.035 ;
        RECT 28.290 126.785 28.460 126.855 ;
        RECT 27.590 126.615 28.460 126.785 ;
        RECT 27.950 126.525 28.460 126.615 ;
        RECT 26.500 126.060 26.805 126.190 ;
        RECT 27.250 126.080 27.780 126.445 ;
        RECT 26.120 125.465 26.385 125.925 ;
        RECT 26.555 125.635 26.805 126.060 ;
        RECT 27.950 125.910 28.120 126.525 ;
        RECT 27.015 125.740 28.120 125.910 ;
        RECT 28.290 125.465 28.460 126.265 ;
        RECT 28.630 125.965 28.800 127.035 ;
        RECT 28.970 126.135 29.160 126.855 ;
        RECT 29.330 126.105 29.650 127.065 ;
        RECT 29.820 127.105 29.990 127.565 ;
        RECT 30.265 127.485 30.475 128.015 ;
        RECT 30.735 127.275 31.065 127.800 ;
        RECT 31.235 127.405 31.405 128.015 ;
        RECT 31.575 127.360 31.905 127.795 ;
        RECT 31.575 127.275 31.955 127.360 ;
        RECT 30.865 127.105 31.065 127.275 ;
        RECT 31.730 127.235 31.955 127.275 ;
        RECT 29.820 126.775 30.695 127.105 ;
        RECT 30.865 126.775 31.615 127.105 ;
        RECT 28.630 125.635 28.880 125.965 ;
        RECT 29.820 125.935 29.990 126.775 ;
        RECT 30.865 126.570 31.055 126.775 ;
        RECT 31.785 126.655 31.955 127.235 ;
        RECT 32.165 127.195 32.395 128.015 ;
        RECT 32.565 127.215 32.895 127.845 ;
        RECT 32.145 126.775 32.475 127.025 ;
        RECT 31.740 126.605 31.955 126.655 ;
        RECT 32.645 126.615 32.895 127.215 ;
        RECT 33.065 127.195 33.275 128.015 ;
        RECT 33.505 127.470 38.850 128.015 ;
        RECT 35.090 126.640 35.430 127.470 ;
        RECT 39.025 127.245 42.535 128.015 ;
        RECT 43.165 127.290 43.455 128.015 ;
        RECT 43.625 127.470 48.970 128.015 ;
        RECT 49.145 127.470 54.490 128.015 ;
        RECT 54.665 127.470 60.010 128.015 ;
        RECT 30.160 126.195 31.055 126.570 ;
        RECT 31.565 126.525 31.955 126.605 ;
        RECT 29.105 125.765 29.990 125.935 ;
        RECT 30.170 125.465 30.485 125.965 ;
        RECT 30.715 125.635 31.055 126.195 ;
        RECT 31.225 125.465 31.395 126.475 ;
        RECT 31.565 125.680 31.895 126.525 ;
        RECT 32.165 125.465 32.395 126.605 ;
        RECT 32.565 125.635 32.895 126.615 ;
        RECT 33.065 125.465 33.275 126.605 ;
        RECT 36.910 125.900 37.260 127.150 ;
        RECT 39.025 126.725 40.675 127.245 ;
        RECT 40.845 126.555 42.535 127.075 ;
        RECT 45.210 126.640 45.550 127.470 ;
        RECT 33.505 125.465 38.850 125.900 ;
        RECT 39.025 125.465 42.535 126.555 ;
        RECT 43.165 125.465 43.455 126.630 ;
        RECT 47.030 125.900 47.380 127.150 ;
        RECT 50.730 126.640 51.070 127.470 ;
        RECT 52.550 125.900 52.900 127.150 ;
        RECT 56.250 126.640 56.590 127.470 ;
        RECT 60.185 127.245 63.695 128.015 ;
        RECT 63.865 127.265 65.075 128.015 ;
        RECT 58.070 125.900 58.420 127.150 ;
        RECT 60.185 126.725 61.835 127.245 ;
        RECT 62.005 126.555 63.695 127.075 ;
        RECT 63.865 126.725 64.385 127.265 ;
        RECT 65.255 127.205 65.525 128.015 ;
        RECT 65.695 127.205 66.025 127.845 ;
        RECT 66.195 127.205 66.435 128.015 ;
        RECT 66.660 127.275 67.275 127.845 ;
        RECT 67.445 127.505 67.660 128.015 ;
        RECT 67.890 127.505 68.170 127.835 ;
        RECT 68.350 127.505 68.590 128.015 ;
        RECT 64.555 126.555 65.075 127.095 ;
        RECT 65.245 126.775 65.595 127.025 ;
        RECT 65.765 126.605 65.935 127.205 ;
        RECT 66.105 126.775 66.455 127.025 ;
        RECT 43.625 125.465 48.970 125.900 ;
        RECT 49.145 125.465 54.490 125.900 ;
        RECT 54.665 125.465 60.010 125.900 ;
        RECT 60.185 125.465 63.695 126.555 ;
        RECT 63.865 125.465 65.075 126.555 ;
        RECT 65.255 125.465 65.585 126.605 ;
        RECT 65.765 126.435 66.445 126.605 ;
        RECT 66.115 125.650 66.445 126.435 ;
        RECT 66.660 126.255 66.975 127.275 ;
        RECT 67.145 126.605 67.315 127.105 ;
        RECT 67.565 126.775 67.830 127.335 ;
        RECT 68.000 126.605 68.170 127.505 ;
        RECT 68.340 126.775 68.695 127.335 ;
        RECT 68.925 127.290 69.215 128.015 ;
        RECT 69.475 127.465 69.645 127.755 ;
        RECT 69.815 127.635 70.145 128.015 ;
        RECT 69.475 127.295 70.140 127.465 ;
        RECT 67.145 126.435 68.570 126.605 ;
        RECT 66.660 125.635 67.195 126.255 ;
        RECT 67.365 125.465 67.695 126.265 ;
        RECT 68.180 126.260 68.570 126.435 ;
        RECT 68.925 125.465 69.215 126.630 ;
        RECT 69.390 126.475 69.740 127.125 ;
        RECT 69.910 126.305 70.140 127.295 ;
        RECT 69.475 126.135 70.140 126.305 ;
        RECT 69.475 125.635 69.645 126.135 ;
        RECT 69.815 125.465 70.145 125.965 ;
        RECT 70.315 125.635 70.500 127.755 ;
        RECT 70.755 127.555 71.005 128.015 ;
        RECT 71.175 127.565 71.510 127.735 ;
        RECT 71.705 127.565 72.380 127.735 ;
        RECT 71.175 127.425 71.345 127.565 ;
        RECT 70.670 126.435 70.950 127.385 ;
        RECT 71.120 127.295 71.345 127.425 ;
        RECT 71.120 126.190 71.290 127.295 ;
        RECT 71.515 127.145 72.040 127.365 ;
        RECT 71.460 126.380 71.700 126.975 ;
        RECT 71.870 126.445 72.040 127.145 ;
        RECT 72.210 126.785 72.380 127.565 ;
        RECT 72.700 127.515 73.070 128.015 ;
        RECT 73.250 127.565 73.655 127.735 ;
        RECT 73.825 127.565 74.610 127.735 ;
        RECT 73.250 127.335 73.420 127.565 ;
        RECT 72.590 127.035 73.420 127.335 ;
        RECT 73.805 127.065 74.270 127.395 ;
        RECT 72.590 127.005 72.790 127.035 ;
        RECT 72.910 126.785 73.080 126.855 ;
        RECT 72.210 126.615 73.080 126.785 ;
        RECT 72.570 126.525 73.080 126.615 ;
        RECT 71.120 126.060 71.425 126.190 ;
        RECT 71.870 126.080 72.400 126.445 ;
        RECT 70.740 125.465 71.005 125.925 ;
        RECT 71.175 125.635 71.425 126.060 ;
        RECT 72.570 125.910 72.740 126.525 ;
        RECT 71.635 125.740 72.740 125.910 ;
        RECT 72.910 125.465 73.080 126.265 ;
        RECT 73.250 125.965 73.420 127.035 ;
        RECT 73.590 126.135 73.780 126.855 ;
        RECT 73.950 126.105 74.270 127.065 ;
        RECT 74.440 127.105 74.610 127.565 ;
        RECT 74.885 127.485 75.095 128.015 ;
        RECT 75.355 127.275 75.685 127.800 ;
        RECT 75.855 127.405 76.025 128.015 ;
        RECT 76.195 127.360 76.525 127.795 ;
        RECT 76.195 127.275 76.575 127.360 ;
        RECT 75.485 127.105 75.685 127.275 ;
        RECT 76.350 127.235 76.575 127.275 ;
        RECT 74.440 126.775 75.315 127.105 ;
        RECT 75.485 126.775 76.235 127.105 ;
        RECT 73.250 125.635 73.500 125.965 ;
        RECT 74.440 125.935 74.610 126.775 ;
        RECT 75.485 126.570 75.675 126.775 ;
        RECT 76.405 126.655 76.575 127.235 ;
        RECT 76.745 127.215 77.440 127.845 ;
        RECT 77.645 127.215 77.955 128.015 ;
        RECT 78.125 127.265 79.335 128.015 ;
        RECT 76.765 126.775 77.100 127.025 ;
        RECT 76.360 126.605 76.575 126.655 ;
        RECT 77.270 126.615 77.440 127.215 ;
        RECT 77.610 126.775 77.945 127.045 ;
        RECT 78.125 126.725 78.645 127.265 ;
        RECT 79.505 127.195 79.765 128.015 ;
        RECT 79.935 127.195 80.265 127.615 ;
        RECT 80.445 127.445 80.705 127.845 ;
        RECT 80.875 127.615 81.205 128.015 ;
        RECT 81.375 127.445 81.545 127.795 ;
        RECT 81.715 127.615 82.090 128.015 ;
        RECT 80.445 127.275 82.110 127.445 ;
        RECT 82.280 127.340 82.555 127.685 ;
        RECT 80.015 127.105 80.265 127.195 ;
        RECT 81.940 127.105 82.110 127.275 ;
        RECT 74.780 126.195 75.675 126.570 ;
        RECT 76.185 126.525 76.575 126.605 ;
        RECT 73.725 125.765 74.610 125.935 ;
        RECT 74.790 125.465 75.105 125.965 ;
        RECT 75.335 125.635 75.675 126.195 ;
        RECT 75.845 125.465 76.015 126.475 ;
        RECT 76.185 125.680 76.515 126.525 ;
        RECT 76.745 125.465 77.005 126.605 ;
        RECT 77.175 125.635 77.505 126.615 ;
        RECT 77.675 125.465 77.955 126.605 ;
        RECT 78.815 126.555 79.335 127.095 ;
        RECT 79.510 126.775 79.845 127.025 ;
        RECT 80.015 126.775 80.730 127.105 ;
        RECT 80.945 126.775 81.770 127.105 ;
        RECT 81.940 126.775 82.215 127.105 ;
        RECT 78.125 125.465 79.335 126.555 ;
        RECT 79.505 125.465 79.765 126.605 ;
        RECT 80.015 126.215 80.185 126.775 ;
        RECT 80.445 126.315 80.775 126.605 ;
        RECT 80.945 126.485 81.190 126.775 ;
        RECT 81.940 126.605 82.110 126.775 ;
        RECT 82.385 126.605 82.555 127.340 ;
        RECT 82.725 127.195 82.985 128.015 ;
        RECT 83.155 127.195 83.485 127.615 ;
        RECT 83.665 127.445 83.925 127.845 ;
        RECT 84.095 127.615 84.425 128.015 ;
        RECT 84.595 127.445 84.765 127.795 ;
        RECT 84.935 127.615 85.310 128.015 ;
        RECT 83.665 127.275 85.330 127.445 ;
        RECT 85.500 127.340 85.775 127.685 ;
        RECT 83.235 127.105 83.485 127.195 ;
        RECT 85.160 127.105 85.330 127.275 ;
        RECT 82.730 126.775 83.065 127.025 ;
        RECT 83.235 126.775 83.950 127.105 ;
        RECT 84.165 126.775 84.990 127.105 ;
        RECT 85.160 126.775 85.435 127.105 ;
        RECT 81.450 126.435 82.110 126.605 ;
        RECT 81.450 126.315 81.620 126.435 ;
        RECT 80.445 126.145 81.620 126.315 ;
        RECT 80.005 125.645 81.620 125.975 ;
        RECT 81.790 125.465 82.070 126.265 ;
        RECT 82.280 125.635 82.555 126.605 ;
        RECT 82.725 125.465 82.985 126.605 ;
        RECT 83.235 126.215 83.405 126.775 ;
        RECT 83.665 126.315 83.995 126.605 ;
        RECT 84.165 126.485 84.410 126.775 ;
        RECT 85.160 126.605 85.330 126.775 ;
        RECT 85.605 126.605 85.775 127.340 ;
        RECT 86.955 127.465 87.125 127.755 ;
        RECT 87.295 127.635 87.625 128.015 ;
        RECT 86.955 127.295 87.620 127.465 ;
        RECT 84.670 126.435 85.330 126.605 ;
        RECT 84.670 126.315 84.840 126.435 ;
        RECT 83.665 126.145 84.840 126.315 ;
        RECT 83.225 125.645 84.840 125.975 ;
        RECT 85.010 125.465 85.290 126.265 ;
        RECT 85.500 125.635 85.775 126.605 ;
        RECT 86.870 126.475 87.220 127.125 ;
        RECT 87.390 126.305 87.620 127.295 ;
        RECT 86.955 126.135 87.620 126.305 ;
        RECT 86.955 125.635 87.125 126.135 ;
        RECT 87.295 125.465 87.625 125.965 ;
        RECT 87.795 125.635 87.980 127.755 ;
        RECT 88.235 127.555 88.485 128.015 ;
        RECT 88.655 127.565 88.990 127.735 ;
        RECT 89.185 127.565 89.860 127.735 ;
        RECT 88.655 127.425 88.825 127.565 ;
        RECT 88.150 126.435 88.430 127.385 ;
        RECT 88.600 127.295 88.825 127.425 ;
        RECT 88.600 126.190 88.770 127.295 ;
        RECT 88.995 127.145 89.520 127.365 ;
        RECT 88.940 126.380 89.180 126.975 ;
        RECT 89.350 126.445 89.520 127.145 ;
        RECT 89.690 126.785 89.860 127.565 ;
        RECT 90.180 127.515 90.550 128.015 ;
        RECT 90.730 127.565 91.135 127.735 ;
        RECT 91.305 127.565 92.090 127.735 ;
        RECT 90.730 127.335 90.900 127.565 ;
        RECT 90.070 127.035 90.900 127.335 ;
        RECT 91.285 127.065 91.750 127.395 ;
        RECT 90.070 127.005 90.270 127.035 ;
        RECT 90.390 126.785 90.560 126.855 ;
        RECT 89.690 126.615 90.560 126.785 ;
        RECT 90.050 126.525 90.560 126.615 ;
        RECT 88.600 126.060 88.905 126.190 ;
        RECT 89.350 126.080 89.880 126.445 ;
        RECT 88.220 125.465 88.485 125.925 ;
        RECT 88.655 125.635 88.905 126.060 ;
        RECT 90.050 125.910 90.220 126.525 ;
        RECT 89.115 125.740 90.220 125.910 ;
        RECT 90.390 125.465 90.560 126.265 ;
        RECT 90.730 125.965 90.900 127.035 ;
        RECT 91.070 126.135 91.260 126.855 ;
        RECT 91.430 126.105 91.750 127.065 ;
        RECT 91.920 127.105 92.090 127.565 ;
        RECT 92.365 127.485 92.575 128.015 ;
        RECT 92.835 127.275 93.165 127.800 ;
        RECT 93.335 127.405 93.505 128.015 ;
        RECT 93.675 127.360 94.005 127.795 ;
        RECT 94.175 127.500 94.345 128.015 ;
        RECT 93.675 127.275 94.055 127.360 ;
        RECT 94.685 127.290 94.975 128.015 ;
        RECT 92.965 127.105 93.165 127.275 ;
        RECT 93.830 127.235 94.055 127.275 ;
        RECT 91.920 126.775 92.795 127.105 ;
        RECT 92.965 126.775 93.715 127.105 ;
        RECT 90.730 125.635 90.980 125.965 ;
        RECT 91.920 125.935 92.090 126.775 ;
        RECT 92.965 126.570 93.155 126.775 ;
        RECT 93.885 126.655 94.055 127.235 ;
        RECT 95.145 127.245 98.655 128.015 ;
        RECT 99.795 127.360 100.125 127.795 ;
        RECT 100.295 127.405 100.465 128.015 ;
        RECT 99.745 127.275 100.125 127.360 ;
        RECT 100.635 127.275 100.965 127.800 ;
        RECT 101.225 127.485 101.435 128.015 ;
        RECT 101.710 127.565 102.495 127.735 ;
        RECT 102.665 127.565 103.070 127.735 ;
        RECT 95.145 126.725 96.795 127.245 ;
        RECT 99.745 127.235 99.970 127.275 ;
        RECT 93.840 126.605 94.055 126.655 ;
        RECT 92.260 126.195 93.155 126.570 ;
        RECT 93.665 126.525 94.055 126.605 ;
        RECT 91.205 125.765 92.090 125.935 ;
        RECT 92.270 125.465 92.585 125.965 ;
        RECT 92.815 125.635 93.155 126.195 ;
        RECT 93.325 125.465 93.495 126.475 ;
        RECT 93.665 125.680 93.995 126.525 ;
        RECT 94.165 125.465 94.335 126.380 ;
        RECT 94.685 125.465 94.975 126.630 ;
        RECT 96.965 126.555 98.655 127.075 ;
        RECT 95.145 125.465 98.655 126.555 ;
        RECT 99.745 126.655 99.915 127.235 ;
        RECT 100.635 127.105 100.835 127.275 ;
        RECT 101.710 127.105 101.880 127.565 ;
        RECT 100.085 126.775 100.835 127.105 ;
        RECT 101.005 126.775 101.880 127.105 ;
        RECT 99.745 126.605 99.960 126.655 ;
        RECT 99.745 126.525 100.135 126.605 ;
        RECT 99.805 125.680 100.135 126.525 ;
        RECT 100.645 126.570 100.835 126.775 ;
        RECT 100.305 125.465 100.475 126.475 ;
        RECT 100.645 126.195 101.540 126.570 ;
        RECT 100.645 125.635 100.985 126.195 ;
        RECT 101.215 125.465 101.530 125.965 ;
        RECT 101.710 125.935 101.880 126.775 ;
        RECT 102.050 127.065 102.515 127.395 ;
        RECT 102.900 127.335 103.070 127.565 ;
        RECT 103.250 127.515 103.620 128.015 ;
        RECT 103.940 127.565 104.615 127.735 ;
        RECT 104.810 127.565 105.145 127.735 ;
        RECT 102.050 126.105 102.370 127.065 ;
        RECT 102.900 127.035 103.730 127.335 ;
        RECT 102.540 126.135 102.730 126.855 ;
        RECT 102.900 125.965 103.070 127.035 ;
        RECT 103.530 127.005 103.730 127.035 ;
        RECT 103.240 126.785 103.410 126.855 ;
        RECT 103.940 126.785 104.110 127.565 ;
        RECT 104.975 127.425 105.145 127.565 ;
        RECT 105.315 127.555 105.565 128.015 ;
        RECT 103.240 126.615 104.110 126.785 ;
        RECT 104.280 127.145 104.805 127.365 ;
        RECT 104.975 127.295 105.200 127.425 ;
        RECT 103.240 126.525 103.750 126.615 ;
        RECT 101.710 125.765 102.595 125.935 ;
        RECT 102.820 125.635 103.070 125.965 ;
        RECT 103.240 125.465 103.410 126.265 ;
        RECT 103.580 125.910 103.750 126.525 ;
        RECT 104.280 126.445 104.450 127.145 ;
        RECT 103.920 126.080 104.450 126.445 ;
        RECT 104.620 126.380 104.860 126.975 ;
        RECT 105.030 126.190 105.200 127.295 ;
        RECT 105.370 126.435 105.650 127.385 ;
        RECT 104.895 126.060 105.200 126.190 ;
        RECT 103.580 125.740 104.685 125.910 ;
        RECT 104.895 125.635 105.145 126.060 ;
        RECT 105.315 125.465 105.580 125.925 ;
        RECT 105.820 125.635 106.005 127.755 ;
        RECT 106.175 127.635 106.505 128.015 ;
        RECT 106.675 127.465 106.845 127.755 ;
        RECT 106.180 127.295 106.845 127.465 ;
        RECT 107.195 127.465 107.365 127.755 ;
        RECT 107.535 127.635 107.865 128.015 ;
        RECT 107.195 127.295 107.860 127.465 ;
        RECT 106.180 126.305 106.410 127.295 ;
        RECT 106.580 126.475 106.930 127.125 ;
        RECT 107.110 126.475 107.460 127.125 ;
        RECT 107.630 126.305 107.860 127.295 ;
        RECT 106.180 126.135 106.845 126.305 ;
        RECT 106.175 125.465 106.505 125.965 ;
        RECT 106.675 125.635 106.845 126.135 ;
        RECT 107.195 126.135 107.860 126.305 ;
        RECT 107.195 125.635 107.365 126.135 ;
        RECT 107.535 125.465 107.865 125.965 ;
        RECT 108.035 125.635 108.220 127.755 ;
        RECT 108.475 127.555 108.725 128.015 ;
        RECT 108.895 127.565 109.230 127.735 ;
        RECT 109.425 127.565 110.100 127.735 ;
        RECT 108.895 127.425 109.065 127.565 ;
        RECT 108.390 126.435 108.670 127.385 ;
        RECT 108.840 127.295 109.065 127.425 ;
        RECT 108.840 126.190 109.010 127.295 ;
        RECT 109.235 127.145 109.760 127.365 ;
        RECT 109.180 126.380 109.420 126.975 ;
        RECT 109.590 126.445 109.760 127.145 ;
        RECT 109.930 126.785 110.100 127.565 ;
        RECT 110.420 127.515 110.790 128.015 ;
        RECT 110.970 127.565 111.375 127.735 ;
        RECT 111.545 127.565 112.330 127.735 ;
        RECT 110.970 127.335 111.140 127.565 ;
        RECT 110.310 127.035 111.140 127.335 ;
        RECT 111.525 127.065 111.990 127.395 ;
        RECT 110.310 127.005 110.510 127.035 ;
        RECT 110.630 126.785 110.800 126.855 ;
        RECT 109.930 126.615 110.800 126.785 ;
        RECT 110.290 126.525 110.800 126.615 ;
        RECT 108.840 126.060 109.145 126.190 ;
        RECT 109.590 126.080 110.120 126.445 ;
        RECT 108.460 125.465 108.725 125.925 ;
        RECT 108.895 125.635 109.145 126.060 ;
        RECT 110.290 125.910 110.460 126.525 ;
        RECT 109.355 125.740 110.460 125.910 ;
        RECT 110.630 125.465 110.800 126.265 ;
        RECT 110.970 125.965 111.140 127.035 ;
        RECT 111.310 126.135 111.500 126.855 ;
        RECT 111.670 126.105 111.990 127.065 ;
        RECT 112.160 127.105 112.330 127.565 ;
        RECT 112.605 127.485 112.815 128.015 ;
        RECT 113.075 127.275 113.405 127.800 ;
        RECT 113.575 127.405 113.745 128.015 ;
        RECT 113.915 127.360 114.245 127.795 ;
        RECT 113.915 127.275 114.295 127.360 ;
        RECT 113.205 127.105 113.405 127.275 ;
        RECT 114.070 127.235 114.295 127.275 ;
        RECT 112.160 126.775 113.035 127.105 ;
        RECT 113.205 126.775 113.955 127.105 ;
        RECT 110.970 125.635 111.220 125.965 ;
        RECT 112.160 125.935 112.330 126.775 ;
        RECT 113.205 126.570 113.395 126.775 ;
        RECT 114.125 126.655 114.295 127.235 ;
        RECT 114.465 127.245 116.135 128.015 ;
        RECT 114.465 126.725 115.215 127.245 ;
        RECT 114.080 126.605 114.295 126.655 ;
        RECT 112.500 126.195 113.395 126.570 ;
        RECT 113.905 126.525 114.295 126.605 ;
        RECT 115.385 126.555 116.135 127.075 ;
        RECT 111.445 125.765 112.330 125.935 ;
        RECT 112.510 125.465 112.825 125.965 ;
        RECT 113.055 125.635 113.395 126.195 ;
        RECT 113.565 125.465 113.735 126.475 ;
        RECT 113.905 125.680 114.235 126.525 ;
        RECT 114.465 125.465 116.135 126.555 ;
        RECT 116.765 127.070 117.105 127.845 ;
        RECT 117.275 127.555 117.445 128.015 ;
        RECT 117.685 127.580 118.045 127.845 ;
        RECT 117.685 127.575 118.040 127.580 ;
        RECT 117.685 127.565 118.035 127.575 ;
        RECT 117.685 127.560 118.030 127.565 ;
        RECT 117.685 127.550 118.025 127.560 ;
        RECT 118.675 127.555 118.845 128.015 ;
        RECT 117.685 127.545 118.020 127.550 ;
        RECT 117.685 127.535 118.010 127.545 ;
        RECT 117.685 127.525 118.000 127.535 ;
        RECT 117.685 127.385 117.985 127.525 ;
        RECT 117.275 127.195 117.985 127.385 ;
        RECT 118.175 127.385 118.505 127.465 ;
        RECT 119.015 127.385 119.355 127.845 ;
        RECT 118.175 127.195 119.355 127.385 ;
        RECT 120.445 127.290 120.735 128.015 ;
        RECT 120.905 127.275 121.290 127.845 ;
        RECT 121.460 127.555 121.785 128.015 ;
        RECT 122.305 127.385 122.585 127.845 ;
        RECT 116.765 125.635 117.045 127.070 ;
        RECT 117.275 126.625 117.560 127.195 ;
        RECT 117.745 126.795 118.215 127.025 ;
        RECT 118.385 127.005 118.715 127.025 ;
        RECT 118.385 126.825 118.835 127.005 ;
        RECT 119.025 126.825 119.355 127.025 ;
        RECT 117.275 126.410 118.425 126.625 ;
        RECT 117.215 125.465 117.925 126.240 ;
        RECT 118.095 125.635 118.425 126.410 ;
        RECT 118.620 125.710 118.835 126.825 ;
        RECT 119.125 126.485 119.355 126.825 ;
        RECT 119.015 125.465 119.345 126.185 ;
        RECT 120.445 125.465 120.735 126.630 ;
        RECT 120.905 126.605 121.185 127.275 ;
        RECT 121.460 127.215 122.585 127.385 ;
        RECT 121.460 127.105 121.910 127.215 ;
        RECT 121.355 126.775 121.910 127.105 ;
        RECT 122.775 127.045 123.175 127.845 ;
        RECT 123.575 127.555 123.845 128.015 ;
        RECT 124.015 127.385 124.300 127.845 ;
        RECT 120.905 125.635 121.290 126.605 ;
        RECT 121.460 126.315 121.910 126.775 ;
        RECT 122.080 126.485 123.175 127.045 ;
        RECT 121.460 126.095 122.585 126.315 ;
        RECT 121.460 125.465 121.785 125.925 ;
        RECT 122.305 125.635 122.585 126.095 ;
        RECT 122.775 125.635 123.175 126.485 ;
        RECT 123.345 127.215 124.300 127.385 ;
        RECT 124.585 127.275 124.970 127.845 ;
        RECT 125.140 127.555 125.465 128.015 ;
        RECT 125.985 127.385 126.265 127.845 ;
        RECT 123.345 126.315 123.555 127.215 ;
        RECT 123.725 126.485 124.415 127.045 ;
        RECT 124.585 126.605 124.865 127.275 ;
        RECT 125.140 127.215 126.265 127.385 ;
        RECT 125.140 127.105 125.590 127.215 ;
        RECT 125.035 126.775 125.590 127.105 ;
        RECT 126.455 127.045 126.855 127.845 ;
        RECT 127.255 127.555 127.525 128.015 ;
        RECT 127.695 127.385 127.980 127.845 ;
        RECT 123.345 126.095 124.300 126.315 ;
        RECT 123.575 125.465 123.845 125.925 ;
        RECT 124.015 125.635 124.300 126.095 ;
        RECT 124.585 125.635 124.970 126.605 ;
        RECT 125.140 126.315 125.590 126.775 ;
        RECT 125.760 126.485 126.855 127.045 ;
        RECT 125.140 126.095 126.265 126.315 ;
        RECT 125.140 125.465 125.465 125.925 ;
        RECT 125.985 125.635 126.265 126.095 ;
        RECT 126.455 125.635 126.855 126.485 ;
        RECT 127.025 127.215 127.980 127.385 ;
        RECT 127.025 126.315 127.235 127.215 ;
        RECT 127.405 126.485 128.095 127.045 ;
        RECT 128.730 126.415 129.065 127.835 ;
        RECT 129.245 127.645 129.990 128.015 ;
        RECT 130.555 127.475 130.810 127.835 ;
        RECT 130.990 127.645 131.320 128.015 ;
        RECT 131.500 127.475 131.725 127.835 ;
        RECT 129.240 127.285 131.725 127.475 ;
        RECT 129.240 126.595 129.465 127.285 ;
        RECT 132.220 127.205 132.465 127.810 ;
        RECT 132.685 127.480 133.195 128.015 ;
        RECT 129.665 126.775 129.945 127.105 ;
        RECT 130.125 126.775 130.700 127.105 ;
        RECT 130.880 126.775 131.315 127.105 ;
        RECT 131.495 126.775 131.765 127.105 ;
        RECT 131.945 127.035 133.175 127.205 ;
        RECT 129.240 126.415 131.735 126.595 ;
        RECT 127.025 126.095 127.980 126.315 ;
        RECT 127.255 125.465 127.525 125.925 ;
        RECT 127.695 125.635 127.980 126.095 ;
        RECT 128.730 125.645 128.995 126.415 ;
        RECT 129.165 125.465 129.495 126.185 ;
        RECT 129.685 126.005 130.875 126.235 ;
        RECT 129.685 125.645 129.945 126.005 ;
        RECT 130.115 125.465 130.445 125.835 ;
        RECT 130.615 125.645 130.875 126.005 ;
        RECT 131.445 125.645 131.735 126.415 ;
        RECT 131.945 126.225 132.285 127.035 ;
        RECT 132.455 126.470 133.205 126.660 ;
        RECT 131.945 125.815 132.460 126.225 ;
        RECT 132.695 125.465 132.865 126.225 ;
        RECT 133.035 125.805 133.205 126.470 ;
        RECT 133.375 126.485 133.565 127.845 ;
        RECT 133.735 126.995 134.010 127.845 ;
        RECT 134.200 127.480 134.730 127.845 ;
        RECT 135.155 127.615 135.485 128.015 ;
        RECT 134.555 127.445 134.730 127.480 ;
        RECT 133.735 126.825 134.015 126.995 ;
        RECT 133.735 126.685 134.010 126.825 ;
        RECT 134.215 126.485 134.385 127.285 ;
        RECT 133.375 126.315 134.385 126.485 ;
        RECT 134.555 127.275 135.485 127.445 ;
        RECT 135.655 127.275 135.910 127.845 ;
        RECT 136.175 127.465 136.345 127.755 ;
        RECT 136.515 127.635 136.845 128.015 ;
        RECT 136.175 127.295 136.840 127.465 ;
        RECT 134.555 126.145 134.725 127.275 ;
        RECT 135.315 127.105 135.485 127.275 ;
        RECT 133.600 125.975 134.725 126.145 ;
        RECT 134.895 126.775 135.090 127.105 ;
        RECT 135.315 126.775 135.570 127.105 ;
        RECT 134.895 125.805 135.065 126.775 ;
        RECT 135.740 126.605 135.910 127.275 ;
        RECT 133.035 125.635 135.065 125.805 ;
        RECT 135.235 125.465 135.405 126.605 ;
        RECT 135.575 125.635 135.910 126.605 ;
        RECT 136.090 126.475 136.440 127.125 ;
        RECT 136.610 126.305 136.840 127.295 ;
        RECT 136.175 126.135 136.840 126.305 ;
        RECT 136.175 125.635 136.345 126.135 ;
        RECT 136.515 125.465 136.845 125.965 ;
        RECT 137.015 125.635 137.200 127.755 ;
        RECT 137.455 127.555 137.705 128.015 ;
        RECT 137.875 127.565 138.210 127.735 ;
        RECT 138.405 127.565 139.080 127.735 ;
        RECT 137.875 127.425 138.045 127.565 ;
        RECT 137.370 126.435 137.650 127.385 ;
        RECT 137.820 127.295 138.045 127.425 ;
        RECT 137.820 126.190 137.990 127.295 ;
        RECT 138.215 127.145 138.740 127.365 ;
        RECT 138.160 126.380 138.400 126.975 ;
        RECT 138.570 126.445 138.740 127.145 ;
        RECT 138.910 126.785 139.080 127.565 ;
        RECT 139.400 127.515 139.770 128.015 ;
        RECT 139.950 127.565 140.355 127.735 ;
        RECT 140.525 127.565 141.310 127.735 ;
        RECT 139.950 127.335 140.120 127.565 ;
        RECT 139.290 127.035 140.120 127.335 ;
        RECT 140.505 127.065 140.970 127.395 ;
        RECT 139.290 127.005 139.490 127.035 ;
        RECT 139.610 126.785 139.780 126.855 ;
        RECT 138.910 126.615 139.780 126.785 ;
        RECT 139.270 126.525 139.780 126.615 ;
        RECT 137.820 126.060 138.125 126.190 ;
        RECT 138.570 126.080 139.100 126.445 ;
        RECT 137.440 125.465 137.705 125.925 ;
        RECT 137.875 125.635 138.125 126.060 ;
        RECT 139.270 125.910 139.440 126.525 ;
        RECT 138.335 125.740 139.440 125.910 ;
        RECT 139.610 125.465 139.780 126.265 ;
        RECT 139.950 125.965 140.120 127.035 ;
        RECT 140.290 126.135 140.480 126.855 ;
        RECT 140.650 126.105 140.970 127.065 ;
        RECT 141.140 127.105 141.310 127.565 ;
        RECT 141.585 127.485 141.795 128.015 ;
        RECT 142.055 127.275 142.385 127.800 ;
        RECT 142.555 127.405 142.725 128.015 ;
        RECT 142.895 127.360 143.225 127.795 ;
        RECT 143.995 127.465 144.165 127.845 ;
        RECT 144.380 127.635 144.710 128.015 ;
        RECT 142.895 127.275 143.275 127.360 ;
        RECT 143.995 127.295 144.710 127.465 ;
        RECT 142.185 127.105 142.385 127.275 ;
        RECT 143.050 127.235 143.275 127.275 ;
        RECT 141.140 126.775 142.015 127.105 ;
        RECT 142.185 126.775 142.935 127.105 ;
        RECT 139.950 125.635 140.200 125.965 ;
        RECT 141.140 125.935 141.310 126.775 ;
        RECT 142.185 126.570 142.375 126.775 ;
        RECT 143.105 126.655 143.275 127.235 ;
        RECT 143.905 126.745 144.260 127.115 ;
        RECT 144.540 127.105 144.710 127.295 ;
        RECT 144.880 127.270 145.135 127.845 ;
        RECT 144.540 126.775 144.795 127.105 ;
        RECT 143.060 126.605 143.275 126.655 ;
        RECT 141.480 126.195 142.375 126.570 ;
        RECT 142.885 126.525 143.275 126.605 ;
        RECT 144.540 126.565 144.710 126.775 ;
        RECT 140.425 125.765 141.310 125.935 ;
        RECT 141.490 125.465 141.805 125.965 ;
        RECT 142.035 125.635 142.375 126.195 ;
        RECT 142.545 125.465 142.715 126.475 ;
        RECT 142.885 125.680 143.215 126.525 ;
        RECT 143.995 126.395 144.710 126.565 ;
        RECT 144.965 126.540 145.135 127.270 ;
        RECT 145.310 127.175 145.570 128.015 ;
        RECT 145.745 127.265 146.955 128.015 ;
        RECT 143.995 125.635 144.165 126.395 ;
        RECT 144.380 125.465 144.710 126.225 ;
        RECT 144.880 125.635 145.135 126.540 ;
        RECT 145.310 125.465 145.570 126.615 ;
        RECT 145.745 126.555 146.265 127.095 ;
        RECT 146.435 126.725 146.955 127.265 ;
        RECT 145.745 125.465 146.955 126.555 ;
        RECT 17.320 125.295 147.040 125.465 ;
        RECT 17.405 124.205 18.615 125.295 ;
        RECT 19.335 124.625 19.505 125.125 ;
        RECT 19.675 124.795 20.005 125.295 ;
        RECT 19.335 124.455 20.000 124.625 ;
        RECT 17.405 123.495 17.925 124.035 ;
        RECT 18.095 123.665 18.615 124.205 ;
        RECT 19.250 123.635 19.600 124.285 ;
        RECT 17.405 122.745 18.615 123.495 ;
        RECT 19.770 123.465 20.000 124.455 ;
        RECT 19.335 123.295 20.000 123.465 ;
        RECT 19.335 123.005 19.505 123.295 ;
        RECT 19.675 122.745 20.005 123.125 ;
        RECT 20.175 123.005 20.360 125.125 ;
        RECT 20.600 124.835 20.865 125.295 ;
        RECT 21.035 124.700 21.285 125.125 ;
        RECT 21.495 124.850 22.600 125.020 ;
        RECT 20.980 124.570 21.285 124.700 ;
        RECT 20.530 123.375 20.810 124.325 ;
        RECT 20.980 123.465 21.150 124.570 ;
        RECT 21.320 123.785 21.560 124.380 ;
        RECT 21.730 124.315 22.260 124.680 ;
        RECT 21.730 123.615 21.900 124.315 ;
        RECT 22.430 124.235 22.600 124.850 ;
        RECT 22.770 124.495 22.940 125.295 ;
        RECT 23.110 124.795 23.360 125.125 ;
        RECT 23.585 124.825 24.470 124.995 ;
        RECT 22.430 124.145 22.940 124.235 ;
        RECT 20.980 123.335 21.205 123.465 ;
        RECT 21.375 123.395 21.900 123.615 ;
        RECT 22.070 123.975 22.940 124.145 ;
        RECT 20.615 122.745 20.865 123.205 ;
        RECT 21.035 123.195 21.205 123.335 ;
        RECT 22.070 123.195 22.240 123.975 ;
        RECT 22.770 123.905 22.940 123.975 ;
        RECT 22.450 123.725 22.650 123.755 ;
        RECT 23.110 123.725 23.280 124.795 ;
        RECT 23.450 123.905 23.640 124.625 ;
        RECT 22.450 123.425 23.280 123.725 ;
        RECT 23.810 123.695 24.130 124.655 ;
        RECT 21.035 123.025 21.370 123.195 ;
        RECT 21.565 123.025 22.240 123.195 ;
        RECT 22.560 122.745 22.930 123.245 ;
        RECT 23.110 123.195 23.280 123.425 ;
        RECT 23.665 123.365 24.130 123.695 ;
        RECT 24.300 123.985 24.470 124.825 ;
        RECT 24.650 124.795 24.965 125.295 ;
        RECT 25.195 124.565 25.535 125.125 ;
        RECT 24.640 124.190 25.535 124.565 ;
        RECT 25.705 124.285 25.875 125.295 ;
        RECT 25.345 123.985 25.535 124.190 ;
        RECT 26.045 124.235 26.375 125.080 ;
        RECT 27.065 124.495 27.505 125.125 ;
        RECT 26.045 124.155 26.435 124.235 ;
        RECT 26.220 124.105 26.435 124.155 ;
        RECT 24.300 123.655 25.175 123.985 ;
        RECT 25.345 123.655 26.095 123.985 ;
        RECT 24.300 123.195 24.470 123.655 ;
        RECT 25.345 123.485 25.545 123.655 ;
        RECT 26.265 123.525 26.435 124.105 ;
        RECT 26.210 123.485 26.435 123.525 ;
        RECT 23.110 123.025 23.515 123.195 ;
        RECT 23.685 123.025 24.470 123.195 ;
        RECT 24.745 122.745 24.955 123.275 ;
        RECT 25.215 122.960 25.545 123.485 ;
        RECT 26.055 123.400 26.435 123.485 ;
        RECT 27.065 123.485 27.375 124.495 ;
        RECT 27.680 124.445 27.995 125.295 ;
        RECT 28.165 124.955 29.595 125.125 ;
        RECT 28.165 124.275 28.335 124.955 ;
        RECT 27.545 124.105 28.335 124.275 ;
        RECT 27.545 123.655 27.715 124.105 ;
        RECT 28.505 123.985 28.705 124.785 ;
        RECT 27.885 123.655 28.275 123.935 ;
        RECT 28.460 123.655 28.705 123.985 ;
        RECT 28.905 123.655 29.155 124.785 ;
        RECT 29.345 124.325 29.595 124.955 ;
        RECT 29.775 124.495 30.105 125.295 ;
        RECT 29.345 124.155 30.115 124.325 ;
        RECT 29.370 123.655 29.775 123.985 ;
        RECT 29.945 123.485 30.115 124.155 ;
        RECT 30.285 124.130 30.575 125.295 ;
        RECT 30.780 124.505 31.315 125.125 ;
        RECT 25.715 122.745 25.885 123.355 ;
        RECT 26.055 122.965 26.385 123.400 ;
        RECT 27.065 122.925 27.505 123.485 ;
        RECT 27.675 122.745 28.125 123.485 ;
        RECT 28.295 123.315 29.455 123.485 ;
        RECT 28.295 122.915 28.465 123.315 ;
        RECT 28.635 122.745 29.055 123.145 ;
        RECT 29.225 122.915 29.455 123.315 ;
        RECT 29.625 122.915 30.115 123.485 ;
        RECT 30.780 123.485 31.095 124.505 ;
        RECT 31.485 124.495 31.815 125.295 ;
        RECT 32.300 124.325 32.690 124.500 ;
        RECT 31.265 124.155 32.690 124.325 ;
        RECT 33.105 124.155 33.315 125.295 ;
        RECT 31.265 123.655 31.435 124.155 ;
        RECT 30.285 122.745 30.575 123.470 ;
        RECT 30.780 122.915 31.395 123.485 ;
        RECT 31.685 123.425 31.950 123.985 ;
        RECT 32.120 123.255 32.290 124.155 ;
        RECT 33.485 124.145 33.815 125.125 ;
        RECT 33.985 124.155 34.215 125.295 ;
        RECT 34.425 124.860 39.770 125.295 ;
        RECT 39.945 124.860 45.290 125.295 ;
        RECT 45.465 124.860 50.810 125.295 ;
        RECT 32.460 123.425 32.815 123.985 ;
        RECT 31.565 122.745 31.780 123.255 ;
        RECT 32.010 122.925 32.290 123.255 ;
        RECT 32.470 122.745 32.710 123.255 ;
        RECT 33.105 122.745 33.315 123.565 ;
        RECT 33.485 123.545 33.735 124.145 ;
        RECT 33.905 123.735 34.235 123.985 ;
        RECT 33.485 122.915 33.815 123.545 ;
        RECT 33.985 122.745 34.215 123.565 ;
        RECT 36.010 123.290 36.350 124.120 ;
        RECT 37.830 123.610 38.180 124.860 ;
        RECT 41.530 123.290 41.870 124.120 ;
        RECT 43.350 123.610 43.700 124.860 ;
        RECT 47.050 123.290 47.390 124.120 ;
        RECT 48.870 123.610 49.220 124.860 ;
        RECT 50.985 124.205 54.495 125.295 ;
        RECT 54.665 124.205 55.875 125.295 ;
        RECT 50.985 123.515 52.635 124.035 ;
        RECT 52.805 123.685 54.495 124.205 ;
        RECT 34.425 122.745 39.770 123.290 ;
        RECT 39.945 122.745 45.290 123.290 ;
        RECT 45.465 122.745 50.810 123.290 ;
        RECT 50.985 122.745 54.495 123.515 ;
        RECT 54.665 123.495 55.185 124.035 ;
        RECT 55.355 123.665 55.875 124.205 ;
        RECT 56.045 124.130 56.335 125.295 ;
        RECT 56.505 124.860 61.850 125.295 ;
        RECT 54.665 122.745 55.875 123.495 ;
        RECT 56.045 122.745 56.335 123.470 ;
        RECT 58.090 123.290 58.430 124.120 ;
        RECT 59.910 123.610 60.260 124.860 ;
        RECT 62.115 124.625 62.285 125.125 ;
        RECT 62.455 124.795 62.785 125.295 ;
        RECT 62.115 124.455 62.780 124.625 ;
        RECT 62.030 123.635 62.380 124.285 ;
        RECT 62.550 123.465 62.780 124.455 ;
        RECT 62.115 123.295 62.780 123.465 ;
        RECT 56.505 122.745 61.850 123.290 ;
        RECT 62.115 123.005 62.285 123.295 ;
        RECT 62.455 122.745 62.785 123.125 ;
        RECT 62.955 123.005 63.140 125.125 ;
        RECT 63.380 124.835 63.645 125.295 ;
        RECT 63.815 124.700 64.065 125.125 ;
        RECT 64.275 124.850 65.380 125.020 ;
        RECT 63.760 124.570 64.065 124.700 ;
        RECT 63.310 123.375 63.590 124.325 ;
        RECT 63.760 123.465 63.930 124.570 ;
        RECT 64.100 123.785 64.340 124.380 ;
        RECT 64.510 124.315 65.040 124.680 ;
        RECT 64.510 123.615 64.680 124.315 ;
        RECT 65.210 124.235 65.380 124.850 ;
        RECT 65.550 124.495 65.720 125.295 ;
        RECT 65.890 124.795 66.140 125.125 ;
        RECT 66.365 124.825 67.250 124.995 ;
        RECT 65.210 124.145 65.720 124.235 ;
        RECT 63.760 123.335 63.985 123.465 ;
        RECT 64.155 123.395 64.680 123.615 ;
        RECT 64.850 123.975 65.720 124.145 ;
        RECT 63.395 122.745 63.645 123.205 ;
        RECT 63.815 123.195 63.985 123.335 ;
        RECT 64.850 123.195 65.020 123.975 ;
        RECT 65.550 123.905 65.720 123.975 ;
        RECT 65.230 123.725 65.430 123.755 ;
        RECT 65.890 123.725 66.060 124.795 ;
        RECT 66.230 123.905 66.420 124.625 ;
        RECT 65.230 123.425 66.060 123.725 ;
        RECT 66.590 123.695 66.910 124.655 ;
        RECT 63.815 123.025 64.150 123.195 ;
        RECT 64.345 123.025 65.020 123.195 ;
        RECT 65.340 122.745 65.710 123.245 ;
        RECT 65.890 123.195 66.060 123.425 ;
        RECT 66.445 123.365 66.910 123.695 ;
        RECT 67.080 123.985 67.250 124.825 ;
        RECT 67.430 124.795 67.745 125.295 ;
        RECT 67.975 124.565 68.315 125.125 ;
        RECT 67.420 124.190 68.315 124.565 ;
        RECT 68.485 124.285 68.655 125.295 ;
        RECT 68.125 123.985 68.315 124.190 ;
        RECT 68.825 124.235 69.155 125.080 ;
        RECT 69.325 124.380 69.495 125.295 ;
        RECT 69.845 124.575 70.305 125.125 ;
        RECT 70.495 124.575 70.825 125.295 ;
        RECT 68.825 124.155 69.215 124.235 ;
        RECT 69.000 124.105 69.215 124.155 ;
        RECT 67.080 123.655 67.955 123.985 ;
        RECT 68.125 123.655 68.875 123.985 ;
        RECT 67.080 123.195 67.250 123.655 ;
        RECT 68.125 123.485 68.325 123.655 ;
        RECT 69.045 123.525 69.215 124.105 ;
        RECT 68.990 123.485 69.215 123.525 ;
        RECT 65.890 123.025 66.295 123.195 ;
        RECT 66.465 123.025 67.250 123.195 ;
        RECT 67.525 122.745 67.735 123.275 ;
        RECT 67.995 122.960 68.325 123.485 ;
        RECT 68.835 123.400 69.215 123.485 ;
        RECT 68.495 122.745 68.665 123.355 ;
        RECT 68.835 122.965 69.165 123.400 ;
        RECT 69.335 122.745 69.505 123.260 ;
        RECT 69.845 123.205 70.095 124.575 ;
        RECT 71.025 124.405 71.325 124.955 ;
        RECT 71.495 124.625 71.775 125.295 ;
        RECT 72.695 124.625 72.865 125.125 ;
        RECT 73.035 124.795 73.365 125.295 ;
        RECT 72.695 124.455 73.360 124.625 ;
        RECT 70.385 124.235 71.325 124.405 ;
        RECT 70.385 123.985 70.555 124.235 ;
        RECT 71.695 123.985 71.960 124.345 ;
        RECT 70.265 123.655 70.555 123.985 ;
        RECT 70.725 123.735 71.065 123.985 ;
        RECT 71.285 123.735 71.960 123.985 ;
        RECT 70.385 123.565 70.555 123.655 ;
        RECT 72.610 123.635 72.960 124.285 ;
        RECT 70.385 123.375 71.775 123.565 ;
        RECT 73.130 123.465 73.360 124.455 ;
        RECT 69.845 122.915 70.405 123.205 ;
        RECT 70.575 122.745 70.825 123.205 ;
        RECT 71.445 123.015 71.775 123.375 ;
        RECT 72.695 123.295 73.360 123.465 ;
        RECT 72.695 123.005 72.865 123.295 ;
        RECT 73.035 122.745 73.365 123.125 ;
        RECT 73.535 123.005 73.720 125.125 ;
        RECT 73.960 124.835 74.225 125.295 ;
        RECT 74.395 124.700 74.645 125.125 ;
        RECT 74.855 124.850 75.960 125.020 ;
        RECT 74.340 124.570 74.645 124.700 ;
        RECT 73.890 123.375 74.170 124.325 ;
        RECT 74.340 123.465 74.510 124.570 ;
        RECT 74.680 123.785 74.920 124.380 ;
        RECT 75.090 124.315 75.620 124.680 ;
        RECT 75.090 123.615 75.260 124.315 ;
        RECT 75.790 124.235 75.960 124.850 ;
        RECT 76.130 124.495 76.300 125.295 ;
        RECT 76.470 124.795 76.720 125.125 ;
        RECT 76.945 124.825 77.830 124.995 ;
        RECT 75.790 124.145 76.300 124.235 ;
        RECT 74.340 123.335 74.565 123.465 ;
        RECT 74.735 123.395 75.260 123.615 ;
        RECT 75.430 123.975 76.300 124.145 ;
        RECT 73.975 122.745 74.225 123.205 ;
        RECT 74.395 123.195 74.565 123.335 ;
        RECT 75.430 123.195 75.600 123.975 ;
        RECT 76.130 123.905 76.300 123.975 ;
        RECT 75.810 123.725 76.010 123.755 ;
        RECT 76.470 123.725 76.640 124.795 ;
        RECT 76.810 123.905 77.000 124.625 ;
        RECT 75.810 123.425 76.640 123.725 ;
        RECT 77.170 123.695 77.490 124.655 ;
        RECT 74.395 123.025 74.730 123.195 ;
        RECT 74.925 123.025 75.600 123.195 ;
        RECT 75.920 122.745 76.290 123.245 ;
        RECT 76.470 123.195 76.640 123.425 ;
        RECT 77.025 123.365 77.490 123.695 ;
        RECT 77.660 123.985 77.830 124.825 ;
        RECT 78.010 124.795 78.325 125.295 ;
        RECT 78.555 124.565 78.895 125.125 ;
        RECT 78.000 124.190 78.895 124.565 ;
        RECT 79.065 124.285 79.235 125.295 ;
        RECT 78.705 123.985 78.895 124.190 ;
        RECT 79.405 124.235 79.735 125.080 ;
        RECT 79.405 124.155 79.795 124.235 ;
        RECT 79.965 124.205 81.635 125.295 ;
        RECT 79.580 124.105 79.795 124.155 ;
        RECT 77.660 123.655 78.535 123.985 ;
        RECT 78.705 123.655 79.455 123.985 ;
        RECT 77.660 123.195 77.830 123.655 ;
        RECT 78.705 123.485 78.905 123.655 ;
        RECT 79.625 123.525 79.795 124.105 ;
        RECT 79.570 123.485 79.795 123.525 ;
        RECT 76.470 123.025 76.875 123.195 ;
        RECT 77.045 123.025 77.830 123.195 ;
        RECT 78.105 122.745 78.315 123.275 ;
        RECT 78.575 122.960 78.905 123.485 ;
        RECT 79.415 123.400 79.795 123.485 ;
        RECT 79.965 123.515 80.715 124.035 ;
        RECT 80.885 123.685 81.635 124.205 ;
        RECT 81.805 124.130 82.095 125.295 ;
        RECT 82.265 124.205 83.475 125.295 ;
        RECT 79.075 122.745 79.245 123.355 ;
        RECT 79.415 122.965 79.745 123.400 ;
        RECT 79.965 122.745 81.635 123.515 ;
        RECT 82.265 123.495 82.785 124.035 ;
        RECT 82.955 123.665 83.475 124.205 ;
        RECT 83.645 124.535 84.160 124.945 ;
        RECT 84.395 124.535 84.565 125.295 ;
        RECT 84.735 124.955 86.765 125.125 ;
        RECT 83.645 123.725 83.985 124.535 ;
        RECT 84.735 124.290 84.905 124.955 ;
        RECT 85.300 124.615 86.425 124.785 ;
        RECT 84.155 124.100 84.905 124.290 ;
        RECT 85.075 124.275 86.085 124.445 ;
        RECT 83.645 123.555 84.875 123.725 ;
        RECT 81.805 122.745 82.095 123.470 ;
        RECT 82.265 122.745 83.475 123.495 ;
        RECT 83.920 122.950 84.165 123.555 ;
        RECT 84.385 122.745 84.895 123.280 ;
        RECT 85.075 122.915 85.265 124.275 ;
        RECT 85.435 123.935 85.710 124.075 ;
        RECT 85.435 123.765 85.715 123.935 ;
        RECT 85.435 122.915 85.710 123.765 ;
        RECT 85.915 123.475 86.085 124.275 ;
        RECT 86.255 123.485 86.425 124.615 ;
        RECT 86.595 123.985 86.765 124.955 ;
        RECT 86.935 124.155 87.105 125.295 ;
        RECT 87.275 124.155 87.610 125.125 ;
        RECT 87.875 124.625 88.045 125.125 ;
        RECT 88.215 124.795 88.545 125.295 ;
        RECT 87.875 124.455 88.540 124.625 ;
        RECT 86.595 123.655 86.790 123.985 ;
        RECT 87.015 123.655 87.270 123.985 ;
        RECT 87.015 123.485 87.185 123.655 ;
        RECT 87.440 123.485 87.610 124.155 ;
        RECT 87.790 123.635 88.140 124.285 ;
        RECT 86.255 123.315 87.185 123.485 ;
        RECT 86.255 123.280 86.430 123.315 ;
        RECT 85.900 122.915 86.430 123.280 ;
        RECT 86.855 122.745 87.185 123.145 ;
        RECT 87.355 122.915 87.610 123.485 ;
        RECT 88.310 123.465 88.540 124.455 ;
        RECT 87.875 123.295 88.540 123.465 ;
        RECT 87.875 123.005 88.045 123.295 ;
        RECT 88.215 122.745 88.545 123.125 ;
        RECT 88.715 123.005 88.900 125.125 ;
        RECT 89.140 124.835 89.405 125.295 ;
        RECT 89.575 124.700 89.825 125.125 ;
        RECT 90.035 124.850 91.140 125.020 ;
        RECT 89.520 124.570 89.825 124.700 ;
        RECT 89.070 123.375 89.350 124.325 ;
        RECT 89.520 123.465 89.690 124.570 ;
        RECT 89.860 123.785 90.100 124.380 ;
        RECT 90.270 124.315 90.800 124.680 ;
        RECT 90.270 123.615 90.440 124.315 ;
        RECT 90.970 124.235 91.140 124.850 ;
        RECT 91.310 124.495 91.480 125.295 ;
        RECT 91.650 124.795 91.900 125.125 ;
        RECT 92.125 124.825 93.010 124.995 ;
        RECT 90.970 124.145 91.480 124.235 ;
        RECT 89.520 123.335 89.745 123.465 ;
        RECT 89.915 123.395 90.440 123.615 ;
        RECT 90.610 123.975 91.480 124.145 ;
        RECT 89.155 122.745 89.405 123.205 ;
        RECT 89.575 123.195 89.745 123.335 ;
        RECT 90.610 123.195 90.780 123.975 ;
        RECT 91.310 123.905 91.480 123.975 ;
        RECT 90.990 123.725 91.190 123.755 ;
        RECT 91.650 123.725 91.820 124.795 ;
        RECT 91.990 123.905 92.180 124.625 ;
        RECT 90.990 123.425 91.820 123.725 ;
        RECT 92.350 123.695 92.670 124.655 ;
        RECT 89.575 123.025 89.910 123.195 ;
        RECT 90.105 123.025 90.780 123.195 ;
        RECT 91.100 122.745 91.470 123.245 ;
        RECT 91.650 123.195 91.820 123.425 ;
        RECT 92.205 123.365 92.670 123.695 ;
        RECT 92.840 123.985 93.010 124.825 ;
        RECT 93.190 124.795 93.505 125.295 ;
        RECT 93.735 124.565 94.075 125.125 ;
        RECT 93.180 124.190 94.075 124.565 ;
        RECT 94.245 124.285 94.415 125.295 ;
        RECT 93.885 123.985 94.075 124.190 ;
        RECT 94.585 124.235 94.915 125.080 ;
        RECT 95.085 124.380 95.255 125.295 ;
        RECT 94.585 124.155 94.975 124.235 ;
        RECT 94.760 124.105 94.975 124.155 ;
        RECT 92.840 123.655 93.715 123.985 ;
        RECT 93.885 123.655 94.635 123.985 ;
        RECT 92.840 123.195 93.010 123.655 ;
        RECT 93.885 123.485 94.085 123.655 ;
        RECT 94.805 123.525 94.975 124.105 ;
        RECT 94.750 123.485 94.975 123.525 ;
        RECT 91.650 123.025 92.055 123.195 ;
        RECT 92.225 123.025 93.010 123.195 ;
        RECT 93.285 122.745 93.495 123.275 ;
        RECT 93.755 122.960 94.085 123.485 ;
        RECT 94.595 123.400 94.975 123.485 ;
        RECT 95.605 124.155 95.990 125.125 ;
        RECT 96.160 124.835 96.485 125.295 ;
        RECT 97.005 124.665 97.285 125.125 ;
        RECT 96.160 124.445 97.285 124.665 ;
        RECT 95.605 123.485 95.885 124.155 ;
        RECT 96.160 123.985 96.610 124.445 ;
        RECT 97.475 124.275 97.875 125.125 ;
        RECT 98.275 124.835 98.545 125.295 ;
        RECT 98.715 124.665 99.000 125.125 ;
        RECT 96.055 123.655 96.610 123.985 ;
        RECT 96.780 123.715 97.875 124.275 ;
        RECT 96.160 123.545 96.610 123.655 ;
        RECT 94.255 122.745 94.425 123.355 ;
        RECT 94.595 122.965 94.925 123.400 ;
        RECT 95.095 122.745 95.265 123.260 ;
        RECT 95.605 122.915 95.990 123.485 ;
        RECT 96.160 123.375 97.285 123.545 ;
        RECT 96.160 122.745 96.485 123.205 ;
        RECT 97.005 122.915 97.285 123.375 ;
        RECT 97.475 122.915 97.875 123.715 ;
        RECT 98.045 124.445 99.000 124.665 ;
        RECT 99.860 124.665 100.145 125.125 ;
        RECT 100.315 124.835 100.585 125.295 ;
        RECT 99.860 124.445 100.815 124.665 ;
        RECT 98.045 123.545 98.255 124.445 ;
        RECT 98.425 123.715 99.115 124.275 ;
        RECT 99.745 123.715 100.435 124.275 ;
        RECT 100.605 123.545 100.815 124.445 ;
        RECT 98.045 123.375 99.000 123.545 ;
        RECT 98.275 122.745 98.545 123.205 ;
        RECT 98.715 122.915 99.000 123.375 ;
        RECT 99.860 123.375 100.815 123.545 ;
        RECT 100.985 124.275 101.385 125.125 ;
        RECT 101.575 124.665 101.855 125.125 ;
        RECT 102.375 124.835 102.700 125.295 ;
        RECT 101.575 124.445 102.700 124.665 ;
        RECT 100.985 123.715 102.080 124.275 ;
        RECT 102.250 123.985 102.700 124.445 ;
        RECT 102.870 124.155 103.255 125.125 ;
        RECT 99.860 122.915 100.145 123.375 ;
        RECT 100.315 122.745 100.585 123.205 ;
        RECT 100.985 122.915 101.385 123.715 ;
        RECT 102.250 123.655 102.805 123.985 ;
        RECT 102.250 123.545 102.700 123.655 ;
        RECT 101.575 123.375 102.700 123.545 ;
        RECT 102.975 123.485 103.255 124.155 ;
        RECT 103.425 124.535 103.940 124.945 ;
        RECT 104.175 124.535 104.345 125.295 ;
        RECT 104.515 124.955 106.545 125.125 ;
        RECT 103.425 123.725 103.765 124.535 ;
        RECT 104.515 124.290 104.685 124.955 ;
        RECT 105.080 124.615 106.205 124.785 ;
        RECT 103.935 124.100 104.685 124.290 ;
        RECT 104.855 124.275 105.865 124.445 ;
        RECT 103.425 123.555 104.655 123.725 ;
        RECT 101.575 122.915 101.855 123.375 ;
        RECT 102.375 122.745 102.700 123.205 ;
        RECT 102.870 122.915 103.255 123.485 ;
        RECT 103.700 122.950 103.945 123.555 ;
        RECT 104.165 122.745 104.675 123.280 ;
        RECT 104.855 122.915 105.045 124.275 ;
        RECT 105.215 123.595 105.490 124.075 ;
        RECT 105.215 123.425 105.495 123.595 ;
        RECT 105.695 123.475 105.865 124.275 ;
        RECT 106.035 123.485 106.205 124.615 ;
        RECT 106.375 123.985 106.545 124.955 ;
        RECT 106.715 124.155 106.885 125.295 ;
        RECT 107.055 124.155 107.390 125.125 ;
        RECT 106.375 123.655 106.570 123.985 ;
        RECT 106.795 123.655 107.050 123.985 ;
        RECT 106.795 123.485 106.965 123.655 ;
        RECT 107.220 123.485 107.390 124.155 ;
        RECT 107.565 124.130 107.855 125.295 ;
        RECT 108.115 124.625 108.285 125.125 ;
        RECT 108.455 124.795 108.785 125.295 ;
        RECT 108.115 124.455 108.780 124.625 ;
        RECT 108.030 123.635 108.380 124.285 ;
        RECT 105.215 122.915 105.490 123.425 ;
        RECT 106.035 123.315 106.965 123.485 ;
        RECT 106.035 123.280 106.210 123.315 ;
        RECT 105.680 122.915 106.210 123.280 ;
        RECT 106.635 122.745 106.965 123.145 ;
        RECT 107.135 122.915 107.390 123.485 ;
        RECT 107.565 122.745 107.855 123.470 ;
        RECT 108.550 123.465 108.780 124.455 ;
        RECT 108.115 123.295 108.780 123.465 ;
        RECT 108.115 123.005 108.285 123.295 ;
        RECT 108.455 122.745 108.785 123.125 ;
        RECT 108.955 123.005 109.140 125.125 ;
        RECT 109.380 124.835 109.645 125.295 ;
        RECT 109.815 124.700 110.065 125.125 ;
        RECT 110.275 124.850 111.380 125.020 ;
        RECT 109.760 124.570 110.065 124.700 ;
        RECT 109.310 123.375 109.590 124.325 ;
        RECT 109.760 123.465 109.930 124.570 ;
        RECT 110.100 123.785 110.340 124.380 ;
        RECT 110.510 124.315 111.040 124.680 ;
        RECT 110.510 123.615 110.680 124.315 ;
        RECT 111.210 124.235 111.380 124.850 ;
        RECT 111.550 124.495 111.720 125.295 ;
        RECT 111.890 124.795 112.140 125.125 ;
        RECT 112.365 124.825 113.250 124.995 ;
        RECT 111.210 124.145 111.720 124.235 ;
        RECT 109.760 123.335 109.985 123.465 ;
        RECT 110.155 123.395 110.680 123.615 ;
        RECT 110.850 123.975 111.720 124.145 ;
        RECT 109.395 122.745 109.645 123.205 ;
        RECT 109.815 123.195 109.985 123.335 ;
        RECT 110.850 123.195 111.020 123.975 ;
        RECT 111.550 123.905 111.720 123.975 ;
        RECT 111.230 123.725 111.430 123.755 ;
        RECT 111.890 123.725 112.060 124.795 ;
        RECT 112.230 123.905 112.420 124.625 ;
        RECT 111.230 123.425 112.060 123.725 ;
        RECT 112.590 123.695 112.910 124.655 ;
        RECT 109.815 123.025 110.150 123.195 ;
        RECT 110.345 123.025 111.020 123.195 ;
        RECT 111.340 122.745 111.710 123.245 ;
        RECT 111.890 123.195 112.060 123.425 ;
        RECT 112.445 123.365 112.910 123.695 ;
        RECT 113.080 123.985 113.250 124.825 ;
        RECT 113.430 124.795 113.745 125.295 ;
        RECT 113.975 124.565 114.315 125.125 ;
        RECT 113.420 124.190 114.315 124.565 ;
        RECT 114.485 124.285 114.655 125.295 ;
        RECT 114.125 123.985 114.315 124.190 ;
        RECT 114.825 124.235 115.155 125.080 ;
        RECT 115.385 124.860 120.730 125.295 ;
        RECT 114.825 124.155 115.215 124.235 ;
        RECT 115.000 124.105 115.215 124.155 ;
        RECT 113.080 123.655 113.955 123.985 ;
        RECT 114.125 123.655 114.875 123.985 ;
        RECT 113.080 123.195 113.250 123.655 ;
        RECT 114.125 123.485 114.325 123.655 ;
        RECT 115.045 123.525 115.215 124.105 ;
        RECT 114.990 123.485 115.215 123.525 ;
        RECT 111.890 123.025 112.295 123.195 ;
        RECT 112.465 123.025 113.250 123.195 ;
        RECT 113.525 122.745 113.735 123.275 ;
        RECT 113.995 122.960 114.325 123.485 ;
        RECT 114.835 123.400 115.215 123.485 ;
        RECT 114.495 122.745 114.665 123.355 ;
        RECT 114.835 122.965 115.165 123.400 ;
        RECT 116.970 123.290 117.310 124.120 ;
        RECT 118.790 123.610 119.140 124.860 ;
        RECT 120.905 123.690 121.185 125.125 ;
        RECT 121.355 124.520 122.065 125.295 ;
        RECT 122.235 124.350 122.565 125.125 ;
        RECT 121.415 124.135 122.565 124.350 ;
        RECT 115.385 122.745 120.730 123.290 ;
        RECT 120.905 122.915 121.245 123.690 ;
        RECT 121.415 123.565 121.700 124.135 ;
        RECT 121.885 123.735 122.355 123.965 ;
        RECT 122.760 123.935 122.975 125.050 ;
        RECT 123.155 124.575 123.485 125.295 ;
        RECT 123.665 124.860 129.010 125.295 ;
        RECT 123.265 123.935 123.495 124.275 ;
        RECT 122.525 123.755 122.975 123.935 ;
        RECT 122.525 123.735 122.855 123.755 ;
        RECT 123.165 123.735 123.495 123.935 ;
        RECT 121.415 123.375 122.125 123.565 ;
        RECT 121.825 123.235 122.125 123.375 ;
        RECT 122.315 123.375 123.495 123.565 ;
        RECT 122.315 123.295 122.645 123.375 ;
        RECT 121.825 123.225 122.140 123.235 ;
        RECT 121.825 123.215 122.150 123.225 ;
        RECT 121.825 123.210 122.160 123.215 ;
        RECT 121.415 122.745 121.585 123.205 ;
        RECT 121.825 123.200 122.165 123.210 ;
        RECT 121.825 123.195 122.170 123.200 ;
        RECT 121.825 123.185 122.175 123.195 ;
        RECT 121.825 123.180 122.180 123.185 ;
        RECT 121.825 122.915 122.185 123.180 ;
        RECT 122.815 122.745 122.985 123.205 ;
        RECT 123.155 122.915 123.495 123.375 ;
        RECT 125.250 123.290 125.590 124.120 ;
        RECT 127.070 123.610 127.420 124.860 ;
        RECT 129.185 124.205 132.695 125.295 ;
        RECT 129.185 123.515 130.835 124.035 ;
        RECT 131.005 123.685 132.695 124.205 ;
        RECT 133.325 124.130 133.615 125.295 ;
        RECT 133.875 124.675 134.045 125.105 ;
        RECT 134.215 124.845 134.545 125.295 ;
        RECT 133.875 124.445 134.550 124.675 ;
        RECT 123.665 122.745 129.010 123.290 ;
        RECT 129.185 122.745 132.695 123.515 ;
        RECT 133.325 122.745 133.615 123.470 ;
        RECT 133.845 123.425 134.145 124.275 ;
        RECT 134.315 123.795 134.550 124.445 ;
        RECT 134.720 124.135 135.005 125.080 ;
        RECT 135.185 124.825 135.870 125.295 ;
        RECT 135.180 124.305 135.875 124.615 ;
        RECT 136.050 124.240 136.355 125.025 ;
        RECT 136.545 124.860 141.890 125.295 ;
        RECT 134.720 123.985 135.580 124.135 ;
        RECT 134.720 123.965 136.005 123.985 ;
        RECT 134.315 123.465 134.850 123.795 ;
        RECT 135.020 123.605 136.005 123.965 ;
        RECT 134.315 123.315 134.535 123.465 ;
        RECT 133.790 122.745 134.125 123.250 ;
        RECT 134.295 122.940 134.535 123.315 ;
        RECT 135.020 123.270 135.190 123.605 ;
        RECT 136.180 123.435 136.355 124.240 ;
        RECT 134.815 123.075 135.190 123.270 ;
        RECT 134.815 122.930 134.985 123.075 ;
        RECT 135.550 122.745 135.945 123.240 ;
        RECT 136.115 122.915 136.355 123.435 ;
        RECT 138.130 123.290 138.470 124.120 ;
        RECT 139.950 123.610 140.300 124.860 ;
        RECT 142.155 124.365 142.325 125.125 ;
        RECT 142.540 124.535 142.870 125.295 ;
        RECT 142.155 124.195 142.870 124.365 ;
        RECT 143.040 124.220 143.295 125.125 ;
        RECT 142.065 123.645 142.420 124.015 ;
        RECT 142.700 123.985 142.870 124.195 ;
        RECT 142.700 123.655 142.955 123.985 ;
        RECT 142.700 123.465 142.870 123.655 ;
        RECT 143.125 123.490 143.295 124.220 ;
        RECT 143.470 124.145 143.730 125.295 ;
        RECT 143.995 124.365 144.165 125.125 ;
        RECT 144.380 124.535 144.710 125.295 ;
        RECT 143.995 124.195 144.710 124.365 ;
        RECT 144.880 124.220 145.135 125.125 ;
        RECT 143.905 123.645 144.260 124.015 ;
        RECT 144.540 123.985 144.710 124.195 ;
        RECT 144.540 123.655 144.795 123.985 ;
        RECT 142.155 123.295 142.870 123.465 ;
        RECT 136.545 122.745 141.890 123.290 ;
        RECT 142.155 122.915 142.325 123.295 ;
        RECT 142.540 122.745 142.870 123.125 ;
        RECT 143.040 122.915 143.295 123.490 ;
        RECT 143.470 122.745 143.730 123.585 ;
        RECT 144.540 123.465 144.710 123.655 ;
        RECT 144.965 123.490 145.135 124.220 ;
        RECT 145.310 124.145 145.570 125.295 ;
        RECT 145.745 124.205 146.955 125.295 ;
        RECT 145.745 123.665 146.265 124.205 ;
        RECT 143.995 123.295 144.710 123.465 ;
        RECT 143.995 122.915 144.165 123.295 ;
        RECT 144.380 122.745 144.710 123.125 ;
        RECT 144.880 122.915 145.135 123.490 ;
        RECT 145.310 122.745 145.570 123.585 ;
        RECT 146.435 123.495 146.955 124.035 ;
        RECT 145.745 122.745 146.955 123.495 ;
        RECT 17.320 122.575 147.040 122.745 ;
        RECT 17.405 121.825 18.615 122.575 ;
        RECT 17.405 121.285 17.925 121.825 ;
        RECT 18.790 121.735 19.050 122.575 ;
        RECT 19.225 121.830 19.480 122.405 ;
        RECT 19.650 122.195 19.980 122.575 ;
        RECT 20.195 122.025 20.365 122.405 ;
        RECT 19.650 121.855 20.365 122.025 ;
        RECT 18.095 121.115 18.615 121.655 ;
        RECT 17.405 120.025 18.615 121.115 ;
        RECT 18.790 120.025 19.050 121.175 ;
        RECT 19.225 121.100 19.395 121.830 ;
        RECT 19.650 121.665 19.820 121.855 ;
        RECT 20.625 121.825 21.835 122.575 ;
        RECT 22.010 121.835 22.265 122.405 ;
        RECT 22.435 122.175 22.765 122.575 ;
        RECT 23.190 122.040 23.720 122.405 ;
        RECT 23.190 122.005 23.365 122.040 ;
        RECT 22.435 121.835 23.365 122.005 ;
        RECT 23.910 121.895 24.185 122.405 ;
        RECT 19.565 121.335 19.820 121.665 ;
        RECT 19.650 121.125 19.820 121.335 ;
        RECT 20.100 121.305 20.455 121.675 ;
        RECT 20.625 121.285 21.145 121.825 ;
        RECT 19.225 120.195 19.480 121.100 ;
        RECT 19.650 120.955 20.365 121.125 ;
        RECT 21.315 121.115 21.835 121.655 ;
        RECT 19.650 120.025 19.980 120.785 ;
        RECT 20.195 120.195 20.365 120.955 ;
        RECT 20.625 120.025 21.835 121.115 ;
        RECT 22.010 121.165 22.180 121.835 ;
        RECT 22.435 121.665 22.605 121.835 ;
        RECT 22.350 121.335 22.605 121.665 ;
        RECT 22.830 121.335 23.025 121.665 ;
        RECT 22.010 120.195 22.345 121.165 ;
        RECT 22.515 120.025 22.685 121.165 ;
        RECT 22.855 120.365 23.025 121.335 ;
        RECT 23.195 120.705 23.365 121.835 ;
        RECT 23.535 121.045 23.705 121.845 ;
        RECT 23.905 121.725 24.185 121.895 ;
        RECT 23.910 121.245 24.185 121.725 ;
        RECT 24.355 121.045 24.545 122.405 ;
        RECT 24.725 122.040 25.235 122.575 ;
        RECT 25.455 121.765 25.700 122.370 ;
        RECT 26.145 122.030 31.490 122.575 ;
        RECT 31.665 122.030 37.010 122.575 ;
        RECT 37.185 122.030 42.530 122.575 ;
        RECT 24.745 121.595 25.975 121.765 ;
        RECT 23.535 120.875 24.545 121.045 ;
        RECT 24.715 121.030 25.465 121.220 ;
        RECT 23.195 120.535 24.320 120.705 ;
        RECT 24.715 120.365 24.885 121.030 ;
        RECT 25.635 120.785 25.975 121.595 ;
        RECT 27.730 121.200 28.070 122.030 ;
        RECT 22.855 120.195 24.885 120.365 ;
        RECT 25.055 120.025 25.225 120.785 ;
        RECT 25.460 120.375 25.975 120.785 ;
        RECT 29.550 120.460 29.900 121.710 ;
        RECT 33.250 121.200 33.590 122.030 ;
        RECT 35.070 120.460 35.420 121.710 ;
        RECT 38.770 121.200 39.110 122.030 ;
        RECT 43.165 121.850 43.455 122.575 ;
        RECT 43.625 122.030 48.970 122.575 ;
        RECT 49.145 122.030 54.490 122.575 ;
        RECT 54.665 122.030 60.010 122.575 ;
        RECT 60.690 122.115 60.955 122.575 ;
        RECT 40.590 120.460 40.940 121.710 ;
        RECT 45.210 121.200 45.550 122.030 ;
        RECT 26.145 120.025 31.490 120.460 ;
        RECT 31.665 120.025 37.010 120.460 ;
        RECT 37.185 120.025 42.530 120.460 ;
        RECT 43.165 120.025 43.455 121.190 ;
        RECT 47.030 120.460 47.380 121.710 ;
        RECT 50.730 121.200 51.070 122.030 ;
        RECT 52.550 120.460 52.900 121.710 ;
        RECT 56.250 121.200 56.590 122.030 ;
        RECT 61.325 121.935 61.495 122.405 ;
        RECT 61.745 122.115 61.915 122.575 ;
        RECT 62.165 121.935 62.335 122.405 ;
        RECT 62.585 122.115 62.755 122.575 ;
        RECT 63.005 121.935 63.175 122.405 ;
        RECT 63.345 122.110 63.595 122.575 ;
        RECT 63.925 122.115 64.170 122.575 ;
        RECT 61.325 121.755 63.695 121.935 ;
        RECT 58.070 120.460 58.420 121.710 ;
        RECT 60.665 121.335 63.175 121.585 ;
        RECT 63.345 121.165 63.695 121.755 ;
        RECT 63.865 121.335 64.180 121.945 ;
        RECT 64.350 121.585 64.600 122.395 ;
        RECT 64.770 122.050 65.030 122.575 ;
        RECT 65.200 121.925 65.460 122.380 ;
        RECT 65.630 122.095 65.890 122.575 ;
        RECT 66.060 121.925 66.320 122.380 ;
        RECT 66.490 122.095 66.750 122.575 ;
        RECT 66.920 121.925 67.180 122.380 ;
        RECT 67.350 122.095 67.610 122.575 ;
        RECT 67.780 121.925 68.040 122.380 ;
        RECT 68.210 122.095 68.510 122.575 ;
        RECT 65.200 121.755 68.510 121.925 ;
        RECT 68.925 121.850 69.215 122.575 ;
        RECT 69.475 122.025 69.645 122.315 ;
        RECT 69.815 122.195 70.145 122.575 ;
        RECT 69.475 121.855 70.140 122.025 ;
        RECT 64.350 121.335 67.370 121.585 ;
        RECT 43.625 120.025 48.970 120.460 ;
        RECT 49.145 120.025 54.490 120.460 ;
        RECT 54.665 120.025 60.010 120.460 ;
        RECT 60.690 120.025 60.985 121.165 ;
        RECT 61.245 120.995 63.695 121.165 ;
        RECT 61.245 120.195 61.575 120.995 ;
        RECT 61.745 120.025 61.915 120.825 ;
        RECT 62.085 120.195 62.415 120.995 ;
        RECT 62.925 120.975 63.695 120.995 ;
        RECT 62.585 120.025 62.755 120.825 ;
        RECT 62.925 120.195 63.255 120.975 ;
        RECT 63.425 120.025 63.595 120.485 ;
        RECT 63.875 120.025 64.170 121.135 ;
        RECT 64.350 120.200 64.600 121.335 ;
        RECT 67.540 121.165 68.510 121.755 ;
        RECT 64.770 120.025 65.030 121.135 ;
        RECT 65.200 120.925 68.510 121.165 ;
        RECT 65.200 120.200 65.460 120.925 ;
        RECT 65.630 120.025 65.890 120.755 ;
        RECT 66.060 120.200 66.320 120.925 ;
        RECT 66.490 120.025 66.750 120.755 ;
        RECT 66.920 120.200 67.180 120.925 ;
        RECT 67.350 120.025 67.610 120.755 ;
        RECT 67.780 120.200 68.040 120.925 ;
        RECT 68.210 120.025 68.505 120.755 ;
        RECT 68.925 120.025 69.215 121.190 ;
        RECT 69.390 121.035 69.740 121.685 ;
        RECT 69.910 120.865 70.140 121.855 ;
        RECT 69.475 120.695 70.140 120.865 ;
        RECT 69.475 120.195 69.645 120.695 ;
        RECT 69.815 120.025 70.145 120.525 ;
        RECT 70.315 120.195 70.500 122.315 ;
        RECT 70.755 122.115 71.005 122.575 ;
        RECT 71.175 122.125 71.510 122.295 ;
        RECT 71.705 122.125 72.380 122.295 ;
        RECT 71.175 121.985 71.345 122.125 ;
        RECT 70.670 120.995 70.950 121.945 ;
        RECT 71.120 121.855 71.345 121.985 ;
        RECT 71.120 120.750 71.290 121.855 ;
        RECT 71.515 121.705 72.040 121.925 ;
        RECT 71.460 120.940 71.700 121.535 ;
        RECT 71.870 121.005 72.040 121.705 ;
        RECT 72.210 121.345 72.380 122.125 ;
        RECT 72.700 122.075 73.070 122.575 ;
        RECT 73.250 122.125 73.655 122.295 ;
        RECT 73.825 122.125 74.610 122.295 ;
        RECT 73.250 121.895 73.420 122.125 ;
        RECT 72.590 121.595 73.420 121.895 ;
        RECT 73.805 121.625 74.270 121.955 ;
        RECT 72.590 121.565 72.790 121.595 ;
        RECT 72.910 121.345 73.080 121.415 ;
        RECT 72.210 121.175 73.080 121.345 ;
        RECT 72.570 121.085 73.080 121.175 ;
        RECT 71.120 120.620 71.425 120.750 ;
        RECT 71.870 120.640 72.400 121.005 ;
        RECT 70.740 120.025 71.005 120.485 ;
        RECT 71.175 120.195 71.425 120.620 ;
        RECT 72.570 120.470 72.740 121.085 ;
        RECT 71.635 120.300 72.740 120.470 ;
        RECT 72.910 120.025 73.080 120.825 ;
        RECT 73.250 120.525 73.420 121.595 ;
        RECT 73.590 120.695 73.780 121.415 ;
        RECT 73.950 120.665 74.270 121.625 ;
        RECT 74.440 121.665 74.610 122.125 ;
        RECT 74.885 122.045 75.095 122.575 ;
        RECT 75.355 121.835 75.685 122.360 ;
        RECT 75.855 121.965 76.025 122.575 ;
        RECT 76.195 121.920 76.525 122.355 ;
        RECT 76.695 122.060 76.865 122.575 ;
        RECT 77.255 121.920 77.585 122.355 ;
        RECT 77.755 121.965 77.925 122.575 ;
        RECT 76.195 121.835 76.575 121.920 ;
        RECT 75.485 121.665 75.685 121.835 ;
        RECT 76.350 121.795 76.575 121.835 ;
        RECT 74.440 121.335 75.315 121.665 ;
        RECT 75.485 121.335 76.235 121.665 ;
        RECT 73.250 120.195 73.500 120.525 ;
        RECT 74.440 120.495 74.610 121.335 ;
        RECT 75.485 121.130 75.675 121.335 ;
        RECT 76.405 121.215 76.575 121.795 ;
        RECT 76.360 121.165 76.575 121.215 ;
        RECT 74.780 120.755 75.675 121.130 ;
        RECT 76.185 121.085 76.575 121.165 ;
        RECT 77.205 121.835 77.585 121.920 ;
        RECT 78.095 121.835 78.425 122.360 ;
        RECT 78.685 122.045 78.895 122.575 ;
        RECT 79.170 122.125 79.955 122.295 ;
        RECT 80.125 122.125 80.530 122.295 ;
        RECT 77.205 121.795 77.430 121.835 ;
        RECT 77.205 121.215 77.375 121.795 ;
        RECT 78.095 121.665 78.295 121.835 ;
        RECT 79.170 121.665 79.340 122.125 ;
        RECT 77.545 121.335 78.295 121.665 ;
        RECT 78.465 121.335 79.340 121.665 ;
        RECT 77.205 121.165 77.420 121.215 ;
        RECT 77.205 121.085 77.595 121.165 ;
        RECT 73.725 120.325 74.610 120.495 ;
        RECT 74.790 120.025 75.105 120.525 ;
        RECT 75.335 120.195 75.675 120.755 ;
        RECT 75.845 120.025 76.015 121.035 ;
        RECT 76.185 120.240 76.515 121.085 ;
        RECT 76.685 120.025 76.855 120.940 ;
        RECT 77.265 120.240 77.595 121.085 ;
        RECT 78.105 121.130 78.295 121.335 ;
        RECT 77.765 120.025 77.935 121.035 ;
        RECT 78.105 120.755 79.000 121.130 ;
        RECT 78.105 120.195 78.445 120.755 ;
        RECT 78.675 120.025 78.990 120.525 ;
        RECT 79.170 120.495 79.340 121.335 ;
        RECT 79.510 121.625 79.975 121.955 ;
        RECT 80.360 121.895 80.530 122.125 ;
        RECT 80.710 122.075 81.080 122.575 ;
        RECT 81.400 122.125 82.075 122.295 ;
        RECT 82.270 122.125 82.605 122.295 ;
        RECT 79.510 120.665 79.830 121.625 ;
        RECT 80.360 121.595 81.190 121.895 ;
        RECT 80.000 120.695 80.190 121.415 ;
        RECT 80.360 120.525 80.530 121.595 ;
        RECT 80.990 121.565 81.190 121.595 ;
        RECT 80.700 121.345 80.870 121.415 ;
        RECT 81.400 121.345 81.570 122.125 ;
        RECT 82.435 121.985 82.605 122.125 ;
        RECT 82.775 122.115 83.025 122.575 ;
        RECT 80.700 121.175 81.570 121.345 ;
        RECT 81.740 121.705 82.265 121.925 ;
        RECT 82.435 121.855 82.660 121.985 ;
        RECT 80.700 121.085 81.210 121.175 ;
        RECT 79.170 120.325 80.055 120.495 ;
        RECT 80.280 120.195 80.530 120.525 ;
        RECT 80.700 120.025 80.870 120.825 ;
        RECT 81.040 120.470 81.210 121.085 ;
        RECT 81.740 121.005 81.910 121.705 ;
        RECT 81.380 120.640 81.910 121.005 ;
        RECT 82.080 120.940 82.320 121.535 ;
        RECT 82.490 120.750 82.660 121.855 ;
        RECT 82.830 120.995 83.110 121.945 ;
        RECT 82.355 120.620 82.660 120.750 ;
        RECT 81.040 120.300 82.145 120.470 ;
        RECT 82.355 120.195 82.605 120.620 ;
        RECT 82.775 120.025 83.040 120.485 ;
        RECT 83.280 120.195 83.465 122.315 ;
        RECT 83.635 122.195 83.965 122.575 ;
        RECT 84.135 122.025 84.305 122.315 ;
        RECT 83.640 121.855 84.305 122.025 ;
        RECT 85.575 122.025 85.745 122.315 ;
        RECT 85.915 122.195 86.245 122.575 ;
        RECT 85.575 121.855 86.240 122.025 ;
        RECT 83.640 120.865 83.870 121.855 ;
        RECT 84.040 121.035 84.390 121.685 ;
        RECT 85.490 121.035 85.840 121.685 ;
        RECT 86.010 120.865 86.240 121.855 ;
        RECT 83.640 120.695 84.305 120.865 ;
        RECT 83.635 120.025 83.965 120.525 ;
        RECT 84.135 120.195 84.305 120.695 ;
        RECT 85.575 120.695 86.240 120.865 ;
        RECT 85.575 120.195 85.745 120.695 ;
        RECT 85.915 120.025 86.245 120.525 ;
        RECT 86.415 120.195 86.600 122.315 ;
        RECT 86.855 122.115 87.105 122.575 ;
        RECT 87.275 122.125 87.610 122.295 ;
        RECT 87.805 122.125 88.480 122.295 ;
        RECT 87.275 121.985 87.445 122.125 ;
        RECT 86.770 120.995 87.050 121.945 ;
        RECT 87.220 121.855 87.445 121.985 ;
        RECT 87.220 120.750 87.390 121.855 ;
        RECT 87.615 121.705 88.140 121.925 ;
        RECT 87.560 120.940 87.800 121.535 ;
        RECT 87.970 121.005 88.140 121.705 ;
        RECT 88.310 121.345 88.480 122.125 ;
        RECT 88.800 122.075 89.170 122.575 ;
        RECT 89.350 122.125 89.755 122.295 ;
        RECT 89.925 122.125 90.710 122.295 ;
        RECT 89.350 121.895 89.520 122.125 ;
        RECT 88.690 121.595 89.520 121.895 ;
        RECT 89.905 121.625 90.370 121.955 ;
        RECT 88.690 121.565 88.890 121.595 ;
        RECT 89.010 121.345 89.180 121.415 ;
        RECT 88.310 121.175 89.180 121.345 ;
        RECT 88.670 121.085 89.180 121.175 ;
        RECT 87.220 120.620 87.525 120.750 ;
        RECT 87.970 120.640 88.500 121.005 ;
        RECT 86.840 120.025 87.105 120.485 ;
        RECT 87.275 120.195 87.525 120.620 ;
        RECT 88.670 120.470 88.840 121.085 ;
        RECT 87.735 120.300 88.840 120.470 ;
        RECT 89.010 120.025 89.180 120.825 ;
        RECT 89.350 120.525 89.520 121.595 ;
        RECT 89.690 120.695 89.880 121.415 ;
        RECT 90.050 120.665 90.370 121.625 ;
        RECT 90.540 121.665 90.710 122.125 ;
        RECT 90.985 122.045 91.195 122.575 ;
        RECT 91.455 121.835 91.785 122.360 ;
        RECT 91.955 121.965 92.125 122.575 ;
        RECT 92.295 121.920 92.625 122.355 ;
        RECT 92.795 122.060 92.965 122.575 ;
        RECT 92.295 121.835 92.675 121.920 ;
        RECT 91.585 121.665 91.785 121.835 ;
        RECT 92.450 121.795 92.675 121.835 ;
        RECT 90.540 121.335 91.415 121.665 ;
        RECT 91.585 121.335 92.335 121.665 ;
        RECT 89.350 120.195 89.600 120.525 ;
        RECT 90.540 120.495 90.710 121.335 ;
        RECT 91.585 121.130 91.775 121.335 ;
        RECT 92.505 121.215 92.675 121.795 ;
        RECT 93.305 121.825 94.515 122.575 ;
        RECT 94.685 121.850 94.975 122.575 ;
        RECT 93.305 121.285 93.825 121.825 ;
        RECT 95.145 121.805 97.735 122.575 ;
        RECT 98.020 121.945 98.305 122.405 ;
        RECT 98.475 122.115 98.745 122.575 ;
        RECT 92.460 121.165 92.675 121.215 ;
        RECT 90.880 120.755 91.775 121.130 ;
        RECT 92.285 121.085 92.675 121.165 ;
        RECT 93.995 121.115 94.515 121.655 ;
        RECT 95.145 121.285 96.355 121.805 ;
        RECT 98.020 121.775 98.975 121.945 ;
        RECT 89.825 120.325 90.710 120.495 ;
        RECT 90.890 120.025 91.205 120.525 ;
        RECT 91.435 120.195 91.775 120.755 ;
        RECT 91.945 120.025 92.115 121.035 ;
        RECT 92.285 120.240 92.615 121.085 ;
        RECT 92.785 120.025 92.955 120.940 ;
        RECT 93.305 120.025 94.515 121.115 ;
        RECT 94.685 120.025 94.975 121.190 ;
        RECT 96.525 121.115 97.735 121.635 ;
        RECT 95.145 120.025 97.735 121.115 ;
        RECT 97.905 121.045 98.595 121.605 ;
        RECT 98.765 120.875 98.975 121.775 ;
        RECT 98.020 120.655 98.975 120.875 ;
        RECT 99.145 121.605 99.545 122.405 ;
        RECT 99.735 121.945 100.015 122.405 ;
        RECT 100.535 122.115 100.860 122.575 ;
        RECT 99.735 121.775 100.860 121.945 ;
        RECT 101.030 121.835 101.415 122.405 ;
        RECT 100.410 121.665 100.860 121.775 ;
        RECT 99.145 121.045 100.240 121.605 ;
        RECT 100.410 121.335 100.965 121.665 ;
        RECT 98.020 120.195 98.305 120.655 ;
        RECT 98.475 120.025 98.745 120.485 ;
        RECT 99.145 120.195 99.545 121.045 ;
        RECT 100.410 120.875 100.860 121.335 ;
        RECT 101.135 121.165 101.415 121.835 ;
        RECT 101.585 121.805 105.095 122.575 ;
        RECT 105.265 121.825 106.475 122.575 ;
        RECT 106.695 122.035 106.920 122.395 ;
        RECT 107.100 122.205 107.430 122.575 ;
        RECT 107.610 122.035 107.865 122.395 ;
        RECT 108.430 122.205 109.175 122.575 ;
        RECT 106.695 121.845 109.180 122.035 ;
        RECT 101.585 121.285 103.235 121.805 ;
        RECT 99.735 120.655 100.860 120.875 ;
        RECT 99.735 120.195 100.015 120.655 ;
        RECT 100.535 120.025 100.860 120.485 ;
        RECT 101.030 120.195 101.415 121.165 ;
        RECT 103.405 121.115 105.095 121.635 ;
        RECT 105.265 121.285 105.785 121.825 ;
        RECT 105.955 121.115 106.475 121.655 ;
        RECT 106.655 121.335 106.925 121.665 ;
        RECT 107.105 121.335 107.540 121.665 ;
        RECT 107.720 121.335 108.295 121.665 ;
        RECT 108.475 121.335 108.755 121.665 ;
        RECT 108.955 121.155 109.180 121.845 ;
        RECT 101.585 120.025 105.095 121.115 ;
        RECT 105.265 120.025 106.475 121.115 ;
        RECT 106.685 120.975 109.180 121.155 ;
        RECT 109.355 120.975 109.690 122.395 ;
        RECT 109.865 121.805 111.535 122.575 ;
        RECT 111.795 122.025 111.965 122.315 ;
        RECT 112.135 122.195 112.465 122.575 ;
        RECT 111.795 121.855 112.460 122.025 ;
        RECT 109.865 121.285 110.615 121.805 ;
        RECT 110.785 121.115 111.535 121.635 ;
        RECT 106.685 120.205 106.975 120.975 ;
        RECT 107.545 120.565 108.735 120.795 ;
        RECT 107.545 120.205 107.805 120.565 ;
        RECT 107.975 120.025 108.305 120.395 ;
        RECT 108.475 120.205 108.735 120.565 ;
        RECT 108.925 120.025 109.255 120.745 ;
        RECT 109.425 120.205 109.690 120.975 ;
        RECT 109.865 120.025 111.535 121.115 ;
        RECT 111.710 121.035 112.060 121.685 ;
        RECT 112.230 120.865 112.460 121.855 ;
        RECT 111.795 120.695 112.460 120.865 ;
        RECT 111.795 120.195 111.965 120.695 ;
        RECT 112.135 120.025 112.465 120.525 ;
        RECT 112.635 120.195 112.820 122.315 ;
        RECT 113.075 122.115 113.325 122.575 ;
        RECT 113.495 122.125 113.830 122.295 ;
        RECT 114.025 122.125 114.700 122.295 ;
        RECT 113.495 121.985 113.665 122.125 ;
        RECT 112.990 120.995 113.270 121.945 ;
        RECT 113.440 121.855 113.665 121.985 ;
        RECT 113.440 120.750 113.610 121.855 ;
        RECT 113.835 121.705 114.360 121.925 ;
        RECT 113.780 120.940 114.020 121.535 ;
        RECT 114.190 121.005 114.360 121.705 ;
        RECT 114.530 121.345 114.700 122.125 ;
        RECT 115.020 122.075 115.390 122.575 ;
        RECT 115.570 122.125 115.975 122.295 ;
        RECT 116.145 122.125 116.930 122.295 ;
        RECT 115.570 121.895 115.740 122.125 ;
        RECT 114.910 121.595 115.740 121.895 ;
        RECT 116.125 121.625 116.590 121.955 ;
        RECT 114.910 121.565 115.110 121.595 ;
        RECT 115.230 121.345 115.400 121.415 ;
        RECT 114.530 121.175 115.400 121.345 ;
        RECT 114.890 121.085 115.400 121.175 ;
        RECT 113.440 120.620 113.745 120.750 ;
        RECT 114.190 120.640 114.720 121.005 ;
        RECT 113.060 120.025 113.325 120.485 ;
        RECT 113.495 120.195 113.745 120.620 ;
        RECT 114.890 120.470 115.060 121.085 ;
        RECT 113.955 120.300 115.060 120.470 ;
        RECT 115.230 120.025 115.400 120.825 ;
        RECT 115.570 120.525 115.740 121.595 ;
        RECT 115.910 120.695 116.100 121.415 ;
        RECT 116.270 120.665 116.590 121.625 ;
        RECT 116.760 121.665 116.930 122.125 ;
        RECT 117.205 122.045 117.415 122.575 ;
        RECT 117.675 121.835 118.005 122.360 ;
        RECT 118.175 121.965 118.345 122.575 ;
        RECT 118.515 121.920 118.845 122.355 ;
        RECT 118.515 121.835 118.895 121.920 ;
        RECT 117.805 121.665 118.005 121.835 ;
        RECT 118.670 121.795 118.895 121.835 ;
        RECT 116.760 121.335 117.635 121.665 ;
        RECT 117.805 121.335 118.555 121.665 ;
        RECT 115.570 120.195 115.820 120.525 ;
        RECT 116.760 120.495 116.930 121.335 ;
        RECT 117.805 121.130 117.995 121.335 ;
        RECT 118.725 121.215 118.895 121.795 ;
        RECT 119.065 121.825 120.275 122.575 ;
        RECT 120.445 121.850 120.735 122.575 ;
        RECT 120.925 121.885 121.165 122.405 ;
        RECT 121.335 122.080 121.730 122.575 ;
        RECT 122.295 122.245 122.465 122.390 ;
        RECT 122.090 122.050 122.465 122.245 ;
        RECT 119.065 121.285 119.585 121.825 ;
        RECT 118.680 121.165 118.895 121.215 ;
        RECT 117.100 120.755 117.995 121.130 ;
        RECT 118.505 121.085 118.895 121.165 ;
        RECT 119.755 121.115 120.275 121.655 ;
        RECT 116.045 120.325 116.930 120.495 ;
        RECT 117.110 120.025 117.425 120.525 ;
        RECT 117.655 120.195 117.995 120.755 ;
        RECT 118.165 120.025 118.335 121.035 ;
        RECT 118.505 120.240 118.835 121.085 ;
        RECT 119.065 120.025 120.275 121.115 ;
        RECT 120.445 120.025 120.735 121.190 ;
        RECT 120.925 121.080 121.100 121.885 ;
        RECT 122.090 121.715 122.260 122.050 ;
        RECT 122.745 122.005 122.985 122.380 ;
        RECT 123.155 122.070 123.490 122.575 ;
        RECT 123.665 122.030 129.010 122.575 ;
        RECT 129.650 122.070 129.985 122.575 ;
        RECT 122.745 121.855 122.965 122.005 ;
        RECT 121.275 121.355 122.260 121.715 ;
        RECT 122.430 121.525 122.965 121.855 ;
        RECT 121.275 121.335 122.560 121.355 ;
        RECT 121.700 121.185 122.560 121.335 ;
        RECT 120.925 120.295 121.230 121.080 ;
        RECT 121.405 120.705 122.100 121.015 ;
        RECT 121.410 120.025 122.095 120.495 ;
        RECT 122.275 120.240 122.560 121.185 ;
        RECT 122.730 120.875 122.965 121.525 ;
        RECT 123.135 121.045 123.435 121.895 ;
        RECT 125.250 121.200 125.590 122.030 ;
        RECT 130.155 122.005 130.395 122.380 ;
        RECT 130.675 122.245 130.845 122.390 ;
        RECT 130.675 122.050 131.050 122.245 ;
        RECT 131.410 122.080 131.805 122.575 ;
        RECT 122.730 120.645 123.405 120.875 ;
        RECT 122.735 120.025 123.065 120.475 ;
        RECT 123.235 120.215 123.405 120.645 ;
        RECT 127.070 120.460 127.420 121.710 ;
        RECT 129.705 121.045 130.005 121.895 ;
        RECT 130.175 121.855 130.395 122.005 ;
        RECT 130.175 121.525 130.710 121.855 ;
        RECT 130.880 121.715 131.050 122.050 ;
        RECT 131.975 121.885 132.215 122.405 ;
        RECT 130.175 120.875 130.410 121.525 ;
        RECT 130.880 121.355 131.865 121.715 ;
        RECT 129.735 120.645 130.410 120.875 ;
        RECT 130.580 121.335 131.865 121.355 ;
        RECT 130.580 121.185 131.440 121.335 ;
        RECT 123.665 120.025 129.010 120.460 ;
        RECT 129.735 120.215 129.905 120.645 ;
        RECT 130.075 120.025 130.405 120.475 ;
        RECT 130.580 120.240 130.865 121.185 ;
        RECT 132.040 121.080 132.215 121.885 ;
        RECT 132.405 121.805 134.995 122.575 ;
        RECT 135.630 121.835 135.885 122.405 ;
        RECT 136.055 122.175 136.385 122.575 ;
        RECT 136.810 122.040 137.340 122.405 ;
        RECT 137.530 122.235 137.805 122.405 ;
        RECT 137.525 122.065 137.805 122.235 ;
        RECT 136.810 122.005 136.985 122.040 ;
        RECT 136.055 121.835 136.985 122.005 ;
        RECT 132.405 121.285 133.615 121.805 ;
        RECT 133.785 121.115 134.995 121.635 ;
        RECT 131.040 120.705 131.735 121.015 ;
        RECT 131.045 120.025 131.730 120.495 ;
        RECT 131.910 120.295 132.215 121.080 ;
        RECT 132.405 120.025 134.995 121.115 ;
        RECT 135.630 121.165 135.800 121.835 ;
        RECT 136.055 121.665 136.225 121.835 ;
        RECT 135.970 121.335 136.225 121.665 ;
        RECT 136.450 121.335 136.645 121.665 ;
        RECT 135.630 120.195 135.965 121.165 ;
        RECT 136.135 120.025 136.305 121.165 ;
        RECT 136.475 120.365 136.645 121.335 ;
        RECT 136.815 120.705 136.985 121.835 ;
        RECT 137.155 121.045 137.325 121.845 ;
        RECT 137.530 121.245 137.805 122.065 ;
        RECT 137.975 121.045 138.165 122.405 ;
        RECT 138.345 122.040 138.855 122.575 ;
        RECT 139.075 121.765 139.320 122.370 ;
        RECT 139.765 122.030 145.110 122.575 ;
        RECT 138.365 121.595 139.595 121.765 ;
        RECT 137.155 120.875 138.165 121.045 ;
        RECT 138.335 121.030 139.085 121.220 ;
        RECT 136.815 120.535 137.940 120.705 ;
        RECT 138.335 120.365 138.505 121.030 ;
        RECT 139.255 120.785 139.595 121.595 ;
        RECT 141.350 121.200 141.690 122.030 ;
        RECT 145.745 121.825 146.955 122.575 ;
        RECT 136.475 120.195 138.505 120.365 ;
        RECT 138.675 120.025 138.845 120.785 ;
        RECT 139.080 120.375 139.595 120.785 ;
        RECT 143.170 120.460 143.520 121.710 ;
        RECT 145.745 121.115 146.265 121.655 ;
        RECT 146.435 121.285 146.955 121.825 ;
        RECT 139.765 120.025 145.110 120.460 ;
        RECT 145.745 120.025 146.955 121.115 ;
        RECT 17.320 119.855 147.040 120.025 ;
        RECT 17.405 118.765 18.615 119.855 ;
        RECT 17.405 118.055 17.925 118.595 ;
        RECT 18.095 118.225 18.615 118.765 ;
        RECT 18.790 118.705 19.050 119.855 ;
        RECT 19.225 118.780 19.480 119.685 ;
        RECT 19.650 119.095 19.980 119.855 ;
        RECT 20.195 118.925 20.365 119.685 ;
        RECT 17.405 117.305 18.615 118.055 ;
        RECT 18.790 117.305 19.050 118.145 ;
        RECT 19.225 118.050 19.395 118.780 ;
        RECT 19.650 118.755 20.365 118.925 ;
        RECT 19.650 118.545 19.820 118.755 ;
        RECT 20.630 118.705 20.890 119.855 ;
        RECT 21.065 118.780 21.320 119.685 ;
        RECT 21.490 119.095 21.820 119.855 ;
        RECT 22.035 118.925 22.205 119.685 ;
        RECT 19.565 118.215 19.820 118.545 ;
        RECT 19.225 117.475 19.480 118.050 ;
        RECT 19.650 118.025 19.820 118.215 ;
        RECT 20.100 118.205 20.455 118.575 ;
        RECT 19.650 117.855 20.365 118.025 ;
        RECT 19.650 117.305 19.980 117.685 ;
        RECT 20.195 117.475 20.365 117.855 ;
        RECT 20.630 117.305 20.890 118.145 ;
        RECT 21.065 118.050 21.235 118.780 ;
        RECT 21.490 118.755 22.205 118.925 ;
        RECT 22.465 118.765 25.975 119.855 ;
        RECT 21.490 118.545 21.660 118.755 ;
        RECT 21.405 118.215 21.660 118.545 ;
        RECT 21.065 117.475 21.320 118.050 ;
        RECT 21.490 118.025 21.660 118.215 ;
        RECT 21.940 118.205 22.295 118.575 ;
        RECT 22.465 118.075 24.115 118.595 ;
        RECT 24.285 118.245 25.975 118.765 ;
        RECT 26.330 118.885 26.720 119.060 ;
        RECT 27.205 119.055 27.535 119.855 ;
        RECT 27.705 119.065 28.240 119.685 ;
        RECT 26.330 118.715 27.755 118.885 ;
        RECT 21.490 117.855 22.205 118.025 ;
        RECT 21.490 117.305 21.820 117.685 ;
        RECT 22.035 117.475 22.205 117.855 ;
        RECT 22.465 117.305 25.975 118.075 ;
        RECT 26.205 117.985 26.560 118.545 ;
        RECT 26.730 117.815 26.900 118.715 ;
        RECT 27.070 117.985 27.335 118.545 ;
        RECT 27.585 118.215 27.755 118.715 ;
        RECT 27.925 118.045 28.240 119.065 ;
        RECT 28.445 118.765 30.115 119.855 ;
        RECT 26.310 117.305 26.550 117.815 ;
        RECT 26.730 117.485 27.010 117.815 ;
        RECT 27.240 117.305 27.455 117.815 ;
        RECT 27.625 117.475 28.240 118.045 ;
        RECT 28.445 118.075 29.195 118.595 ;
        RECT 29.365 118.245 30.115 118.765 ;
        RECT 30.285 118.690 30.575 119.855 ;
        RECT 30.745 119.420 36.090 119.855 ;
        RECT 36.265 119.420 41.610 119.855 ;
        RECT 41.785 119.420 47.130 119.855 ;
        RECT 47.305 119.420 52.650 119.855 ;
        RECT 28.445 117.305 30.115 118.075 ;
        RECT 30.285 117.305 30.575 118.030 ;
        RECT 32.330 117.850 32.670 118.680 ;
        RECT 34.150 118.170 34.500 119.420 ;
        RECT 37.850 117.850 38.190 118.680 ;
        RECT 39.670 118.170 40.020 119.420 ;
        RECT 43.370 117.850 43.710 118.680 ;
        RECT 45.190 118.170 45.540 119.420 ;
        RECT 48.890 117.850 49.230 118.680 ;
        RECT 50.710 118.170 51.060 119.420 ;
        RECT 52.825 118.765 55.415 119.855 ;
        RECT 52.825 118.075 54.035 118.595 ;
        RECT 54.205 118.245 55.415 118.765 ;
        RECT 56.045 118.690 56.335 119.855 ;
        RECT 56.505 119.420 61.850 119.855 ;
        RECT 30.745 117.305 36.090 117.850 ;
        RECT 36.265 117.305 41.610 117.850 ;
        RECT 41.785 117.305 47.130 117.850 ;
        RECT 47.305 117.305 52.650 117.850 ;
        RECT 52.825 117.305 55.415 118.075 ;
        RECT 56.045 117.305 56.335 118.030 ;
        RECT 58.090 117.850 58.430 118.680 ;
        RECT 59.910 118.170 60.260 119.420 ;
        RECT 62.025 118.765 64.615 119.855 ;
        RECT 62.025 118.075 63.235 118.595 ;
        RECT 63.405 118.245 64.615 118.765 ;
        RECT 64.790 118.715 65.125 119.685 ;
        RECT 65.295 118.715 65.465 119.855 ;
        RECT 65.635 119.515 67.665 119.685 ;
        RECT 56.505 117.305 61.850 117.850 ;
        RECT 62.025 117.305 64.615 118.075 ;
        RECT 64.790 118.045 64.960 118.715 ;
        RECT 65.635 118.545 65.805 119.515 ;
        RECT 65.130 118.215 65.385 118.545 ;
        RECT 65.610 118.215 65.805 118.545 ;
        RECT 65.975 119.175 67.100 119.345 ;
        RECT 65.215 118.045 65.385 118.215 ;
        RECT 65.975 118.045 66.145 119.175 ;
        RECT 64.790 117.475 65.045 118.045 ;
        RECT 65.215 117.875 66.145 118.045 ;
        RECT 66.315 118.835 67.325 119.005 ;
        RECT 66.315 118.035 66.485 118.835 ;
        RECT 65.970 117.840 66.145 117.875 ;
        RECT 65.215 117.305 65.545 117.705 ;
        RECT 65.970 117.475 66.500 117.840 ;
        RECT 66.690 117.815 66.965 118.635 ;
        RECT 66.685 117.645 66.965 117.815 ;
        RECT 66.690 117.475 66.965 117.645 ;
        RECT 67.135 117.475 67.325 118.835 ;
        RECT 67.495 118.850 67.665 119.515 ;
        RECT 67.835 119.095 68.005 119.855 ;
        RECT 68.240 119.095 68.755 119.505 ;
        RECT 67.495 118.660 68.245 118.850 ;
        RECT 68.415 118.285 68.755 119.095 ;
        RECT 68.925 118.765 71.515 119.855 ;
        RECT 67.525 118.115 68.755 118.285 ;
        RECT 67.505 117.305 68.015 117.840 ;
        RECT 68.235 117.510 68.480 118.115 ;
        RECT 68.925 118.075 70.135 118.595 ;
        RECT 70.305 118.245 71.515 118.765 ;
        RECT 71.690 118.715 72.025 119.685 ;
        RECT 72.195 118.715 72.365 119.855 ;
        RECT 72.535 119.515 74.565 119.685 ;
        RECT 68.925 117.305 71.515 118.075 ;
        RECT 71.690 118.045 71.860 118.715 ;
        RECT 72.535 118.545 72.705 119.515 ;
        RECT 72.030 118.215 72.285 118.545 ;
        RECT 72.510 118.215 72.705 118.545 ;
        RECT 72.875 119.175 74.000 119.345 ;
        RECT 72.115 118.045 72.285 118.215 ;
        RECT 72.875 118.045 73.045 119.175 ;
        RECT 71.690 117.475 71.945 118.045 ;
        RECT 72.115 117.875 73.045 118.045 ;
        RECT 73.215 118.835 74.225 119.005 ;
        RECT 73.215 118.035 73.385 118.835 ;
        RECT 73.590 118.155 73.865 118.635 ;
        RECT 73.585 117.985 73.865 118.155 ;
        RECT 72.870 117.840 73.045 117.875 ;
        RECT 72.115 117.305 72.445 117.705 ;
        RECT 72.870 117.475 73.400 117.840 ;
        RECT 73.590 117.475 73.865 117.985 ;
        RECT 74.035 117.475 74.225 118.835 ;
        RECT 74.395 118.850 74.565 119.515 ;
        RECT 74.735 119.095 74.905 119.855 ;
        RECT 75.140 119.095 75.655 119.505 ;
        RECT 75.825 119.420 81.170 119.855 ;
        RECT 74.395 118.660 75.145 118.850 ;
        RECT 75.315 118.285 75.655 119.095 ;
        RECT 74.425 118.115 75.655 118.285 ;
        RECT 74.405 117.305 74.915 117.840 ;
        RECT 75.135 117.510 75.380 118.115 ;
        RECT 77.410 117.850 77.750 118.680 ;
        RECT 79.230 118.170 79.580 119.420 ;
        RECT 81.805 118.690 82.095 119.855 ;
        RECT 82.270 118.715 82.605 119.685 ;
        RECT 82.775 118.715 82.945 119.855 ;
        RECT 83.115 119.515 85.145 119.685 ;
        RECT 82.270 118.045 82.440 118.715 ;
        RECT 83.115 118.545 83.285 119.515 ;
        RECT 82.610 118.215 82.865 118.545 ;
        RECT 83.090 118.215 83.285 118.545 ;
        RECT 83.455 119.175 84.580 119.345 ;
        RECT 82.695 118.045 82.865 118.215 ;
        RECT 83.455 118.045 83.625 119.175 ;
        RECT 75.825 117.305 81.170 117.850 ;
        RECT 81.805 117.305 82.095 118.030 ;
        RECT 82.270 117.475 82.525 118.045 ;
        RECT 82.695 117.875 83.625 118.045 ;
        RECT 83.795 118.835 84.805 119.005 ;
        RECT 83.795 118.035 83.965 118.835 ;
        RECT 84.170 118.495 84.445 118.635 ;
        RECT 84.165 118.325 84.445 118.495 ;
        RECT 83.450 117.840 83.625 117.875 ;
        RECT 82.695 117.305 83.025 117.705 ;
        RECT 83.450 117.475 83.980 117.840 ;
        RECT 84.170 117.475 84.445 118.325 ;
        RECT 84.615 117.475 84.805 118.835 ;
        RECT 84.975 118.850 85.145 119.515 ;
        RECT 85.315 119.095 85.485 119.855 ;
        RECT 85.720 119.095 86.235 119.505 ;
        RECT 84.975 118.660 85.725 118.850 ;
        RECT 85.895 118.285 86.235 119.095 ;
        RECT 86.405 118.765 89.915 119.855 ;
        RECT 90.085 118.765 91.295 119.855 ;
        RECT 91.715 119.125 92.010 119.855 ;
        RECT 92.180 118.955 92.440 119.680 ;
        RECT 92.610 119.125 92.870 119.855 ;
        RECT 93.040 118.955 93.300 119.680 ;
        RECT 93.470 119.125 93.730 119.855 ;
        RECT 93.900 118.955 94.160 119.680 ;
        RECT 94.330 119.125 94.590 119.855 ;
        RECT 94.760 118.955 95.020 119.680 ;
        RECT 85.005 118.115 86.235 118.285 ;
        RECT 84.985 117.305 85.495 117.840 ;
        RECT 85.715 117.510 85.960 118.115 ;
        RECT 86.405 118.075 88.055 118.595 ;
        RECT 88.225 118.245 89.915 118.765 ;
        RECT 86.405 117.305 89.915 118.075 ;
        RECT 90.085 118.055 90.605 118.595 ;
        RECT 90.775 118.225 91.295 118.765 ;
        RECT 91.710 118.715 95.020 118.955 ;
        RECT 95.190 118.745 95.450 119.855 ;
        RECT 91.710 118.125 92.680 118.715 ;
        RECT 95.620 118.545 95.870 119.680 ;
        RECT 96.050 118.745 96.345 119.855 ;
        RECT 96.530 118.715 96.865 119.685 ;
        RECT 97.035 118.715 97.205 119.855 ;
        RECT 97.375 119.515 99.405 119.685 ;
        RECT 92.850 118.295 95.870 118.545 ;
        RECT 90.085 117.305 91.295 118.055 ;
        RECT 91.710 117.955 95.020 118.125 ;
        RECT 91.710 117.305 92.010 117.785 ;
        RECT 92.180 117.500 92.440 117.955 ;
        RECT 92.610 117.305 92.870 117.785 ;
        RECT 93.040 117.500 93.300 117.955 ;
        RECT 93.470 117.305 93.730 117.785 ;
        RECT 93.900 117.500 94.160 117.955 ;
        RECT 94.330 117.305 94.590 117.785 ;
        RECT 94.760 117.500 95.020 117.955 ;
        RECT 95.190 117.305 95.450 117.830 ;
        RECT 95.620 117.485 95.870 118.295 ;
        RECT 96.040 117.935 96.355 118.545 ;
        RECT 96.530 118.045 96.700 118.715 ;
        RECT 97.375 118.545 97.545 119.515 ;
        RECT 96.870 118.215 97.125 118.545 ;
        RECT 97.350 118.215 97.545 118.545 ;
        RECT 97.715 119.175 98.840 119.345 ;
        RECT 96.955 118.045 97.125 118.215 ;
        RECT 97.715 118.045 97.885 119.175 ;
        RECT 96.050 117.305 96.295 117.765 ;
        RECT 96.530 117.475 96.785 118.045 ;
        RECT 96.955 117.875 97.885 118.045 ;
        RECT 98.055 118.835 99.065 119.005 ;
        RECT 98.055 118.035 98.225 118.835 ;
        RECT 98.430 118.155 98.705 118.635 ;
        RECT 98.425 117.985 98.705 118.155 ;
        RECT 97.710 117.840 97.885 117.875 ;
        RECT 96.955 117.305 97.285 117.705 ;
        RECT 97.710 117.475 98.240 117.840 ;
        RECT 98.430 117.475 98.705 117.985 ;
        RECT 98.875 117.475 99.065 118.835 ;
        RECT 99.235 118.850 99.405 119.515 ;
        RECT 99.575 119.095 99.745 119.855 ;
        RECT 99.980 119.095 100.495 119.505 ;
        RECT 99.235 118.660 99.985 118.850 ;
        RECT 100.155 118.285 100.495 119.095 ;
        RECT 99.265 118.115 100.495 118.285 ;
        RECT 100.670 118.715 101.005 119.685 ;
        RECT 101.175 118.715 101.345 119.855 ;
        RECT 101.515 119.515 103.545 119.685 ;
        RECT 99.245 117.305 99.755 117.840 ;
        RECT 99.975 117.510 100.220 118.115 ;
        RECT 100.670 118.045 100.840 118.715 ;
        RECT 101.515 118.545 101.685 119.515 ;
        RECT 101.010 118.215 101.265 118.545 ;
        RECT 101.490 118.215 101.685 118.545 ;
        RECT 101.855 119.175 102.980 119.345 ;
        RECT 101.095 118.045 101.265 118.215 ;
        RECT 101.855 118.045 102.025 119.175 ;
        RECT 100.670 117.475 100.925 118.045 ;
        RECT 101.095 117.875 102.025 118.045 ;
        RECT 102.195 118.835 103.205 119.005 ;
        RECT 102.195 118.035 102.365 118.835 ;
        RECT 102.570 118.155 102.845 118.635 ;
        RECT 102.565 117.985 102.845 118.155 ;
        RECT 101.850 117.840 102.025 117.875 ;
        RECT 101.095 117.305 101.425 117.705 ;
        RECT 101.850 117.475 102.380 117.840 ;
        RECT 102.570 117.475 102.845 117.985 ;
        RECT 103.015 117.475 103.205 118.835 ;
        RECT 103.375 118.850 103.545 119.515 ;
        RECT 103.715 119.095 103.885 119.855 ;
        RECT 104.120 119.095 104.635 119.505 ;
        RECT 103.375 118.660 104.125 118.850 ;
        RECT 104.295 118.285 104.635 119.095 ;
        RECT 104.805 118.765 107.395 119.855 ;
        RECT 103.405 118.115 104.635 118.285 ;
        RECT 103.385 117.305 103.895 117.840 ;
        RECT 104.115 117.510 104.360 118.115 ;
        RECT 104.805 118.075 106.015 118.595 ;
        RECT 106.185 118.245 107.395 118.765 ;
        RECT 107.565 118.690 107.855 119.855 ;
        RECT 109.035 119.235 109.205 119.665 ;
        RECT 109.375 119.405 109.705 119.855 ;
        RECT 109.035 119.005 109.710 119.235 ;
        RECT 104.805 117.305 107.395 118.075 ;
        RECT 107.565 117.305 107.855 118.030 ;
        RECT 109.005 117.985 109.305 118.835 ;
        RECT 109.475 118.355 109.710 119.005 ;
        RECT 109.880 118.695 110.165 119.640 ;
        RECT 110.345 119.385 111.030 119.855 ;
        RECT 110.340 118.865 111.035 119.175 ;
        RECT 111.210 118.800 111.515 119.585 ;
        RECT 109.880 118.545 110.740 118.695 ;
        RECT 109.880 118.525 111.165 118.545 ;
        RECT 109.475 118.025 110.010 118.355 ;
        RECT 110.180 118.165 111.165 118.525 ;
        RECT 109.475 117.875 109.695 118.025 ;
        RECT 108.950 117.305 109.285 117.810 ;
        RECT 109.455 117.500 109.695 117.875 ;
        RECT 110.180 117.830 110.350 118.165 ;
        RECT 111.340 117.995 111.515 118.800 ;
        RECT 109.975 117.635 110.350 117.830 ;
        RECT 109.975 117.490 110.145 117.635 ;
        RECT 110.710 117.305 111.105 117.800 ;
        RECT 111.275 117.475 111.515 117.995 ;
        RECT 111.710 118.715 112.045 119.685 ;
        RECT 112.215 118.715 112.385 119.855 ;
        RECT 112.555 119.515 114.585 119.685 ;
        RECT 111.710 118.045 111.880 118.715 ;
        RECT 112.555 118.545 112.725 119.515 ;
        RECT 112.050 118.215 112.305 118.545 ;
        RECT 112.530 118.215 112.725 118.545 ;
        RECT 112.895 119.175 114.020 119.345 ;
        RECT 112.135 118.045 112.305 118.215 ;
        RECT 112.895 118.045 113.065 119.175 ;
        RECT 111.710 117.475 111.965 118.045 ;
        RECT 112.135 117.875 113.065 118.045 ;
        RECT 113.235 118.835 114.245 119.005 ;
        RECT 113.235 118.035 113.405 118.835 ;
        RECT 113.610 118.155 113.885 118.635 ;
        RECT 113.605 117.985 113.885 118.155 ;
        RECT 112.890 117.840 113.065 117.875 ;
        RECT 112.135 117.305 112.465 117.705 ;
        RECT 112.890 117.475 113.420 117.840 ;
        RECT 113.610 117.475 113.885 117.985 ;
        RECT 114.055 117.475 114.245 118.835 ;
        RECT 114.415 118.850 114.585 119.515 ;
        RECT 114.755 119.095 114.925 119.855 ;
        RECT 115.160 119.095 115.675 119.505 ;
        RECT 114.415 118.660 115.165 118.850 ;
        RECT 115.335 118.285 115.675 119.095 ;
        RECT 115.845 118.765 117.515 119.855 ;
        RECT 114.445 118.115 115.675 118.285 ;
        RECT 114.425 117.305 114.935 117.840 ;
        RECT 115.155 117.510 115.400 118.115 ;
        RECT 115.845 118.075 116.595 118.595 ;
        RECT 116.765 118.245 117.515 118.765 ;
        RECT 117.690 118.905 117.955 119.675 ;
        RECT 118.125 119.135 118.455 119.855 ;
        RECT 118.645 119.315 118.905 119.675 ;
        RECT 119.075 119.485 119.405 119.855 ;
        RECT 119.575 119.315 119.835 119.675 ;
        RECT 118.645 119.085 119.835 119.315 ;
        RECT 120.405 118.905 120.695 119.675 ;
        RECT 120.995 119.185 121.165 119.685 ;
        RECT 121.335 119.355 121.665 119.855 ;
        RECT 120.995 119.015 121.660 119.185 ;
        RECT 115.845 117.305 117.515 118.075 ;
        RECT 117.690 117.485 118.025 118.905 ;
        RECT 118.200 118.725 120.695 118.905 ;
        RECT 118.200 118.035 118.425 118.725 ;
        RECT 118.625 118.215 118.905 118.545 ;
        RECT 119.085 118.215 119.660 118.545 ;
        RECT 119.840 118.215 120.275 118.545 ;
        RECT 120.455 118.215 120.725 118.545 ;
        RECT 120.910 118.195 121.260 118.845 ;
        RECT 118.200 117.845 120.685 118.035 ;
        RECT 121.430 118.025 121.660 119.015 ;
        RECT 118.205 117.305 118.950 117.675 ;
        RECT 119.515 117.485 119.770 117.845 ;
        RECT 119.950 117.305 120.280 117.675 ;
        RECT 120.460 117.485 120.685 117.845 ;
        RECT 120.995 117.855 121.660 118.025 ;
        RECT 120.995 117.565 121.165 117.855 ;
        RECT 121.335 117.305 121.665 117.685 ;
        RECT 121.835 117.565 122.020 119.685 ;
        RECT 122.260 119.395 122.525 119.855 ;
        RECT 122.695 119.260 122.945 119.685 ;
        RECT 123.155 119.410 124.260 119.580 ;
        RECT 122.640 119.130 122.945 119.260 ;
        RECT 122.190 117.935 122.470 118.885 ;
        RECT 122.640 118.025 122.810 119.130 ;
        RECT 122.980 118.345 123.220 118.940 ;
        RECT 123.390 118.875 123.920 119.240 ;
        RECT 123.390 118.175 123.560 118.875 ;
        RECT 124.090 118.795 124.260 119.410 ;
        RECT 124.430 119.055 124.600 119.855 ;
        RECT 124.770 119.355 125.020 119.685 ;
        RECT 125.245 119.385 126.130 119.555 ;
        RECT 124.090 118.705 124.600 118.795 ;
        RECT 122.640 117.895 122.865 118.025 ;
        RECT 123.035 117.955 123.560 118.175 ;
        RECT 123.730 118.535 124.600 118.705 ;
        RECT 122.275 117.305 122.525 117.765 ;
        RECT 122.695 117.755 122.865 117.895 ;
        RECT 123.730 117.755 123.900 118.535 ;
        RECT 124.430 118.465 124.600 118.535 ;
        RECT 124.110 118.285 124.310 118.315 ;
        RECT 124.770 118.285 124.940 119.355 ;
        RECT 125.110 118.465 125.300 119.185 ;
        RECT 124.110 117.985 124.940 118.285 ;
        RECT 125.470 118.255 125.790 119.215 ;
        RECT 122.695 117.585 123.030 117.755 ;
        RECT 123.225 117.585 123.900 117.755 ;
        RECT 124.220 117.305 124.590 117.805 ;
        RECT 124.770 117.755 124.940 117.985 ;
        RECT 125.325 117.925 125.790 118.255 ;
        RECT 125.960 118.545 126.130 119.385 ;
        RECT 126.310 119.355 126.625 119.855 ;
        RECT 126.855 119.125 127.195 119.685 ;
        RECT 126.300 118.750 127.195 119.125 ;
        RECT 127.365 118.845 127.535 119.855 ;
        RECT 127.005 118.545 127.195 118.750 ;
        RECT 127.705 118.795 128.035 119.640 ;
        RECT 127.705 118.715 128.095 118.795 ;
        RECT 128.265 118.765 129.935 119.855 ;
        RECT 130.655 119.235 130.825 119.665 ;
        RECT 130.995 119.405 131.325 119.855 ;
        RECT 130.655 119.005 131.330 119.235 ;
        RECT 127.880 118.665 128.095 118.715 ;
        RECT 125.960 118.215 126.835 118.545 ;
        RECT 127.005 118.215 127.755 118.545 ;
        RECT 125.960 117.755 126.130 118.215 ;
        RECT 127.005 118.045 127.205 118.215 ;
        RECT 127.925 118.085 128.095 118.665 ;
        RECT 127.870 118.045 128.095 118.085 ;
        RECT 124.770 117.585 125.175 117.755 ;
        RECT 125.345 117.585 126.130 117.755 ;
        RECT 126.405 117.305 126.615 117.835 ;
        RECT 126.875 117.520 127.205 118.045 ;
        RECT 127.715 117.960 128.095 118.045 ;
        RECT 128.265 118.075 129.015 118.595 ;
        RECT 129.185 118.245 129.935 118.765 ;
        RECT 127.375 117.305 127.545 117.915 ;
        RECT 127.715 117.525 128.045 117.960 ;
        RECT 128.265 117.305 129.935 118.075 ;
        RECT 130.625 117.985 130.925 118.835 ;
        RECT 131.095 118.355 131.330 119.005 ;
        RECT 131.500 118.695 131.785 119.640 ;
        RECT 131.965 119.385 132.650 119.855 ;
        RECT 131.960 118.865 132.655 119.175 ;
        RECT 132.830 118.800 133.135 119.585 ;
        RECT 131.500 118.545 132.360 118.695 ;
        RECT 131.500 118.525 132.785 118.545 ;
        RECT 131.095 118.025 131.630 118.355 ;
        RECT 131.800 118.165 132.785 118.525 ;
        RECT 131.095 117.875 131.315 118.025 ;
        RECT 130.570 117.305 130.905 117.810 ;
        RECT 131.075 117.500 131.315 117.875 ;
        RECT 131.800 117.830 131.970 118.165 ;
        RECT 132.960 117.995 133.135 118.800 ;
        RECT 133.325 118.690 133.615 119.855 ;
        RECT 133.790 118.905 134.055 119.675 ;
        RECT 134.225 119.135 134.555 119.855 ;
        RECT 134.745 119.315 135.005 119.675 ;
        RECT 135.175 119.485 135.505 119.855 ;
        RECT 135.675 119.315 135.935 119.675 ;
        RECT 134.745 119.085 135.935 119.315 ;
        RECT 136.505 118.905 136.795 119.675 ;
        RECT 137.555 119.185 137.725 119.685 ;
        RECT 137.895 119.355 138.225 119.855 ;
        RECT 137.555 119.015 138.220 119.185 ;
        RECT 131.595 117.635 131.970 117.830 ;
        RECT 131.595 117.490 131.765 117.635 ;
        RECT 132.330 117.305 132.725 117.800 ;
        RECT 132.895 117.475 133.135 117.995 ;
        RECT 133.325 117.305 133.615 118.030 ;
        RECT 133.790 117.485 134.125 118.905 ;
        RECT 134.300 118.725 136.795 118.905 ;
        RECT 134.300 118.035 134.525 118.725 ;
        RECT 134.725 118.215 135.005 118.545 ;
        RECT 135.185 118.215 135.760 118.545 ;
        RECT 135.940 118.215 136.375 118.545 ;
        RECT 136.555 118.215 136.825 118.545 ;
        RECT 137.470 118.195 137.820 118.845 ;
        RECT 134.300 117.845 136.785 118.035 ;
        RECT 137.990 118.025 138.220 119.015 ;
        RECT 134.305 117.305 135.050 117.675 ;
        RECT 135.615 117.485 135.870 117.845 ;
        RECT 136.050 117.305 136.380 117.675 ;
        RECT 136.560 117.485 136.785 117.845 ;
        RECT 137.555 117.855 138.220 118.025 ;
        RECT 137.555 117.565 137.725 117.855 ;
        RECT 137.895 117.305 138.225 117.685 ;
        RECT 138.395 117.565 138.580 119.685 ;
        RECT 138.820 119.395 139.085 119.855 ;
        RECT 139.255 119.260 139.505 119.685 ;
        RECT 139.715 119.410 140.820 119.580 ;
        RECT 139.200 119.130 139.505 119.260 ;
        RECT 138.750 117.935 139.030 118.885 ;
        RECT 139.200 118.025 139.370 119.130 ;
        RECT 139.540 118.345 139.780 118.940 ;
        RECT 139.950 118.875 140.480 119.240 ;
        RECT 139.950 118.175 140.120 118.875 ;
        RECT 140.650 118.795 140.820 119.410 ;
        RECT 140.990 119.055 141.160 119.855 ;
        RECT 141.330 119.355 141.580 119.685 ;
        RECT 141.805 119.385 142.690 119.555 ;
        RECT 140.650 118.705 141.160 118.795 ;
        RECT 139.200 117.895 139.425 118.025 ;
        RECT 139.595 117.955 140.120 118.175 ;
        RECT 140.290 118.535 141.160 118.705 ;
        RECT 138.835 117.305 139.085 117.765 ;
        RECT 139.255 117.755 139.425 117.895 ;
        RECT 140.290 117.755 140.460 118.535 ;
        RECT 140.990 118.465 141.160 118.535 ;
        RECT 140.670 118.285 140.870 118.315 ;
        RECT 141.330 118.285 141.500 119.355 ;
        RECT 141.670 118.465 141.860 119.185 ;
        RECT 140.670 117.985 141.500 118.285 ;
        RECT 142.030 118.255 142.350 119.215 ;
        RECT 139.255 117.585 139.590 117.755 ;
        RECT 139.785 117.585 140.460 117.755 ;
        RECT 140.780 117.305 141.150 117.805 ;
        RECT 141.330 117.755 141.500 117.985 ;
        RECT 141.885 117.925 142.350 118.255 ;
        RECT 142.520 118.545 142.690 119.385 ;
        RECT 142.870 119.355 143.185 119.855 ;
        RECT 143.415 119.125 143.755 119.685 ;
        RECT 142.860 118.750 143.755 119.125 ;
        RECT 143.925 118.845 144.095 119.855 ;
        RECT 143.565 118.545 143.755 118.750 ;
        RECT 144.265 118.795 144.595 119.640 ;
        RECT 144.265 118.715 144.655 118.795 ;
        RECT 144.440 118.665 144.655 118.715 ;
        RECT 142.520 118.215 143.395 118.545 ;
        RECT 143.565 118.215 144.315 118.545 ;
        RECT 142.520 117.755 142.690 118.215 ;
        RECT 143.565 118.045 143.765 118.215 ;
        RECT 144.485 118.085 144.655 118.665 ;
        RECT 145.745 118.765 146.955 119.855 ;
        RECT 145.745 118.225 146.265 118.765 ;
        RECT 144.430 118.045 144.655 118.085 ;
        RECT 146.435 118.055 146.955 118.595 ;
        RECT 141.330 117.585 141.735 117.755 ;
        RECT 141.905 117.585 142.690 117.755 ;
        RECT 142.965 117.305 143.175 117.835 ;
        RECT 143.435 117.520 143.765 118.045 ;
        RECT 144.275 117.960 144.655 118.045 ;
        RECT 143.935 117.305 144.105 117.915 ;
        RECT 144.275 117.525 144.605 117.960 ;
        RECT 145.745 117.305 146.955 118.055 ;
        RECT 17.320 117.135 147.040 117.305 ;
        RECT 17.405 116.385 18.615 117.135 ;
        RECT 19.705 116.635 19.965 116.965 ;
        RECT 20.175 116.655 20.450 117.135 ;
        RECT 17.405 115.845 17.925 116.385 ;
        RECT 18.095 115.675 18.615 116.215 ;
        RECT 17.405 114.585 18.615 115.675 ;
        RECT 19.705 115.725 19.875 116.635 ;
        RECT 20.660 116.565 20.865 116.965 ;
        RECT 21.035 116.735 21.370 117.135 ;
        RECT 20.045 115.895 20.405 116.475 ;
        RECT 20.660 116.395 21.345 116.565 ;
        RECT 20.585 115.725 20.835 116.225 ;
        RECT 19.705 115.555 20.835 115.725 ;
        RECT 19.705 114.785 19.975 115.555 ;
        RECT 21.005 115.365 21.345 116.395 ;
        RECT 21.545 116.385 22.755 117.135 ;
        RECT 22.975 116.480 23.305 116.915 ;
        RECT 23.475 116.525 23.645 117.135 ;
        RECT 22.925 116.395 23.305 116.480 ;
        RECT 23.815 116.395 24.145 116.920 ;
        RECT 24.405 116.605 24.615 117.135 ;
        RECT 24.890 116.685 25.675 116.855 ;
        RECT 25.845 116.685 26.250 116.855 ;
        RECT 21.545 115.845 22.065 116.385 ;
        RECT 22.925 116.355 23.150 116.395 ;
        RECT 22.235 115.675 22.755 116.215 ;
        RECT 20.145 114.585 20.475 115.365 ;
        RECT 20.680 115.190 21.345 115.365 ;
        RECT 20.680 114.785 20.865 115.190 ;
        RECT 21.035 114.585 21.370 115.010 ;
        RECT 21.545 114.585 22.755 115.675 ;
        RECT 22.925 115.775 23.095 116.355 ;
        RECT 23.815 116.225 24.015 116.395 ;
        RECT 24.890 116.225 25.060 116.685 ;
        RECT 23.265 115.895 24.015 116.225 ;
        RECT 24.185 115.895 25.060 116.225 ;
        RECT 22.925 115.725 23.140 115.775 ;
        RECT 22.925 115.645 23.315 115.725 ;
        RECT 22.985 114.800 23.315 115.645 ;
        RECT 23.825 115.690 24.015 115.895 ;
        RECT 23.485 114.585 23.655 115.595 ;
        RECT 23.825 115.315 24.720 115.690 ;
        RECT 23.825 114.755 24.165 115.315 ;
        RECT 24.395 114.585 24.710 115.085 ;
        RECT 24.890 115.055 25.060 115.895 ;
        RECT 25.230 116.185 25.695 116.515 ;
        RECT 26.080 116.455 26.250 116.685 ;
        RECT 26.430 116.635 26.800 117.135 ;
        RECT 27.120 116.685 27.795 116.855 ;
        RECT 27.990 116.685 28.325 116.855 ;
        RECT 25.230 115.225 25.550 116.185 ;
        RECT 26.080 116.155 26.910 116.455 ;
        RECT 25.720 115.255 25.910 115.975 ;
        RECT 26.080 115.085 26.250 116.155 ;
        RECT 26.710 116.125 26.910 116.155 ;
        RECT 26.420 115.905 26.590 115.975 ;
        RECT 27.120 115.905 27.290 116.685 ;
        RECT 28.155 116.545 28.325 116.685 ;
        RECT 28.495 116.675 28.745 117.135 ;
        RECT 26.420 115.735 27.290 115.905 ;
        RECT 27.460 116.265 27.985 116.485 ;
        RECT 28.155 116.415 28.380 116.545 ;
        RECT 26.420 115.645 26.930 115.735 ;
        RECT 24.890 114.885 25.775 115.055 ;
        RECT 26.000 114.755 26.250 115.085 ;
        RECT 26.420 114.585 26.590 115.385 ;
        RECT 26.760 115.030 26.930 115.645 ;
        RECT 27.460 115.565 27.630 116.265 ;
        RECT 27.100 115.200 27.630 115.565 ;
        RECT 27.800 115.500 28.040 116.095 ;
        RECT 28.210 115.310 28.380 116.415 ;
        RECT 28.550 115.555 28.830 116.505 ;
        RECT 28.075 115.180 28.380 115.310 ;
        RECT 26.760 114.860 27.865 115.030 ;
        RECT 28.075 114.755 28.325 115.180 ;
        RECT 28.495 114.585 28.760 115.045 ;
        RECT 29.000 114.755 29.185 116.875 ;
        RECT 29.355 116.755 29.685 117.135 ;
        RECT 29.855 116.585 30.025 116.875 ;
        RECT 29.360 116.415 30.025 116.585 ;
        RECT 29.360 115.425 29.590 116.415 ;
        RECT 30.285 116.335 30.625 116.965 ;
        RECT 30.915 116.675 31.085 117.135 ;
        RECT 31.355 116.505 31.685 116.950 ;
        RECT 29.760 115.595 30.110 116.245 ;
        RECT 30.285 115.765 30.555 116.335 ;
        RECT 30.935 116.315 31.685 116.505 ;
        RECT 31.855 116.485 32.025 116.805 ;
        RECT 32.250 116.675 32.580 117.135 ;
        RECT 32.780 116.485 33.110 116.965 ;
        RECT 33.325 116.675 33.655 117.135 ;
        RECT 33.825 116.485 34.155 116.965 ;
        RECT 34.425 116.590 39.770 117.135 ;
        RECT 31.855 116.315 34.155 116.485 ;
        RECT 30.935 116.145 31.305 116.315 ;
        RECT 30.725 115.935 31.305 116.145 ;
        RECT 31.475 115.935 31.895 116.145 ;
        RECT 31.045 115.765 31.305 115.935 ;
        RECT 29.360 115.255 30.025 115.425 ;
        RECT 29.355 114.585 29.685 115.085 ;
        RECT 29.855 114.755 30.025 115.255 ;
        RECT 30.285 114.755 30.810 115.765 ;
        RECT 31.045 115.475 31.795 115.765 ;
        RECT 31.045 114.585 31.375 115.305 ;
        RECT 31.545 114.755 31.795 115.475 ;
        RECT 32.065 114.830 32.395 116.145 ;
        RECT 32.605 114.830 32.935 116.145 ;
        RECT 33.105 114.830 33.475 116.145 ;
        RECT 33.685 115.895 34.195 116.145 ;
        RECT 36.010 115.760 36.350 116.590 ;
        RECT 39.945 116.365 42.535 117.135 ;
        RECT 43.165 116.410 43.455 117.135 ;
        RECT 43.625 116.590 48.970 117.135 ;
        RECT 49.145 116.590 54.490 117.135 ;
        RECT 54.665 116.590 60.010 117.135 ;
        RECT 60.185 116.590 65.530 117.135 ;
        RECT 33.805 114.585 34.135 115.705 ;
        RECT 37.830 115.020 38.180 116.270 ;
        RECT 39.945 115.845 41.155 116.365 ;
        RECT 41.325 115.675 42.535 116.195 ;
        RECT 45.210 115.760 45.550 116.590 ;
        RECT 34.425 114.585 39.770 115.020 ;
        RECT 39.945 114.585 42.535 115.675 ;
        RECT 43.165 114.585 43.455 115.750 ;
        RECT 47.030 115.020 47.380 116.270 ;
        RECT 50.730 115.760 51.070 116.590 ;
        RECT 52.550 115.020 52.900 116.270 ;
        RECT 56.250 115.760 56.590 116.590 ;
        RECT 58.070 115.020 58.420 116.270 ;
        RECT 61.770 115.760 62.110 116.590 ;
        RECT 65.705 116.365 68.295 117.135 ;
        RECT 68.925 116.410 69.215 117.135 ;
        RECT 69.385 116.590 74.730 117.135 ;
        RECT 74.905 116.590 80.250 117.135 ;
        RECT 80.425 116.590 85.770 117.135 ;
        RECT 86.875 116.645 87.205 117.135 ;
        RECT 63.590 115.020 63.940 116.270 ;
        RECT 65.705 115.845 66.915 116.365 ;
        RECT 67.085 115.675 68.295 116.195 ;
        RECT 70.970 115.760 71.310 116.590 ;
        RECT 43.625 114.585 48.970 115.020 ;
        RECT 49.145 114.585 54.490 115.020 ;
        RECT 54.665 114.585 60.010 115.020 ;
        RECT 60.185 114.585 65.530 115.020 ;
        RECT 65.705 114.585 68.295 115.675 ;
        RECT 68.925 114.585 69.215 115.750 ;
        RECT 72.790 115.020 73.140 116.270 ;
        RECT 76.490 115.760 76.830 116.590 ;
        RECT 78.310 115.020 78.660 116.270 ;
        RECT 82.010 115.760 82.350 116.590 ;
        RECT 87.375 116.540 87.995 116.965 ;
        RECT 83.830 115.020 84.180 116.270 ;
        RECT 86.865 115.895 87.205 116.475 ;
        RECT 87.375 116.205 87.735 116.540 ;
        RECT 88.455 116.445 88.785 117.135 ;
        RECT 89.685 116.675 89.930 117.135 ;
        RECT 87.375 115.925 88.795 116.205 ;
        RECT 69.385 114.585 74.730 115.020 ;
        RECT 74.905 114.585 80.250 115.020 ;
        RECT 80.425 114.585 85.770 115.020 ;
        RECT 86.875 114.585 87.205 115.725 ;
        RECT 87.375 114.755 87.735 115.925 ;
        RECT 87.935 114.585 88.265 115.755 ;
        RECT 88.465 114.755 88.795 115.925 ;
        RECT 89.625 115.895 89.940 116.505 ;
        RECT 90.110 116.145 90.360 116.955 ;
        RECT 90.530 116.610 90.790 117.135 ;
        RECT 90.960 116.485 91.220 116.940 ;
        RECT 91.390 116.655 91.650 117.135 ;
        RECT 91.820 116.485 92.080 116.940 ;
        RECT 92.250 116.655 92.510 117.135 ;
        RECT 92.680 116.485 92.940 116.940 ;
        RECT 93.110 116.655 93.370 117.135 ;
        RECT 93.540 116.485 93.800 116.940 ;
        RECT 93.970 116.655 94.270 117.135 ;
        RECT 90.960 116.315 94.270 116.485 ;
        RECT 94.685 116.410 94.975 117.135 ;
        RECT 95.235 116.585 95.405 116.875 ;
        RECT 95.575 116.755 95.905 117.135 ;
        RECT 95.235 116.415 95.900 116.585 ;
        RECT 90.110 115.895 93.130 116.145 ;
        RECT 88.995 114.585 89.325 115.755 ;
        RECT 89.635 114.585 89.930 115.695 ;
        RECT 90.110 114.760 90.360 115.895 ;
        RECT 93.300 115.725 94.270 116.315 ;
        RECT 90.530 114.585 90.790 115.695 ;
        RECT 90.960 115.485 94.270 115.725 ;
        RECT 90.960 114.760 91.220 115.485 ;
        RECT 91.390 114.585 91.650 115.315 ;
        RECT 91.820 114.760 92.080 115.485 ;
        RECT 92.250 114.585 92.510 115.315 ;
        RECT 92.680 114.760 92.940 115.485 ;
        RECT 93.110 114.585 93.370 115.315 ;
        RECT 93.540 114.760 93.800 115.485 ;
        RECT 93.970 114.585 94.265 115.315 ;
        RECT 94.685 114.585 94.975 115.750 ;
        RECT 95.150 115.595 95.500 116.245 ;
        RECT 95.670 115.425 95.900 116.415 ;
        RECT 95.235 115.255 95.900 115.425 ;
        RECT 95.235 114.755 95.405 115.255 ;
        RECT 95.575 114.585 95.905 115.085 ;
        RECT 96.075 114.755 96.260 116.875 ;
        RECT 96.515 116.675 96.765 117.135 ;
        RECT 96.935 116.685 97.270 116.855 ;
        RECT 97.465 116.685 98.140 116.855 ;
        RECT 96.935 116.545 97.105 116.685 ;
        RECT 96.430 115.555 96.710 116.505 ;
        RECT 96.880 116.415 97.105 116.545 ;
        RECT 96.880 115.310 97.050 116.415 ;
        RECT 97.275 116.265 97.800 116.485 ;
        RECT 97.220 115.500 97.460 116.095 ;
        RECT 97.630 115.565 97.800 116.265 ;
        RECT 97.970 115.905 98.140 116.685 ;
        RECT 98.460 116.635 98.830 117.135 ;
        RECT 99.010 116.685 99.415 116.855 ;
        RECT 99.585 116.685 100.370 116.855 ;
        RECT 99.010 116.455 99.180 116.685 ;
        RECT 98.350 116.155 99.180 116.455 ;
        RECT 99.565 116.185 100.030 116.515 ;
        RECT 98.350 116.125 98.550 116.155 ;
        RECT 98.670 115.905 98.840 115.975 ;
        RECT 97.970 115.735 98.840 115.905 ;
        RECT 98.330 115.645 98.840 115.735 ;
        RECT 96.880 115.180 97.185 115.310 ;
        RECT 97.630 115.200 98.160 115.565 ;
        RECT 96.500 114.585 96.765 115.045 ;
        RECT 96.935 114.755 97.185 115.180 ;
        RECT 98.330 115.030 98.500 115.645 ;
        RECT 97.395 114.860 98.500 115.030 ;
        RECT 98.670 114.585 98.840 115.385 ;
        RECT 99.010 115.085 99.180 116.155 ;
        RECT 99.350 115.255 99.540 115.975 ;
        RECT 99.710 115.225 100.030 116.185 ;
        RECT 100.200 116.225 100.370 116.685 ;
        RECT 100.645 116.605 100.855 117.135 ;
        RECT 101.115 116.395 101.445 116.920 ;
        RECT 101.615 116.525 101.785 117.135 ;
        RECT 101.955 116.480 102.285 116.915 ;
        RECT 102.575 116.735 102.905 117.135 ;
        RECT 103.075 116.565 103.245 116.835 ;
        RECT 103.415 116.735 103.745 117.135 ;
        RECT 103.915 116.565 104.170 116.835 ;
        RECT 104.345 116.590 109.690 117.135 ;
        RECT 101.955 116.395 102.335 116.480 ;
        RECT 101.245 116.225 101.445 116.395 ;
        RECT 102.110 116.355 102.335 116.395 ;
        RECT 100.200 115.895 101.075 116.225 ;
        RECT 101.245 115.895 101.995 116.225 ;
        RECT 99.010 114.755 99.260 115.085 ;
        RECT 100.200 115.055 100.370 115.895 ;
        RECT 101.245 115.690 101.435 115.895 ;
        RECT 102.165 115.775 102.335 116.355 ;
        RECT 102.120 115.725 102.335 115.775 ;
        RECT 100.540 115.315 101.435 115.690 ;
        RECT 101.945 115.645 102.335 115.725 ;
        RECT 99.485 114.885 100.370 115.055 ;
        RECT 100.550 114.585 100.865 115.085 ;
        RECT 101.095 114.755 101.435 115.315 ;
        RECT 101.605 114.585 101.775 115.595 ;
        RECT 101.945 114.800 102.275 115.645 ;
        RECT 102.505 115.555 102.775 116.565 ;
        RECT 102.945 116.395 104.170 116.565 ;
        RECT 102.945 115.725 103.115 116.395 ;
        RECT 103.285 115.895 103.665 116.225 ;
        RECT 103.835 115.895 104.170 116.225 ;
        RECT 102.945 115.555 103.260 115.725 ;
        RECT 102.510 114.585 102.825 115.385 ;
        RECT 103.090 114.940 103.260 115.555 ;
        RECT 103.430 115.215 103.665 115.895 ;
        RECT 105.930 115.760 106.270 116.590 ;
        RECT 109.865 116.365 113.375 117.135 ;
        RECT 114.010 116.395 114.265 116.965 ;
        RECT 114.435 116.735 114.765 117.135 ;
        RECT 115.190 116.600 115.720 116.965 ;
        RECT 115.910 116.795 116.185 116.965 ;
        RECT 115.905 116.625 116.185 116.795 ;
        RECT 115.190 116.565 115.365 116.600 ;
        RECT 114.435 116.395 115.365 116.565 ;
        RECT 103.835 114.940 104.170 115.725 ;
        RECT 107.750 115.020 108.100 116.270 ;
        RECT 109.865 115.845 111.515 116.365 ;
        RECT 111.685 115.675 113.375 116.195 ;
        RECT 103.090 114.770 104.170 114.940 ;
        RECT 104.345 114.585 109.690 115.020 ;
        RECT 109.865 114.585 113.375 115.675 ;
        RECT 114.010 115.725 114.180 116.395 ;
        RECT 114.435 116.225 114.605 116.395 ;
        RECT 114.350 115.895 114.605 116.225 ;
        RECT 114.830 115.895 115.025 116.225 ;
        RECT 114.010 114.755 114.345 115.725 ;
        RECT 114.515 114.585 114.685 115.725 ;
        RECT 114.855 114.925 115.025 115.895 ;
        RECT 115.195 115.265 115.365 116.395 ;
        RECT 115.535 115.605 115.705 116.405 ;
        RECT 115.910 115.805 116.185 116.625 ;
        RECT 116.355 115.605 116.545 116.965 ;
        RECT 116.725 116.600 117.235 117.135 ;
        RECT 117.455 116.325 117.700 116.930 ;
        RECT 118.145 116.365 119.815 117.135 ;
        RECT 120.445 116.410 120.735 117.135 ;
        RECT 121.885 116.675 122.130 117.135 ;
        RECT 116.745 116.155 117.975 116.325 ;
        RECT 115.535 115.435 116.545 115.605 ;
        RECT 116.715 115.590 117.465 115.780 ;
        RECT 115.195 115.095 116.320 115.265 ;
        RECT 116.715 114.925 116.885 115.590 ;
        RECT 117.635 115.345 117.975 116.155 ;
        RECT 118.145 115.845 118.895 116.365 ;
        RECT 119.065 115.675 119.815 116.195 ;
        RECT 121.825 115.895 122.140 116.505 ;
        RECT 122.310 116.145 122.560 116.955 ;
        RECT 122.730 116.610 122.990 117.135 ;
        RECT 123.160 116.485 123.420 116.940 ;
        RECT 123.590 116.655 123.850 117.135 ;
        RECT 124.020 116.485 124.280 116.940 ;
        RECT 124.450 116.655 124.710 117.135 ;
        RECT 124.880 116.485 125.140 116.940 ;
        RECT 125.310 116.655 125.570 117.135 ;
        RECT 125.740 116.485 126.000 116.940 ;
        RECT 126.170 116.655 126.470 117.135 ;
        RECT 123.160 116.315 126.470 116.485 ;
        RECT 122.310 115.895 125.330 116.145 ;
        RECT 114.855 114.755 116.885 114.925 ;
        RECT 117.055 114.585 117.225 115.345 ;
        RECT 117.460 114.935 117.975 115.345 ;
        RECT 118.145 114.585 119.815 115.675 ;
        RECT 120.445 114.585 120.735 115.750 ;
        RECT 121.835 114.585 122.130 115.695 ;
        RECT 122.310 114.760 122.560 115.895 ;
        RECT 125.500 115.725 126.470 116.315 ;
        RECT 122.730 114.585 122.990 115.695 ;
        RECT 123.160 115.485 126.470 115.725 ;
        RECT 126.890 116.395 127.145 116.965 ;
        RECT 127.315 116.735 127.645 117.135 ;
        RECT 128.070 116.600 128.600 116.965 ;
        RECT 128.790 116.795 129.065 116.965 ;
        RECT 128.785 116.625 129.065 116.795 ;
        RECT 128.070 116.565 128.245 116.600 ;
        RECT 127.315 116.395 128.245 116.565 ;
        RECT 126.890 115.725 127.060 116.395 ;
        RECT 127.315 116.225 127.485 116.395 ;
        RECT 127.230 115.895 127.485 116.225 ;
        RECT 127.710 115.895 127.905 116.225 ;
        RECT 123.160 114.760 123.420 115.485 ;
        RECT 123.590 114.585 123.850 115.315 ;
        RECT 124.020 114.760 124.280 115.485 ;
        RECT 124.450 114.585 124.710 115.315 ;
        RECT 124.880 114.760 125.140 115.485 ;
        RECT 125.310 114.585 125.570 115.315 ;
        RECT 125.740 114.760 126.000 115.485 ;
        RECT 126.170 114.585 126.465 115.315 ;
        RECT 126.890 114.755 127.225 115.725 ;
        RECT 127.395 114.585 127.565 115.725 ;
        RECT 127.735 114.925 127.905 115.895 ;
        RECT 128.075 115.265 128.245 116.395 ;
        RECT 128.415 115.605 128.585 116.405 ;
        RECT 128.790 115.805 129.065 116.625 ;
        RECT 129.235 115.605 129.425 116.965 ;
        RECT 129.605 116.600 130.115 117.135 ;
        RECT 130.335 116.325 130.580 116.930 ;
        RECT 131.025 116.385 132.235 117.135 ;
        RECT 132.495 116.585 132.665 116.875 ;
        RECT 132.835 116.755 133.165 117.135 ;
        RECT 132.495 116.415 133.160 116.585 ;
        RECT 129.625 116.155 130.855 116.325 ;
        RECT 128.415 115.435 129.425 115.605 ;
        RECT 129.595 115.590 130.345 115.780 ;
        RECT 128.075 115.095 129.200 115.265 ;
        RECT 129.595 114.925 129.765 115.590 ;
        RECT 130.515 115.345 130.855 116.155 ;
        RECT 131.025 115.845 131.545 116.385 ;
        RECT 131.715 115.675 132.235 116.215 ;
        RECT 127.735 114.755 129.765 114.925 ;
        RECT 129.935 114.585 130.105 115.345 ;
        RECT 130.340 114.935 130.855 115.345 ;
        RECT 131.025 114.585 132.235 115.675 ;
        RECT 132.410 115.595 132.760 116.245 ;
        RECT 132.930 115.425 133.160 116.415 ;
        RECT 132.495 115.255 133.160 115.425 ;
        RECT 132.495 114.755 132.665 115.255 ;
        RECT 132.835 114.585 133.165 115.085 ;
        RECT 133.335 114.755 133.520 116.875 ;
        RECT 133.775 116.675 134.025 117.135 ;
        RECT 134.195 116.685 134.530 116.855 ;
        RECT 134.725 116.685 135.400 116.855 ;
        RECT 134.195 116.545 134.365 116.685 ;
        RECT 133.690 115.555 133.970 116.505 ;
        RECT 134.140 116.415 134.365 116.545 ;
        RECT 134.140 115.310 134.310 116.415 ;
        RECT 134.535 116.265 135.060 116.485 ;
        RECT 134.480 115.500 134.720 116.095 ;
        RECT 134.890 115.565 135.060 116.265 ;
        RECT 135.230 115.905 135.400 116.685 ;
        RECT 135.720 116.635 136.090 117.135 ;
        RECT 136.270 116.685 136.675 116.855 ;
        RECT 136.845 116.685 137.630 116.855 ;
        RECT 136.270 116.455 136.440 116.685 ;
        RECT 135.610 116.155 136.440 116.455 ;
        RECT 136.825 116.185 137.290 116.515 ;
        RECT 135.610 116.125 135.810 116.155 ;
        RECT 135.930 115.905 136.100 115.975 ;
        RECT 135.230 115.735 136.100 115.905 ;
        RECT 135.590 115.645 136.100 115.735 ;
        RECT 134.140 115.180 134.445 115.310 ;
        RECT 134.890 115.200 135.420 115.565 ;
        RECT 133.760 114.585 134.025 115.045 ;
        RECT 134.195 114.755 134.445 115.180 ;
        RECT 135.590 115.030 135.760 115.645 ;
        RECT 134.655 114.860 135.760 115.030 ;
        RECT 135.930 114.585 136.100 115.385 ;
        RECT 136.270 115.085 136.440 116.155 ;
        RECT 136.610 115.255 136.800 115.975 ;
        RECT 136.970 115.225 137.290 116.185 ;
        RECT 137.460 116.225 137.630 116.685 ;
        RECT 137.905 116.605 138.115 117.135 ;
        RECT 138.375 116.395 138.705 116.920 ;
        RECT 138.875 116.525 139.045 117.135 ;
        RECT 139.215 116.480 139.545 116.915 ;
        RECT 139.215 116.395 139.595 116.480 ;
        RECT 138.505 116.225 138.705 116.395 ;
        RECT 139.370 116.355 139.595 116.395 ;
        RECT 137.460 115.895 138.335 116.225 ;
        RECT 138.505 115.895 139.255 116.225 ;
        RECT 136.270 114.755 136.520 115.085 ;
        RECT 137.460 115.055 137.630 115.895 ;
        RECT 138.505 115.690 138.695 115.895 ;
        RECT 139.425 115.775 139.595 116.355 ;
        RECT 139.765 116.365 141.435 117.135 ;
        RECT 142.155 116.585 142.325 116.965 ;
        RECT 142.540 116.755 142.870 117.135 ;
        RECT 142.155 116.415 142.870 116.585 ;
        RECT 139.765 115.845 140.515 116.365 ;
        RECT 139.380 115.725 139.595 115.775 ;
        RECT 137.800 115.315 138.695 115.690 ;
        RECT 139.205 115.645 139.595 115.725 ;
        RECT 140.685 115.675 141.435 116.195 ;
        RECT 142.065 115.865 142.420 116.235 ;
        RECT 142.700 116.225 142.870 116.415 ;
        RECT 143.040 116.390 143.295 116.965 ;
        RECT 142.700 115.895 142.955 116.225 ;
        RECT 142.700 115.685 142.870 115.895 ;
        RECT 136.745 114.885 137.630 115.055 ;
        RECT 137.810 114.585 138.125 115.085 ;
        RECT 138.355 114.755 138.695 115.315 ;
        RECT 138.865 114.585 139.035 115.595 ;
        RECT 139.205 114.800 139.535 115.645 ;
        RECT 139.765 114.585 141.435 115.675 ;
        RECT 142.155 115.515 142.870 115.685 ;
        RECT 143.125 115.660 143.295 116.390 ;
        RECT 143.470 116.295 143.730 117.135 ;
        RECT 143.995 116.585 144.165 116.965 ;
        RECT 144.380 116.755 144.710 117.135 ;
        RECT 143.995 116.415 144.710 116.585 ;
        RECT 143.905 115.865 144.260 116.235 ;
        RECT 144.540 116.225 144.710 116.415 ;
        RECT 144.880 116.390 145.135 116.965 ;
        RECT 144.540 115.895 144.795 116.225 ;
        RECT 142.155 114.755 142.325 115.515 ;
        RECT 142.540 114.585 142.870 115.345 ;
        RECT 143.040 114.755 143.295 115.660 ;
        RECT 143.470 114.585 143.730 115.735 ;
        RECT 144.540 115.685 144.710 115.895 ;
        RECT 143.995 115.515 144.710 115.685 ;
        RECT 144.965 115.660 145.135 116.390 ;
        RECT 145.310 116.295 145.570 117.135 ;
        RECT 145.745 116.385 146.955 117.135 ;
        RECT 143.995 114.755 144.165 115.515 ;
        RECT 144.380 114.585 144.710 115.345 ;
        RECT 144.880 114.755 145.135 115.660 ;
        RECT 145.310 114.585 145.570 115.735 ;
        RECT 145.745 115.675 146.265 116.215 ;
        RECT 146.435 115.845 146.955 116.385 ;
        RECT 145.745 114.585 146.955 115.675 ;
        RECT 17.320 114.415 147.040 114.585 ;
        RECT 17.405 113.325 18.615 114.415 ;
        RECT 19.335 113.745 19.505 114.245 ;
        RECT 19.675 113.915 20.005 114.415 ;
        RECT 19.335 113.575 20.000 113.745 ;
        RECT 17.405 112.615 17.925 113.155 ;
        RECT 18.095 112.785 18.615 113.325 ;
        RECT 19.250 112.755 19.600 113.405 ;
        RECT 17.405 111.865 18.615 112.615 ;
        RECT 19.770 112.585 20.000 113.575 ;
        RECT 19.335 112.415 20.000 112.585 ;
        RECT 19.335 112.125 19.505 112.415 ;
        RECT 19.675 111.865 20.005 112.245 ;
        RECT 20.175 112.125 20.360 114.245 ;
        RECT 20.600 113.955 20.865 114.415 ;
        RECT 21.035 113.820 21.285 114.245 ;
        RECT 21.495 113.970 22.600 114.140 ;
        RECT 20.980 113.690 21.285 113.820 ;
        RECT 20.530 112.495 20.810 113.445 ;
        RECT 20.980 112.585 21.150 113.690 ;
        RECT 21.320 112.905 21.560 113.500 ;
        RECT 21.730 113.435 22.260 113.800 ;
        RECT 21.730 112.735 21.900 113.435 ;
        RECT 22.430 113.355 22.600 113.970 ;
        RECT 22.770 113.615 22.940 114.415 ;
        RECT 23.110 113.915 23.360 114.245 ;
        RECT 23.585 113.945 24.470 114.115 ;
        RECT 22.430 113.265 22.940 113.355 ;
        RECT 20.980 112.455 21.205 112.585 ;
        RECT 21.375 112.515 21.900 112.735 ;
        RECT 22.070 113.095 22.940 113.265 ;
        RECT 20.615 111.865 20.865 112.325 ;
        RECT 21.035 112.315 21.205 112.455 ;
        RECT 22.070 112.315 22.240 113.095 ;
        RECT 22.770 113.025 22.940 113.095 ;
        RECT 22.450 112.845 22.650 112.875 ;
        RECT 23.110 112.845 23.280 113.915 ;
        RECT 23.450 113.025 23.640 113.745 ;
        RECT 22.450 112.545 23.280 112.845 ;
        RECT 23.810 112.815 24.130 113.775 ;
        RECT 21.035 112.145 21.370 112.315 ;
        RECT 21.565 112.145 22.240 112.315 ;
        RECT 22.560 111.865 22.930 112.365 ;
        RECT 23.110 112.315 23.280 112.545 ;
        RECT 23.665 112.485 24.130 112.815 ;
        RECT 24.300 113.105 24.470 113.945 ;
        RECT 24.650 113.915 24.965 114.415 ;
        RECT 25.195 113.685 25.535 114.245 ;
        RECT 24.640 113.310 25.535 113.685 ;
        RECT 25.705 113.405 25.875 114.415 ;
        RECT 25.345 113.105 25.535 113.310 ;
        RECT 26.045 113.355 26.375 114.200 ;
        RECT 27.065 113.460 27.335 114.415 ;
        RECT 27.520 113.360 27.825 114.145 ;
        RECT 28.005 113.945 28.690 114.415 ;
        RECT 28.000 113.425 28.695 113.735 ;
        RECT 26.045 113.275 26.435 113.355 ;
        RECT 26.220 113.225 26.435 113.275 ;
        RECT 24.300 112.775 25.175 113.105 ;
        RECT 25.345 112.775 26.095 113.105 ;
        RECT 24.300 112.315 24.470 112.775 ;
        RECT 25.345 112.605 25.545 112.775 ;
        RECT 26.265 112.645 26.435 113.225 ;
        RECT 26.210 112.605 26.435 112.645 ;
        RECT 23.110 112.145 23.515 112.315 ;
        RECT 23.685 112.145 24.470 112.315 ;
        RECT 24.745 111.865 24.955 112.395 ;
        RECT 25.215 112.080 25.545 112.605 ;
        RECT 26.055 112.520 26.435 112.605 ;
        RECT 27.520 112.555 27.695 113.360 ;
        RECT 28.870 113.255 29.155 114.200 ;
        RECT 29.355 113.965 29.685 114.415 ;
        RECT 29.855 113.795 30.025 114.225 ;
        RECT 28.295 113.105 29.155 113.255 ;
        RECT 27.865 113.085 29.155 113.105 ;
        RECT 29.345 113.565 30.025 113.795 ;
        RECT 27.865 112.725 28.855 113.085 ;
        RECT 29.345 112.915 29.580 113.565 ;
        RECT 25.715 111.865 25.885 112.475 ;
        RECT 26.055 112.085 26.385 112.520 ;
        RECT 27.065 111.865 27.335 112.500 ;
        RECT 27.520 112.035 27.755 112.555 ;
        RECT 28.685 112.390 28.855 112.725 ;
        RECT 29.025 112.585 29.580 112.915 ;
        RECT 29.365 112.435 29.580 112.585 ;
        RECT 29.750 112.715 30.050 113.395 ;
        RECT 30.285 113.250 30.575 114.415 ;
        RECT 30.835 113.745 31.005 114.245 ;
        RECT 31.175 113.915 31.505 114.415 ;
        RECT 30.835 113.575 31.500 113.745 ;
        RECT 30.750 112.755 31.100 113.405 ;
        RECT 29.750 112.545 30.055 112.715 ;
        RECT 27.925 111.865 28.325 112.360 ;
        RECT 28.685 112.195 29.085 112.390 ;
        RECT 28.915 112.050 29.085 112.195 ;
        RECT 29.365 112.060 29.605 112.435 ;
        RECT 29.775 111.865 30.105 112.370 ;
        RECT 30.285 111.865 30.575 112.590 ;
        RECT 31.270 112.585 31.500 113.575 ;
        RECT 30.835 112.415 31.500 112.585 ;
        RECT 30.835 112.125 31.005 112.415 ;
        RECT 31.175 111.865 31.505 112.245 ;
        RECT 31.675 112.125 31.860 114.245 ;
        RECT 32.100 113.955 32.365 114.415 ;
        RECT 32.535 113.820 32.785 114.245 ;
        RECT 32.995 113.970 34.100 114.140 ;
        RECT 32.480 113.690 32.785 113.820 ;
        RECT 32.030 112.495 32.310 113.445 ;
        RECT 32.480 112.585 32.650 113.690 ;
        RECT 32.820 112.905 33.060 113.500 ;
        RECT 33.230 113.435 33.760 113.800 ;
        RECT 33.230 112.735 33.400 113.435 ;
        RECT 33.930 113.355 34.100 113.970 ;
        RECT 34.270 113.615 34.440 114.415 ;
        RECT 34.610 113.915 34.860 114.245 ;
        RECT 35.085 113.945 35.970 114.115 ;
        RECT 33.930 113.265 34.440 113.355 ;
        RECT 32.480 112.455 32.705 112.585 ;
        RECT 32.875 112.515 33.400 112.735 ;
        RECT 33.570 113.095 34.440 113.265 ;
        RECT 32.115 111.865 32.365 112.325 ;
        RECT 32.535 112.315 32.705 112.455 ;
        RECT 33.570 112.315 33.740 113.095 ;
        RECT 34.270 113.025 34.440 113.095 ;
        RECT 33.950 112.845 34.150 112.875 ;
        RECT 34.610 112.845 34.780 113.915 ;
        RECT 34.950 113.025 35.140 113.745 ;
        RECT 33.950 112.545 34.780 112.845 ;
        RECT 35.310 112.815 35.630 113.775 ;
        RECT 32.535 112.145 32.870 112.315 ;
        RECT 33.065 112.145 33.740 112.315 ;
        RECT 34.060 111.865 34.430 112.365 ;
        RECT 34.610 112.315 34.780 112.545 ;
        RECT 35.165 112.485 35.630 112.815 ;
        RECT 35.800 113.105 35.970 113.945 ;
        RECT 36.150 113.915 36.465 114.415 ;
        RECT 36.695 113.685 37.035 114.245 ;
        RECT 36.140 113.310 37.035 113.685 ;
        RECT 37.205 113.405 37.375 114.415 ;
        RECT 36.845 113.105 37.035 113.310 ;
        RECT 37.545 113.355 37.875 114.200 ;
        RECT 38.105 113.980 43.450 114.415 ;
        RECT 43.625 113.980 48.970 114.415 ;
        RECT 49.145 113.980 54.490 114.415 ;
        RECT 37.545 113.275 37.935 113.355 ;
        RECT 37.720 113.225 37.935 113.275 ;
        RECT 35.800 112.775 36.675 113.105 ;
        RECT 36.845 112.775 37.595 113.105 ;
        RECT 35.800 112.315 35.970 112.775 ;
        RECT 36.845 112.605 37.045 112.775 ;
        RECT 37.765 112.645 37.935 113.225 ;
        RECT 37.710 112.605 37.935 112.645 ;
        RECT 34.610 112.145 35.015 112.315 ;
        RECT 35.185 112.145 35.970 112.315 ;
        RECT 36.245 111.865 36.455 112.395 ;
        RECT 36.715 112.080 37.045 112.605 ;
        RECT 37.555 112.520 37.935 112.605 ;
        RECT 37.215 111.865 37.385 112.475 ;
        RECT 37.555 112.085 37.885 112.520 ;
        RECT 39.690 112.410 40.030 113.240 ;
        RECT 41.510 112.730 41.860 113.980 ;
        RECT 45.210 112.410 45.550 113.240 ;
        RECT 47.030 112.730 47.380 113.980 ;
        RECT 50.730 112.410 51.070 113.240 ;
        RECT 52.550 112.730 52.900 113.980 ;
        RECT 54.665 113.325 55.875 114.415 ;
        RECT 54.665 112.615 55.185 113.155 ;
        RECT 55.355 112.785 55.875 113.325 ;
        RECT 56.045 113.250 56.335 114.415 ;
        RECT 56.505 113.980 61.850 114.415 ;
        RECT 62.025 113.980 67.370 114.415 ;
        RECT 67.545 113.980 72.890 114.415 ;
        RECT 73.065 113.980 78.410 114.415 ;
        RECT 38.105 111.865 43.450 112.410 ;
        RECT 43.625 111.865 48.970 112.410 ;
        RECT 49.145 111.865 54.490 112.410 ;
        RECT 54.665 111.865 55.875 112.615 ;
        RECT 56.045 111.865 56.335 112.590 ;
        RECT 58.090 112.410 58.430 113.240 ;
        RECT 59.910 112.730 60.260 113.980 ;
        RECT 63.610 112.410 63.950 113.240 ;
        RECT 65.430 112.730 65.780 113.980 ;
        RECT 69.130 112.410 69.470 113.240 ;
        RECT 70.950 112.730 71.300 113.980 ;
        RECT 74.650 112.410 74.990 113.240 ;
        RECT 76.470 112.730 76.820 113.980 ;
        RECT 78.585 113.325 81.175 114.415 ;
        RECT 78.585 112.635 79.795 113.155 ;
        RECT 79.965 112.805 81.175 113.325 ;
        RECT 81.805 113.250 82.095 114.415 ;
        RECT 82.265 113.325 85.775 114.415 ;
        RECT 86.955 113.795 87.125 114.225 ;
        RECT 87.295 113.965 87.625 114.415 ;
        RECT 86.955 113.565 87.630 113.795 ;
        RECT 82.265 112.635 83.915 113.155 ;
        RECT 84.085 112.805 85.775 113.325 ;
        RECT 56.505 111.865 61.850 112.410 ;
        RECT 62.025 111.865 67.370 112.410 ;
        RECT 67.545 111.865 72.890 112.410 ;
        RECT 73.065 111.865 78.410 112.410 ;
        RECT 78.585 111.865 81.175 112.635 ;
        RECT 81.805 111.865 82.095 112.590 ;
        RECT 82.265 111.865 85.775 112.635 ;
        RECT 86.925 112.545 87.225 113.395 ;
        RECT 87.395 112.915 87.630 113.565 ;
        RECT 87.800 113.255 88.085 114.200 ;
        RECT 88.265 113.945 88.950 114.415 ;
        RECT 88.260 113.425 88.955 113.735 ;
        RECT 89.130 113.360 89.435 114.145 ;
        RECT 87.800 113.105 88.660 113.255 ;
        RECT 87.800 113.085 89.085 113.105 ;
        RECT 87.395 112.585 87.930 112.915 ;
        RECT 88.100 112.725 89.085 113.085 ;
        RECT 87.395 112.435 87.615 112.585 ;
        RECT 86.870 111.865 87.205 112.370 ;
        RECT 87.375 112.060 87.615 112.435 ;
        RECT 88.100 112.390 88.270 112.725 ;
        RECT 89.260 112.555 89.435 113.360 ;
        RECT 90.215 113.245 90.545 114.415 ;
        RECT 90.745 113.075 91.075 114.245 ;
        RECT 91.275 113.245 91.605 114.415 ;
        RECT 91.805 113.075 92.165 114.245 ;
        RECT 92.335 113.275 92.665 114.415 ;
        RECT 93.395 113.745 93.565 114.245 ;
        RECT 93.735 113.915 94.065 114.415 ;
        RECT 93.395 113.575 94.060 113.745 ;
        RECT 90.745 112.795 92.165 113.075 ;
        RECT 87.895 112.195 88.270 112.390 ;
        RECT 87.895 112.050 88.065 112.195 ;
        RECT 88.630 111.865 89.025 112.360 ;
        RECT 89.195 112.035 89.435 112.555 ;
        RECT 90.755 111.865 91.085 112.555 ;
        RECT 91.805 112.460 92.165 112.795 ;
        RECT 92.335 112.525 92.675 113.105 ;
        RECT 93.310 112.755 93.660 113.405 ;
        RECT 93.830 112.585 94.060 113.575 ;
        RECT 91.545 112.035 92.165 112.460 ;
        RECT 93.395 112.415 94.060 112.585 ;
        RECT 92.335 111.865 92.665 112.355 ;
        RECT 93.395 112.125 93.565 112.415 ;
        RECT 93.735 111.865 94.065 112.245 ;
        RECT 94.235 112.125 94.420 114.245 ;
        RECT 94.660 113.955 94.925 114.415 ;
        RECT 95.095 113.820 95.345 114.245 ;
        RECT 95.555 113.970 96.660 114.140 ;
        RECT 95.040 113.690 95.345 113.820 ;
        RECT 94.590 112.495 94.870 113.445 ;
        RECT 95.040 112.585 95.210 113.690 ;
        RECT 95.380 112.905 95.620 113.500 ;
        RECT 95.790 113.435 96.320 113.800 ;
        RECT 95.790 112.735 95.960 113.435 ;
        RECT 96.490 113.355 96.660 113.970 ;
        RECT 96.830 113.615 97.000 114.415 ;
        RECT 97.170 113.915 97.420 114.245 ;
        RECT 97.645 113.945 98.530 114.115 ;
        RECT 96.490 113.265 97.000 113.355 ;
        RECT 95.040 112.455 95.265 112.585 ;
        RECT 95.435 112.515 95.960 112.735 ;
        RECT 96.130 113.095 97.000 113.265 ;
        RECT 94.675 111.865 94.925 112.325 ;
        RECT 95.095 112.315 95.265 112.455 ;
        RECT 96.130 112.315 96.300 113.095 ;
        RECT 96.830 113.025 97.000 113.095 ;
        RECT 96.510 112.845 96.710 112.875 ;
        RECT 97.170 112.845 97.340 113.915 ;
        RECT 97.510 113.025 97.700 113.745 ;
        RECT 96.510 112.545 97.340 112.845 ;
        RECT 97.870 112.815 98.190 113.775 ;
        RECT 95.095 112.145 95.430 112.315 ;
        RECT 95.625 112.145 96.300 112.315 ;
        RECT 96.620 111.865 96.990 112.365 ;
        RECT 97.170 112.315 97.340 112.545 ;
        RECT 97.725 112.485 98.190 112.815 ;
        RECT 98.360 113.105 98.530 113.945 ;
        RECT 98.710 113.915 99.025 114.415 ;
        RECT 99.255 113.685 99.595 114.245 ;
        RECT 98.700 113.310 99.595 113.685 ;
        RECT 99.765 113.405 99.935 114.415 ;
        RECT 99.405 113.105 99.595 113.310 ;
        RECT 100.105 113.355 100.435 114.200 ;
        RECT 100.105 113.275 100.495 113.355 ;
        RECT 100.715 113.320 100.965 114.415 ;
        RECT 101.700 114.075 103.765 114.245 ;
        RECT 100.280 113.225 100.495 113.275 ;
        RECT 101.135 113.235 101.490 113.650 ;
        RECT 101.700 113.235 101.945 114.075 ;
        RECT 98.360 112.775 99.235 113.105 ;
        RECT 99.405 112.775 100.155 113.105 ;
        RECT 98.360 112.315 98.530 112.775 ;
        RECT 99.405 112.605 99.605 112.775 ;
        RECT 100.325 112.645 100.495 113.225 ;
        RECT 101.320 113.065 101.490 113.235 ;
        RECT 100.665 112.855 101.150 113.065 ;
        RECT 101.320 112.855 101.945 113.065 ;
        RECT 101.320 112.685 101.490 112.855 ;
        RECT 102.115 112.685 102.365 113.905 ;
        RECT 102.535 113.235 102.805 114.075 ;
        RECT 103.095 113.405 103.345 113.905 ;
        RECT 103.515 113.575 103.765 114.075 ;
        RECT 103.935 113.405 104.185 114.245 ;
        RECT 104.355 113.575 104.605 114.415 ;
        RECT 104.775 113.405 105.090 114.245 ;
        RECT 105.270 113.990 105.605 114.415 ;
        RECT 105.775 113.810 105.960 114.215 ;
        RECT 103.095 113.235 105.090 113.405 ;
        RECT 105.295 113.635 105.960 113.810 ;
        RECT 106.165 113.635 106.495 114.415 ;
        RECT 102.540 112.855 104.045 113.065 ;
        RECT 104.215 112.855 105.070 113.065 ;
        RECT 100.270 112.605 100.495 112.645 ;
        RECT 97.170 112.145 97.575 112.315 ;
        RECT 97.745 112.145 98.530 112.315 ;
        RECT 98.805 111.865 99.015 112.395 ;
        RECT 99.275 112.080 99.605 112.605 ;
        RECT 100.115 112.520 100.495 112.605 ;
        RECT 99.775 111.865 99.945 112.475 ;
        RECT 100.115 112.085 100.445 112.520 ;
        RECT 100.675 111.865 100.965 112.605 ;
        RECT 101.135 112.160 101.490 112.685 ;
        RECT 101.700 111.865 101.905 112.675 ;
        RECT 102.075 112.505 104.645 112.685 ;
        RECT 102.075 112.035 102.405 112.505 ;
        RECT 102.575 111.865 103.305 112.335 ;
        RECT 103.475 112.035 103.805 112.505 ;
        RECT 103.975 111.865 104.145 112.335 ;
        RECT 104.315 112.035 104.645 112.505 ;
        RECT 104.815 111.865 105.090 112.685 ;
        RECT 105.295 112.605 105.635 113.635 ;
        RECT 106.665 113.445 106.935 114.215 ;
        RECT 105.805 113.275 106.935 113.445 ;
        RECT 105.805 112.775 106.055 113.275 ;
        RECT 105.295 112.435 105.980 112.605 ;
        RECT 106.235 112.525 106.595 113.105 ;
        RECT 105.270 111.865 105.605 112.265 ;
        RECT 105.775 112.035 105.980 112.435 ;
        RECT 106.765 112.365 106.935 113.275 ;
        RECT 107.565 113.250 107.855 114.415 ;
        RECT 108.030 113.465 108.295 114.235 ;
        RECT 108.465 113.695 108.795 114.415 ;
        RECT 108.985 113.875 109.245 114.235 ;
        RECT 109.415 114.045 109.745 114.415 ;
        RECT 109.915 113.875 110.175 114.235 ;
        RECT 108.985 113.645 110.175 113.875 ;
        RECT 110.745 113.465 111.035 114.235 ;
        RECT 106.190 111.865 106.465 112.345 ;
        RECT 106.675 112.035 106.935 112.365 ;
        RECT 107.565 111.865 107.855 112.590 ;
        RECT 108.030 112.045 108.365 113.465 ;
        RECT 108.540 113.285 111.035 113.465 ;
        RECT 111.245 113.325 112.915 114.415 ;
        RECT 113.635 113.745 113.805 114.245 ;
        RECT 113.975 113.915 114.305 114.415 ;
        RECT 113.635 113.575 114.300 113.745 ;
        RECT 108.540 112.595 108.765 113.285 ;
        RECT 108.965 112.775 109.245 113.105 ;
        RECT 109.425 112.775 110.000 113.105 ;
        RECT 110.180 112.775 110.615 113.105 ;
        RECT 110.795 112.775 111.065 113.105 ;
        RECT 111.245 112.635 111.995 113.155 ;
        RECT 112.165 112.805 112.915 113.325 ;
        RECT 113.550 112.755 113.900 113.405 ;
        RECT 108.540 112.405 111.025 112.595 ;
        RECT 108.545 111.865 109.290 112.235 ;
        RECT 109.855 112.045 110.110 112.405 ;
        RECT 110.290 111.865 110.620 112.235 ;
        RECT 110.800 112.045 111.025 112.405 ;
        RECT 111.245 111.865 112.915 112.635 ;
        RECT 114.070 112.585 114.300 113.575 ;
        RECT 113.635 112.415 114.300 112.585 ;
        RECT 113.635 112.125 113.805 112.415 ;
        RECT 113.975 111.865 114.305 112.245 ;
        RECT 114.475 112.125 114.660 114.245 ;
        RECT 114.900 113.955 115.165 114.415 ;
        RECT 115.335 113.820 115.585 114.245 ;
        RECT 115.795 113.970 116.900 114.140 ;
        RECT 115.280 113.690 115.585 113.820 ;
        RECT 114.830 112.495 115.110 113.445 ;
        RECT 115.280 112.585 115.450 113.690 ;
        RECT 115.620 112.905 115.860 113.500 ;
        RECT 116.030 113.435 116.560 113.800 ;
        RECT 116.030 112.735 116.200 113.435 ;
        RECT 116.730 113.355 116.900 113.970 ;
        RECT 117.070 113.615 117.240 114.415 ;
        RECT 117.410 113.915 117.660 114.245 ;
        RECT 117.885 113.945 118.770 114.115 ;
        RECT 116.730 113.265 117.240 113.355 ;
        RECT 115.280 112.455 115.505 112.585 ;
        RECT 115.675 112.515 116.200 112.735 ;
        RECT 116.370 113.095 117.240 113.265 ;
        RECT 114.915 111.865 115.165 112.325 ;
        RECT 115.335 112.315 115.505 112.455 ;
        RECT 116.370 112.315 116.540 113.095 ;
        RECT 117.070 113.025 117.240 113.095 ;
        RECT 116.750 112.845 116.950 112.875 ;
        RECT 117.410 112.845 117.580 113.915 ;
        RECT 117.750 113.025 117.940 113.745 ;
        RECT 116.750 112.545 117.580 112.845 ;
        RECT 118.110 112.815 118.430 113.775 ;
        RECT 115.335 112.145 115.670 112.315 ;
        RECT 115.865 112.145 116.540 112.315 ;
        RECT 116.860 111.865 117.230 112.365 ;
        RECT 117.410 112.315 117.580 112.545 ;
        RECT 117.965 112.485 118.430 112.815 ;
        RECT 118.600 113.105 118.770 113.945 ;
        RECT 118.950 113.915 119.265 114.415 ;
        RECT 119.495 113.685 119.835 114.245 ;
        RECT 118.940 113.310 119.835 113.685 ;
        RECT 120.005 113.405 120.175 114.415 ;
        RECT 119.645 113.105 119.835 113.310 ;
        RECT 120.345 113.355 120.675 114.200 ;
        RECT 120.345 113.275 120.735 113.355 ;
        RECT 120.915 113.305 121.210 114.415 ;
        RECT 120.520 113.225 120.735 113.275 ;
        RECT 118.600 112.775 119.475 113.105 ;
        RECT 119.645 112.775 120.395 113.105 ;
        RECT 118.600 112.315 118.770 112.775 ;
        RECT 119.645 112.605 119.845 112.775 ;
        RECT 120.565 112.645 120.735 113.225 ;
        RECT 121.390 113.105 121.640 114.240 ;
        RECT 121.810 113.305 122.070 114.415 ;
        RECT 122.240 113.515 122.500 114.240 ;
        RECT 122.670 113.685 122.930 114.415 ;
        RECT 123.100 113.515 123.360 114.240 ;
        RECT 123.530 113.685 123.790 114.415 ;
        RECT 123.960 113.515 124.220 114.240 ;
        RECT 124.390 113.685 124.650 114.415 ;
        RECT 124.820 113.515 125.080 114.240 ;
        RECT 125.250 113.685 125.545 114.415 ;
        RECT 122.240 113.275 125.550 113.515 ;
        RECT 125.965 113.325 129.475 114.415 ;
        RECT 120.510 112.605 120.735 112.645 ;
        RECT 117.410 112.145 117.815 112.315 ;
        RECT 117.985 112.145 118.770 112.315 ;
        RECT 119.045 111.865 119.255 112.395 ;
        RECT 119.515 112.080 119.845 112.605 ;
        RECT 120.355 112.520 120.735 112.605 ;
        RECT 120.015 111.865 120.185 112.475 ;
        RECT 120.355 112.085 120.685 112.520 ;
        RECT 120.905 112.495 121.220 113.105 ;
        RECT 121.390 112.855 124.410 113.105 ;
        RECT 120.965 111.865 121.210 112.325 ;
        RECT 121.390 112.045 121.640 112.855 ;
        RECT 124.580 112.685 125.550 113.275 ;
        RECT 122.240 112.515 125.550 112.685 ;
        RECT 125.965 112.635 127.615 113.155 ;
        RECT 127.785 112.805 129.475 113.325 ;
        RECT 129.735 113.405 129.905 114.245 ;
        RECT 130.075 114.075 131.245 114.245 ;
        RECT 130.075 113.575 130.405 114.075 ;
        RECT 130.915 114.035 131.245 114.075 ;
        RECT 131.435 113.995 131.790 114.415 ;
        RECT 130.575 113.815 130.805 113.905 ;
        RECT 131.960 113.815 132.210 114.245 ;
        RECT 130.575 113.575 132.210 113.815 ;
        RECT 132.380 113.655 132.710 114.415 ;
        RECT 132.880 113.575 133.135 114.245 ;
        RECT 129.735 113.235 132.795 113.405 ;
        RECT 129.650 112.855 130.000 113.065 ;
        RECT 130.170 112.855 130.615 113.055 ;
        RECT 130.785 112.855 131.260 113.055 ;
        RECT 121.810 111.865 122.070 112.390 ;
        RECT 122.240 112.060 122.500 112.515 ;
        RECT 122.670 111.865 122.930 112.345 ;
        RECT 123.100 112.060 123.360 112.515 ;
        RECT 123.530 111.865 123.790 112.345 ;
        RECT 123.960 112.060 124.220 112.515 ;
        RECT 124.390 111.865 124.650 112.345 ;
        RECT 124.820 112.060 125.080 112.515 ;
        RECT 125.250 111.865 125.550 112.345 ;
        RECT 125.965 111.865 129.475 112.635 ;
        RECT 129.735 112.515 130.800 112.685 ;
        RECT 129.735 112.035 129.905 112.515 ;
        RECT 130.075 111.865 130.405 112.345 ;
        RECT 130.630 112.285 130.800 112.515 ;
        RECT 130.980 112.455 131.260 112.855 ;
        RECT 131.530 112.855 131.860 113.055 ;
        RECT 132.030 112.855 132.395 113.055 ;
        RECT 131.530 112.455 131.815 112.855 ;
        RECT 132.625 112.685 132.795 113.235 ;
        RECT 131.995 112.515 132.795 112.685 ;
        RECT 131.995 112.285 132.165 112.515 ;
        RECT 132.965 112.445 133.135 113.575 ;
        RECT 133.325 113.250 133.615 114.415 ;
        RECT 133.790 113.275 134.125 114.245 ;
        RECT 134.295 113.275 134.465 114.415 ;
        RECT 134.635 114.075 136.665 114.245 ;
        RECT 133.790 112.605 133.960 113.275 ;
        RECT 134.635 113.105 134.805 114.075 ;
        RECT 134.130 112.775 134.385 113.105 ;
        RECT 134.610 112.775 134.805 113.105 ;
        RECT 134.975 113.735 136.100 113.905 ;
        RECT 134.215 112.605 134.385 112.775 ;
        RECT 134.975 112.605 135.145 113.735 ;
        RECT 132.950 112.365 133.135 112.445 ;
        RECT 130.630 112.035 132.165 112.285 ;
        RECT 132.335 111.865 132.665 112.345 ;
        RECT 132.880 112.035 133.135 112.365 ;
        RECT 133.325 111.865 133.615 112.590 ;
        RECT 133.790 112.035 134.045 112.605 ;
        RECT 134.215 112.435 135.145 112.605 ;
        RECT 135.315 113.395 136.325 113.565 ;
        RECT 135.315 112.595 135.485 113.395 ;
        RECT 135.690 113.055 135.965 113.195 ;
        RECT 135.685 112.885 135.965 113.055 ;
        RECT 134.970 112.400 135.145 112.435 ;
        RECT 134.215 111.865 134.545 112.265 ;
        RECT 134.970 112.035 135.500 112.400 ;
        RECT 135.690 112.035 135.965 112.885 ;
        RECT 136.135 112.035 136.325 113.395 ;
        RECT 136.495 113.410 136.665 114.075 ;
        RECT 136.835 113.655 137.005 114.415 ;
        RECT 137.240 113.655 137.755 114.065 ;
        RECT 136.495 113.220 137.245 113.410 ;
        RECT 137.415 112.845 137.755 113.655 ;
        RECT 137.925 113.325 141.435 114.415 ;
        RECT 136.525 112.675 137.755 112.845 ;
        RECT 136.505 111.865 137.015 112.400 ;
        RECT 137.235 112.070 137.480 112.675 ;
        RECT 137.925 112.635 139.575 113.155 ;
        RECT 139.745 112.805 141.435 113.325 ;
        RECT 142.155 113.485 142.325 114.245 ;
        RECT 142.540 113.655 142.870 114.415 ;
        RECT 142.155 113.315 142.870 113.485 ;
        RECT 143.040 113.340 143.295 114.245 ;
        RECT 142.065 112.765 142.420 113.135 ;
        RECT 142.700 113.105 142.870 113.315 ;
        RECT 142.700 112.775 142.955 113.105 ;
        RECT 137.925 111.865 141.435 112.635 ;
        RECT 142.700 112.585 142.870 112.775 ;
        RECT 143.125 112.610 143.295 113.340 ;
        RECT 143.470 113.265 143.730 114.415 ;
        RECT 143.995 113.485 144.165 114.245 ;
        RECT 144.380 113.655 144.710 114.415 ;
        RECT 143.995 113.315 144.710 113.485 ;
        RECT 144.880 113.340 145.135 114.245 ;
        RECT 143.905 112.765 144.260 113.135 ;
        RECT 144.540 113.105 144.710 113.315 ;
        RECT 144.540 112.775 144.795 113.105 ;
        RECT 142.155 112.415 142.870 112.585 ;
        RECT 142.155 112.035 142.325 112.415 ;
        RECT 142.540 111.865 142.870 112.245 ;
        RECT 143.040 112.035 143.295 112.610 ;
        RECT 143.470 111.865 143.730 112.705 ;
        RECT 144.540 112.585 144.710 112.775 ;
        RECT 144.965 112.610 145.135 113.340 ;
        RECT 145.310 113.265 145.570 114.415 ;
        RECT 145.745 113.325 146.955 114.415 ;
        RECT 145.745 112.785 146.265 113.325 ;
        RECT 143.995 112.415 144.710 112.585 ;
        RECT 143.995 112.035 144.165 112.415 ;
        RECT 144.380 111.865 144.710 112.245 ;
        RECT 144.880 112.035 145.135 112.610 ;
        RECT 145.310 111.865 145.570 112.705 ;
        RECT 146.435 112.615 146.955 113.155 ;
        RECT 145.745 111.865 146.955 112.615 ;
        RECT 17.320 111.695 147.040 111.865 ;
        RECT 17.405 110.945 18.615 111.695 ;
        RECT 18.875 111.145 19.045 111.525 ;
        RECT 19.225 111.315 19.555 111.695 ;
        RECT 18.875 110.975 19.540 111.145 ;
        RECT 19.735 111.020 19.995 111.525 ;
        RECT 17.405 110.405 17.925 110.945 ;
        RECT 18.095 110.235 18.615 110.775 ;
        RECT 18.805 110.425 19.145 110.795 ;
        RECT 19.370 110.720 19.540 110.975 ;
        RECT 19.370 110.390 19.645 110.720 ;
        RECT 19.370 110.245 19.540 110.390 ;
        RECT 17.405 109.145 18.615 110.235 ;
        RECT 18.865 110.075 19.540 110.245 ;
        RECT 19.815 110.220 19.995 111.020 ;
        RECT 20.255 111.145 20.425 111.525 ;
        RECT 20.605 111.315 20.935 111.695 ;
        RECT 20.255 110.975 20.920 111.145 ;
        RECT 21.115 111.020 21.375 111.525 ;
        RECT 20.185 110.425 20.525 110.795 ;
        RECT 20.750 110.720 20.920 110.975 ;
        RECT 20.750 110.390 21.025 110.720 ;
        RECT 20.750 110.245 20.920 110.390 ;
        RECT 18.865 109.315 19.045 110.075 ;
        RECT 19.225 109.145 19.555 109.905 ;
        RECT 19.725 109.315 19.995 110.220 ;
        RECT 20.245 110.075 20.920 110.245 ;
        RECT 21.195 110.220 21.375 111.020 ;
        RECT 20.245 109.315 20.425 110.075 ;
        RECT 20.605 109.145 20.935 109.905 ;
        RECT 21.105 109.315 21.375 110.220 ;
        RECT 21.550 110.955 21.805 111.525 ;
        RECT 21.975 111.295 22.305 111.695 ;
        RECT 22.730 111.160 23.260 111.525 ;
        RECT 23.450 111.355 23.725 111.525 ;
        RECT 23.445 111.185 23.725 111.355 ;
        RECT 22.730 111.125 22.905 111.160 ;
        RECT 21.975 110.955 22.905 111.125 ;
        RECT 21.550 110.285 21.720 110.955 ;
        RECT 21.975 110.785 22.145 110.955 ;
        RECT 21.890 110.455 22.145 110.785 ;
        RECT 22.370 110.455 22.565 110.785 ;
        RECT 21.550 109.315 21.885 110.285 ;
        RECT 22.055 109.145 22.225 110.285 ;
        RECT 22.395 109.485 22.565 110.455 ;
        RECT 22.735 109.825 22.905 110.955 ;
        RECT 23.075 110.165 23.245 110.965 ;
        RECT 23.450 110.365 23.725 111.185 ;
        RECT 23.895 110.165 24.085 111.525 ;
        RECT 24.265 111.160 24.775 111.695 ;
        RECT 24.995 110.885 25.240 111.490 ;
        RECT 26.235 111.145 26.405 111.435 ;
        RECT 26.575 111.315 26.905 111.695 ;
        RECT 26.235 110.975 26.900 111.145 ;
        RECT 24.285 110.715 25.515 110.885 ;
        RECT 23.075 109.995 24.085 110.165 ;
        RECT 24.255 110.150 25.005 110.340 ;
        RECT 22.735 109.655 23.860 109.825 ;
        RECT 24.255 109.485 24.425 110.150 ;
        RECT 25.175 109.905 25.515 110.715 ;
        RECT 26.150 110.155 26.500 110.805 ;
        RECT 26.670 109.985 26.900 110.975 ;
        RECT 22.395 109.315 24.425 109.485 ;
        RECT 24.595 109.145 24.765 109.905 ;
        RECT 25.000 109.495 25.515 109.905 ;
        RECT 26.235 109.815 26.900 109.985 ;
        RECT 26.235 109.315 26.405 109.815 ;
        RECT 26.575 109.145 26.905 109.645 ;
        RECT 27.075 109.315 27.260 111.435 ;
        RECT 27.515 111.235 27.765 111.695 ;
        RECT 27.935 111.245 28.270 111.415 ;
        RECT 28.465 111.245 29.140 111.415 ;
        RECT 27.935 111.105 28.105 111.245 ;
        RECT 27.430 110.115 27.710 111.065 ;
        RECT 27.880 110.975 28.105 111.105 ;
        RECT 27.880 109.870 28.050 110.975 ;
        RECT 28.275 110.825 28.800 111.045 ;
        RECT 28.220 110.060 28.460 110.655 ;
        RECT 28.630 110.125 28.800 110.825 ;
        RECT 28.970 110.465 29.140 111.245 ;
        RECT 29.460 111.195 29.830 111.695 ;
        RECT 30.010 111.245 30.415 111.415 ;
        RECT 30.585 111.245 31.370 111.415 ;
        RECT 30.010 111.015 30.180 111.245 ;
        RECT 29.350 110.715 30.180 111.015 ;
        RECT 30.565 110.745 31.030 111.075 ;
        RECT 29.350 110.685 29.550 110.715 ;
        RECT 29.670 110.465 29.840 110.535 ;
        RECT 28.970 110.295 29.840 110.465 ;
        RECT 29.330 110.205 29.840 110.295 ;
        RECT 27.880 109.740 28.185 109.870 ;
        RECT 28.630 109.760 29.160 110.125 ;
        RECT 27.500 109.145 27.765 109.605 ;
        RECT 27.935 109.315 28.185 109.740 ;
        RECT 29.330 109.590 29.500 110.205 ;
        RECT 28.395 109.420 29.500 109.590 ;
        RECT 29.670 109.145 29.840 109.945 ;
        RECT 30.010 109.645 30.180 110.715 ;
        RECT 30.350 109.815 30.540 110.535 ;
        RECT 30.710 109.785 31.030 110.745 ;
        RECT 31.200 110.785 31.370 111.245 ;
        RECT 31.645 111.165 31.855 111.695 ;
        RECT 32.115 110.955 32.445 111.480 ;
        RECT 32.615 111.085 32.785 111.695 ;
        RECT 32.955 111.040 33.285 111.475 ;
        RECT 33.515 111.190 33.845 111.695 ;
        RECT 34.015 111.125 34.255 111.500 ;
        RECT 34.535 111.365 34.705 111.510 ;
        RECT 34.535 111.170 34.935 111.365 ;
        RECT 35.295 111.200 35.695 111.695 ;
        RECT 32.955 110.955 33.335 111.040 ;
        RECT 32.245 110.785 32.445 110.955 ;
        RECT 33.110 110.915 33.335 110.955 ;
        RECT 31.200 110.455 32.075 110.785 ;
        RECT 32.245 110.455 32.995 110.785 ;
        RECT 30.010 109.315 30.260 109.645 ;
        RECT 31.200 109.615 31.370 110.455 ;
        RECT 32.245 110.250 32.435 110.455 ;
        RECT 33.165 110.335 33.335 110.915 ;
        RECT 33.565 110.845 33.870 111.015 ;
        RECT 33.120 110.285 33.335 110.335 ;
        RECT 31.540 109.875 32.435 110.250 ;
        RECT 32.945 110.205 33.335 110.285 ;
        RECT 30.485 109.445 31.370 109.615 ;
        RECT 31.550 109.145 31.865 109.645 ;
        RECT 32.095 109.315 32.435 109.875 ;
        RECT 32.605 109.145 32.775 110.155 ;
        RECT 32.945 109.360 33.275 110.205 ;
        RECT 33.570 110.165 33.870 110.845 ;
        RECT 34.040 110.975 34.255 111.125 ;
        RECT 34.040 110.645 34.595 110.975 ;
        RECT 34.765 110.835 34.935 111.170 ;
        RECT 35.865 111.005 36.100 111.525 ;
        RECT 36.285 111.060 36.555 111.695 ;
        RECT 36.725 111.150 42.070 111.695 ;
        RECT 34.040 109.995 34.275 110.645 ;
        RECT 34.765 110.475 35.755 110.835 ;
        RECT 33.595 109.765 34.275 109.995 ;
        RECT 34.465 110.455 35.755 110.475 ;
        RECT 34.465 110.305 35.325 110.455 ;
        RECT 33.595 109.335 33.765 109.765 ;
        RECT 33.935 109.145 34.265 109.595 ;
        RECT 34.465 109.360 34.750 110.305 ;
        RECT 35.925 110.200 36.100 111.005 ;
        RECT 38.310 110.320 38.650 111.150 ;
        RECT 43.165 110.970 43.455 111.695 ;
        RECT 43.625 111.150 48.970 111.695 ;
        RECT 49.145 111.150 54.490 111.695 ;
        RECT 54.665 111.150 60.010 111.695 ;
        RECT 60.185 111.150 65.530 111.695 ;
        RECT 34.925 109.825 35.620 110.135 ;
        RECT 34.930 109.145 35.615 109.615 ;
        RECT 35.795 109.415 36.100 110.200 ;
        RECT 36.285 109.145 36.555 110.100 ;
        RECT 40.130 109.580 40.480 110.830 ;
        RECT 45.210 110.320 45.550 111.150 ;
        RECT 36.725 109.145 42.070 109.580 ;
        RECT 43.165 109.145 43.455 110.310 ;
        RECT 47.030 109.580 47.380 110.830 ;
        RECT 50.730 110.320 51.070 111.150 ;
        RECT 52.550 109.580 52.900 110.830 ;
        RECT 56.250 110.320 56.590 111.150 ;
        RECT 58.070 109.580 58.420 110.830 ;
        RECT 61.770 110.320 62.110 111.150 ;
        RECT 65.705 110.925 68.295 111.695 ;
        RECT 68.925 110.970 69.215 111.695 ;
        RECT 69.385 110.925 72.895 111.695 ;
        RECT 73.990 111.190 74.325 111.695 ;
        RECT 74.495 111.125 74.735 111.500 ;
        RECT 75.015 111.365 75.185 111.510 ;
        RECT 75.015 111.170 75.390 111.365 ;
        RECT 75.750 111.200 76.145 111.695 ;
        RECT 63.590 109.580 63.940 110.830 ;
        RECT 65.705 110.405 66.915 110.925 ;
        RECT 67.085 110.235 68.295 110.755 ;
        RECT 69.385 110.405 71.035 110.925 ;
        RECT 43.625 109.145 48.970 109.580 ;
        RECT 49.145 109.145 54.490 109.580 ;
        RECT 54.665 109.145 60.010 109.580 ;
        RECT 60.185 109.145 65.530 109.580 ;
        RECT 65.705 109.145 68.295 110.235 ;
        RECT 68.925 109.145 69.215 110.310 ;
        RECT 71.205 110.235 72.895 110.755 ;
        RECT 69.385 109.145 72.895 110.235 ;
        RECT 74.045 110.165 74.345 111.015 ;
        RECT 74.515 110.975 74.735 111.125 ;
        RECT 74.515 110.645 75.050 110.975 ;
        RECT 75.220 110.835 75.390 111.170 ;
        RECT 76.315 111.005 76.555 111.525 ;
        RECT 74.515 109.995 74.750 110.645 ;
        RECT 75.220 110.475 76.205 110.835 ;
        RECT 74.075 109.765 74.750 109.995 ;
        RECT 74.920 110.455 76.205 110.475 ;
        RECT 74.920 110.305 75.780 110.455 ;
        RECT 74.075 109.335 74.245 109.765 ;
        RECT 74.415 109.145 74.745 109.595 ;
        RECT 74.920 109.360 75.205 110.305 ;
        RECT 76.380 110.200 76.555 111.005 ;
        RECT 76.745 110.945 77.955 111.695 ;
        RECT 78.130 110.955 78.385 111.525 ;
        RECT 78.555 111.295 78.885 111.695 ;
        RECT 79.310 111.160 79.840 111.525 ;
        RECT 80.030 111.355 80.305 111.525 ;
        RECT 80.025 111.185 80.305 111.355 ;
        RECT 79.310 111.125 79.485 111.160 ;
        RECT 78.555 110.955 79.485 111.125 ;
        RECT 76.745 110.405 77.265 110.945 ;
        RECT 77.435 110.235 77.955 110.775 ;
        RECT 75.380 109.825 76.075 110.135 ;
        RECT 75.385 109.145 76.070 109.615 ;
        RECT 76.250 109.415 76.555 110.200 ;
        RECT 76.745 109.145 77.955 110.235 ;
        RECT 78.130 110.285 78.300 110.955 ;
        RECT 78.555 110.785 78.725 110.955 ;
        RECT 78.470 110.455 78.725 110.785 ;
        RECT 78.950 110.455 79.145 110.785 ;
        RECT 78.130 109.315 78.465 110.285 ;
        RECT 78.635 109.145 78.805 110.285 ;
        RECT 78.975 109.485 79.145 110.455 ;
        RECT 79.315 109.825 79.485 110.955 ;
        RECT 79.655 110.165 79.825 110.965 ;
        RECT 80.030 110.365 80.305 111.185 ;
        RECT 80.475 110.165 80.665 111.525 ;
        RECT 80.845 111.160 81.355 111.695 ;
        RECT 81.575 110.885 81.820 111.490 ;
        RECT 82.265 110.925 83.935 111.695 ;
        RECT 84.570 110.955 84.825 111.525 ;
        RECT 84.995 111.295 85.325 111.695 ;
        RECT 85.750 111.160 86.280 111.525 ;
        RECT 86.470 111.355 86.745 111.525 ;
        RECT 86.465 111.185 86.745 111.355 ;
        RECT 85.750 111.125 85.925 111.160 ;
        RECT 84.995 110.955 85.925 111.125 ;
        RECT 80.865 110.715 82.095 110.885 ;
        RECT 79.655 109.995 80.665 110.165 ;
        RECT 80.835 110.150 81.585 110.340 ;
        RECT 79.315 109.655 80.440 109.825 ;
        RECT 80.835 109.485 81.005 110.150 ;
        RECT 81.755 109.905 82.095 110.715 ;
        RECT 82.265 110.405 83.015 110.925 ;
        RECT 83.185 110.235 83.935 110.755 ;
        RECT 78.975 109.315 81.005 109.485 ;
        RECT 81.175 109.145 81.345 109.905 ;
        RECT 81.580 109.495 82.095 109.905 ;
        RECT 82.265 109.145 83.935 110.235 ;
        RECT 84.570 110.285 84.740 110.955 ;
        RECT 84.995 110.785 85.165 110.955 ;
        RECT 84.910 110.455 85.165 110.785 ;
        RECT 85.390 110.455 85.585 110.785 ;
        RECT 84.570 109.315 84.905 110.285 ;
        RECT 85.075 109.145 85.245 110.285 ;
        RECT 85.415 109.485 85.585 110.455 ;
        RECT 85.755 109.825 85.925 110.955 ;
        RECT 86.095 110.165 86.265 110.965 ;
        RECT 86.470 110.365 86.745 111.185 ;
        RECT 86.915 110.165 87.105 111.525 ;
        RECT 87.285 111.160 87.795 111.695 ;
        RECT 88.015 110.885 88.260 111.490 ;
        RECT 88.705 110.925 90.375 111.695 ;
        RECT 90.550 111.065 90.885 111.525 ;
        RECT 91.055 111.235 91.225 111.695 ;
        RECT 91.395 111.065 91.725 111.525 ;
        RECT 91.895 111.235 92.065 111.695 ;
        RECT 92.235 111.315 94.245 111.525 ;
        RECT 92.235 111.065 92.485 111.315 ;
        RECT 87.305 110.715 88.535 110.885 ;
        RECT 86.095 109.995 87.105 110.165 ;
        RECT 87.275 110.150 88.025 110.340 ;
        RECT 85.755 109.655 86.880 109.825 ;
        RECT 87.275 109.485 87.445 110.150 ;
        RECT 88.195 109.905 88.535 110.715 ;
        RECT 88.705 110.405 89.455 110.925 ;
        RECT 90.550 110.875 92.485 111.065 ;
        RECT 92.655 110.975 93.825 111.145 ;
        RECT 89.625 110.235 90.375 110.755 ;
        RECT 92.655 110.705 92.905 110.975 ;
        RECT 93.995 110.895 94.245 111.315 ;
        RECT 94.685 110.970 94.975 111.695 ;
        RECT 96.070 110.855 96.330 111.695 ;
        RECT 96.505 110.950 96.760 111.525 ;
        RECT 96.930 111.315 97.260 111.695 ;
        RECT 97.475 111.145 97.645 111.525 ;
        RECT 96.930 110.975 97.645 111.145 ;
        RECT 90.570 110.455 92.190 110.705 ;
        RECT 92.370 110.285 92.905 110.705 ;
        RECT 93.075 110.455 94.515 110.705 ;
        RECT 85.415 109.315 87.445 109.485 ;
        RECT 87.615 109.145 87.785 109.905 ;
        RECT 88.020 109.495 88.535 109.905 ;
        RECT 88.705 109.145 90.375 110.235 ;
        RECT 90.550 109.145 90.805 110.285 ;
        RECT 90.975 110.115 93.825 110.285 ;
        RECT 90.975 109.315 91.305 110.115 ;
        RECT 91.475 109.145 91.645 109.945 ;
        RECT 91.815 109.315 92.145 110.115 ;
        RECT 92.315 109.145 92.485 109.945 ;
        RECT 92.655 109.315 92.985 110.115 ;
        RECT 93.155 109.145 93.325 109.945 ;
        RECT 93.495 109.315 93.825 110.115 ;
        RECT 93.995 109.145 94.245 109.945 ;
        RECT 94.685 109.145 94.975 110.310 ;
        RECT 96.070 109.145 96.330 110.295 ;
        RECT 96.505 110.220 96.675 110.950 ;
        RECT 96.930 110.785 97.100 110.975 ;
        RECT 97.910 110.875 98.185 111.695 ;
        RECT 98.355 111.055 98.685 111.525 ;
        RECT 98.855 111.225 99.025 111.695 ;
        RECT 99.195 111.055 99.525 111.525 ;
        RECT 99.695 111.225 100.425 111.695 ;
        RECT 100.595 111.055 100.925 111.525 ;
        RECT 98.355 110.875 100.925 111.055 ;
        RECT 101.095 110.885 101.300 111.695 ;
        RECT 101.510 110.875 101.865 111.400 ;
        RECT 102.035 110.955 102.325 111.695 ;
        RECT 102.570 111.425 103.055 111.525 ;
        RECT 102.570 111.235 104.020 111.425 ;
        RECT 104.200 111.335 104.530 111.695 ;
        RECT 105.065 111.335 105.395 111.695 ;
        RECT 102.570 110.975 103.055 111.235 ;
        RECT 103.840 111.165 104.020 111.235 ;
        RECT 104.705 111.165 104.895 111.265 ;
        RECT 105.565 111.165 105.755 111.525 ;
        RECT 105.925 111.335 106.255 111.695 ;
        RECT 100.635 110.845 100.895 110.875 ;
        RECT 96.845 110.455 97.100 110.785 ;
        RECT 96.930 110.245 97.100 110.455 ;
        RECT 97.380 110.425 97.735 110.795 ;
        RECT 97.930 110.495 98.785 110.705 ;
        RECT 98.955 110.495 100.460 110.705 ;
        RECT 96.505 109.315 96.760 110.220 ;
        RECT 96.930 110.075 97.645 110.245 ;
        RECT 96.930 109.145 97.260 109.905 ;
        RECT 97.475 109.315 97.645 110.075 ;
        RECT 97.910 110.155 99.905 110.325 ;
        RECT 97.910 109.315 98.225 110.155 ;
        RECT 98.395 109.145 98.645 109.985 ;
        RECT 98.815 109.315 99.065 110.155 ;
        RECT 99.235 109.485 99.485 109.985 ;
        RECT 99.655 109.655 99.905 110.155 ;
        RECT 100.195 109.485 100.465 110.325 ;
        RECT 100.635 109.655 100.885 110.845 ;
        RECT 101.510 110.705 101.680 110.875 ;
        RECT 101.055 110.495 101.680 110.705 ;
        RECT 101.850 110.495 102.335 110.705 ;
        RECT 101.510 110.325 101.680 110.495 ;
        RECT 101.055 109.485 101.300 110.325 ;
        RECT 101.510 109.910 101.865 110.325 ;
        RECT 102.570 110.285 102.790 110.975 ;
        RECT 102.960 110.455 103.270 110.785 ;
        RECT 99.235 109.315 101.300 109.485 ;
        RECT 102.035 109.145 102.285 110.240 ;
        RECT 102.570 109.615 102.930 110.285 ;
        RECT 103.100 109.905 103.270 110.455 ;
        RECT 103.440 110.440 103.655 111.055 ;
        RECT 103.840 110.975 104.535 111.165 ;
        RECT 103.945 110.440 104.135 110.785 ;
        RECT 104.305 110.760 104.535 110.975 ;
        RECT 104.705 110.935 105.955 111.165 ;
        RECT 104.305 110.425 105.520 110.760 ;
        RECT 104.305 110.255 104.475 110.425 ;
        RECT 103.700 110.085 104.475 110.255 ;
        RECT 105.690 110.245 105.955 110.935 ;
        RECT 104.645 110.075 105.955 110.245 ;
        RECT 106.135 110.075 106.415 111.165 ;
        RECT 106.585 109.905 106.865 111.355 ;
        RECT 107.840 110.885 108.085 111.490 ;
        RECT 108.305 111.160 108.815 111.695 ;
        RECT 103.100 109.675 106.865 109.905 ;
        RECT 107.565 110.715 108.795 110.885 ;
        RECT 107.565 109.905 107.905 110.715 ;
        RECT 108.075 110.150 108.825 110.340 ;
        RECT 103.150 109.145 103.600 109.505 ;
        RECT 104.165 109.145 104.495 109.505 ;
        RECT 105.065 109.145 105.400 109.505 ;
        RECT 105.925 109.145 106.255 109.505 ;
        RECT 107.565 109.495 108.080 109.905 ;
        RECT 108.315 109.145 108.485 109.905 ;
        RECT 108.655 109.485 108.825 110.150 ;
        RECT 108.995 110.165 109.185 111.525 ;
        RECT 109.355 111.355 109.630 111.525 ;
        RECT 109.355 111.185 109.635 111.355 ;
        RECT 109.355 110.365 109.630 111.185 ;
        RECT 109.820 111.160 110.350 111.525 ;
        RECT 110.775 111.295 111.105 111.695 ;
        RECT 110.175 111.125 110.350 111.160 ;
        RECT 109.835 110.165 110.005 110.965 ;
        RECT 108.995 109.995 110.005 110.165 ;
        RECT 110.175 110.955 111.105 111.125 ;
        RECT 111.275 110.955 111.530 111.525 ;
        RECT 112.630 111.190 112.965 111.695 ;
        RECT 113.135 111.125 113.375 111.500 ;
        RECT 113.655 111.365 113.825 111.510 ;
        RECT 113.655 111.170 114.030 111.365 ;
        RECT 114.390 111.200 114.785 111.695 ;
        RECT 110.175 109.825 110.345 110.955 ;
        RECT 110.935 110.785 111.105 110.955 ;
        RECT 109.220 109.655 110.345 109.825 ;
        RECT 110.515 110.455 110.710 110.785 ;
        RECT 110.935 110.455 111.190 110.785 ;
        RECT 110.515 109.485 110.685 110.455 ;
        RECT 111.360 110.285 111.530 110.955 ;
        RECT 108.655 109.315 110.685 109.485 ;
        RECT 110.855 109.145 111.025 110.285 ;
        RECT 111.195 109.315 111.530 110.285 ;
        RECT 112.685 110.165 112.985 111.015 ;
        RECT 113.155 110.975 113.375 111.125 ;
        RECT 113.155 110.645 113.690 110.975 ;
        RECT 113.860 110.835 114.030 111.170 ;
        RECT 114.955 111.005 115.195 111.525 ;
        RECT 113.155 109.995 113.390 110.645 ;
        RECT 113.860 110.475 114.845 110.835 ;
        RECT 112.715 109.765 113.390 109.995 ;
        RECT 113.560 110.455 114.845 110.475 ;
        RECT 113.560 110.305 114.420 110.455 ;
        RECT 112.715 109.335 112.885 109.765 ;
        RECT 113.055 109.145 113.385 109.595 ;
        RECT 113.560 109.360 113.845 110.305 ;
        RECT 115.020 110.200 115.195 111.005 ;
        RECT 115.385 110.925 118.895 111.695 ;
        RECT 119.065 110.945 120.275 111.695 ;
        RECT 120.445 110.970 120.735 111.695 ;
        RECT 121.455 111.145 121.625 111.435 ;
        RECT 121.795 111.315 122.125 111.695 ;
        RECT 121.455 110.975 122.120 111.145 ;
        RECT 115.385 110.405 117.035 110.925 ;
        RECT 117.205 110.235 118.895 110.755 ;
        RECT 119.065 110.405 119.585 110.945 ;
        RECT 119.755 110.235 120.275 110.775 ;
        RECT 114.020 109.825 114.715 110.135 ;
        RECT 114.025 109.145 114.710 109.615 ;
        RECT 114.890 109.415 115.195 110.200 ;
        RECT 115.385 109.145 118.895 110.235 ;
        RECT 119.065 109.145 120.275 110.235 ;
        RECT 120.445 109.145 120.735 110.310 ;
        RECT 121.370 110.155 121.720 110.805 ;
        RECT 121.890 109.985 122.120 110.975 ;
        RECT 121.455 109.815 122.120 109.985 ;
        RECT 121.455 109.315 121.625 109.815 ;
        RECT 121.795 109.145 122.125 109.645 ;
        RECT 122.295 109.315 122.480 111.435 ;
        RECT 122.735 111.235 122.985 111.695 ;
        RECT 123.155 111.245 123.490 111.415 ;
        RECT 123.685 111.245 124.360 111.415 ;
        RECT 123.155 111.105 123.325 111.245 ;
        RECT 122.650 110.115 122.930 111.065 ;
        RECT 123.100 110.975 123.325 111.105 ;
        RECT 123.100 109.870 123.270 110.975 ;
        RECT 123.495 110.825 124.020 111.045 ;
        RECT 123.440 110.060 123.680 110.655 ;
        RECT 123.850 110.125 124.020 110.825 ;
        RECT 124.190 110.465 124.360 111.245 ;
        RECT 124.680 111.195 125.050 111.695 ;
        RECT 125.230 111.245 125.635 111.415 ;
        RECT 125.805 111.245 126.590 111.415 ;
        RECT 125.230 111.015 125.400 111.245 ;
        RECT 124.570 110.715 125.400 111.015 ;
        RECT 125.785 110.745 126.250 111.075 ;
        RECT 124.570 110.685 124.770 110.715 ;
        RECT 124.890 110.465 125.060 110.535 ;
        RECT 124.190 110.295 125.060 110.465 ;
        RECT 124.550 110.205 125.060 110.295 ;
        RECT 123.100 109.740 123.405 109.870 ;
        RECT 123.850 109.760 124.380 110.125 ;
        RECT 122.720 109.145 122.985 109.605 ;
        RECT 123.155 109.315 123.405 109.740 ;
        RECT 124.550 109.590 124.720 110.205 ;
        RECT 123.615 109.420 124.720 109.590 ;
        RECT 124.890 109.145 125.060 109.945 ;
        RECT 125.230 109.645 125.400 110.715 ;
        RECT 125.570 109.815 125.760 110.535 ;
        RECT 125.930 109.785 126.250 110.745 ;
        RECT 126.420 110.785 126.590 111.245 ;
        RECT 126.865 111.165 127.075 111.695 ;
        RECT 127.335 110.955 127.665 111.480 ;
        RECT 127.835 111.085 128.005 111.695 ;
        RECT 128.175 111.040 128.505 111.475 ;
        RECT 128.175 110.955 128.555 111.040 ;
        RECT 127.465 110.785 127.665 110.955 ;
        RECT 128.330 110.915 128.555 110.955 ;
        RECT 126.420 110.455 127.295 110.785 ;
        RECT 127.465 110.455 128.215 110.785 ;
        RECT 125.230 109.315 125.480 109.645 ;
        RECT 126.420 109.615 126.590 110.455 ;
        RECT 127.465 110.250 127.655 110.455 ;
        RECT 128.385 110.335 128.555 110.915 ;
        RECT 128.340 110.285 128.555 110.335 ;
        RECT 126.760 109.875 127.655 110.250 ;
        RECT 128.165 110.205 128.555 110.285 ;
        RECT 128.730 110.955 128.985 111.525 ;
        RECT 129.155 111.295 129.485 111.695 ;
        RECT 129.910 111.160 130.440 111.525 ;
        RECT 129.910 111.125 130.085 111.160 ;
        RECT 129.155 110.955 130.085 111.125 ;
        RECT 128.730 110.285 128.900 110.955 ;
        RECT 129.155 110.785 129.325 110.955 ;
        RECT 129.070 110.455 129.325 110.785 ;
        RECT 129.550 110.455 129.745 110.785 ;
        RECT 125.705 109.445 126.590 109.615 ;
        RECT 126.770 109.145 127.085 109.645 ;
        RECT 127.315 109.315 127.655 109.875 ;
        RECT 127.825 109.145 127.995 110.155 ;
        RECT 128.165 109.360 128.495 110.205 ;
        RECT 128.730 109.315 129.065 110.285 ;
        RECT 129.235 109.145 129.405 110.285 ;
        RECT 129.575 109.485 129.745 110.455 ;
        RECT 129.915 109.825 130.085 110.955 ;
        RECT 130.255 110.165 130.425 110.965 ;
        RECT 130.630 110.675 130.905 111.525 ;
        RECT 130.625 110.505 130.905 110.675 ;
        RECT 130.630 110.365 130.905 110.505 ;
        RECT 131.075 110.165 131.265 111.525 ;
        RECT 131.445 111.160 131.955 111.695 ;
        RECT 132.175 110.885 132.420 111.490 ;
        RECT 132.865 110.925 134.535 111.695 ;
        RECT 134.710 111.190 135.045 111.695 ;
        RECT 135.215 111.125 135.455 111.500 ;
        RECT 135.735 111.365 135.905 111.510 ;
        RECT 135.735 111.170 136.110 111.365 ;
        RECT 136.470 111.200 136.865 111.695 ;
        RECT 131.465 110.715 132.695 110.885 ;
        RECT 130.255 109.995 131.265 110.165 ;
        RECT 131.435 110.150 132.185 110.340 ;
        RECT 129.915 109.655 131.040 109.825 ;
        RECT 131.435 109.485 131.605 110.150 ;
        RECT 132.355 109.905 132.695 110.715 ;
        RECT 132.865 110.405 133.615 110.925 ;
        RECT 133.785 110.235 134.535 110.755 ;
        RECT 129.575 109.315 131.605 109.485 ;
        RECT 131.775 109.145 131.945 109.905 ;
        RECT 132.180 109.495 132.695 109.905 ;
        RECT 132.865 109.145 134.535 110.235 ;
        RECT 134.765 110.165 135.065 111.015 ;
        RECT 135.235 110.975 135.455 111.125 ;
        RECT 135.235 110.645 135.770 110.975 ;
        RECT 135.940 110.835 136.110 111.170 ;
        RECT 137.035 111.005 137.275 111.525 ;
        RECT 135.235 109.995 135.470 110.645 ;
        RECT 135.940 110.475 136.925 110.835 ;
        RECT 134.795 109.765 135.470 109.995 ;
        RECT 135.640 110.455 136.925 110.475 ;
        RECT 135.640 110.305 136.500 110.455 ;
        RECT 134.795 109.335 134.965 109.765 ;
        RECT 135.135 109.145 135.465 109.595 ;
        RECT 135.640 109.360 135.925 110.305 ;
        RECT 137.100 110.200 137.275 111.005 ;
        RECT 137.555 111.145 137.725 111.435 ;
        RECT 137.895 111.315 138.225 111.695 ;
        RECT 137.555 110.975 138.220 111.145 ;
        RECT 136.100 109.825 136.795 110.135 ;
        RECT 136.105 109.145 136.790 109.615 ;
        RECT 136.970 109.415 137.275 110.200 ;
        RECT 137.470 110.155 137.820 110.805 ;
        RECT 137.990 109.985 138.220 110.975 ;
        RECT 137.555 109.815 138.220 109.985 ;
        RECT 137.555 109.315 137.725 109.815 ;
        RECT 137.895 109.145 138.225 109.645 ;
        RECT 138.395 109.315 138.580 111.435 ;
        RECT 138.835 111.235 139.085 111.695 ;
        RECT 139.255 111.245 139.590 111.415 ;
        RECT 139.785 111.245 140.460 111.415 ;
        RECT 139.255 111.105 139.425 111.245 ;
        RECT 138.750 110.115 139.030 111.065 ;
        RECT 139.200 110.975 139.425 111.105 ;
        RECT 139.200 109.870 139.370 110.975 ;
        RECT 139.595 110.825 140.120 111.045 ;
        RECT 139.540 110.060 139.780 110.655 ;
        RECT 139.950 110.125 140.120 110.825 ;
        RECT 140.290 110.465 140.460 111.245 ;
        RECT 140.780 111.195 141.150 111.695 ;
        RECT 141.330 111.245 141.735 111.415 ;
        RECT 141.905 111.245 142.690 111.415 ;
        RECT 141.330 111.015 141.500 111.245 ;
        RECT 140.670 110.715 141.500 111.015 ;
        RECT 141.885 110.745 142.350 111.075 ;
        RECT 140.670 110.685 140.870 110.715 ;
        RECT 140.990 110.465 141.160 110.535 ;
        RECT 140.290 110.295 141.160 110.465 ;
        RECT 140.650 110.205 141.160 110.295 ;
        RECT 139.200 109.740 139.505 109.870 ;
        RECT 139.950 109.760 140.480 110.125 ;
        RECT 138.820 109.145 139.085 109.605 ;
        RECT 139.255 109.315 139.505 109.740 ;
        RECT 140.650 109.590 140.820 110.205 ;
        RECT 139.715 109.420 140.820 109.590 ;
        RECT 140.990 109.145 141.160 109.945 ;
        RECT 141.330 109.645 141.500 110.715 ;
        RECT 141.670 109.815 141.860 110.535 ;
        RECT 142.030 109.785 142.350 110.745 ;
        RECT 142.520 110.785 142.690 111.245 ;
        RECT 142.965 111.165 143.175 111.695 ;
        RECT 143.435 110.955 143.765 111.480 ;
        RECT 143.935 111.085 144.105 111.695 ;
        RECT 144.275 111.040 144.605 111.475 ;
        RECT 144.275 110.955 144.655 111.040 ;
        RECT 143.565 110.785 143.765 110.955 ;
        RECT 144.430 110.915 144.655 110.955 ;
        RECT 145.745 110.945 146.955 111.695 ;
        RECT 142.520 110.455 143.395 110.785 ;
        RECT 143.565 110.455 144.315 110.785 ;
        RECT 141.330 109.315 141.580 109.645 ;
        RECT 142.520 109.615 142.690 110.455 ;
        RECT 143.565 110.250 143.755 110.455 ;
        RECT 144.485 110.335 144.655 110.915 ;
        RECT 144.440 110.285 144.655 110.335 ;
        RECT 142.860 109.875 143.755 110.250 ;
        RECT 144.265 110.205 144.655 110.285 ;
        RECT 145.745 110.235 146.265 110.775 ;
        RECT 146.435 110.405 146.955 110.945 ;
        RECT 141.805 109.445 142.690 109.615 ;
        RECT 142.870 109.145 143.185 109.645 ;
        RECT 143.415 109.315 143.755 109.875 ;
        RECT 143.925 109.145 144.095 110.155 ;
        RECT 144.265 109.360 144.595 110.205 ;
        RECT 145.745 109.145 146.955 110.235 ;
        RECT 17.320 108.975 147.040 109.145 ;
        RECT 17.405 107.885 18.615 108.975 ;
        RECT 18.785 108.540 24.130 108.975 ;
        RECT 17.405 107.175 17.925 107.715 ;
        RECT 18.095 107.345 18.615 107.885 ;
        RECT 17.405 106.425 18.615 107.175 ;
        RECT 20.370 106.970 20.710 107.800 ;
        RECT 22.190 107.290 22.540 108.540 ;
        RECT 24.305 107.885 27.815 108.975 ;
        RECT 24.305 107.195 25.955 107.715 ;
        RECT 26.125 107.365 27.815 107.885 ;
        RECT 28.915 107.835 29.245 108.975 ;
        RECT 29.775 108.005 30.105 108.790 ;
        RECT 29.425 107.835 30.105 108.005 ;
        RECT 28.905 107.415 29.255 107.665 ;
        RECT 29.425 107.235 29.595 107.835 ;
        RECT 30.285 107.810 30.575 108.975 ;
        RECT 30.745 108.540 36.090 108.975 ;
        RECT 36.265 108.540 41.610 108.975 ;
        RECT 41.785 108.540 47.130 108.975 ;
        RECT 47.305 108.540 52.650 108.975 ;
        RECT 29.765 107.415 30.115 107.665 ;
        RECT 18.785 106.425 24.130 106.970 ;
        RECT 24.305 106.425 27.815 107.195 ;
        RECT 28.915 106.425 29.185 107.235 ;
        RECT 29.355 106.595 29.685 107.235 ;
        RECT 29.855 106.425 30.095 107.235 ;
        RECT 30.285 106.425 30.575 107.150 ;
        RECT 32.330 106.970 32.670 107.800 ;
        RECT 34.150 107.290 34.500 108.540 ;
        RECT 37.850 106.970 38.190 107.800 ;
        RECT 39.670 107.290 40.020 108.540 ;
        RECT 43.370 106.970 43.710 107.800 ;
        RECT 45.190 107.290 45.540 108.540 ;
        RECT 48.890 106.970 49.230 107.800 ;
        RECT 50.710 107.290 51.060 108.540 ;
        RECT 52.825 107.885 55.415 108.975 ;
        RECT 52.825 107.195 54.035 107.715 ;
        RECT 54.205 107.365 55.415 107.885 ;
        RECT 56.045 107.810 56.335 108.975 ;
        RECT 56.505 108.540 61.850 108.975 ;
        RECT 62.025 108.540 67.370 108.975 ;
        RECT 30.745 106.425 36.090 106.970 ;
        RECT 36.265 106.425 41.610 106.970 ;
        RECT 41.785 106.425 47.130 106.970 ;
        RECT 47.305 106.425 52.650 106.970 ;
        RECT 52.825 106.425 55.415 107.195 ;
        RECT 56.045 106.425 56.335 107.150 ;
        RECT 58.090 106.970 58.430 107.800 ;
        RECT 59.910 107.290 60.260 108.540 ;
        RECT 63.610 106.970 63.950 107.800 ;
        RECT 65.430 107.290 65.780 108.540 ;
        RECT 67.545 107.885 71.055 108.975 ;
        RECT 71.315 108.355 71.485 108.785 ;
        RECT 71.655 108.525 71.985 108.975 ;
        RECT 71.315 108.125 71.990 108.355 ;
        RECT 67.545 107.195 69.195 107.715 ;
        RECT 69.365 107.365 71.055 107.885 ;
        RECT 56.505 106.425 61.850 106.970 ;
        RECT 62.025 106.425 67.370 106.970 ;
        RECT 67.545 106.425 71.055 107.195 ;
        RECT 71.285 107.105 71.585 107.955 ;
        RECT 71.755 107.475 71.990 108.125 ;
        RECT 72.160 107.815 72.445 108.760 ;
        RECT 72.625 108.505 73.310 108.975 ;
        RECT 72.620 107.985 73.315 108.295 ;
        RECT 73.490 107.920 73.795 108.705 ;
        RECT 74.075 108.305 74.245 108.805 ;
        RECT 74.415 108.475 74.745 108.975 ;
        RECT 74.075 108.135 74.740 108.305 ;
        RECT 72.160 107.665 73.020 107.815 ;
        RECT 72.160 107.645 73.445 107.665 ;
        RECT 71.755 107.145 72.290 107.475 ;
        RECT 72.460 107.285 73.445 107.645 ;
        RECT 71.755 106.995 71.975 107.145 ;
        RECT 71.230 106.425 71.565 106.930 ;
        RECT 71.735 106.620 71.975 106.995 ;
        RECT 72.460 106.950 72.630 107.285 ;
        RECT 73.620 107.115 73.795 107.920 ;
        RECT 73.990 107.315 74.340 107.965 ;
        RECT 74.510 107.145 74.740 108.135 ;
        RECT 72.255 106.755 72.630 106.950 ;
        RECT 72.255 106.610 72.425 106.755 ;
        RECT 72.990 106.425 73.385 106.920 ;
        RECT 73.555 106.595 73.795 107.115 ;
        RECT 74.075 106.975 74.740 107.145 ;
        RECT 74.075 106.685 74.245 106.975 ;
        RECT 74.415 106.425 74.745 106.805 ;
        RECT 74.915 106.685 75.100 108.805 ;
        RECT 75.340 108.515 75.605 108.975 ;
        RECT 75.775 108.380 76.025 108.805 ;
        RECT 76.235 108.530 77.340 108.700 ;
        RECT 75.720 108.250 76.025 108.380 ;
        RECT 75.270 107.055 75.550 108.005 ;
        RECT 75.720 107.145 75.890 108.250 ;
        RECT 76.060 107.465 76.300 108.060 ;
        RECT 76.470 107.995 77.000 108.360 ;
        RECT 76.470 107.295 76.640 107.995 ;
        RECT 77.170 107.915 77.340 108.530 ;
        RECT 77.510 108.175 77.680 108.975 ;
        RECT 77.850 108.475 78.100 108.805 ;
        RECT 78.325 108.505 79.210 108.675 ;
        RECT 77.170 107.825 77.680 107.915 ;
        RECT 75.720 107.015 75.945 107.145 ;
        RECT 76.115 107.075 76.640 107.295 ;
        RECT 76.810 107.655 77.680 107.825 ;
        RECT 75.355 106.425 75.605 106.885 ;
        RECT 75.775 106.875 75.945 107.015 ;
        RECT 76.810 106.875 76.980 107.655 ;
        RECT 77.510 107.585 77.680 107.655 ;
        RECT 77.190 107.405 77.390 107.435 ;
        RECT 77.850 107.405 78.020 108.475 ;
        RECT 78.190 107.585 78.380 108.305 ;
        RECT 77.190 107.105 78.020 107.405 ;
        RECT 78.550 107.375 78.870 108.335 ;
        RECT 75.775 106.705 76.110 106.875 ;
        RECT 76.305 106.705 76.980 106.875 ;
        RECT 77.300 106.425 77.670 106.925 ;
        RECT 77.850 106.875 78.020 107.105 ;
        RECT 78.405 107.045 78.870 107.375 ;
        RECT 79.040 107.665 79.210 108.505 ;
        RECT 79.390 108.475 79.705 108.975 ;
        RECT 79.935 108.245 80.275 108.805 ;
        RECT 79.380 107.870 80.275 108.245 ;
        RECT 80.445 107.965 80.615 108.975 ;
        RECT 80.085 107.665 80.275 107.870 ;
        RECT 80.785 107.915 81.115 108.760 ;
        RECT 80.785 107.835 81.175 107.915 ;
        RECT 80.960 107.785 81.175 107.835 ;
        RECT 81.805 107.810 82.095 108.975 ;
        RECT 82.355 108.305 82.525 108.805 ;
        RECT 82.695 108.475 83.025 108.975 ;
        RECT 82.355 108.135 83.020 108.305 ;
        RECT 79.040 107.335 79.915 107.665 ;
        RECT 80.085 107.335 80.835 107.665 ;
        RECT 79.040 106.875 79.210 107.335 ;
        RECT 80.085 107.165 80.285 107.335 ;
        RECT 81.005 107.205 81.175 107.785 ;
        RECT 82.270 107.315 82.620 107.965 ;
        RECT 80.950 107.165 81.175 107.205 ;
        RECT 77.850 106.705 78.255 106.875 ;
        RECT 78.425 106.705 79.210 106.875 ;
        RECT 79.485 106.425 79.695 106.955 ;
        RECT 79.955 106.640 80.285 107.165 ;
        RECT 80.795 107.080 81.175 107.165 ;
        RECT 80.455 106.425 80.625 107.035 ;
        RECT 80.795 106.645 81.125 107.080 ;
        RECT 81.805 106.425 82.095 107.150 ;
        RECT 82.790 107.145 83.020 108.135 ;
        RECT 82.355 106.975 83.020 107.145 ;
        RECT 82.355 106.685 82.525 106.975 ;
        RECT 82.695 106.425 83.025 106.805 ;
        RECT 83.195 106.685 83.380 108.805 ;
        RECT 83.620 108.515 83.885 108.975 ;
        RECT 84.055 108.380 84.305 108.805 ;
        RECT 84.515 108.530 85.620 108.700 ;
        RECT 84.000 108.250 84.305 108.380 ;
        RECT 83.550 107.055 83.830 108.005 ;
        RECT 84.000 107.145 84.170 108.250 ;
        RECT 84.340 107.465 84.580 108.060 ;
        RECT 84.750 107.995 85.280 108.360 ;
        RECT 84.750 107.295 84.920 107.995 ;
        RECT 85.450 107.915 85.620 108.530 ;
        RECT 85.790 108.175 85.960 108.975 ;
        RECT 86.130 108.475 86.380 108.805 ;
        RECT 86.605 108.505 87.490 108.675 ;
        RECT 85.450 107.825 85.960 107.915 ;
        RECT 84.000 107.015 84.225 107.145 ;
        RECT 84.395 107.075 84.920 107.295 ;
        RECT 85.090 107.655 85.960 107.825 ;
        RECT 83.635 106.425 83.885 106.885 ;
        RECT 84.055 106.875 84.225 107.015 ;
        RECT 85.090 106.875 85.260 107.655 ;
        RECT 85.790 107.585 85.960 107.655 ;
        RECT 85.470 107.405 85.670 107.435 ;
        RECT 86.130 107.405 86.300 108.475 ;
        RECT 86.470 107.585 86.660 108.305 ;
        RECT 85.470 107.105 86.300 107.405 ;
        RECT 86.830 107.375 87.150 108.335 ;
        RECT 84.055 106.705 84.390 106.875 ;
        RECT 84.585 106.705 85.260 106.875 ;
        RECT 85.580 106.425 85.950 106.925 ;
        RECT 86.130 106.875 86.300 107.105 ;
        RECT 86.685 107.045 87.150 107.375 ;
        RECT 87.320 107.665 87.490 108.505 ;
        RECT 87.670 108.475 87.985 108.975 ;
        RECT 88.215 108.245 88.555 108.805 ;
        RECT 87.660 107.870 88.555 108.245 ;
        RECT 88.725 107.965 88.895 108.975 ;
        RECT 88.365 107.665 88.555 107.870 ;
        RECT 89.065 107.915 89.395 108.760 ;
        RECT 89.065 107.835 89.455 107.915 ;
        RECT 89.240 107.785 89.455 107.835 ;
        RECT 87.320 107.335 88.195 107.665 ;
        RECT 88.365 107.335 89.115 107.665 ;
        RECT 87.320 106.875 87.490 107.335 ;
        RECT 88.365 107.165 88.565 107.335 ;
        RECT 89.285 107.205 89.455 107.785 ;
        RECT 89.230 107.165 89.455 107.205 ;
        RECT 86.130 106.705 86.535 106.875 ;
        RECT 86.705 106.705 87.490 106.875 ;
        RECT 87.765 106.425 87.975 106.955 ;
        RECT 88.235 106.640 88.565 107.165 ;
        RECT 89.075 107.080 89.455 107.165 ;
        RECT 90.550 107.835 90.885 108.805 ;
        RECT 91.055 107.835 91.225 108.975 ;
        RECT 91.395 108.635 93.425 108.805 ;
        RECT 90.550 107.165 90.720 107.835 ;
        RECT 91.395 107.665 91.565 108.635 ;
        RECT 90.890 107.335 91.145 107.665 ;
        RECT 91.370 107.335 91.565 107.665 ;
        RECT 91.735 108.295 92.860 108.465 ;
        RECT 90.975 107.165 91.145 107.335 ;
        RECT 91.735 107.165 91.905 108.295 ;
        RECT 88.735 106.425 88.905 107.035 ;
        RECT 89.075 106.645 89.405 107.080 ;
        RECT 90.550 106.595 90.805 107.165 ;
        RECT 90.975 106.995 91.905 107.165 ;
        RECT 92.075 107.955 93.085 108.125 ;
        RECT 92.075 107.155 92.245 107.955 ;
        RECT 91.730 106.960 91.905 106.995 ;
        RECT 90.975 106.425 91.305 106.825 ;
        RECT 91.730 106.595 92.260 106.960 ;
        RECT 92.450 106.935 92.725 107.755 ;
        RECT 92.445 106.765 92.725 106.935 ;
        RECT 92.450 106.595 92.725 106.765 ;
        RECT 92.895 106.595 93.085 107.955 ;
        RECT 93.255 107.970 93.425 108.635 ;
        RECT 93.595 108.215 93.765 108.975 ;
        RECT 94.000 108.215 94.515 108.625 ;
        RECT 93.255 107.780 94.005 107.970 ;
        RECT 94.175 107.405 94.515 108.215 ;
        RECT 94.690 107.835 94.945 108.975 ;
        RECT 95.115 108.005 95.445 108.805 ;
        RECT 95.615 108.175 95.785 108.975 ;
        RECT 95.955 108.005 96.285 108.805 ;
        RECT 96.455 108.175 96.625 108.975 ;
        RECT 96.795 108.005 97.125 108.805 ;
        RECT 97.295 108.175 97.465 108.975 ;
        RECT 97.635 108.005 97.965 108.805 ;
        RECT 98.135 108.175 98.385 108.975 ;
        RECT 99.095 108.175 99.345 108.975 ;
        RECT 95.115 107.835 97.965 108.005 ;
        RECT 99.515 108.005 99.845 108.805 ;
        RECT 100.015 108.175 100.185 108.975 ;
        RECT 100.355 108.005 100.685 108.805 ;
        RECT 100.855 108.175 101.025 108.975 ;
        RECT 101.195 108.005 101.525 108.805 ;
        RECT 101.695 108.175 101.865 108.975 ;
        RECT 102.035 108.005 102.365 108.805 ;
        RECT 99.515 107.835 102.365 108.005 ;
        RECT 102.535 107.835 102.790 108.975 ;
        RECT 103.430 107.835 103.765 108.805 ;
        RECT 103.935 107.835 104.105 108.975 ;
        RECT 104.275 108.635 106.305 108.805 ;
        RECT 94.710 107.415 96.330 107.665 ;
        RECT 96.510 107.415 97.045 107.835 ;
        RECT 97.215 107.415 98.655 107.665 ;
        RECT 98.825 107.415 100.265 107.665 ;
        RECT 100.435 107.415 100.970 107.835 ;
        RECT 101.150 107.415 102.770 107.665 ;
        RECT 93.285 107.235 94.515 107.405 ;
        RECT 93.265 106.425 93.775 106.960 ;
        RECT 93.995 106.630 94.240 107.235 ;
        RECT 94.690 107.055 96.625 107.245 ;
        RECT 94.690 106.595 95.025 107.055 ;
        RECT 95.195 106.425 95.365 106.885 ;
        RECT 95.535 106.595 95.865 107.055 ;
        RECT 96.035 106.425 96.205 106.885 ;
        RECT 96.375 106.805 96.625 107.055 ;
        RECT 96.795 107.145 97.045 107.415 ;
        RECT 96.795 106.975 97.965 107.145 ;
        RECT 98.135 106.805 98.385 107.225 ;
        RECT 96.375 106.595 98.385 106.805 ;
        RECT 99.095 106.805 99.345 107.225 ;
        RECT 100.435 107.145 100.685 107.415 ;
        RECT 99.515 106.975 100.685 107.145 ;
        RECT 100.855 107.055 102.790 107.245 ;
        RECT 100.855 106.805 101.105 107.055 ;
        RECT 99.095 106.595 101.105 106.805 ;
        RECT 101.275 106.425 101.445 106.885 ;
        RECT 101.615 106.595 101.945 107.055 ;
        RECT 102.115 106.425 102.285 106.885 ;
        RECT 102.455 106.595 102.790 107.055 ;
        RECT 103.430 107.165 103.600 107.835 ;
        RECT 104.275 107.665 104.445 108.635 ;
        RECT 103.770 107.335 104.025 107.665 ;
        RECT 104.250 107.335 104.445 107.665 ;
        RECT 104.615 108.295 105.740 108.465 ;
        RECT 103.855 107.165 104.025 107.335 ;
        RECT 104.615 107.165 104.785 108.295 ;
        RECT 103.430 106.595 103.685 107.165 ;
        RECT 103.855 106.995 104.785 107.165 ;
        RECT 104.955 107.955 105.965 108.125 ;
        RECT 104.955 107.155 105.125 107.955 ;
        RECT 105.330 107.615 105.605 107.755 ;
        RECT 105.325 107.445 105.605 107.615 ;
        RECT 104.610 106.960 104.785 106.995 ;
        RECT 103.855 106.425 104.185 106.825 ;
        RECT 104.610 106.595 105.140 106.960 ;
        RECT 105.330 106.595 105.605 107.445 ;
        RECT 105.775 106.595 105.965 107.955 ;
        RECT 106.135 107.970 106.305 108.635 ;
        RECT 106.475 108.215 106.645 108.975 ;
        RECT 106.880 108.215 107.395 108.625 ;
        RECT 106.135 107.780 106.885 107.970 ;
        RECT 107.055 107.405 107.395 108.215 ;
        RECT 107.565 107.810 107.855 108.975 ;
        RECT 108.085 107.915 108.415 108.760 ;
        RECT 108.585 107.965 108.755 108.975 ;
        RECT 108.925 108.245 109.265 108.805 ;
        RECT 109.495 108.475 109.810 108.975 ;
        RECT 109.990 108.505 110.875 108.675 ;
        RECT 108.025 107.835 108.415 107.915 ;
        RECT 108.925 107.870 109.820 108.245 ;
        RECT 106.165 107.235 107.395 107.405 ;
        RECT 108.025 107.785 108.240 107.835 ;
        RECT 106.145 106.425 106.655 106.960 ;
        RECT 106.875 106.630 107.120 107.235 ;
        RECT 108.025 107.205 108.195 107.785 ;
        RECT 108.925 107.665 109.115 107.870 ;
        RECT 109.990 107.665 110.160 108.505 ;
        RECT 111.100 108.475 111.350 108.805 ;
        RECT 108.365 107.335 109.115 107.665 ;
        RECT 109.285 107.335 110.160 107.665 ;
        RECT 108.025 107.165 108.250 107.205 ;
        RECT 108.915 107.165 109.115 107.335 ;
        RECT 107.565 106.425 107.855 107.150 ;
        RECT 108.025 107.080 108.405 107.165 ;
        RECT 108.075 106.645 108.405 107.080 ;
        RECT 108.575 106.425 108.745 107.035 ;
        RECT 108.915 106.640 109.245 107.165 ;
        RECT 109.505 106.425 109.715 106.955 ;
        RECT 109.990 106.875 110.160 107.335 ;
        RECT 110.330 107.375 110.650 108.335 ;
        RECT 110.820 107.585 111.010 108.305 ;
        RECT 111.180 107.405 111.350 108.475 ;
        RECT 111.520 108.175 111.690 108.975 ;
        RECT 111.860 108.530 112.965 108.700 ;
        RECT 111.860 107.915 112.030 108.530 ;
        RECT 113.175 108.380 113.425 108.805 ;
        RECT 113.595 108.515 113.860 108.975 ;
        RECT 112.200 107.995 112.730 108.360 ;
        RECT 113.175 108.250 113.480 108.380 ;
        RECT 111.520 107.825 112.030 107.915 ;
        RECT 111.520 107.655 112.390 107.825 ;
        RECT 111.520 107.585 111.690 107.655 ;
        RECT 111.810 107.405 112.010 107.435 ;
        RECT 110.330 107.045 110.795 107.375 ;
        RECT 111.180 107.105 112.010 107.405 ;
        RECT 111.180 106.875 111.350 107.105 ;
        RECT 109.990 106.705 110.775 106.875 ;
        RECT 110.945 106.705 111.350 106.875 ;
        RECT 111.530 106.425 111.900 106.925 ;
        RECT 112.220 106.875 112.390 107.655 ;
        RECT 112.560 107.295 112.730 107.995 ;
        RECT 112.900 107.465 113.140 108.060 ;
        RECT 112.560 107.075 113.085 107.295 ;
        RECT 113.310 107.145 113.480 108.250 ;
        RECT 113.255 107.015 113.480 107.145 ;
        RECT 113.650 107.055 113.930 108.005 ;
        RECT 113.255 106.875 113.425 107.015 ;
        RECT 112.220 106.705 112.895 106.875 ;
        RECT 113.090 106.705 113.425 106.875 ;
        RECT 113.595 106.425 113.845 106.885 ;
        RECT 114.100 106.685 114.285 108.805 ;
        RECT 114.455 108.475 114.785 108.975 ;
        RECT 114.955 108.305 115.125 108.805 ;
        RECT 115.385 108.540 120.730 108.975 ;
        RECT 114.460 108.135 115.125 108.305 ;
        RECT 114.460 107.145 114.690 108.135 ;
        RECT 114.860 107.315 115.210 107.965 ;
        RECT 114.460 106.975 115.125 107.145 ;
        RECT 114.455 106.425 114.785 106.805 ;
        RECT 114.955 106.685 115.125 106.975 ;
        RECT 116.970 106.970 117.310 107.800 ;
        RECT 118.790 107.290 119.140 108.540 ;
        RECT 121.455 108.355 121.625 108.785 ;
        RECT 121.795 108.525 122.125 108.975 ;
        RECT 121.455 108.125 122.130 108.355 ;
        RECT 121.425 107.105 121.725 107.955 ;
        RECT 121.895 107.475 122.130 108.125 ;
        RECT 122.300 107.815 122.585 108.760 ;
        RECT 122.765 108.505 123.450 108.975 ;
        RECT 122.760 107.985 123.455 108.295 ;
        RECT 123.630 107.920 123.935 108.705 ;
        RECT 122.300 107.665 123.160 107.815 ;
        RECT 122.300 107.645 123.585 107.665 ;
        RECT 121.895 107.145 122.430 107.475 ;
        RECT 122.600 107.285 123.585 107.645 ;
        RECT 121.895 106.995 122.115 107.145 ;
        RECT 115.385 106.425 120.730 106.970 ;
        RECT 121.370 106.425 121.705 106.930 ;
        RECT 121.875 106.620 122.115 106.995 ;
        RECT 122.600 106.950 122.770 107.285 ;
        RECT 123.760 107.115 123.935 107.920 ;
        RECT 122.395 106.755 122.770 106.950 ;
        RECT 122.395 106.610 122.565 106.755 ;
        RECT 123.130 106.425 123.525 106.920 ;
        RECT 123.695 106.595 123.935 107.115 ;
        RECT 124.145 107.920 124.450 108.705 ;
        RECT 124.630 108.505 125.315 108.975 ;
        RECT 124.625 107.985 125.320 108.295 ;
        RECT 124.145 107.115 124.320 107.920 ;
        RECT 125.495 107.815 125.780 108.760 ;
        RECT 125.955 108.525 126.285 108.975 ;
        RECT 126.455 108.355 126.625 108.785 ;
        RECT 126.885 108.540 132.230 108.975 ;
        RECT 124.920 107.665 125.780 107.815 ;
        RECT 124.495 107.645 125.780 107.665 ;
        RECT 125.950 108.125 126.625 108.355 ;
        RECT 124.495 107.285 125.480 107.645 ;
        RECT 125.950 107.475 126.185 108.125 ;
        RECT 124.145 106.595 124.385 107.115 ;
        RECT 125.310 106.950 125.480 107.285 ;
        RECT 125.650 107.145 126.185 107.475 ;
        RECT 125.965 106.995 126.185 107.145 ;
        RECT 126.355 107.105 126.655 107.955 ;
        RECT 124.555 106.425 124.950 106.920 ;
        RECT 125.310 106.755 125.685 106.950 ;
        RECT 125.515 106.610 125.685 106.755 ;
        RECT 125.965 106.620 126.205 106.995 ;
        RECT 128.470 106.970 128.810 107.800 ;
        RECT 130.290 107.290 130.640 108.540 ;
        RECT 133.325 107.810 133.615 108.975 ;
        RECT 133.785 107.885 136.375 108.975 ;
        RECT 133.785 107.195 134.995 107.715 ;
        RECT 135.165 107.365 136.375 107.885 ;
        RECT 136.550 107.835 136.885 108.805 ;
        RECT 137.055 107.835 137.225 108.975 ;
        RECT 137.395 108.635 139.425 108.805 ;
        RECT 126.375 106.425 126.710 106.930 ;
        RECT 126.885 106.425 132.230 106.970 ;
        RECT 133.325 106.425 133.615 107.150 ;
        RECT 133.785 106.425 136.375 107.195 ;
        RECT 136.550 107.165 136.720 107.835 ;
        RECT 137.395 107.665 137.565 108.635 ;
        RECT 136.890 107.335 137.145 107.665 ;
        RECT 137.370 107.335 137.565 107.665 ;
        RECT 137.735 108.295 138.860 108.465 ;
        RECT 136.975 107.165 137.145 107.335 ;
        RECT 137.735 107.165 137.905 108.295 ;
        RECT 136.550 106.595 136.805 107.165 ;
        RECT 136.975 106.995 137.905 107.165 ;
        RECT 138.075 107.955 139.085 108.125 ;
        RECT 138.075 107.155 138.245 107.955 ;
        RECT 138.450 107.615 138.725 107.755 ;
        RECT 138.445 107.445 138.725 107.615 ;
        RECT 137.730 106.960 137.905 106.995 ;
        RECT 136.975 106.425 137.305 106.825 ;
        RECT 137.730 106.595 138.260 106.960 ;
        RECT 138.450 106.595 138.725 107.445 ;
        RECT 138.895 106.595 139.085 107.955 ;
        RECT 139.255 107.970 139.425 108.635 ;
        RECT 139.595 108.215 139.765 108.975 ;
        RECT 140.000 108.215 140.515 108.625 ;
        RECT 139.255 107.780 140.005 107.970 ;
        RECT 140.175 107.405 140.515 108.215 ;
        RECT 139.285 107.235 140.515 107.405 ;
        RECT 140.705 108.135 140.960 108.805 ;
        RECT 141.130 108.215 141.460 108.975 ;
        RECT 141.630 108.375 141.880 108.805 ;
        RECT 142.050 108.555 142.405 108.975 ;
        RECT 142.595 108.635 143.765 108.805 ;
        RECT 142.595 108.595 142.925 108.635 ;
        RECT 143.035 108.375 143.265 108.465 ;
        RECT 141.630 108.135 143.265 108.375 ;
        RECT 143.435 108.135 143.765 108.635 ;
        RECT 139.265 106.425 139.775 106.960 ;
        RECT 139.995 106.630 140.240 107.235 ;
        RECT 140.705 107.005 140.875 108.135 ;
        RECT 143.935 107.965 144.105 108.805 ;
        RECT 141.045 107.795 144.105 107.965 ;
        RECT 144.365 107.885 145.575 108.975 ;
        RECT 141.045 107.245 141.215 107.795 ;
        RECT 141.445 107.415 141.810 107.615 ;
        RECT 141.980 107.415 142.310 107.615 ;
        RECT 141.045 107.075 141.845 107.245 ;
        RECT 140.705 106.935 140.890 107.005 ;
        RECT 140.705 106.925 140.915 106.935 ;
        RECT 140.705 106.595 140.960 106.925 ;
        RECT 141.175 106.425 141.505 106.905 ;
        RECT 141.675 106.845 141.845 107.075 ;
        RECT 142.025 107.015 142.310 107.415 ;
        RECT 142.580 107.415 143.055 107.615 ;
        RECT 143.225 107.415 143.670 107.615 ;
        RECT 143.840 107.415 144.190 107.625 ;
        RECT 142.580 107.015 142.860 107.415 ;
        RECT 143.040 107.075 144.105 107.245 ;
        RECT 143.040 106.845 143.210 107.075 ;
        RECT 141.675 106.595 143.210 106.845 ;
        RECT 143.435 106.425 143.765 106.905 ;
        RECT 143.935 106.595 144.105 107.075 ;
        RECT 144.365 107.175 144.885 107.715 ;
        RECT 145.055 107.345 145.575 107.885 ;
        RECT 145.745 107.885 146.955 108.975 ;
        RECT 145.745 107.345 146.265 107.885 ;
        RECT 146.435 107.175 146.955 107.715 ;
        RECT 144.365 106.425 145.575 107.175 ;
        RECT 145.745 106.425 146.955 107.175 ;
        RECT 17.320 106.255 147.040 106.425 ;
        RECT 17.405 105.505 18.615 106.255 ;
        RECT 17.405 104.965 17.925 105.505 ;
        RECT 18.790 105.415 19.050 106.255 ;
        RECT 19.225 105.510 19.480 106.085 ;
        RECT 19.650 105.875 19.980 106.255 ;
        RECT 20.195 105.705 20.365 106.085 ;
        RECT 19.650 105.535 20.365 105.705 ;
        RECT 18.095 104.795 18.615 105.335 ;
        RECT 17.405 103.705 18.615 104.795 ;
        RECT 18.790 103.705 19.050 104.855 ;
        RECT 19.225 104.780 19.395 105.510 ;
        RECT 19.650 105.345 19.820 105.535 ;
        RECT 20.625 105.485 22.295 106.255 ;
        RECT 19.565 105.015 19.820 105.345 ;
        RECT 19.650 104.805 19.820 105.015 ;
        RECT 20.100 104.985 20.455 105.355 ;
        RECT 20.625 104.965 21.375 105.485 ;
        RECT 22.740 105.445 22.985 106.050 ;
        RECT 23.205 105.720 23.715 106.255 ;
        RECT 19.225 103.875 19.480 104.780 ;
        RECT 19.650 104.635 20.365 104.805 ;
        RECT 21.545 104.795 22.295 105.315 ;
        RECT 19.650 103.705 19.980 104.465 ;
        RECT 20.195 103.875 20.365 104.635 ;
        RECT 20.625 103.705 22.295 104.795 ;
        RECT 22.465 105.275 23.695 105.445 ;
        RECT 22.465 104.465 22.805 105.275 ;
        RECT 22.975 104.710 23.725 104.900 ;
        RECT 22.465 104.055 22.980 104.465 ;
        RECT 23.215 103.705 23.385 104.465 ;
        RECT 23.555 104.045 23.725 104.710 ;
        RECT 23.895 104.725 24.085 106.085 ;
        RECT 24.255 105.235 24.530 106.085 ;
        RECT 24.720 105.720 25.250 106.085 ;
        RECT 25.675 105.855 26.005 106.255 ;
        RECT 25.075 105.685 25.250 105.720 ;
        RECT 24.255 105.065 24.535 105.235 ;
        RECT 24.255 104.925 24.530 105.065 ;
        RECT 24.735 104.725 24.905 105.525 ;
        RECT 23.895 104.555 24.905 104.725 ;
        RECT 25.075 105.515 26.005 105.685 ;
        RECT 26.175 105.515 26.430 106.085 ;
        RECT 27.155 105.705 27.325 105.995 ;
        RECT 27.495 105.875 27.825 106.255 ;
        RECT 27.155 105.535 27.820 105.705 ;
        RECT 25.075 104.385 25.245 105.515 ;
        RECT 25.835 105.345 26.005 105.515 ;
        RECT 24.120 104.215 25.245 104.385 ;
        RECT 25.415 105.015 25.610 105.345 ;
        RECT 25.835 105.015 26.090 105.345 ;
        RECT 25.415 104.045 25.585 105.015 ;
        RECT 26.260 104.845 26.430 105.515 ;
        RECT 23.555 103.875 25.585 104.045 ;
        RECT 25.755 103.705 25.925 104.845 ;
        RECT 26.095 103.875 26.430 104.845 ;
        RECT 27.070 104.715 27.420 105.365 ;
        RECT 27.590 104.545 27.820 105.535 ;
        RECT 27.155 104.375 27.820 104.545 ;
        RECT 27.155 103.875 27.325 104.375 ;
        RECT 27.495 103.705 27.825 104.205 ;
        RECT 27.995 103.875 28.180 105.995 ;
        RECT 28.435 105.795 28.685 106.255 ;
        RECT 28.855 105.805 29.190 105.975 ;
        RECT 29.385 105.805 30.060 105.975 ;
        RECT 28.855 105.665 29.025 105.805 ;
        RECT 28.350 104.675 28.630 105.625 ;
        RECT 28.800 105.535 29.025 105.665 ;
        RECT 28.800 104.430 28.970 105.535 ;
        RECT 29.195 105.385 29.720 105.605 ;
        RECT 29.140 104.620 29.380 105.215 ;
        RECT 29.550 104.685 29.720 105.385 ;
        RECT 29.890 105.025 30.060 105.805 ;
        RECT 30.380 105.755 30.750 106.255 ;
        RECT 30.930 105.805 31.335 105.975 ;
        RECT 31.505 105.805 32.290 105.975 ;
        RECT 30.930 105.575 31.100 105.805 ;
        RECT 30.270 105.275 31.100 105.575 ;
        RECT 31.485 105.305 31.950 105.635 ;
        RECT 30.270 105.245 30.470 105.275 ;
        RECT 30.590 105.025 30.760 105.095 ;
        RECT 29.890 104.855 30.760 105.025 ;
        RECT 30.250 104.765 30.760 104.855 ;
        RECT 28.800 104.300 29.105 104.430 ;
        RECT 29.550 104.320 30.080 104.685 ;
        RECT 28.420 103.705 28.685 104.165 ;
        RECT 28.855 103.875 29.105 104.300 ;
        RECT 30.250 104.150 30.420 104.765 ;
        RECT 29.315 103.980 30.420 104.150 ;
        RECT 30.590 103.705 30.760 104.505 ;
        RECT 30.930 104.205 31.100 105.275 ;
        RECT 31.270 104.375 31.460 105.095 ;
        RECT 31.630 104.345 31.950 105.305 ;
        RECT 32.120 105.345 32.290 105.805 ;
        RECT 32.565 105.725 32.775 106.255 ;
        RECT 33.035 105.515 33.365 106.040 ;
        RECT 33.535 105.645 33.705 106.255 ;
        RECT 33.875 105.600 34.205 106.035 ;
        RECT 34.425 105.710 39.770 106.255 ;
        RECT 33.875 105.515 34.255 105.600 ;
        RECT 33.165 105.345 33.365 105.515 ;
        RECT 34.030 105.475 34.255 105.515 ;
        RECT 32.120 105.015 32.995 105.345 ;
        RECT 33.165 105.015 33.915 105.345 ;
        RECT 30.930 103.875 31.180 104.205 ;
        RECT 32.120 104.175 32.290 105.015 ;
        RECT 33.165 104.810 33.355 105.015 ;
        RECT 34.085 104.895 34.255 105.475 ;
        RECT 34.040 104.845 34.255 104.895 ;
        RECT 36.010 104.880 36.350 105.710 ;
        RECT 39.945 105.485 42.535 106.255 ;
        RECT 43.165 105.530 43.455 106.255 ;
        RECT 43.625 105.710 48.970 106.255 ;
        RECT 49.145 105.710 54.490 106.255 ;
        RECT 54.665 105.710 60.010 106.255 ;
        RECT 60.185 105.710 65.530 106.255 ;
        RECT 32.460 104.435 33.355 104.810 ;
        RECT 33.865 104.765 34.255 104.845 ;
        RECT 31.405 104.005 32.290 104.175 ;
        RECT 32.470 103.705 32.785 104.205 ;
        RECT 33.015 103.875 33.355 104.435 ;
        RECT 33.525 103.705 33.695 104.715 ;
        RECT 33.865 103.920 34.195 104.765 ;
        RECT 37.830 104.140 38.180 105.390 ;
        RECT 39.945 104.965 41.155 105.485 ;
        RECT 41.325 104.795 42.535 105.315 ;
        RECT 45.210 104.880 45.550 105.710 ;
        RECT 34.425 103.705 39.770 104.140 ;
        RECT 39.945 103.705 42.535 104.795 ;
        RECT 43.165 103.705 43.455 104.870 ;
        RECT 47.030 104.140 47.380 105.390 ;
        RECT 50.730 104.880 51.070 105.710 ;
        RECT 52.550 104.140 52.900 105.390 ;
        RECT 56.250 104.880 56.590 105.710 ;
        RECT 58.070 104.140 58.420 105.390 ;
        RECT 61.770 104.880 62.110 105.710 ;
        RECT 65.705 105.485 68.295 106.255 ;
        RECT 68.925 105.530 69.215 106.255 ;
        RECT 69.385 105.485 71.055 106.255 ;
        RECT 71.315 105.705 71.485 105.995 ;
        RECT 71.655 105.875 71.985 106.255 ;
        RECT 71.315 105.535 71.980 105.705 ;
        RECT 63.590 104.140 63.940 105.390 ;
        RECT 65.705 104.965 66.915 105.485 ;
        RECT 67.085 104.795 68.295 105.315 ;
        RECT 69.385 104.965 70.135 105.485 ;
        RECT 43.625 103.705 48.970 104.140 ;
        RECT 49.145 103.705 54.490 104.140 ;
        RECT 54.665 103.705 60.010 104.140 ;
        RECT 60.185 103.705 65.530 104.140 ;
        RECT 65.705 103.705 68.295 104.795 ;
        RECT 68.925 103.705 69.215 104.870 ;
        RECT 70.305 104.795 71.055 105.315 ;
        RECT 69.385 103.705 71.055 104.795 ;
        RECT 71.230 104.715 71.580 105.365 ;
        RECT 71.750 104.545 71.980 105.535 ;
        RECT 71.315 104.375 71.980 104.545 ;
        RECT 71.315 103.875 71.485 104.375 ;
        RECT 71.655 103.705 71.985 104.205 ;
        RECT 72.155 103.875 72.340 105.995 ;
        RECT 72.595 105.795 72.845 106.255 ;
        RECT 73.015 105.805 73.350 105.975 ;
        RECT 73.545 105.805 74.220 105.975 ;
        RECT 73.015 105.665 73.185 105.805 ;
        RECT 72.510 104.675 72.790 105.625 ;
        RECT 72.960 105.535 73.185 105.665 ;
        RECT 72.960 104.430 73.130 105.535 ;
        RECT 73.355 105.385 73.880 105.605 ;
        RECT 73.300 104.620 73.540 105.215 ;
        RECT 73.710 104.685 73.880 105.385 ;
        RECT 74.050 105.025 74.220 105.805 ;
        RECT 74.540 105.755 74.910 106.255 ;
        RECT 75.090 105.805 75.495 105.975 ;
        RECT 75.665 105.805 76.450 105.975 ;
        RECT 75.090 105.575 75.260 105.805 ;
        RECT 74.430 105.275 75.260 105.575 ;
        RECT 75.645 105.305 76.110 105.635 ;
        RECT 74.430 105.245 74.630 105.275 ;
        RECT 74.750 105.025 74.920 105.095 ;
        RECT 74.050 104.855 74.920 105.025 ;
        RECT 74.410 104.765 74.920 104.855 ;
        RECT 72.960 104.300 73.265 104.430 ;
        RECT 73.710 104.320 74.240 104.685 ;
        RECT 72.580 103.705 72.845 104.165 ;
        RECT 73.015 103.875 73.265 104.300 ;
        RECT 74.410 104.150 74.580 104.765 ;
        RECT 73.475 103.980 74.580 104.150 ;
        RECT 74.750 103.705 74.920 104.505 ;
        RECT 75.090 104.205 75.260 105.275 ;
        RECT 75.430 104.375 75.620 105.095 ;
        RECT 75.790 104.345 76.110 105.305 ;
        RECT 76.280 105.345 76.450 105.805 ;
        RECT 76.725 105.725 76.935 106.255 ;
        RECT 77.195 105.515 77.525 106.040 ;
        RECT 77.695 105.645 77.865 106.255 ;
        RECT 78.035 105.600 78.365 106.035 ;
        RECT 78.035 105.515 78.415 105.600 ;
        RECT 77.325 105.345 77.525 105.515 ;
        RECT 78.190 105.475 78.415 105.515 ;
        RECT 76.280 105.015 77.155 105.345 ;
        RECT 77.325 105.015 78.075 105.345 ;
        RECT 75.090 103.875 75.340 104.205 ;
        RECT 76.280 104.175 76.450 105.015 ;
        RECT 77.325 104.810 77.515 105.015 ;
        RECT 78.245 104.895 78.415 105.475 ;
        RECT 78.200 104.845 78.415 104.895 ;
        RECT 76.620 104.435 77.515 104.810 ;
        RECT 78.025 104.765 78.415 104.845 ;
        RECT 78.590 105.515 78.845 106.085 ;
        RECT 79.015 105.855 79.345 106.255 ;
        RECT 79.770 105.720 80.300 106.085 ;
        RECT 79.770 105.685 79.945 105.720 ;
        RECT 79.015 105.515 79.945 105.685 ;
        RECT 80.490 105.575 80.765 106.085 ;
        RECT 78.590 104.845 78.760 105.515 ;
        RECT 79.015 105.345 79.185 105.515 ;
        RECT 78.930 105.015 79.185 105.345 ;
        RECT 79.410 105.015 79.605 105.345 ;
        RECT 75.565 104.005 76.450 104.175 ;
        RECT 76.630 103.705 76.945 104.205 ;
        RECT 77.175 103.875 77.515 104.435 ;
        RECT 77.685 103.705 77.855 104.715 ;
        RECT 78.025 103.920 78.355 104.765 ;
        RECT 78.590 103.875 78.925 104.845 ;
        RECT 79.095 103.705 79.265 104.845 ;
        RECT 79.435 104.045 79.605 105.015 ;
        RECT 79.775 104.385 79.945 105.515 ;
        RECT 80.115 104.725 80.285 105.525 ;
        RECT 80.485 105.405 80.765 105.575 ;
        RECT 80.490 104.925 80.765 105.405 ;
        RECT 80.935 104.725 81.125 106.085 ;
        RECT 81.305 105.720 81.815 106.255 ;
        RECT 82.035 105.445 82.280 106.050 ;
        RECT 82.815 105.605 82.985 106.085 ;
        RECT 83.155 105.775 83.485 106.255 ;
        RECT 83.710 105.835 85.245 106.085 ;
        RECT 83.710 105.605 83.880 105.835 ;
        RECT 81.325 105.275 82.555 105.445 ;
        RECT 82.815 105.435 83.880 105.605 ;
        RECT 80.115 104.555 81.125 104.725 ;
        RECT 81.295 104.710 82.045 104.900 ;
        RECT 79.775 104.215 80.900 104.385 ;
        RECT 81.295 104.045 81.465 104.710 ;
        RECT 82.215 104.465 82.555 105.275 ;
        RECT 84.060 105.265 84.340 105.665 ;
        RECT 82.730 105.055 83.080 105.265 ;
        RECT 83.250 105.065 83.695 105.265 ;
        RECT 83.865 105.065 84.340 105.265 ;
        RECT 84.610 105.265 84.895 105.665 ;
        RECT 85.075 105.605 85.245 105.835 ;
        RECT 85.415 105.775 85.745 106.255 ;
        RECT 85.960 105.755 86.215 106.085 ;
        RECT 86.005 105.745 86.215 105.755 ;
        RECT 86.030 105.675 86.215 105.745 ;
        RECT 85.075 105.435 85.875 105.605 ;
        RECT 84.610 105.065 84.940 105.265 ;
        RECT 85.110 105.065 85.475 105.265 ;
        RECT 85.705 104.885 85.875 105.435 ;
        RECT 79.435 103.875 81.465 104.045 ;
        RECT 81.635 103.705 81.805 104.465 ;
        RECT 82.040 104.055 82.555 104.465 ;
        RECT 82.815 104.715 85.875 104.885 ;
        RECT 82.815 103.875 82.985 104.715 ;
        RECT 86.045 104.545 86.215 105.675 ;
        RECT 86.955 105.705 87.125 105.995 ;
        RECT 87.295 105.875 87.625 106.255 ;
        RECT 86.955 105.535 87.620 105.705 ;
        RECT 86.870 104.715 87.220 105.365 ;
        RECT 87.390 104.545 87.620 105.535 ;
        RECT 83.155 104.045 83.485 104.545 ;
        RECT 83.655 104.305 85.290 104.545 ;
        RECT 83.655 104.215 83.885 104.305 ;
        RECT 83.995 104.045 84.325 104.085 ;
        RECT 83.155 103.875 84.325 104.045 ;
        RECT 84.515 103.705 84.870 104.125 ;
        RECT 85.040 103.875 85.290 104.305 ;
        RECT 85.460 103.705 85.790 104.465 ;
        RECT 85.960 103.875 86.215 104.545 ;
        RECT 86.955 104.375 87.620 104.545 ;
        RECT 86.955 103.875 87.125 104.375 ;
        RECT 87.295 103.705 87.625 104.205 ;
        RECT 87.795 103.875 87.980 105.995 ;
        RECT 88.235 105.795 88.485 106.255 ;
        RECT 88.655 105.805 88.990 105.975 ;
        RECT 89.185 105.805 89.860 105.975 ;
        RECT 88.655 105.665 88.825 105.805 ;
        RECT 88.150 104.675 88.430 105.625 ;
        RECT 88.600 105.535 88.825 105.665 ;
        RECT 88.600 104.430 88.770 105.535 ;
        RECT 88.995 105.385 89.520 105.605 ;
        RECT 88.940 104.620 89.180 105.215 ;
        RECT 89.350 104.685 89.520 105.385 ;
        RECT 89.690 105.025 89.860 105.805 ;
        RECT 90.180 105.755 90.550 106.255 ;
        RECT 90.730 105.805 91.135 105.975 ;
        RECT 91.305 105.805 92.090 105.975 ;
        RECT 90.730 105.575 90.900 105.805 ;
        RECT 90.070 105.275 90.900 105.575 ;
        RECT 91.285 105.305 91.750 105.635 ;
        RECT 90.070 105.245 90.270 105.275 ;
        RECT 90.390 105.025 90.560 105.095 ;
        RECT 89.690 104.855 90.560 105.025 ;
        RECT 90.050 104.765 90.560 104.855 ;
        RECT 88.600 104.300 88.905 104.430 ;
        RECT 89.350 104.320 89.880 104.685 ;
        RECT 88.220 103.705 88.485 104.165 ;
        RECT 88.655 103.875 88.905 104.300 ;
        RECT 90.050 104.150 90.220 104.765 ;
        RECT 89.115 103.980 90.220 104.150 ;
        RECT 90.390 103.705 90.560 104.505 ;
        RECT 90.730 104.205 90.900 105.275 ;
        RECT 91.070 104.375 91.260 105.095 ;
        RECT 91.430 104.345 91.750 105.305 ;
        RECT 91.920 105.345 92.090 105.805 ;
        RECT 92.365 105.725 92.575 106.255 ;
        RECT 92.835 105.515 93.165 106.040 ;
        RECT 93.335 105.645 93.505 106.255 ;
        RECT 93.675 105.600 94.005 106.035 ;
        RECT 93.675 105.515 94.055 105.600 ;
        RECT 94.685 105.530 94.975 106.255 ;
        RECT 95.415 105.875 97.425 106.085 ;
        RECT 92.965 105.345 93.165 105.515 ;
        RECT 93.830 105.475 94.055 105.515 ;
        RECT 91.920 105.015 92.795 105.345 ;
        RECT 92.965 105.015 93.715 105.345 ;
        RECT 90.730 103.875 90.980 104.205 ;
        RECT 91.920 104.175 92.090 105.015 ;
        RECT 92.965 104.810 93.155 105.015 ;
        RECT 93.885 104.895 94.055 105.475 ;
        RECT 95.415 105.455 95.665 105.875 ;
        RECT 95.835 105.535 97.005 105.705 ;
        RECT 96.755 105.265 97.005 105.535 ;
        RECT 97.175 105.625 97.425 105.875 ;
        RECT 97.595 105.795 97.765 106.255 ;
        RECT 97.935 105.625 98.265 106.085 ;
        RECT 98.435 105.795 98.605 106.255 ;
        RECT 98.775 105.625 99.110 106.085 ;
        RECT 97.175 105.435 99.110 105.625 ;
        RECT 99.285 105.505 100.495 106.255 ;
        RECT 100.670 105.855 101.005 106.255 ;
        RECT 101.175 105.685 101.380 106.085 ;
        RECT 101.590 105.775 101.865 106.255 ;
        RECT 102.075 105.755 102.335 106.085 ;
        RECT 100.695 105.515 101.380 105.685 ;
        RECT 95.145 105.015 96.585 105.265 ;
        RECT 93.840 104.845 94.055 104.895 ;
        RECT 92.260 104.435 93.155 104.810 ;
        RECT 93.665 104.765 94.055 104.845 ;
        RECT 91.205 104.005 92.090 104.175 ;
        RECT 92.270 103.705 92.585 104.205 ;
        RECT 92.815 103.875 93.155 104.435 ;
        RECT 93.325 103.705 93.495 104.715 ;
        RECT 93.665 103.920 93.995 104.765 ;
        RECT 94.685 103.705 94.975 104.870 ;
        RECT 96.755 104.845 97.290 105.265 ;
        RECT 97.470 105.015 99.090 105.265 ;
        RECT 99.285 104.965 99.805 105.505 ;
        RECT 95.835 104.675 98.685 104.845 ;
        RECT 95.415 103.705 95.665 104.505 ;
        RECT 95.835 103.875 96.165 104.675 ;
        RECT 96.335 103.705 96.505 104.505 ;
        RECT 96.675 103.875 97.005 104.675 ;
        RECT 97.175 103.705 97.345 104.505 ;
        RECT 97.515 103.875 97.845 104.675 ;
        RECT 98.015 103.705 98.185 104.505 ;
        RECT 98.355 103.875 98.685 104.675 ;
        RECT 98.855 103.705 99.110 104.845 ;
        RECT 99.975 104.795 100.495 105.335 ;
        RECT 99.285 103.705 100.495 104.795 ;
        RECT 100.695 104.485 101.035 105.515 ;
        RECT 101.205 104.845 101.455 105.345 ;
        RECT 101.635 105.015 101.995 105.595 ;
        RECT 102.165 104.845 102.335 105.755 ;
        RECT 102.595 105.705 102.765 105.995 ;
        RECT 102.935 105.875 103.265 106.255 ;
        RECT 102.595 105.535 103.260 105.705 ;
        RECT 101.205 104.675 102.335 104.845 ;
        RECT 102.510 104.715 102.860 105.365 ;
        RECT 100.695 104.310 101.360 104.485 ;
        RECT 100.670 103.705 101.005 104.130 ;
        RECT 101.175 103.905 101.360 104.310 ;
        RECT 101.565 103.705 101.895 104.485 ;
        RECT 102.065 103.905 102.335 104.675 ;
        RECT 103.030 104.545 103.260 105.535 ;
        RECT 102.595 104.375 103.260 104.545 ;
        RECT 102.595 103.875 102.765 104.375 ;
        RECT 102.935 103.705 103.265 104.205 ;
        RECT 103.435 103.875 103.620 105.995 ;
        RECT 103.875 105.795 104.125 106.255 ;
        RECT 104.295 105.805 104.630 105.975 ;
        RECT 104.825 105.805 105.500 105.975 ;
        RECT 104.295 105.665 104.465 105.805 ;
        RECT 103.790 104.675 104.070 105.625 ;
        RECT 104.240 105.535 104.465 105.665 ;
        RECT 104.240 104.430 104.410 105.535 ;
        RECT 104.635 105.385 105.160 105.605 ;
        RECT 104.580 104.620 104.820 105.215 ;
        RECT 104.990 104.685 105.160 105.385 ;
        RECT 105.330 105.025 105.500 105.805 ;
        RECT 105.820 105.755 106.190 106.255 ;
        RECT 106.370 105.805 106.775 105.975 ;
        RECT 106.945 105.805 107.730 105.975 ;
        RECT 106.370 105.575 106.540 105.805 ;
        RECT 105.710 105.275 106.540 105.575 ;
        RECT 106.925 105.305 107.390 105.635 ;
        RECT 105.710 105.245 105.910 105.275 ;
        RECT 106.030 105.025 106.200 105.095 ;
        RECT 105.330 104.855 106.200 105.025 ;
        RECT 105.690 104.765 106.200 104.855 ;
        RECT 104.240 104.300 104.545 104.430 ;
        RECT 104.990 104.320 105.520 104.685 ;
        RECT 103.860 103.705 104.125 104.165 ;
        RECT 104.295 103.875 104.545 104.300 ;
        RECT 105.690 104.150 105.860 104.765 ;
        RECT 104.755 103.980 105.860 104.150 ;
        RECT 106.030 103.705 106.200 104.505 ;
        RECT 106.370 104.205 106.540 105.275 ;
        RECT 106.710 104.375 106.900 105.095 ;
        RECT 107.070 104.345 107.390 105.305 ;
        RECT 107.560 105.345 107.730 105.805 ;
        RECT 108.005 105.725 108.215 106.255 ;
        RECT 108.475 105.515 108.805 106.040 ;
        RECT 108.975 105.645 109.145 106.255 ;
        RECT 109.315 105.600 109.645 106.035 ;
        RECT 109.315 105.515 109.695 105.600 ;
        RECT 108.605 105.345 108.805 105.515 ;
        RECT 109.470 105.475 109.695 105.515 ;
        RECT 109.870 105.490 110.325 106.255 ;
        RECT 110.600 105.875 111.900 106.085 ;
        RECT 112.155 105.895 112.485 106.255 ;
        RECT 111.730 105.725 111.900 105.875 ;
        RECT 112.655 105.755 112.915 106.085 ;
        RECT 112.685 105.745 112.915 105.755 ;
        RECT 107.560 105.015 108.435 105.345 ;
        RECT 108.605 105.015 109.355 105.345 ;
        RECT 106.370 103.875 106.620 104.205 ;
        RECT 107.560 104.175 107.730 105.015 ;
        RECT 108.605 104.810 108.795 105.015 ;
        RECT 109.525 104.895 109.695 105.475 ;
        RECT 110.800 105.265 111.020 105.665 ;
        RECT 109.865 105.065 110.355 105.265 ;
        RECT 110.545 105.055 111.020 105.265 ;
        RECT 111.265 105.265 111.475 105.665 ;
        RECT 111.730 105.600 112.485 105.725 ;
        RECT 111.730 105.555 112.575 105.600 ;
        RECT 112.305 105.435 112.575 105.555 ;
        RECT 111.265 105.055 111.595 105.265 ;
        RECT 111.765 104.995 112.175 105.300 ;
        RECT 109.480 104.845 109.695 104.895 ;
        RECT 107.900 104.435 108.795 104.810 ;
        RECT 109.305 104.765 109.695 104.845 ;
        RECT 109.870 104.825 111.045 104.885 ;
        RECT 112.405 104.860 112.575 105.435 ;
        RECT 112.375 104.825 112.575 104.860 ;
        RECT 106.845 104.005 107.730 104.175 ;
        RECT 107.910 103.705 108.225 104.205 ;
        RECT 108.455 103.875 108.795 104.435 ;
        RECT 108.965 103.705 109.135 104.715 ;
        RECT 109.305 103.920 109.635 104.765 ;
        RECT 109.870 104.715 112.575 104.825 ;
        RECT 109.870 104.095 110.125 104.715 ;
        RECT 110.715 104.655 112.515 104.715 ;
        RECT 110.715 104.625 111.045 104.655 ;
        RECT 112.745 104.555 112.915 105.745 ;
        RECT 113.085 105.710 118.430 106.255 ;
        RECT 114.670 104.880 115.010 105.710 ;
        RECT 118.605 105.485 120.275 106.255 ;
        RECT 120.445 105.530 120.735 106.255 ;
        RECT 120.905 105.505 122.115 106.255 ;
        RECT 122.375 105.705 122.545 105.995 ;
        RECT 122.715 105.875 123.045 106.255 ;
        RECT 122.375 105.535 123.040 105.705 ;
        RECT 110.375 104.455 110.560 104.545 ;
        RECT 111.150 104.455 111.985 104.465 ;
        RECT 110.375 104.255 111.985 104.455 ;
        RECT 110.375 104.215 110.605 104.255 ;
        RECT 109.870 103.875 110.205 104.095 ;
        RECT 111.210 103.705 111.565 104.085 ;
        RECT 111.735 103.875 111.985 104.255 ;
        RECT 112.235 103.705 112.485 104.485 ;
        RECT 112.655 103.875 112.915 104.555 ;
        RECT 116.490 104.140 116.840 105.390 ;
        RECT 118.605 104.965 119.355 105.485 ;
        RECT 119.525 104.795 120.275 105.315 ;
        RECT 120.905 104.965 121.425 105.505 ;
        RECT 113.085 103.705 118.430 104.140 ;
        RECT 118.605 103.705 120.275 104.795 ;
        RECT 120.445 103.705 120.735 104.870 ;
        RECT 121.595 104.795 122.115 105.335 ;
        RECT 120.905 103.705 122.115 104.795 ;
        RECT 122.290 104.715 122.640 105.365 ;
        RECT 122.810 104.545 123.040 105.535 ;
        RECT 122.375 104.375 123.040 104.545 ;
        RECT 122.375 103.875 122.545 104.375 ;
        RECT 122.715 103.705 123.045 104.205 ;
        RECT 123.215 103.875 123.400 105.995 ;
        RECT 123.655 105.795 123.905 106.255 ;
        RECT 124.075 105.805 124.410 105.975 ;
        RECT 124.605 105.805 125.280 105.975 ;
        RECT 124.075 105.665 124.245 105.805 ;
        RECT 123.570 104.675 123.850 105.625 ;
        RECT 124.020 105.535 124.245 105.665 ;
        RECT 124.020 104.430 124.190 105.535 ;
        RECT 124.415 105.385 124.940 105.605 ;
        RECT 124.360 104.620 124.600 105.215 ;
        RECT 124.770 104.685 124.940 105.385 ;
        RECT 125.110 105.025 125.280 105.805 ;
        RECT 125.600 105.755 125.970 106.255 ;
        RECT 126.150 105.805 126.555 105.975 ;
        RECT 126.725 105.805 127.510 105.975 ;
        RECT 126.150 105.575 126.320 105.805 ;
        RECT 125.490 105.275 126.320 105.575 ;
        RECT 126.705 105.305 127.170 105.635 ;
        RECT 125.490 105.245 125.690 105.275 ;
        RECT 125.810 105.025 125.980 105.095 ;
        RECT 125.110 104.855 125.980 105.025 ;
        RECT 125.470 104.765 125.980 104.855 ;
        RECT 124.020 104.300 124.325 104.430 ;
        RECT 124.770 104.320 125.300 104.685 ;
        RECT 123.640 103.705 123.905 104.165 ;
        RECT 124.075 103.875 124.325 104.300 ;
        RECT 125.470 104.150 125.640 104.765 ;
        RECT 124.535 103.980 125.640 104.150 ;
        RECT 125.810 103.705 125.980 104.505 ;
        RECT 126.150 104.205 126.320 105.275 ;
        RECT 126.490 104.375 126.680 105.095 ;
        RECT 126.850 104.345 127.170 105.305 ;
        RECT 127.340 105.345 127.510 105.805 ;
        RECT 127.785 105.725 127.995 106.255 ;
        RECT 128.255 105.515 128.585 106.040 ;
        RECT 128.755 105.645 128.925 106.255 ;
        RECT 129.095 105.600 129.425 106.035 ;
        RECT 129.095 105.515 129.475 105.600 ;
        RECT 128.385 105.345 128.585 105.515 ;
        RECT 129.250 105.475 129.475 105.515 ;
        RECT 127.340 105.015 128.215 105.345 ;
        RECT 128.385 105.015 129.135 105.345 ;
        RECT 126.150 103.875 126.400 104.205 ;
        RECT 127.340 104.175 127.510 105.015 ;
        RECT 128.385 104.810 128.575 105.015 ;
        RECT 129.305 104.895 129.475 105.475 ;
        RECT 129.260 104.845 129.475 104.895 ;
        RECT 127.680 104.435 128.575 104.810 ;
        RECT 129.085 104.765 129.475 104.845 ;
        RECT 129.650 105.515 129.905 106.085 ;
        RECT 130.075 105.855 130.405 106.255 ;
        RECT 130.830 105.720 131.360 106.085 ;
        RECT 131.550 105.915 131.825 106.085 ;
        RECT 131.545 105.745 131.825 105.915 ;
        RECT 130.830 105.685 131.005 105.720 ;
        RECT 130.075 105.515 131.005 105.685 ;
        RECT 129.650 104.845 129.820 105.515 ;
        RECT 130.075 105.345 130.245 105.515 ;
        RECT 129.990 105.015 130.245 105.345 ;
        RECT 130.470 105.015 130.665 105.345 ;
        RECT 126.625 104.005 127.510 104.175 ;
        RECT 127.690 103.705 128.005 104.205 ;
        RECT 128.235 103.875 128.575 104.435 ;
        RECT 128.745 103.705 128.915 104.715 ;
        RECT 129.085 103.920 129.415 104.765 ;
        RECT 129.650 103.875 129.985 104.845 ;
        RECT 130.155 103.705 130.325 104.845 ;
        RECT 130.495 104.045 130.665 105.015 ;
        RECT 130.835 104.385 131.005 105.515 ;
        RECT 131.175 104.725 131.345 105.525 ;
        RECT 131.550 104.925 131.825 105.745 ;
        RECT 131.995 104.725 132.185 106.085 ;
        RECT 132.365 105.720 132.875 106.255 ;
        RECT 133.095 105.445 133.340 106.050 ;
        RECT 133.785 105.485 135.455 106.255 ;
        RECT 135.630 105.515 135.885 106.085 ;
        RECT 136.055 105.855 136.385 106.255 ;
        RECT 136.810 105.720 137.340 106.085 ;
        RECT 137.530 105.915 137.805 106.085 ;
        RECT 137.525 105.745 137.805 105.915 ;
        RECT 136.810 105.685 136.985 105.720 ;
        RECT 136.055 105.515 136.985 105.685 ;
        RECT 132.385 105.275 133.615 105.445 ;
        RECT 131.175 104.555 132.185 104.725 ;
        RECT 132.355 104.710 133.105 104.900 ;
        RECT 130.835 104.215 131.960 104.385 ;
        RECT 132.355 104.045 132.525 104.710 ;
        RECT 133.275 104.465 133.615 105.275 ;
        RECT 133.785 104.965 134.535 105.485 ;
        RECT 134.705 104.795 135.455 105.315 ;
        RECT 130.495 103.875 132.525 104.045 ;
        RECT 132.695 103.705 132.865 104.465 ;
        RECT 133.100 104.055 133.615 104.465 ;
        RECT 133.785 103.705 135.455 104.795 ;
        RECT 135.630 104.845 135.800 105.515 ;
        RECT 136.055 105.345 136.225 105.515 ;
        RECT 135.970 105.015 136.225 105.345 ;
        RECT 136.450 105.015 136.645 105.345 ;
        RECT 135.630 103.875 135.965 104.845 ;
        RECT 136.135 103.705 136.305 104.845 ;
        RECT 136.475 104.045 136.645 105.015 ;
        RECT 136.815 104.385 136.985 105.515 ;
        RECT 137.155 104.725 137.325 105.525 ;
        RECT 137.530 104.925 137.805 105.745 ;
        RECT 137.975 104.725 138.165 106.085 ;
        RECT 138.345 105.720 138.855 106.255 ;
        RECT 139.075 105.445 139.320 106.050 ;
        RECT 139.770 105.515 140.025 106.085 ;
        RECT 140.195 105.855 140.525 106.255 ;
        RECT 140.950 105.720 141.480 106.085 ;
        RECT 140.950 105.685 141.125 105.720 ;
        RECT 140.195 105.515 141.125 105.685 ;
        RECT 138.365 105.275 139.595 105.445 ;
        RECT 137.155 104.555 138.165 104.725 ;
        RECT 138.335 104.710 139.085 104.900 ;
        RECT 136.815 104.215 137.940 104.385 ;
        RECT 138.335 104.045 138.505 104.710 ;
        RECT 139.255 104.465 139.595 105.275 ;
        RECT 136.475 103.875 138.505 104.045 ;
        RECT 138.675 103.705 138.845 104.465 ;
        RECT 139.080 104.055 139.595 104.465 ;
        RECT 139.770 104.845 139.940 105.515 ;
        RECT 140.195 105.345 140.365 105.515 ;
        RECT 140.110 105.015 140.365 105.345 ;
        RECT 140.590 105.015 140.785 105.345 ;
        RECT 139.770 103.875 140.105 104.845 ;
        RECT 140.275 103.705 140.445 104.845 ;
        RECT 140.615 104.045 140.785 105.015 ;
        RECT 140.955 104.385 141.125 105.515 ;
        RECT 141.295 104.725 141.465 105.525 ;
        RECT 141.670 105.235 141.945 106.085 ;
        RECT 141.665 105.065 141.945 105.235 ;
        RECT 141.670 104.925 141.945 105.065 ;
        RECT 142.115 104.725 142.305 106.085 ;
        RECT 142.485 105.720 142.995 106.255 ;
        RECT 143.215 105.445 143.460 106.050 ;
        RECT 143.995 105.705 144.165 106.085 ;
        RECT 144.380 105.875 144.710 106.255 ;
        RECT 143.995 105.535 144.710 105.705 ;
        RECT 142.505 105.275 143.735 105.445 ;
        RECT 141.295 104.555 142.305 104.725 ;
        RECT 142.475 104.710 143.225 104.900 ;
        RECT 140.955 104.215 142.080 104.385 ;
        RECT 142.475 104.045 142.645 104.710 ;
        RECT 143.395 104.465 143.735 105.275 ;
        RECT 143.905 104.985 144.260 105.355 ;
        RECT 144.540 105.345 144.710 105.535 ;
        RECT 144.880 105.510 145.135 106.085 ;
        RECT 144.540 105.015 144.795 105.345 ;
        RECT 144.540 104.805 144.710 105.015 ;
        RECT 140.615 103.875 142.645 104.045 ;
        RECT 142.815 103.705 142.985 104.465 ;
        RECT 143.220 104.055 143.735 104.465 ;
        RECT 143.995 104.635 144.710 104.805 ;
        RECT 144.965 104.780 145.135 105.510 ;
        RECT 145.310 105.415 145.570 106.255 ;
        RECT 145.745 105.505 146.955 106.255 ;
        RECT 143.995 103.875 144.165 104.635 ;
        RECT 144.380 103.705 144.710 104.465 ;
        RECT 144.880 103.875 145.135 104.780 ;
        RECT 145.310 103.705 145.570 104.855 ;
        RECT 145.745 104.795 146.265 105.335 ;
        RECT 146.435 104.965 146.955 105.505 ;
        RECT 145.745 103.705 146.955 104.795 ;
        RECT 17.320 103.535 147.040 103.705 ;
        RECT 17.405 102.445 18.615 103.535 ;
        RECT 19.305 102.475 19.635 103.320 ;
        RECT 19.805 102.525 19.975 103.535 ;
        RECT 20.145 102.805 20.485 103.365 ;
        RECT 20.715 103.035 21.030 103.535 ;
        RECT 21.210 103.065 22.095 103.235 ;
        RECT 17.405 101.735 17.925 102.275 ;
        RECT 18.095 101.905 18.615 102.445 ;
        RECT 19.245 102.395 19.635 102.475 ;
        RECT 20.145 102.430 21.040 102.805 ;
        RECT 19.245 102.345 19.460 102.395 ;
        RECT 19.245 101.765 19.415 102.345 ;
        RECT 20.145 102.225 20.335 102.430 ;
        RECT 21.210 102.225 21.380 103.065 ;
        RECT 22.320 103.035 22.570 103.365 ;
        RECT 19.585 101.895 20.335 102.225 ;
        RECT 20.505 101.895 21.380 102.225 ;
        RECT 17.405 100.985 18.615 101.735 ;
        RECT 19.245 101.725 19.470 101.765 ;
        RECT 20.135 101.725 20.335 101.895 ;
        RECT 19.245 101.640 19.625 101.725 ;
        RECT 19.295 101.205 19.625 101.640 ;
        RECT 19.795 100.985 19.965 101.595 ;
        RECT 20.135 101.200 20.465 101.725 ;
        RECT 20.725 100.985 20.935 101.515 ;
        RECT 21.210 101.435 21.380 101.895 ;
        RECT 21.550 101.935 21.870 102.895 ;
        RECT 22.040 102.145 22.230 102.865 ;
        RECT 22.400 101.965 22.570 103.035 ;
        RECT 22.740 102.735 22.910 103.535 ;
        RECT 23.080 103.090 24.185 103.260 ;
        RECT 23.080 102.475 23.250 103.090 ;
        RECT 24.395 102.940 24.645 103.365 ;
        RECT 24.815 103.075 25.080 103.535 ;
        RECT 23.420 102.555 23.950 102.920 ;
        RECT 24.395 102.810 24.700 102.940 ;
        RECT 22.740 102.385 23.250 102.475 ;
        RECT 22.740 102.215 23.610 102.385 ;
        RECT 22.740 102.145 22.910 102.215 ;
        RECT 23.030 101.965 23.230 101.995 ;
        RECT 21.550 101.605 22.015 101.935 ;
        RECT 22.400 101.665 23.230 101.965 ;
        RECT 22.400 101.435 22.570 101.665 ;
        RECT 21.210 101.265 21.995 101.435 ;
        RECT 22.165 101.265 22.570 101.435 ;
        RECT 22.750 100.985 23.120 101.485 ;
        RECT 23.440 101.435 23.610 102.215 ;
        RECT 23.780 101.855 23.950 102.555 ;
        RECT 24.120 102.025 24.360 102.620 ;
        RECT 23.780 101.635 24.305 101.855 ;
        RECT 24.530 101.705 24.700 102.810 ;
        RECT 24.475 101.575 24.700 101.705 ;
        RECT 24.870 101.615 25.150 102.565 ;
        RECT 24.475 101.435 24.645 101.575 ;
        RECT 23.440 101.265 24.115 101.435 ;
        RECT 24.310 101.265 24.645 101.435 ;
        RECT 24.815 100.985 25.065 101.445 ;
        RECT 25.320 101.245 25.505 103.365 ;
        RECT 25.675 103.035 26.005 103.535 ;
        RECT 26.175 102.865 26.345 103.365 ;
        RECT 25.680 102.695 26.345 102.865 ;
        RECT 25.680 101.705 25.910 102.695 ;
        RECT 26.080 101.875 26.430 102.525 ;
        RECT 26.605 102.445 30.115 103.535 ;
        RECT 26.605 101.755 28.255 102.275 ;
        RECT 28.425 101.925 30.115 102.445 ;
        RECT 30.285 102.370 30.575 103.535 ;
        RECT 30.750 102.395 31.085 103.365 ;
        RECT 31.255 102.395 31.425 103.535 ;
        RECT 31.595 103.195 33.625 103.365 ;
        RECT 25.680 101.535 26.345 101.705 ;
        RECT 25.675 100.985 26.005 101.365 ;
        RECT 26.175 101.245 26.345 101.535 ;
        RECT 26.605 100.985 30.115 101.755 ;
        RECT 30.750 101.725 30.920 102.395 ;
        RECT 31.595 102.225 31.765 103.195 ;
        RECT 31.090 101.895 31.345 102.225 ;
        RECT 31.570 101.895 31.765 102.225 ;
        RECT 31.935 102.855 33.060 103.025 ;
        RECT 31.175 101.725 31.345 101.895 ;
        RECT 31.935 101.725 32.105 102.855 ;
        RECT 30.285 100.985 30.575 101.710 ;
        RECT 30.750 101.155 31.005 101.725 ;
        RECT 31.175 101.555 32.105 101.725 ;
        RECT 32.275 102.515 33.285 102.685 ;
        RECT 32.275 101.715 32.445 102.515 ;
        RECT 32.650 102.175 32.925 102.315 ;
        RECT 32.645 102.005 32.925 102.175 ;
        RECT 31.930 101.520 32.105 101.555 ;
        RECT 31.175 100.985 31.505 101.385 ;
        RECT 31.930 101.155 32.460 101.520 ;
        RECT 32.650 101.155 32.925 102.005 ;
        RECT 33.095 101.155 33.285 102.515 ;
        RECT 33.455 102.530 33.625 103.195 ;
        RECT 33.795 102.775 33.965 103.535 ;
        RECT 34.200 102.775 34.715 103.185 ;
        RECT 34.885 103.100 40.230 103.535 ;
        RECT 40.405 103.100 45.750 103.535 ;
        RECT 45.925 103.100 51.270 103.535 ;
        RECT 33.455 102.340 34.205 102.530 ;
        RECT 34.375 101.965 34.715 102.775 ;
        RECT 33.485 101.795 34.715 101.965 ;
        RECT 33.465 100.985 33.975 101.520 ;
        RECT 34.195 101.190 34.440 101.795 ;
        RECT 36.470 101.530 36.810 102.360 ;
        RECT 38.290 101.850 38.640 103.100 ;
        RECT 41.990 101.530 42.330 102.360 ;
        RECT 43.810 101.850 44.160 103.100 ;
        RECT 47.510 101.530 47.850 102.360 ;
        RECT 49.330 101.850 49.680 103.100 ;
        RECT 51.445 102.445 54.955 103.535 ;
        RECT 51.445 101.755 53.095 102.275 ;
        RECT 53.265 101.925 54.955 102.445 ;
        RECT 56.045 102.370 56.335 103.535 ;
        RECT 56.505 103.100 61.850 103.535 ;
        RECT 34.885 100.985 40.230 101.530 ;
        RECT 40.405 100.985 45.750 101.530 ;
        RECT 45.925 100.985 51.270 101.530 ;
        RECT 51.445 100.985 54.955 101.755 ;
        RECT 56.045 100.985 56.335 101.710 ;
        RECT 58.090 101.530 58.430 102.360 ;
        RECT 59.910 101.850 60.260 103.100 ;
        RECT 62.025 102.445 63.235 103.535 ;
        RECT 63.495 102.865 63.665 103.365 ;
        RECT 63.835 103.035 64.165 103.535 ;
        RECT 63.495 102.695 64.160 102.865 ;
        RECT 62.025 101.735 62.545 102.275 ;
        RECT 62.715 101.905 63.235 102.445 ;
        RECT 63.410 101.875 63.760 102.525 ;
        RECT 56.505 100.985 61.850 101.530 ;
        RECT 62.025 100.985 63.235 101.735 ;
        RECT 63.930 101.705 64.160 102.695 ;
        RECT 63.495 101.535 64.160 101.705 ;
        RECT 63.495 101.245 63.665 101.535 ;
        RECT 63.835 100.985 64.165 101.365 ;
        RECT 64.335 101.245 64.520 103.365 ;
        RECT 64.760 103.075 65.025 103.535 ;
        RECT 65.195 102.940 65.445 103.365 ;
        RECT 65.655 103.090 66.760 103.260 ;
        RECT 65.140 102.810 65.445 102.940 ;
        RECT 64.690 101.615 64.970 102.565 ;
        RECT 65.140 101.705 65.310 102.810 ;
        RECT 65.480 102.025 65.720 102.620 ;
        RECT 65.890 102.555 66.420 102.920 ;
        RECT 65.890 101.855 66.060 102.555 ;
        RECT 66.590 102.475 66.760 103.090 ;
        RECT 66.930 102.735 67.100 103.535 ;
        RECT 67.270 103.035 67.520 103.365 ;
        RECT 67.745 103.065 68.630 103.235 ;
        RECT 66.590 102.385 67.100 102.475 ;
        RECT 65.140 101.575 65.365 101.705 ;
        RECT 65.535 101.635 66.060 101.855 ;
        RECT 66.230 102.215 67.100 102.385 ;
        RECT 64.775 100.985 65.025 101.445 ;
        RECT 65.195 101.435 65.365 101.575 ;
        RECT 66.230 101.435 66.400 102.215 ;
        RECT 66.930 102.145 67.100 102.215 ;
        RECT 66.610 101.965 66.810 101.995 ;
        RECT 67.270 101.965 67.440 103.035 ;
        RECT 67.610 102.145 67.800 102.865 ;
        RECT 66.610 101.665 67.440 101.965 ;
        RECT 67.970 101.935 68.290 102.895 ;
        RECT 65.195 101.265 65.530 101.435 ;
        RECT 65.725 101.265 66.400 101.435 ;
        RECT 66.720 100.985 67.090 101.485 ;
        RECT 67.270 101.435 67.440 101.665 ;
        RECT 67.825 101.605 68.290 101.935 ;
        RECT 68.460 102.225 68.630 103.065 ;
        RECT 68.810 103.035 69.125 103.535 ;
        RECT 69.355 102.805 69.695 103.365 ;
        RECT 68.800 102.430 69.695 102.805 ;
        RECT 69.865 102.525 70.035 103.535 ;
        RECT 69.505 102.225 69.695 102.430 ;
        RECT 70.205 102.475 70.535 103.320 ;
        RECT 70.205 102.395 70.595 102.475 ;
        RECT 70.380 102.345 70.595 102.395 ;
        RECT 68.460 101.895 69.335 102.225 ;
        RECT 69.505 101.895 70.255 102.225 ;
        RECT 68.460 101.435 68.630 101.895 ;
        RECT 69.505 101.725 69.705 101.895 ;
        RECT 70.425 101.765 70.595 102.345 ;
        RECT 70.370 101.725 70.595 101.765 ;
        RECT 67.270 101.265 67.675 101.435 ;
        RECT 67.845 101.265 68.630 101.435 ;
        RECT 68.905 100.985 69.115 101.515 ;
        RECT 69.375 101.200 69.705 101.725 ;
        RECT 70.215 101.640 70.595 101.725 ;
        RECT 70.770 102.395 71.105 103.365 ;
        RECT 71.275 102.395 71.445 103.535 ;
        RECT 71.615 103.195 73.645 103.365 ;
        RECT 70.770 101.725 70.940 102.395 ;
        RECT 71.615 102.225 71.785 103.195 ;
        RECT 71.110 101.895 71.365 102.225 ;
        RECT 71.590 101.895 71.785 102.225 ;
        RECT 71.955 102.855 73.080 103.025 ;
        RECT 71.195 101.725 71.365 101.895 ;
        RECT 71.955 101.725 72.125 102.855 ;
        RECT 69.875 100.985 70.045 101.595 ;
        RECT 70.215 101.205 70.545 101.640 ;
        RECT 70.770 101.155 71.025 101.725 ;
        RECT 71.195 101.555 72.125 101.725 ;
        RECT 72.295 102.515 73.305 102.685 ;
        RECT 72.295 101.715 72.465 102.515 ;
        RECT 72.670 102.175 72.945 102.315 ;
        RECT 72.665 102.005 72.945 102.175 ;
        RECT 71.950 101.520 72.125 101.555 ;
        RECT 71.195 100.985 71.525 101.385 ;
        RECT 71.950 101.155 72.480 101.520 ;
        RECT 72.670 101.155 72.945 102.005 ;
        RECT 73.115 101.155 73.305 102.515 ;
        RECT 73.475 102.530 73.645 103.195 ;
        RECT 73.815 102.775 73.985 103.535 ;
        RECT 74.220 102.775 74.735 103.185 ;
        RECT 74.905 103.100 80.250 103.535 ;
        RECT 73.475 102.340 74.225 102.530 ;
        RECT 74.395 101.965 74.735 102.775 ;
        RECT 73.505 101.795 74.735 101.965 ;
        RECT 73.485 100.985 73.995 101.520 ;
        RECT 74.215 101.190 74.460 101.795 ;
        RECT 76.490 101.530 76.830 102.360 ;
        RECT 78.310 101.850 78.660 103.100 ;
        RECT 80.425 102.445 81.635 103.535 ;
        RECT 80.425 101.735 80.945 102.275 ;
        RECT 81.115 101.905 81.635 102.445 ;
        RECT 81.805 102.370 82.095 103.535 ;
        RECT 82.355 102.915 82.525 103.345 ;
        RECT 82.695 103.085 83.025 103.535 ;
        RECT 82.355 102.685 83.030 102.915 ;
        RECT 74.905 100.985 80.250 101.530 ;
        RECT 80.425 100.985 81.635 101.735 ;
        RECT 81.805 100.985 82.095 101.710 ;
        RECT 82.325 101.665 82.625 102.515 ;
        RECT 82.795 102.035 83.030 102.685 ;
        RECT 83.200 102.375 83.485 103.320 ;
        RECT 83.665 103.065 84.350 103.535 ;
        RECT 83.660 102.545 84.355 102.855 ;
        RECT 84.530 102.480 84.835 103.265 ;
        RECT 83.200 102.225 84.060 102.375 ;
        RECT 83.200 102.205 84.485 102.225 ;
        RECT 82.795 101.705 83.330 102.035 ;
        RECT 83.500 101.845 84.485 102.205 ;
        RECT 82.795 101.555 83.015 101.705 ;
        RECT 82.270 100.985 82.605 101.490 ;
        RECT 82.775 101.180 83.015 101.555 ;
        RECT 83.500 101.510 83.670 101.845 ;
        RECT 84.660 101.675 84.835 102.480 ;
        RECT 85.025 102.445 88.535 103.535 ;
        RECT 83.295 101.315 83.670 101.510 ;
        RECT 83.295 101.170 83.465 101.315 ;
        RECT 84.030 100.985 84.425 101.480 ;
        RECT 84.595 101.155 84.835 101.675 ;
        RECT 85.025 101.755 86.675 102.275 ;
        RECT 86.845 101.925 88.535 102.445 ;
        RECT 88.705 102.685 88.965 103.365 ;
        RECT 89.135 102.755 89.385 103.535 ;
        RECT 89.635 102.985 89.885 103.365 ;
        RECT 90.055 103.155 90.410 103.535 ;
        RECT 91.415 103.145 91.750 103.365 ;
        RECT 91.015 102.985 91.245 103.025 ;
        RECT 89.635 102.785 91.245 102.985 ;
        RECT 89.635 102.775 90.470 102.785 ;
        RECT 91.060 102.695 91.245 102.785 ;
        RECT 85.025 100.985 88.535 101.755 ;
        RECT 88.705 101.485 88.875 102.685 ;
        RECT 90.575 102.585 90.905 102.615 ;
        RECT 89.105 102.525 90.905 102.585 ;
        RECT 91.495 102.525 91.750 103.145 ;
        RECT 91.925 103.100 97.270 103.535 ;
        RECT 97.445 103.100 102.790 103.535 ;
        RECT 89.045 102.415 91.750 102.525 ;
        RECT 89.045 102.380 89.245 102.415 ;
        RECT 89.045 101.805 89.215 102.380 ;
        RECT 90.575 102.355 91.750 102.415 ;
        RECT 89.445 101.940 89.855 102.245 ;
        RECT 90.025 101.975 90.355 102.185 ;
        RECT 89.045 101.685 89.315 101.805 ;
        RECT 89.045 101.640 89.890 101.685 ;
        RECT 89.135 101.515 89.890 101.640 ;
        RECT 90.145 101.575 90.355 101.975 ;
        RECT 90.600 101.975 91.075 102.185 ;
        RECT 91.265 101.975 91.755 102.175 ;
        RECT 90.600 101.575 90.820 101.975 ;
        RECT 88.705 101.155 88.965 101.485 ;
        RECT 89.720 101.365 89.890 101.515 ;
        RECT 89.135 100.985 89.465 101.345 ;
        RECT 89.720 101.155 91.020 101.365 ;
        RECT 91.295 100.985 91.750 101.750 ;
        RECT 93.510 101.530 93.850 102.360 ;
        RECT 95.330 101.850 95.680 103.100 ;
        RECT 99.030 101.530 99.370 102.360 ;
        RECT 100.850 101.850 101.200 103.100 ;
        RECT 102.985 102.480 103.290 103.265 ;
        RECT 103.470 103.065 104.155 103.535 ;
        RECT 103.465 102.545 104.160 102.855 ;
        RECT 102.985 101.675 103.160 102.480 ;
        RECT 104.335 102.375 104.620 103.320 ;
        RECT 104.795 103.085 105.125 103.535 ;
        RECT 105.295 102.915 105.465 103.345 ;
        RECT 103.760 102.225 104.620 102.375 ;
        RECT 103.335 102.205 104.620 102.225 ;
        RECT 104.790 102.685 105.465 102.915 ;
        RECT 103.335 101.845 104.320 102.205 ;
        RECT 104.790 102.035 105.025 102.685 ;
        RECT 91.925 100.985 97.270 101.530 ;
        RECT 97.445 100.985 102.790 101.530 ;
        RECT 102.985 101.155 103.225 101.675 ;
        RECT 104.150 101.510 104.320 101.845 ;
        RECT 104.490 101.705 105.025 102.035 ;
        RECT 104.805 101.555 105.025 101.705 ;
        RECT 105.195 101.665 105.495 102.515 ;
        RECT 105.725 102.445 107.395 103.535 ;
        RECT 105.725 101.755 106.475 102.275 ;
        RECT 106.645 101.925 107.395 102.445 ;
        RECT 107.565 102.370 107.855 103.535 ;
        RECT 108.115 102.915 108.285 103.345 ;
        RECT 108.455 103.085 108.785 103.535 ;
        RECT 108.115 102.685 108.790 102.915 ;
        RECT 103.395 100.985 103.790 101.480 ;
        RECT 104.150 101.315 104.525 101.510 ;
        RECT 104.355 101.170 104.525 101.315 ;
        RECT 104.805 101.180 105.045 101.555 ;
        RECT 105.215 100.985 105.550 101.490 ;
        RECT 105.725 100.985 107.395 101.755 ;
        RECT 107.565 100.985 107.855 101.710 ;
        RECT 108.085 101.665 108.385 102.515 ;
        RECT 108.555 102.035 108.790 102.685 ;
        RECT 108.960 102.375 109.245 103.320 ;
        RECT 109.425 103.065 110.110 103.535 ;
        RECT 109.420 102.545 110.115 102.855 ;
        RECT 110.290 102.480 110.595 103.265 ;
        RECT 108.960 102.225 109.820 102.375 ;
        RECT 108.960 102.205 110.245 102.225 ;
        RECT 108.555 101.705 109.090 102.035 ;
        RECT 109.260 101.845 110.245 102.205 ;
        RECT 108.555 101.555 108.775 101.705 ;
        RECT 108.030 100.985 108.365 101.490 ;
        RECT 108.535 101.180 108.775 101.555 ;
        RECT 109.260 101.510 109.430 101.845 ;
        RECT 110.420 101.675 110.595 102.480 ;
        RECT 110.785 102.445 112.455 103.535 ;
        RECT 109.055 101.315 109.430 101.510 ;
        RECT 109.055 101.170 109.225 101.315 ;
        RECT 109.790 100.985 110.185 101.480 ;
        RECT 110.355 101.155 110.595 101.675 ;
        RECT 110.785 101.755 111.535 102.275 ;
        RECT 111.705 101.925 112.455 102.445 ;
        RECT 113.085 102.775 113.600 103.185 ;
        RECT 113.835 102.775 114.005 103.535 ;
        RECT 114.175 103.195 116.205 103.365 ;
        RECT 113.085 101.965 113.425 102.775 ;
        RECT 114.175 102.530 114.345 103.195 ;
        RECT 114.740 102.855 115.865 103.025 ;
        RECT 113.595 102.340 114.345 102.530 ;
        RECT 114.515 102.515 115.525 102.685 ;
        RECT 113.085 101.795 114.315 101.965 ;
        RECT 110.785 100.985 112.455 101.755 ;
        RECT 113.360 101.190 113.605 101.795 ;
        RECT 113.825 100.985 114.335 101.520 ;
        RECT 114.515 101.155 114.705 102.515 ;
        RECT 114.875 102.175 115.150 102.315 ;
        RECT 114.875 102.005 115.155 102.175 ;
        RECT 114.875 101.155 115.150 102.005 ;
        RECT 115.355 101.715 115.525 102.515 ;
        RECT 115.695 101.725 115.865 102.855 ;
        RECT 116.035 102.225 116.205 103.195 ;
        RECT 116.375 102.395 116.545 103.535 ;
        RECT 116.715 102.395 117.050 103.365 ;
        RECT 117.315 102.865 117.485 103.365 ;
        RECT 117.655 103.035 117.985 103.535 ;
        RECT 117.315 102.695 117.980 102.865 ;
        RECT 116.035 101.895 116.230 102.225 ;
        RECT 116.455 101.895 116.710 102.225 ;
        RECT 116.455 101.725 116.625 101.895 ;
        RECT 116.880 101.725 117.050 102.395 ;
        RECT 117.230 101.875 117.580 102.525 ;
        RECT 115.695 101.555 116.625 101.725 ;
        RECT 115.695 101.520 115.870 101.555 ;
        RECT 115.340 101.155 115.870 101.520 ;
        RECT 116.295 100.985 116.625 101.385 ;
        RECT 116.795 101.155 117.050 101.725 ;
        RECT 117.750 101.705 117.980 102.695 ;
        RECT 117.315 101.535 117.980 101.705 ;
        RECT 117.315 101.245 117.485 101.535 ;
        RECT 117.655 100.985 117.985 101.365 ;
        RECT 118.155 101.245 118.340 103.365 ;
        RECT 118.580 103.075 118.845 103.535 ;
        RECT 119.015 102.940 119.265 103.365 ;
        RECT 119.475 103.090 120.580 103.260 ;
        RECT 118.960 102.810 119.265 102.940 ;
        RECT 118.510 101.615 118.790 102.565 ;
        RECT 118.960 101.705 119.130 102.810 ;
        RECT 119.300 102.025 119.540 102.620 ;
        RECT 119.710 102.555 120.240 102.920 ;
        RECT 119.710 101.855 119.880 102.555 ;
        RECT 120.410 102.475 120.580 103.090 ;
        RECT 120.750 102.735 120.920 103.535 ;
        RECT 121.090 103.035 121.340 103.365 ;
        RECT 121.565 103.065 122.450 103.235 ;
        RECT 120.410 102.385 120.920 102.475 ;
        RECT 118.960 101.575 119.185 101.705 ;
        RECT 119.355 101.635 119.880 101.855 ;
        RECT 120.050 102.215 120.920 102.385 ;
        RECT 118.595 100.985 118.845 101.445 ;
        RECT 119.015 101.435 119.185 101.575 ;
        RECT 120.050 101.435 120.220 102.215 ;
        RECT 120.750 102.145 120.920 102.215 ;
        RECT 120.430 101.965 120.630 101.995 ;
        RECT 121.090 101.965 121.260 103.035 ;
        RECT 121.430 102.145 121.620 102.865 ;
        RECT 120.430 101.665 121.260 101.965 ;
        RECT 121.790 101.935 122.110 102.895 ;
        RECT 119.015 101.265 119.350 101.435 ;
        RECT 119.545 101.265 120.220 101.435 ;
        RECT 120.540 100.985 120.910 101.485 ;
        RECT 121.090 101.435 121.260 101.665 ;
        RECT 121.645 101.605 122.110 101.935 ;
        RECT 122.280 102.225 122.450 103.065 ;
        RECT 122.630 103.035 122.945 103.535 ;
        RECT 123.175 102.805 123.515 103.365 ;
        RECT 122.620 102.430 123.515 102.805 ;
        RECT 123.685 102.525 123.855 103.535 ;
        RECT 123.325 102.225 123.515 102.430 ;
        RECT 124.025 102.475 124.355 103.320 ;
        RECT 124.585 103.100 129.930 103.535 ;
        RECT 124.025 102.395 124.415 102.475 ;
        RECT 124.200 102.345 124.415 102.395 ;
        RECT 122.280 101.895 123.155 102.225 ;
        RECT 123.325 101.895 124.075 102.225 ;
        RECT 122.280 101.435 122.450 101.895 ;
        RECT 123.325 101.725 123.525 101.895 ;
        RECT 124.245 101.765 124.415 102.345 ;
        RECT 124.190 101.725 124.415 101.765 ;
        RECT 121.090 101.265 121.495 101.435 ;
        RECT 121.665 101.265 122.450 101.435 ;
        RECT 122.725 100.985 122.935 101.515 ;
        RECT 123.195 101.200 123.525 101.725 ;
        RECT 124.035 101.640 124.415 101.725 ;
        RECT 123.695 100.985 123.865 101.595 ;
        RECT 124.035 101.205 124.365 101.640 ;
        RECT 126.170 101.530 126.510 102.360 ;
        RECT 127.990 101.850 128.340 103.100 ;
        RECT 130.655 102.915 130.825 103.345 ;
        RECT 130.995 103.085 131.325 103.535 ;
        RECT 130.655 102.685 131.330 102.915 ;
        RECT 130.625 101.665 130.925 102.515 ;
        RECT 131.095 102.035 131.330 102.685 ;
        RECT 131.500 102.375 131.785 103.320 ;
        RECT 131.965 103.065 132.650 103.535 ;
        RECT 131.960 102.545 132.655 102.855 ;
        RECT 132.830 102.480 133.135 103.265 ;
        RECT 131.500 102.225 132.360 102.375 ;
        RECT 131.500 102.205 132.785 102.225 ;
        RECT 131.095 101.705 131.630 102.035 ;
        RECT 131.800 101.845 132.785 102.205 ;
        RECT 131.095 101.555 131.315 101.705 ;
        RECT 124.585 100.985 129.930 101.530 ;
        RECT 130.570 100.985 130.905 101.490 ;
        RECT 131.075 101.180 131.315 101.555 ;
        RECT 131.800 101.510 131.970 101.845 ;
        RECT 132.960 101.675 133.135 102.480 ;
        RECT 133.325 102.370 133.615 103.535 ;
        RECT 133.785 102.445 135.455 103.535 ;
        RECT 136.175 102.865 136.345 103.365 ;
        RECT 136.515 103.035 136.845 103.535 ;
        RECT 136.175 102.695 136.840 102.865 ;
        RECT 133.785 101.755 134.535 102.275 ;
        RECT 134.705 101.925 135.455 102.445 ;
        RECT 136.090 101.875 136.440 102.525 ;
        RECT 131.595 101.315 131.970 101.510 ;
        RECT 131.595 101.170 131.765 101.315 ;
        RECT 132.330 100.985 132.725 101.480 ;
        RECT 132.895 101.155 133.135 101.675 ;
        RECT 133.325 100.985 133.615 101.710 ;
        RECT 133.785 100.985 135.455 101.755 ;
        RECT 136.610 101.705 136.840 102.695 ;
        RECT 136.175 101.535 136.840 101.705 ;
        RECT 136.175 101.245 136.345 101.535 ;
        RECT 136.515 100.985 136.845 101.365 ;
        RECT 137.015 101.245 137.200 103.365 ;
        RECT 137.440 103.075 137.705 103.535 ;
        RECT 137.875 102.940 138.125 103.365 ;
        RECT 138.335 103.090 139.440 103.260 ;
        RECT 137.820 102.810 138.125 102.940 ;
        RECT 137.370 101.615 137.650 102.565 ;
        RECT 137.820 101.705 137.990 102.810 ;
        RECT 138.160 102.025 138.400 102.620 ;
        RECT 138.570 102.555 139.100 102.920 ;
        RECT 138.570 101.855 138.740 102.555 ;
        RECT 139.270 102.475 139.440 103.090 ;
        RECT 139.610 102.735 139.780 103.535 ;
        RECT 139.950 103.035 140.200 103.365 ;
        RECT 140.425 103.065 141.310 103.235 ;
        RECT 139.270 102.385 139.780 102.475 ;
        RECT 137.820 101.575 138.045 101.705 ;
        RECT 138.215 101.635 138.740 101.855 ;
        RECT 138.910 102.215 139.780 102.385 ;
        RECT 137.455 100.985 137.705 101.445 ;
        RECT 137.875 101.435 138.045 101.575 ;
        RECT 138.910 101.435 139.080 102.215 ;
        RECT 139.610 102.145 139.780 102.215 ;
        RECT 139.290 101.965 139.490 101.995 ;
        RECT 139.950 101.965 140.120 103.035 ;
        RECT 140.290 102.145 140.480 102.865 ;
        RECT 139.290 101.665 140.120 101.965 ;
        RECT 140.650 101.935 140.970 102.895 ;
        RECT 137.875 101.265 138.210 101.435 ;
        RECT 138.405 101.265 139.080 101.435 ;
        RECT 139.400 100.985 139.770 101.485 ;
        RECT 139.950 101.435 140.120 101.665 ;
        RECT 140.505 101.605 140.970 101.935 ;
        RECT 141.140 102.225 141.310 103.065 ;
        RECT 141.490 103.035 141.805 103.535 ;
        RECT 142.035 102.805 142.375 103.365 ;
        RECT 141.480 102.430 142.375 102.805 ;
        RECT 142.545 102.525 142.715 103.535 ;
        RECT 142.185 102.225 142.375 102.430 ;
        RECT 142.885 102.475 143.215 103.320 ;
        RECT 143.995 102.605 144.165 103.365 ;
        RECT 144.380 102.775 144.710 103.535 ;
        RECT 142.885 102.395 143.275 102.475 ;
        RECT 143.995 102.435 144.710 102.605 ;
        RECT 144.880 102.460 145.135 103.365 ;
        RECT 143.060 102.345 143.275 102.395 ;
        RECT 141.140 101.895 142.015 102.225 ;
        RECT 142.185 101.895 142.935 102.225 ;
        RECT 141.140 101.435 141.310 101.895 ;
        RECT 142.185 101.725 142.385 101.895 ;
        RECT 143.105 101.765 143.275 102.345 ;
        RECT 143.905 101.885 144.260 102.255 ;
        RECT 144.540 102.225 144.710 102.435 ;
        RECT 144.540 101.895 144.795 102.225 ;
        RECT 143.050 101.725 143.275 101.765 ;
        RECT 139.950 101.265 140.355 101.435 ;
        RECT 140.525 101.265 141.310 101.435 ;
        RECT 141.585 100.985 141.795 101.515 ;
        RECT 142.055 101.200 142.385 101.725 ;
        RECT 142.895 101.640 143.275 101.725 ;
        RECT 144.540 101.705 144.710 101.895 ;
        RECT 144.965 101.730 145.135 102.460 ;
        RECT 145.310 102.385 145.570 103.535 ;
        RECT 145.745 102.445 146.955 103.535 ;
        RECT 145.745 101.905 146.265 102.445 ;
        RECT 142.555 100.985 142.725 101.595 ;
        RECT 142.895 101.205 143.225 101.640 ;
        RECT 143.995 101.535 144.710 101.705 ;
        RECT 143.995 101.155 144.165 101.535 ;
        RECT 144.380 100.985 144.710 101.365 ;
        RECT 144.880 101.155 145.135 101.730 ;
        RECT 145.310 100.985 145.570 101.825 ;
        RECT 146.435 101.735 146.955 102.275 ;
        RECT 145.745 100.985 146.955 101.735 ;
        RECT 17.320 100.815 147.040 100.985 ;
        RECT 17.405 100.065 18.615 100.815 ;
        RECT 17.405 99.525 17.925 100.065 ;
        RECT 18.790 99.975 19.050 100.815 ;
        RECT 19.225 100.070 19.480 100.645 ;
        RECT 19.650 100.435 19.980 100.815 ;
        RECT 20.195 100.265 20.365 100.645 ;
        RECT 19.650 100.095 20.365 100.265 ;
        RECT 21.135 100.160 21.465 100.595 ;
        RECT 21.635 100.205 21.805 100.815 ;
        RECT 18.095 99.355 18.615 99.895 ;
        RECT 17.405 98.265 18.615 99.355 ;
        RECT 18.790 98.265 19.050 99.415 ;
        RECT 19.225 99.340 19.395 100.070 ;
        RECT 19.650 99.905 19.820 100.095 ;
        RECT 21.085 100.075 21.465 100.160 ;
        RECT 21.975 100.075 22.305 100.600 ;
        RECT 22.565 100.285 22.775 100.815 ;
        RECT 23.050 100.365 23.835 100.535 ;
        RECT 24.005 100.365 24.410 100.535 ;
        RECT 21.085 100.035 21.310 100.075 ;
        RECT 19.565 99.575 19.820 99.905 ;
        RECT 19.650 99.365 19.820 99.575 ;
        RECT 20.100 99.545 20.455 99.915 ;
        RECT 21.085 99.455 21.255 100.035 ;
        RECT 21.975 99.905 22.175 100.075 ;
        RECT 23.050 99.905 23.220 100.365 ;
        RECT 21.425 99.575 22.175 99.905 ;
        RECT 22.345 99.575 23.220 99.905 ;
        RECT 21.085 99.405 21.300 99.455 ;
        RECT 19.225 98.435 19.480 99.340 ;
        RECT 19.650 99.195 20.365 99.365 ;
        RECT 21.085 99.325 21.475 99.405 ;
        RECT 19.650 98.265 19.980 99.025 ;
        RECT 20.195 98.435 20.365 99.195 ;
        RECT 21.145 98.480 21.475 99.325 ;
        RECT 21.985 99.370 22.175 99.575 ;
        RECT 21.645 98.265 21.815 99.275 ;
        RECT 21.985 98.995 22.880 99.370 ;
        RECT 21.985 98.435 22.325 98.995 ;
        RECT 22.555 98.265 22.870 98.765 ;
        RECT 23.050 98.735 23.220 99.575 ;
        RECT 23.390 99.865 23.855 100.195 ;
        RECT 24.240 100.135 24.410 100.365 ;
        RECT 24.590 100.315 24.960 100.815 ;
        RECT 25.280 100.365 25.955 100.535 ;
        RECT 26.150 100.365 26.485 100.535 ;
        RECT 23.390 98.905 23.710 99.865 ;
        RECT 24.240 99.835 25.070 100.135 ;
        RECT 23.880 98.935 24.070 99.655 ;
        RECT 24.240 98.765 24.410 99.835 ;
        RECT 24.870 99.805 25.070 99.835 ;
        RECT 24.580 99.585 24.750 99.655 ;
        RECT 25.280 99.585 25.450 100.365 ;
        RECT 26.315 100.225 26.485 100.365 ;
        RECT 26.655 100.355 26.905 100.815 ;
        RECT 24.580 99.415 25.450 99.585 ;
        RECT 25.620 99.945 26.145 100.165 ;
        RECT 26.315 100.095 26.540 100.225 ;
        RECT 24.580 99.325 25.090 99.415 ;
        RECT 23.050 98.565 23.935 98.735 ;
        RECT 24.160 98.435 24.410 98.765 ;
        RECT 24.580 98.265 24.750 99.065 ;
        RECT 24.920 98.710 25.090 99.325 ;
        RECT 25.620 99.245 25.790 99.945 ;
        RECT 25.260 98.880 25.790 99.245 ;
        RECT 25.960 99.180 26.200 99.775 ;
        RECT 26.370 98.990 26.540 100.095 ;
        RECT 26.710 99.235 26.990 100.185 ;
        RECT 26.235 98.860 26.540 98.990 ;
        RECT 24.920 98.540 26.025 98.710 ;
        RECT 26.235 98.435 26.485 98.860 ;
        RECT 26.655 98.265 26.920 98.725 ;
        RECT 27.160 98.435 27.345 100.555 ;
        RECT 27.515 100.435 27.845 100.815 ;
        RECT 28.015 100.265 28.185 100.555 ;
        RECT 27.520 100.095 28.185 100.265 ;
        RECT 27.520 99.105 27.750 100.095 ;
        RECT 28.450 100.075 28.705 100.645 ;
        RECT 28.875 100.415 29.205 100.815 ;
        RECT 29.630 100.280 30.160 100.645 ;
        RECT 29.630 100.245 29.805 100.280 ;
        RECT 28.875 100.075 29.805 100.245 ;
        RECT 30.350 100.135 30.625 100.645 ;
        RECT 27.920 99.275 28.270 99.925 ;
        RECT 28.450 99.405 28.620 100.075 ;
        RECT 28.875 99.905 29.045 100.075 ;
        RECT 28.790 99.575 29.045 99.905 ;
        RECT 29.270 99.575 29.465 99.905 ;
        RECT 27.520 98.935 28.185 99.105 ;
        RECT 27.515 98.265 27.845 98.765 ;
        RECT 28.015 98.435 28.185 98.935 ;
        RECT 28.450 98.435 28.785 99.405 ;
        RECT 28.955 98.265 29.125 99.405 ;
        RECT 29.295 98.605 29.465 99.575 ;
        RECT 29.635 98.945 29.805 100.075 ;
        RECT 29.975 99.285 30.145 100.085 ;
        RECT 30.345 99.965 30.625 100.135 ;
        RECT 30.350 99.485 30.625 99.965 ;
        RECT 30.795 99.285 30.985 100.645 ;
        RECT 31.165 100.280 31.675 100.815 ;
        RECT 31.895 100.005 32.140 100.610 ;
        RECT 32.585 100.270 37.930 100.815 ;
        RECT 31.185 99.835 32.415 100.005 ;
        RECT 29.975 99.115 30.985 99.285 ;
        RECT 31.155 99.270 31.905 99.460 ;
        RECT 29.635 98.775 30.760 98.945 ;
        RECT 31.155 98.605 31.325 99.270 ;
        RECT 32.075 99.025 32.415 99.835 ;
        RECT 34.170 99.440 34.510 100.270 ;
        RECT 38.105 100.045 41.615 100.815 ;
        RECT 41.785 100.065 42.995 100.815 ;
        RECT 43.165 100.090 43.455 100.815 ;
        RECT 43.625 100.270 48.970 100.815 ;
        RECT 49.145 100.270 54.490 100.815 ;
        RECT 54.665 100.270 60.010 100.815 ;
        RECT 29.295 98.435 31.325 98.605 ;
        RECT 31.495 98.265 31.665 99.025 ;
        RECT 31.900 98.615 32.415 99.025 ;
        RECT 35.990 98.700 36.340 99.950 ;
        RECT 38.105 99.525 39.755 100.045 ;
        RECT 39.925 99.355 41.615 99.875 ;
        RECT 41.785 99.525 42.305 100.065 ;
        RECT 42.475 99.355 42.995 99.895 ;
        RECT 45.210 99.440 45.550 100.270 ;
        RECT 32.585 98.265 37.930 98.700 ;
        RECT 38.105 98.265 41.615 99.355 ;
        RECT 41.785 98.265 42.995 99.355 ;
        RECT 43.165 98.265 43.455 99.430 ;
        RECT 47.030 98.700 47.380 99.950 ;
        RECT 50.730 99.440 51.070 100.270 ;
        RECT 52.550 98.700 52.900 99.950 ;
        RECT 56.250 99.440 56.590 100.270 ;
        RECT 60.185 100.045 63.695 100.815 ;
        RECT 64.345 100.125 64.585 100.645 ;
        RECT 64.755 100.320 65.150 100.815 ;
        RECT 65.715 100.485 65.885 100.630 ;
        RECT 65.510 100.290 65.885 100.485 ;
        RECT 58.070 98.700 58.420 99.950 ;
        RECT 60.185 99.525 61.835 100.045 ;
        RECT 62.005 99.355 63.695 99.875 ;
        RECT 43.625 98.265 48.970 98.700 ;
        RECT 49.145 98.265 54.490 98.700 ;
        RECT 54.665 98.265 60.010 98.700 ;
        RECT 60.185 98.265 63.695 99.355 ;
        RECT 64.345 99.320 64.520 100.125 ;
        RECT 65.510 99.955 65.680 100.290 ;
        RECT 66.165 100.245 66.405 100.620 ;
        RECT 66.575 100.310 66.910 100.815 ;
        RECT 66.165 100.095 66.385 100.245 ;
        RECT 64.695 99.595 65.680 99.955 ;
        RECT 65.850 99.765 66.385 100.095 ;
        RECT 64.695 99.575 65.980 99.595 ;
        RECT 65.120 99.425 65.980 99.575 ;
        RECT 64.345 98.535 64.650 99.320 ;
        RECT 64.825 98.945 65.520 99.255 ;
        RECT 64.830 98.265 65.515 98.735 ;
        RECT 65.695 98.480 65.980 99.425 ;
        RECT 66.150 99.115 66.385 99.765 ;
        RECT 66.555 99.285 66.855 100.135 ;
        RECT 67.085 100.045 68.755 100.815 ;
        RECT 68.925 100.090 69.215 100.815 ;
        RECT 69.385 100.270 74.730 100.815 ;
        RECT 74.905 100.270 80.250 100.815 ;
        RECT 80.425 100.270 85.770 100.815 ;
        RECT 85.945 100.270 91.290 100.815 ;
        RECT 67.085 99.525 67.835 100.045 ;
        RECT 68.005 99.355 68.755 99.875 ;
        RECT 70.970 99.440 71.310 100.270 ;
        RECT 66.150 98.885 66.825 99.115 ;
        RECT 66.155 98.265 66.485 98.715 ;
        RECT 66.655 98.455 66.825 98.885 ;
        RECT 67.085 98.265 68.755 99.355 ;
        RECT 68.925 98.265 69.215 99.430 ;
        RECT 72.790 98.700 73.140 99.950 ;
        RECT 76.490 99.440 76.830 100.270 ;
        RECT 78.310 98.700 78.660 99.950 ;
        RECT 82.010 99.440 82.350 100.270 ;
        RECT 83.830 98.700 84.180 99.950 ;
        RECT 87.530 99.440 87.870 100.270 ;
        RECT 91.465 100.045 94.055 100.815 ;
        RECT 94.685 100.090 94.975 100.815 ;
        RECT 95.145 100.270 100.490 100.815 ;
        RECT 100.665 100.270 106.010 100.815 ;
        RECT 107.110 100.310 107.445 100.815 ;
        RECT 89.350 98.700 89.700 99.950 ;
        RECT 91.465 99.525 92.675 100.045 ;
        RECT 92.845 99.355 94.055 99.875 ;
        RECT 96.730 99.440 97.070 100.270 ;
        RECT 69.385 98.265 74.730 98.700 ;
        RECT 74.905 98.265 80.250 98.700 ;
        RECT 80.425 98.265 85.770 98.700 ;
        RECT 85.945 98.265 91.290 98.700 ;
        RECT 91.465 98.265 94.055 99.355 ;
        RECT 94.685 98.265 94.975 99.430 ;
        RECT 98.550 98.700 98.900 99.950 ;
        RECT 102.250 99.440 102.590 100.270 ;
        RECT 107.615 100.245 107.855 100.620 ;
        RECT 108.135 100.485 108.305 100.630 ;
        RECT 108.135 100.290 108.510 100.485 ;
        RECT 108.870 100.320 109.265 100.815 ;
        RECT 104.070 98.700 104.420 99.950 ;
        RECT 107.165 99.285 107.465 100.135 ;
        RECT 107.635 100.095 107.855 100.245 ;
        RECT 107.635 99.765 108.170 100.095 ;
        RECT 108.340 99.955 108.510 100.290 ;
        RECT 109.435 100.125 109.675 100.645 ;
        RECT 109.865 100.270 115.210 100.815 ;
        RECT 116.310 100.310 116.645 100.815 ;
        RECT 107.635 99.115 107.870 99.765 ;
        RECT 108.340 99.595 109.325 99.955 ;
        RECT 107.195 98.885 107.870 99.115 ;
        RECT 108.040 99.575 109.325 99.595 ;
        RECT 108.040 99.425 108.900 99.575 ;
        RECT 95.145 98.265 100.490 98.700 ;
        RECT 100.665 98.265 106.010 98.700 ;
        RECT 107.195 98.455 107.365 98.885 ;
        RECT 107.535 98.265 107.865 98.715 ;
        RECT 108.040 98.480 108.325 99.425 ;
        RECT 109.500 99.320 109.675 100.125 ;
        RECT 111.450 99.440 111.790 100.270 ;
        RECT 116.815 100.245 117.055 100.620 ;
        RECT 117.335 100.485 117.505 100.630 ;
        RECT 117.335 100.290 117.710 100.485 ;
        RECT 118.070 100.320 118.465 100.815 ;
        RECT 108.500 98.945 109.195 99.255 ;
        RECT 108.505 98.265 109.190 98.735 ;
        RECT 109.370 98.535 109.675 99.320 ;
        RECT 113.270 98.700 113.620 99.950 ;
        RECT 116.365 99.285 116.665 100.135 ;
        RECT 116.835 100.095 117.055 100.245 ;
        RECT 116.835 99.765 117.370 100.095 ;
        RECT 117.540 99.955 117.710 100.290 ;
        RECT 118.635 100.125 118.875 100.645 ;
        RECT 116.835 99.115 117.070 99.765 ;
        RECT 117.540 99.595 118.525 99.955 ;
        RECT 116.395 98.885 117.070 99.115 ;
        RECT 117.240 99.575 118.525 99.595 ;
        RECT 117.240 99.425 118.100 99.575 ;
        RECT 109.865 98.265 115.210 98.700 ;
        RECT 116.395 98.455 116.565 98.885 ;
        RECT 116.735 98.265 117.065 98.715 ;
        RECT 117.240 98.480 117.525 99.425 ;
        RECT 118.700 99.320 118.875 100.125 ;
        RECT 119.065 100.065 120.275 100.815 ;
        RECT 120.445 100.090 120.735 100.815 ;
        RECT 120.905 100.270 126.250 100.815 ;
        RECT 126.425 100.270 131.770 100.815 ;
        RECT 119.065 99.525 119.585 100.065 ;
        RECT 119.755 99.355 120.275 99.895 ;
        RECT 122.490 99.440 122.830 100.270 ;
        RECT 117.700 98.945 118.395 99.255 ;
        RECT 117.705 98.265 118.390 98.735 ;
        RECT 118.570 98.535 118.875 99.320 ;
        RECT 119.065 98.265 120.275 99.355 ;
        RECT 120.445 98.265 120.735 99.430 ;
        RECT 124.310 98.700 124.660 99.950 ;
        RECT 128.010 99.440 128.350 100.270 ;
        RECT 131.945 100.045 133.615 100.815 ;
        RECT 133.790 100.310 134.125 100.815 ;
        RECT 134.295 100.245 134.535 100.620 ;
        RECT 134.815 100.485 134.985 100.630 ;
        RECT 134.815 100.290 135.190 100.485 ;
        RECT 135.550 100.320 135.945 100.815 ;
        RECT 129.830 98.700 130.180 99.950 ;
        RECT 131.945 99.525 132.695 100.045 ;
        RECT 132.865 99.355 133.615 99.875 ;
        RECT 120.905 98.265 126.250 98.700 ;
        RECT 126.425 98.265 131.770 98.700 ;
        RECT 131.945 98.265 133.615 99.355 ;
        RECT 133.845 99.285 134.145 100.135 ;
        RECT 134.315 100.095 134.535 100.245 ;
        RECT 134.315 99.765 134.850 100.095 ;
        RECT 135.020 99.955 135.190 100.290 ;
        RECT 136.115 100.125 136.355 100.645 ;
        RECT 134.315 99.115 134.550 99.765 ;
        RECT 135.020 99.595 136.005 99.955 ;
        RECT 133.875 98.885 134.550 99.115 ;
        RECT 134.720 99.575 136.005 99.595 ;
        RECT 134.720 99.425 135.580 99.575 ;
        RECT 133.875 98.455 134.045 98.885 ;
        RECT 134.215 98.265 134.545 98.715 ;
        RECT 134.720 98.480 135.005 99.425 ;
        RECT 136.180 99.320 136.355 100.125 ;
        RECT 136.635 100.265 136.805 100.555 ;
        RECT 136.975 100.435 137.305 100.815 ;
        RECT 136.635 100.095 137.300 100.265 ;
        RECT 135.180 98.945 135.875 99.255 ;
        RECT 135.185 98.265 135.870 98.735 ;
        RECT 136.050 98.535 136.355 99.320 ;
        RECT 136.550 99.275 136.900 99.925 ;
        RECT 137.070 99.105 137.300 100.095 ;
        RECT 136.635 98.935 137.300 99.105 ;
        RECT 136.635 98.435 136.805 98.935 ;
        RECT 136.975 98.265 137.305 98.765 ;
        RECT 137.475 98.435 137.660 100.555 ;
        RECT 137.915 100.355 138.165 100.815 ;
        RECT 138.335 100.365 138.670 100.535 ;
        RECT 138.865 100.365 139.540 100.535 ;
        RECT 138.335 100.225 138.505 100.365 ;
        RECT 137.830 99.235 138.110 100.185 ;
        RECT 138.280 100.095 138.505 100.225 ;
        RECT 138.280 98.990 138.450 100.095 ;
        RECT 138.675 99.945 139.200 100.165 ;
        RECT 138.620 99.180 138.860 99.775 ;
        RECT 139.030 99.245 139.200 99.945 ;
        RECT 139.370 99.585 139.540 100.365 ;
        RECT 139.860 100.315 140.230 100.815 ;
        RECT 140.410 100.365 140.815 100.535 ;
        RECT 140.985 100.365 141.770 100.535 ;
        RECT 140.410 100.135 140.580 100.365 ;
        RECT 139.750 99.835 140.580 100.135 ;
        RECT 140.965 99.865 141.430 100.195 ;
        RECT 139.750 99.805 139.950 99.835 ;
        RECT 140.070 99.585 140.240 99.655 ;
        RECT 139.370 99.415 140.240 99.585 ;
        RECT 139.730 99.325 140.240 99.415 ;
        RECT 138.280 98.860 138.585 98.990 ;
        RECT 139.030 98.880 139.560 99.245 ;
        RECT 137.900 98.265 138.165 98.725 ;
        RECT 138.335 98.435 138.585 98.860 ;
        RECT 139.730 98.710 139.900 99.325 ;
        RECT 138.795 98.540 139.900 98.710 ;
        RECT 140.070 98.265 140.240 99.065 ;
        RECT 140.410 98.765 140.580 99.835 ;
        RECT 140.750 98.935 140.940 99.655 ;
        RECT 141.110 98.905 141.430 99.865 ;
        RECT 141.600 99.905 141.770 100.365 ;
        RECT 142.045 100.285 142.255 100.815 ;
        RECT 142.515 100.075 142.845 100.600 ;
        RECT 143.015 100.205 143.185 100.815 ;
        RECT 143.355 100.160 143.685 100.595 ;
        RECT 143.995 100.265 144.165 100.645 ;
        RECT 144.380 100.435 144.710 100.815 ;
        RECT 143.355 100.075 143.735 100.160 ;
        RECT 143.995 100.095 144.710 100.265 ;
        RECT 142.645 99.905 142.845 100.075 ;
        RECT 143.510 100.035 143.735 100.075 ;
        RECT 141.600 99.575 142.475 99.905 ;
        RECT 142.645 99.575 143.395 99.905 ;
        RECT 140.410 98.435 140.660 98.765 ;
        RECT 141.600 98.735 141.770 99.575 ;
        RECT 142.645 99.370 142.835 99.575 ;
        RECT 143.565 99.455 143.735 100.035 ;
        RECT 143.905 99.545 144.260 99.915 ;
        RECT 144.540 99.905 144.710 100.095 ;
        RECT 144.880 100.070 145.135 100.645 ;
        RECT 144.540 99.575 144.795 99.905 ;
        RECT 143.520 99.405 143.735 99.455 ;
        RECT 141.940 98.995 142.835 99.370 ;
        RECT 143.345 99.325 143.735 99.405 ;
        RECT 144.540 99.365 144.710 99.575 ;
        RECT 140.885 98.565 141.770 98.735 ;
        RECT 141.950 98.265 142.265 98.765 ;
        RECT 142.495 98.435 142.835 98.995 ;
        RECT 143.005 98.265 143.175 99.275 ;
        RECT 143.345 98.480 143.675 99.325 ;
        RECT 143.995 99.195 144.710 99.365 ;
        RECT 144.965 99.340 145.135 100.070 ;
        RECT 145.310 99.975 145.570 100.815 ;
        RECT 145.745 100.065 146.955 100.815 ;
        RECT 143.995 98.435 144.165 99.195 ;
        RECT 144.380 98.265 144.710 99.025 ;
        RECT 144.880 98.435 145.135 99.340 ;
        RECT 145.310 98.265 145.570 99.415 ;
        RECT 145.745 99.355 146.265 99.895 ;
        RECT 146.435 99.525 146.955 100.065 ;
        RECT 145.745 98.265 146.955 99.355 ;
        RECT 17.320 98.095 147.040 98.265 ;
        RECT 17.405 97.005 18.615 98.095 ;
        RECT 19.305 97.035 19.635 97.880 ;
        RECT 19.805 97.085 19.975 98.095 ;
        RECT 20.145 97.365 20.485 97.925 ;
        RECT 20.715 97.595 21.030 98.095 ;
        RECT 21.210 97.625 22.095 97.795 ;
        RECT 17.405 96.295 17.925 96.835 ;
        RECT 18.095 96.465 18.615 97.005 ;
        RECT 19.245 96.955 19.635 97.035 ;
        RECT 20.145 96.990 21.040 97.365 ;
        RECT 19.245 96.905 19.460 96.955 ;
        RECT 19.245 96.325 19.415 96.905 ;
        RECT 20.145 96.785 20.335 96.990 ;
        RECT 21.210 96.785 21.380 97.625 ;
        RECT 22.320 97.595 22.570 97.925 ;
        RECT 19.585 96.455 20.335 96.785 ;
        RECT 20.505 96.455 21.380 96.785 ;
        RECT 17.405 95.545 18.615 96.295 ;
        RECT 19.245 96.285 19.470 96.325 ;
        RECT 20.135 96.285 20.335 96.455 ;
        RECT 19.245 96.200 19.625 96.285 ;
        RECT 19.295 95.765 19.625 96.200 ;
        RECT 19.795 95.545 19.965 96.155 ;
        RECT 20.135 95.760 20.465 96.285 ;
        RECT 20.725 95.545 20.935 96.075 ;
        RECT 21.210 95.995 21.380 96.455 ;
        RECT 21.550 96.495 21.870 97.455 ;
        RECT 22.040 96.705 22.230 97.425 ;
        RECT 22.400 96.525 22.570 97.595 ;
        RECT 22.740 97.295 22.910 98.095 ;
        RECT 23.080 97.650 24.185 97.820 ;
        RECT 23.080 97.035 23.250 97.650 ;
        RECT 24.395 97.500 24.645 97.925 ;
        RECT 24.815 97.635 25.080 98.095 ;
        RECT 23.420 97.115 23.950 97.480 ;
        RECT 24.395 97.370 24.700 97.500 ;
        RECT 22.740 96.945 23.250 97.035 ;
        RECT 22.740 96.775 23.610 96.945 ;
        RECT 22.740 96.705 22.910 96.775 ;
        RECT 23.030 96.525 23.230 96.555 ;
        RECT 21.550 96.165 22.015 96.495 ;
        RECT 22.400 96.225 23.230 96.525 ;
        RECT 22.400 95.995 22.570 96.225 ;
        RECT 21.210 95.825 21.995 95.995 ;
        RECT 22.165 95.825 22.570 95.995 ;
        RECT 22.750 95.545 23.120 96.045 ;
        RECT 23.440 95.995 23.610 96.775 ;
        RECT 23.780 96.415 23.950 97.115 ;
        RECT 24.120 96.585 24.360 97.180 ;
        RECT 23.780 96.195 24.305 96.415 ;
        RECT 24.530 96.265 24.700 97.370 ;
        RECT 24.475 96.135 24.700 96.265 ;
        RECT 24.870 96.175 25.150 97.125 ;
        RECT 24.475 95.995 24.645 96.135 ;
        RECT 23.440 95.825 24.115 95.995 ;
        RECT 24.310 95.825 24.645 95.995 ;
        RECT 24.815 95.545 25.065 96.005 ;
        RECT 25.320 95.805 25.505 97.925 ;
        RECT 25.675 97.595 26.005 98.095 ;
        RECT 26.175 97.425 26.345 97.925 ;
        RECT 25.680 97.255 26.345 97.425 ;
        RECT 25.680 96.265 25.910 97.255 ;
        RECT 26.080 96.435 26.430 97.085 ;
        RECT 26.605 97.005 27.815 98.095 ;
        RECT 26.605 96.295 27.125 96.835 ;
        RECT 27.295 96.465 27.815 97.005 ;
        RECT 27.990 96.955 28.265 97.925 ;
        RECT 28.475 97.295 28.755 98.095 ;
        RECT 28.925 97.585 30.115 97.875 ;
        RECT 28.925 97.245 30.095 97.415 ;
        RECT 28.925 97.125 29.095 97.245 ;
        RECT 28.435 96.955 29.095 97.125 ;
        RECT 25.680 96.095 26.345 96.265 ;
        RECT 25.675 95.545 26.005 95.925 ;
        RECT 26.175 95.805 26.345 96.095 ;
        RECT 26.605 95.545 27.815 96.295 ;
        RECT 27.990 96.220 28.160 96.955 ;
        RECT 28.435 96.785 28.605 96.955 ;
        RECT 29.405 96.785 29.600 97.075 ;
        RECT 29.770 96.955 30.095 97.245 ;
        RECT 30.285 96.930 30.575 98.095 ;
        RECT 30.745 96.940 31.085 97.925 ;
        RECT 31.255 97.665 31.665 98.095 ;
        RECT 32.410 97.675 32.740 98.095 ;
        RECT 32.910 97.495 33.235 97.925 ;
        RECT 31.255 97.325 33.235 97.495 ;
        RECT 28.330 96.455 28.605 96.785 ;
        RECT 28.775 96.455 29.600 96.785 ;
        RECT 29.770 96.455 30.115 96.785 ;
        RECT 28.435 96.285 28.605 96.455 ;
        RECT 30.745 96.285 31.000 96.940 ;
        RECT 31.255 96.785 31.520 97.325 ;
        RECT 31.735 96.985 32.360 97.155 ;
        RECT 31.170 96.455 31.520 96.785 ;
        RECT 31.690 96.455 32.020 96.785 ;
        RECT 32.190 96.285 32.360 96.985 ;
        RECT 27.990 95.875 28.265 96.220 ;
        RECT 28.435 96.115 30.100 96.285 ;
        RECT 28.455 95.545 28.835 95.945 ;
        RECT 29.005 95.765 29.175 96.115 ;
        RECT 29.345 95.545 29.675 95.945 ;
        RECT 29.845 95.765 30.100 96.115 ;
        RECT 30.285 95.545 30.575 96.270 ;
        RECT 30.745 95.910 31.105 96.285 ;
        RECT 31.370 95.545 31.540 96.285 ;
        RECT 31.820 96.115 32.360 96.285 ;
        RECT 32.530 96.915 33.235 97.325 ;
        RECT 33.710 96.995 34.040 98.095 ;
        RECT 34.430 97.585 36.085 97.875 ;
        RECT 34.430 97.245 36.020 97.415 ;
        RECT 36.255 97.295 36.535 98.095 ;
        RECT 34.430 96.955 34.750 97.245 ;
        RECT 35.850 97.125 36.020 97.245 ;
        RECT 31.820 95.910 31.990 96.115 ;
        RECT 32.530 95.715 32.700 96.915 ;
        RECT 34.945 96.905 35.660 97.075 ;
        RECT 35.850 96.955 36.575 97.125 ;
        RECT 36.745 96.955 37.015 97.925 ;
        RECT 37.185 97.660 42.530 98.095 ;
        RECT 42.705 97.660 48.050 98.095 ;
        RECT 48.225 97.660 53.570 98.095 ;
        RECT 32.870 96.535 33.440 96.745 ;
        RECT 33.610 96.535 34.255 96.745 ;
        RECT 32.930 96.195 34.100 96.365 ;
        RECT 34.430 96.215 34.780 96.785 ;
        RECT 34.950 96.455 35.660 96.905 ;
        RECT 36.405 96.785 36.575 96.955 ;
        RECT 35.830 96.455 36.235 96.785 ;
        RECT 36.405 96.455 36.675 96.785 ;
        RECT 36.405 96.285 36.575 96.455 ;
        RECT 32.930 95.715 33.260 96.195 ;
        RECT 33.430 95.545 33.600 96.015 ;
        RECT 33.770 95.730 34.100 96.195 ;
        RECT 34.965 96.115 36.575 96.285 ;
        RECT 36.845 96.220 37.015 96.955 ;
        RECT 34.435 95.545 34.765 96.045 ;
        RECT 34.965 95.765 35.135 96.115 ;
        RECT 35.335 95.545 35.665 95.945 ;
        RECT 35.835 95.765 36.005 96.115 ;
        RECT 36.175 95.545 36.555 95.945 ;
        RECT 36.745 95.875 37.015 96.220 ;
        RECT 38.770 96.090 39.110 96.920 ;
        RECT 40.590 96.410 40.940 97.660 ;
        RECT 44.290 96.090 44.630 96.920 ;
        RECT 46.110 96.410 46.460 97.660 ;
        RECT 49.810 96.090 50.150 96.920 ;
        RECT 51.630 96.410 51.980 97.660 ;
        RECT 53.745 97.005 55.415 98.095 ;
        RECT 53.745 96.315 54.495 96.835 ;
        RECT 54.665 96.485 55.415 97.005 ;
        RECT 56.045 96.930 56.335 98.095 ;
        RECT 56.505 97.660 61.850 98.095 ;
        RECT 37.185 95.545 42.530 96.090 ;
        RECT 42.705 95.545 48.050 96.090 ;
        RECT 48.225 95.545 53.570 96.090 ;
        RECT 53.745 95.545 55.415 96.315 ;
        RECT 56.045 95.545 56.335 96.270 ;
        RECT 58.090 96.090 58.430 96.920 ;
        RECT 59.910 96.410 60.260 97.660 ;
        RECT 62.115 97.475 62.285 97.905 ;
        RECT 62.455 97.645 62.785 98.095 ;
        RECT 62.115 97.245 62.790 97.475 ;
        RECT 62.085 96.225 62.385 97.075 ;
        RECT 62.555 96.595 62.790 97.245 ;
        RECT 62.960 96.935 63.245 97.880 ;
        RECT 63.425 97.625 64.110 98.095 ;
        RECT 63.420 97.105 64.115 97.415 ;
        RECT 64.290 97.040 64.595 97.825 ;
        RECT 62.960 96.785 63.820 96.935 ;
        RECT 62.960 96.765 64.245 96.785 ;
        RECT 62.555 96.265 63.090 96.595 ;
        RECT 63.260 96.405 64.245 96.765 ;
        RECT 62.555 96.115 62.775 96.265 ;
        RECT 56.505 95.545 61.850 96.090 ;
        RECT 62.030 95.545 62.365 96.050 ;
        RECT 62.535 95.740 62.775 96.115 ;
        RECT 63.260 96.070 63.430 96.405 ;
        RECT 64.420 96.235 64.595 97.040 ;
        RECT 64.785 97.005 67.375 98.095 ;
        RECT 63.055 95.875 63.430 96.070 ;
        RECT 63.055 95.730 63.225 95.875 ;
        RECT 63.790 95.545 64.185 96.040 ;
        RECT 64.355 95.715 64.595 96.235 ;
        RECT 64.785 96.315 65.995 96.835 ;
        RECT 66.165 96.485 67.375 97.005 ;
        RECT 67.550 96.955 67.885 97.925 ;
        RECT 68.055 96.955 68.225 98.095 ;
        RECT 68.395 97.755 70.425 97.925 ;
        RECT 64.785 95.545 67.375 96.315 ;
        RECT 67.550 96.285 67.720 96.955 ;
        RECT 68.395 96.785 68.565 97.755 ;
        RECT 67.890 96.455 68.145 96.785 ;
        RECT 68.370 96.455 68.565 96.785 ;
        RECT 68.735 97.415 69.860 97.585 ;
        RECT 67.975 96.285 68.145 96.455 ;
        RECT 68.735 96.285 68.905 97.415 ;
        RECT 67.550 95.715 67.805 96.285 ;
        RECT 67.975 96.115 68.905 96.285 ;
        RECT 69.075 97.075 70.085 97.245 ;
        RECT 69.075 96.275 69.245 97.075 ;
        RECT 69.450 96.395 69.725 96.875 ;
        RECT 69.445 96.225 69.725 96.395 ;
        RECT 68.730 96.080 68.905 96.115 ;
        RECT 67.975 95.545 68.305 95.945 ;
        RECT 68.730 95.715 69.260 96.080 ;
        RECT 69.450 95.715 69.725 96.225 ;
        RECT 69.895 95.715 70.085 97.075 ;
        RECT 70.255 97.090 70.425 97.755 ;
        RECT 70.595 97.335 70.765 98.095 ;
        RECT 71.000 97.335 71.515 97.745 ;
        RECT 70.255 96.900 71.005 97.090 ;
        RECT 71.175 96.525 71.515 97.335 ;
        RECT 71.690 97.705 72.025 97.925 ;
        RECT 73.030 97.715 73.385 98.095 ;
        RECT 71.690 97.085 71.945 97.705 ;
        RECT 72.195 97.545 72.425 97.585 ;
        RECT 73.555 97.545 73.805 97.925 ;
        RECT 72.195 97.345 73.805 97.545 ;
        RECT 72.195 97.255 72.380 97.345 ;
        RECT 72.970 97.335 73.805 97.345 ;
        RECT 74.055 97.315 74.305 98.095 ;
        RECT 74.475 97.245 74.735 97.925 ;
        RECT 72.535 97.145 72.865 97.175 ;
        RECT 72.535 97.085 74.335 97.145 ;
        RECT 71.690 96.975 74.395 97.085 ;
        RECT 71.690 96.915 72.865 96.975 ;
        RECT 74.195 96.940 74.395 96.975 ;
        RECT 71.685 96.535 72.175 96.735 ;
        RECT 72.365 96.535 72.840 96.745 ;
        RECT 70.285 96.355 71.515 96.525 ;
        RECT 70.265 95.545 70.775 96.080 ;
        RECT 70.995 95.750 71.240 96.355 ;
        RECT 71.690 95.545 72.145 96.310 ;
        RECT 72.620 96.135 72.840 96.535 ;
        RECT 73.085 96.535 73.415 96.745 ;
        RECT 73.085 96.135 73.295 96.535 ;
        RECT 73.585 96.500 73.995 96.805 ;
        RECT 74.225 96.365 74.395 96.940 ;
        RECT 74.125 96.245 74.395 96.365 ;
        RECT 73.550 96.200 74.395 96.245 ;
        RECT 73.550 96.075 74.305 96.200 ;
        RECT 73.550 95.925 73.720 96.075 ;
        RECT 74.565 96.045 74.735 97.245 ;
        RECT 74.905 97.005 78.415 98.095 ;
        RECT 79.135 97.475 79.305 97.905 ;
        RECT 79.475 97.645 79.805 98.095 ;
        RECT 79.135 97.245 79.810 97.475 ;
        RECT 72.420 95.715 73.720 95.925 ;
        RECT 73.975 95.545 74.305 95.905 ;
        RECT 74.475 95.715 74.735 96.045 ;
        RECT 74.905 96.315 76.555 96.835 ;
        RECT 76.725 96.485 78.415 97.005 ;
        RECT 74.905 95.545 78.415 96.315 ;
        RECT 79.105 96.225 79.405 97.075 ;
        RECT 79.575 96.595 79.810 97.245 ;
        RECT 79.980 96.935 80.265 97.880 ;
        RECT 80.445 97.625 81.130 98.095 ;
        RECT 80.440 97.105 81.135 97.415 ;
        RECT 81.310 97.040 81.615 97.825 ;
        RECT 79.980 96.785 80.840 96.935 ;
        RECT 79.980 96.765 81.265 96.785 ;
        RECT 79.575 96.265 80.110 96.595 ;
        RECT 80.280 96.405 81.265 96.765 ;
        RECT 79.575 96.115 79.795 96.265 ;
        RECT 79.050 95.545 79.385 96.050 ;
        RECT 79.555 95.740 79.795 96.115 ;
        RECT 80.280 96.070 80.450 96.405 ;
        RECT 81.440 96.235 81.615 97.040 ;
        RECT 81.805 96.930 82.095 98.095 ;
        RECT 82.265 97.005 83.935 98.095 ;
        RECT 82.265 96.315 83.015 96.835 ;
        RECT 83.185 96.485 83.935 97.005 ;
        RECT 84.110 96.955 84.445 97.925 ;
        RECT 84.615 96.955 84.785 98.095 ;
        RECT 84.955 97.755 86.985 97.925 ;
        RECT 80.075 95.875 80.450 96.070 ;
        RECT 80.075 95.730 80.245 95.875 ;
        RECT 80.810 95.545 81.205 96.040 ;
        RECT 81.375 95.715 81.615 96.235 ;
        RECT 81.805 95.545 82.095 96.270 ;
        RECT 82.265 95.545 83.935 96.315 ;
        RECT 84.110 96.285 84.280 96.955 ;
        RECT 84.955 96.785 85.125 97.755 ;
        RECT 84.450 96.455 84.705 96.785 ;
        RECT 84.930 96.455 85.125 96.785 ;
        RECT 85.295 97.415 86.420 97.585 ;
        RECT 84.535 96.285 84.705 96.455 ;
        RECT 85.295 96.285 85.465 97.415 ;
        RECT 84.110 95.715 84.365 96.285 ;
        RECT 84.535 96.115 85.465 96.285 ;
        RECT 85.635 97.075 86.645 97.245 ;
        RECT 85.635 96.275 85.805 97.075 ;
        RECT 85.290 96.080 85.465 96.115 ;
        RECT 84.535 95.545 84.865 95.945 ;
        RECT 85.290 95.715 85.820 96.080 ;
        RECT 86.010 96.055 86.285 96.875 ;
        RECT 86.005 95.885 86.285 96.055 ;
        RECT 86.010 95.715 86.285 95.885 ;
        RECT 86.455 95.715 86.645 97.075 ;
        RECT 86.815 97.090 86.985 97.755 ;
        RECT 87.155 97.335 87.325 98.095 ;
        RECT 87.560 97.335 88.075 97.745 ;
        RECT 86.815 96.900 87.565 97.090 ;
        RECT 87.735 96.525 88.075 97.335 ;
        RECT 88.245 97.005 89.915 98.095 ;
        RECT 86.845 96.355 88.075 96.525 ;
        RECT 86.825 95.545 87.335 96.080 ;
        RECT 87.555 95.750 87.800 96.355 ;
        RECT 88.245 96.315 88.995 96.835 ;
        RECT 89.165 96.485 89.915 97.005 ;
        RECT 90.635 97.085 90.805 97.925 ;
        RECT 90.975 97.755 92.145 97.925 ;
        RECT 90.975 97.255 91.305 97.755 ;
        RECT 91.815 97.715 92.145 97.755 ;
        RECT 92.335 97.675 92.690 98.095 ;
        RECT 91.475 97.495 91.705 97.585 ;
        RECT 92.860 97.495 93.110 97.925 ;
        RECT 91.475 97.255 93.110 97.495 ;
        RECT 93.280 97.335 93.610 98.095 ;
        RECT 93.780 97.255 94.035 97.925 ;
        RECT 90.635 96.915 93.695 97.085 ;
        RECT 90.550 96.535 90.900 96.745 ;
        RECT 91.070 96.535 91.515 96.735 ;
        RECT 91.685 96.535 92.160 96.735 ;
        RECT 88.245 95.545 89.915 96.315 ;
        RECT 90.635 96.195 91.700 96.365 ;
        RECT 90.635 95.715 90.805 96.195 ;
        RECT 90.975 95.545 91.305 96.025 ;
        RECT 91.530 95.965 91.700 96.195 ;
        RECT 91.880 96.135 92.160 96.535 ;
        RECT 92.430 96.535 92.760 96.735 ;
        RECT 92.930 96.535 93.295 96.735 ;
        RECT 92.430 96.135 92.715 96.535 ;
        RECT 93.525 96.365 93.695 96.915 ;
        RECT 92.895 96.195 93.695 96.365 ;
        RECT 92.895 95.965 93.065 96.195 ;
        RECT 93.865 96.125 94.035 97.255 ;
        RECT 94.225 97.005 95.435 98.095 ;
        RECT 93.850 96.055 94.035 96.125 ;
        RECT 93.825 96.045 94.035 96.055 ;
        RECT 91.530 95.715 93.065 95.965 ;
        RECT 93.235 95.545 93.565 96.025 ;
        RECT 93.780 95.715 94.035 96.045 ;
        RECT 94.225 96.295 94.745 96.835 ;
        RECT 94.915 96.465 95.435 97.005 ;
        RECT 95.605 97.125 95.875 97.895 ;
        RECT 96.045 97.315 96.375 98.095 ;
        RECT 96.580 97.490 96.765 97.895 ;
        RECT 96.935 97.670 97.270 98.095 ;
        RECT 96.580 97.315 97.245 97.490 ;
        RECT 95.605 96.955 96.735 97.125 ;
        RECT 94.225 95.545 95.435 96.295 ;
        RECT 95.605 96.045 95.775 96.955 ;
        RECT 95.945 96.205 96.305 96.785 ;
        RECT 96.485 96.455 96.735 96.955 ;
        RECT 96.905 96.285 97.245 97.315 ;
        RECT 96.560 96.115 97.245 96.285 ;
        RECT 97.445 96.955 97.705 97.925 ;
        RECT 97.875 97.670 98.260 98.095 ;
        RECT 98.430 97.500 98.685 97.925 ;
        RECT 97.875 97.305 98.685 97.500 ;
        RECT 97.445 96.285 97.630 96.955 ;
        RECT 97.875 96.785 98.225 97.305 ;
        RECT 98.875 97.135 99.120 97.925 ;
        RECT 99.290 97.670 99.675 98.095 ;
        RECT 99.845 97.500 100.120 97.925 ;
        RECT 97.800 96.455 98.225 96.785 ;
        RECT 98.395 96.955 99.120 97.135 ;
        RECT 99.290 97.305 100.120 97.500 ;
        RECT 98.395 96.455 99.045 96.955 ;
        RECT 99.290 96.785 99.640 97.305 ;
        RECT 100.290 97.135 100.715 97.925 ;
        RECT 100.885 97.670 101.270 98.095 ;
        RECT 101.440 97.500 101.875 97.925 ;
        RECT 99.215 96.455 99.640 96.785 ;
        RECT 99.810 96.955 100.715 97.135 ;
        RECT 100.885 97.330 101.875 97.500 ;
        RECT 99.810 96.455 100.640 96.955 ;
        RECT 100.885 96.785 101.220 97.330 ;
        RECT 100.810 96.455 101.220 96.785 ;
        RECT 101.390 96.455 101.875 97.160 ;
        RECT 102.050 96.955 102.385 97.925 ;
        RECT 102.555 96.955 102.725 98.095 ;
        RECT 102.895 97.755 104.925 97.925 ;
        RECT 97.875 96.285 98.225 96.455 ;
        RECT 98.875 96.285 99.045 96.455 ;
        RECT 99.290 96.285 99.640 96.455 ;
        RECT 100.290 96.285 100.640 96.455 ;
        RECT 100.885 96.285 101.220 96.455 ;
        RECT 102.050 96.285 102.220 96.955 ;
        RECT 102.895 96.785 103.065 97.755 ;
        RECT 102.390 96.455 102.645 96.785 ;
        RECT 102.870 96.455 103.065 96.785 ;
        RECT 103.235 97.415 104.360 97.585 ;
        RECT 102.475 96.285 102.645 96.455 ;
        RECT 103.235 96.285 103.405 97.415 ;
        RECT 95.605 95.715 95.865 96.045 ;
        RECT 96.075 95.545 96.350 96.025 ;
        RECT 96.560 95.715 96.765 96.115 ;
        RECT 96.935 95.545 97.270 95.945 ;
        RECT 97.445 95.715 97.705 96.285 ;
        RECT 97.875 96.115 98.685 96.285 ;
        RECT 97.875 95.545 98.260 95.945 ;
        RECT 98.430 95.715 98.685 96.115 ;
        RECT 98.875 95.715 99.120 96.285 ;
        RECT 99.290 96.115 100.100 96.285 ;
        RECT 99.290 95.545 99.675 95.945 ;
        RECT 99.845 95.715 100.100 96.115 ;
        RECT 100.290 95.715 100.715 96.285 ;
        RECT 100.885 96.115 101.875 96.285 ;
        RECT 100.885 95.545 101.270 95.945 ;
        RECT 101.440 95.715 101.875 96.115 ;
        RECT 102.050 95.715 102.305 96.285 ;
        RECT 102.475 96.115 103.405 96.285 ;
        RECT 103.575 97.075 104.585 97.245 ;
        RECT 103.575 96.275 103.745 97.075 ;
        RECT 103.950 96.395 104.225 96.875 ;
        RECT 103.945 96.225 104.225 96.395 ;
        RECT 103.230 96.080 103.405 96.115 ;
        RECT 102.475 95.545 102.805 95.945 ;
        RECT 103.230 95.715 103.760 96.080 ;
        RECT 103.950 95.715 104.225 96.225 ;
        RECT 104.395 95.715 104.585 97.075 ;
        RECT 104.755 97.090 104.925 97.755 ;
        RECT 105.095 97.335 105.265 98.095 ;
        RECT 105.500 97.335 106.015 97.745 ;
        RECT 104.755 96.900 105.505 97.090 ;
        RECT 105.675 96.525 106.015 97.335 ;
        RECT 106.185 97.005 107.395 98.095 ;
        RECT 104.785 96.355 106.015 96.525 ;
        RECT 104.765 95.545 105.275 96.080 ;
        RECT 105.495 95.750 105.740 96.355 ;
        RECT 106.185 96.295 106.705 96.835 ;
        RECT 106.875 96.465 107.395 97.005 ;
        RECT 107.565 96.930 107.855 98.095 ;
        RECT 108.490 96.955 108.825 97.925 ;
        RECT 108.995 96.955 109.165 98.095 ;
        RECT 109.335 97.755 111.365 97.925 ;
        RECT 106.185 95.545 107.395 96.295 ;
        RECT 108.490 96.285 108.660 96.955 ;
        RECT 109.335 96.785 109.505 97.755 ;
        RECT 108.830 96.455 109.085 96.785 ;
        RECT 109.310 96.455 109.505 96.785 ;
        RECT 109.675 97.415 110.800 97.585 ;
        RECT 108.915 96.285 109.085 96.455 ;
        RECT 109.675 96.285 109.845 97.415 ;
        RECT 107.565 95.545 107.855 96.270 ;
        RECT 108.490 95.715 108.745 96.285 ;
        RECT 108.915 96.115 109.845 96.285 ;
        RECT 110.015 97.075 111.025 97.245 ;
        RECT 110.015 96.275 110.185 97.075 ;
        RECT 109.670 96.080 109.845 96.115 ;
        RECT 108.915 95.545 109.245 95.945 ;
        RECT 109.670 95.715 110.200 96.080 ;
        RECT 110.390 96.055 110.665 96.875 ;
        RECT 110.385 95.885 110.665 96.055 ;
        RECT 110.390 95.715 110.665 95.885 ;
        RECT 110.835 95.715 111.025 97.075 ;
        RECT 111.195 97.090 111.365 97.755 ;
        RECT 111.535 97.335 111.705 98.095 ;
        RECT 111.940 97.335 112.455 97.745 ;
        RECT 111.195 96.900 111.945 97.090 ;
        RECT 112.115 96.525 112.455 97.335 ;
        RECT 112.625 97.005 114.295 98.095 ;
        RECT 111.225 96.355 112.455 96.525 ;
        RECT 111.205 95.545 111.715 96.080 ;
        RECT 111.935 95.750 112.180 96.355 ;
        RECT 112.625 96.315 113.375 96.835 ;
        RECT 113.545 96.485 114.295 97.005 ;
        RECT 114.555 97.085 114.725 97.925 ;
        RECT 114.895 97.755 116.065 97.925 ;
        RECT 114.895 97.255 115.225 97.755 ;
        RECT 115.735 97.715 116.065 97.755 ;
        RECT 116.255 97.675 116.610 98.095 ;
        RECT 115.395 97.495 115.625 97.585 ;
        RECT 116.780 97.495 117.030 97.925 ;
        RECT 115.395 97.255 117.030 97.495 ;
        RECT 117.200 97.335 117.530 98.095 ;
        RECT 117.700 97.255 117.955 97.925 ;
        RECT 118.145 97.660 123.490 98.095 ;
        RECT 114.555 96.915 117.615 97.085 ;
        RECT 114.470 96.535 114.820 96.745 ;
        RECT 114.990 96.535 115.435 96.735 ;
        RECT 115.605 96.535 116.080 96.735 ;
        RECT 112.625 95.545 114.295 96.315 ;
        RECT 114.555 96.195 115.620 96.365 ;
        RECT 114.555 95.715 114.725 96.195 ;
        RECT 114.895 95.545 115.225 96.025 ;
        RECT 115.450 95.965 115.620 96.195 ;
        RECT 115.800 96.135 116.080 96.535 ;
        RECT 116.350 96.535 116.680 96.735 ;
        RECT 116.850 96.535 117.215 96.735 ;
        RECT 116.350 96.135 116.635 96.535 ;
        RECT 117.445 96.365 117.615 96.915 ;
        RECT 116.815 96.195 117.615 96.365 ;
        RECT 116.815 95.965 116.985 96.195 ;
        RECT 117.785 96.125 117.955 97.255 ;
        RECT 117.770 96.045 117.955 96.125 ;
        RECT 119.730 96.090 120.070 96.920 ;
        RECT 121.550 96.410 121.900 97.660 ;
        RECT 123.665 97.005 126.255 98.095 ;
        RECT 126.515 97.475 126.685 97.905 ;
        RECT 126.855 97.645 127.185 98.095 ;
        RECT 126.515 97.245 127.190 97.475 ;
        RECT 123.665 96.315 124.875 96.835 ;
        RECT 125.045 96.485 126.255 97.005 ;
        RECT 115.450 95.715 116.985 95.965 ;
        RECT 117.155 95.545 117.485 96.025 ;
        RECT 117.700 95.715 117.955 96.045 ;
        RECT 118.145 95.545 123.490 96.090 ;
        RECT 123.665 95.545 126.255 96.315 ;
        RECT 126.485 96.225 126.785 97.075 ;
        RECT 126.955 96.595 127.190 97.245 ;
        RECT 127.360 96.935 127.645 97.880 ;
        RECT 127.825 97.625 128.510 98.095 ;
        RECT 127.820 97.105 128.515 97.415 ;
        RECT 128.690 97.040 128.995 97.825 ;
        RECT 127.360 96.785 128.220 96.935 ;
        RECT 127.360 96.765 128.645 96.785 ;
        RECT 126.955 96.265 127.490 96.595 ;
        RECT 127.660 96.405 128.645 96.765 ;
        RECT 126.955 96.115 127.175 96.265 ;
        RECT 126.430 95.545 126.765 96.050 ;
        RECT 126.935 95.740 127.175 96.115 ;
        RECT 127.660 96.070 127.830 96.405 ;
        RECT 128.820 96.235 128.995 97.040 ;
        RECT 127.455 95.875 127.830 96.070 ;
        RECT 127.455 95.730 127.625 95.875 ;
        RECT 128.190 95.545 128.585 96.040 ;
        RECT 128.755 95.715 128.995 96.235 ;
        RECT 129.185 97.125 129.455 97.895 ;
        RECT 129.625 97.315 129.955 98.095 ;
        RECT 130.160 97.490 130.345 97.895 ;
        RECT 130.515 97.670 130.850 98.095 ;
        RECT 131.030 97.670 131.365 98.095 ;
        RECT 131.535 97.490 131.720 97.895 ;
        RECT 130.160 97.315 130.825 97.490 ;
        RECT 129.185 96.955 130.315 97.125 ;
        RECT 129.185 96.045 129.355 96.955 ;
        RECT 129.525 96.205 129.885 96.785 ;
        RECT 130.065 96.455 130.315 96.955 ;
        RECT 130.485 96.285 130.825 97.315 ;
        RECT 130.140 96.115 130.825 96.285 ;
        RECT 131.055 97.315 131.720 97.490 ;
        RECT 131.925 97.315 132.255 98.095 ;
        RECT 131.055 96.285 131.395 97.315 ;
        RECT 132.425 97.125 132.695 97.895 ;
        RECT 131.565 96.955 132.695 97.125 ;
        RECT 131.565 96.455 131.815 96.955 ;
        RECT 131.055 96.115 131.740 96.285 ;
        RECT 131.995 96.205 132.355 96.785 ;
        RECT 129.185 95.715 129.445 96.045 ;
        RECT 129.655 95.545 129.930 96.025 ;
        RECT 130.140 95.715 130.345 96.115 ;
        RECT 130.515 95.545 130.850 95.945 ;
        RECT 131.030 95.545 131.365 95.945 ;
        RECT 131.535 95.715 131.740 96.115 ;
        RECT 132.525 96.045 132.695 96.955 ;
        RECT 133.325 96.930 133.615 98.095 ;
        RECT 133.875 97.475 134.045 97.905 ;
        RECT 134.215 97.645 134.545 98.095 ;
        RECT 133.875 97.245 134.550 97.475 ;
        RECT 131.950 95.545 132.225 96.025 ;
        RECT 132.435 95.715 132.695 96.045 ;
        RECT 133.325 95.545 133.615 96.270 ;
        RECT 133.845 96.225 134.145 97.075 ;
        RECT 134.315 96.595 134.550 97.245 ;
        RECT 134.720 96.935 135.005 97.880 ;
        RECT 135.185 97.625 135.870 98.095 ;
        RECT 135.180 97.105 135.875 97.415 ;
        RECT 136.050 97.040 136.355 97.825 ;
        RECT 134.720 96.785 135.580 96.935 ;
        RECT 136.145 96.905 136.355 97.040 ;
        RECT 134.720 96.765 136.005 96.785 ;
        RECT 134.315 96.265 134.850 96.595 ;
        RECT 135.020 96.405 136.005 96.765 ;
        RECT 134.315 96.115 134.535 96.265 ;
        RECT 133.790 95.545 134.125 96.050 ;
        RECT 134.295 95.740 134.535 96.115 ;
        RECT 135.020 96.070 135.190 96.405 ;
        RECT 136.180 96.235 136.355 96.905 ;
        RECT 134.815 95.875 135.190 96.070 ;
        RECT 134.815 95.730 134.985 95.875 ;
        RECT 135.550 95.545 135.945 96.040 ;
        RECT 136.115 95.715 136.355 96.235 ;
        RECT 136.545 97.245 136.805 97.925 ;
        RECT 136.975 97.315 137.225 98.095 ;
        RECT 137.475 97.545 137.725 97.925 ;
        RECT 137.895 97.715 138.250 98.095 ;
        RECT 139.255 97.705 139.590 97.925 ;
        RECT 138.855 97.545 139.085 97.585 ;
        RECT 137.475 97.345 139.085 97.545 ;
        RECT 137.475 97.335 138.310 97.345 ;
        RECT 138.900 97.255 139.085 97.345 ;
        RECT 136.545 96.055 136.715 97.245 ;
        RECT 138.415 97.145 138.745 97.175 ;
        RECT 136.945 97.085 138.745 97.145 ;
        RECT 139.335 97.085 139.590 97.705 ;
        RECT 136.885 96.975 139.590 97.085 ;
        RECT 139.765 97.005 141.435 98.095 ;
        RECT 136.885 96.940 137.085 96.975 ;
        RECT 136.885 96.365 137.055 96.940 ;
        RECT 138.415 96.915 139.590 96.975 ;
        RECT 137.285 96.500 137.695 96.805 ;
        RECT 137.865 96.535 138.195 96.745 ;
        RECT 136.885 96.245 137.155 96.365 ;
        RECT 136.885 96.200 137.730 96.245 ;
        RECT 136.975 96.075 137.730 96.200 ;
        RECT 137.985 96.135 138.195 96.535 ;
        RECT 138.440 96.535 138.915 96.745 ;
        RECT 139.105 96.535 139.595 96.735 ;
        RECT 138.440 96.135 138.660 96.535 ;
        RECT 139.765 96.315 140.515 96.835 ;
        RECT 140.685 96.485 141.435 97.005 ;
        RECT 142.155 97.165 142.325 97.925 ;
        RECT 142.540 97.335 142.870 98.095 ;
        RECT 142.155 96.995 142.870 97.165 ;
        RECT 143.040 97.020 143.295 97.925 ;
        RECT 142.065 96.445 142.420 96.815 ;
        RECT 142.700 96.785 142.870 96.995 ;
        RECT 142.700 96.455 142.955 96.785 ;
        RECT 136.545 96.045 136.775 96.055 ;
        RECT 136.545 95.715 136.805 96.045 ;
        RECT 137.560 95.925 137.730 96.075 ;
        RECT 136.975 95.545 137.305 95.905 ;
        RECT 137.560 95.715 138.860 95.925 ;
        RECT 139.135 95.545 139.590 96.310 ;
        RECT 139.765 95.545 141.435 96.315 ;
        RECT 142.700 96.265 142.870 96.455 ;
        RECT 143.125 96.290 143.295 97.020 ;
        RECT 143.470 96.945 143.730 98.095 ;
        RECT 143.995 97.165 144.165 97.925 ;
        RECT 144.380 97.335 144.710 98.095 ;
        RECT 143.995 96.995 144.710 97.165 ;
        RECT 144.880 97.020 145.135 97.925 ;
        RECT 143.905 96.445 144.260 96.815 ;
        RECT 144.540 96.785 144.710 96.995 ;
        RECT 144.540 96.455 144.795 96.785 ;
        RECT 142.155 96.095 142.870 96.265 ;
        RECT 142.155 95.715 142.325 96.095 ;
        RECT 142.540 95.545 142.870 95.925 ;
        RECT 143.040 95.715 143.295 96.290 ;
        RECT 143.470 95.545 143.730 96.385 ;
        RECT 144.540 96.265 144.710 96.455 ;
        RECT 144.965 96.290 145.135 97.020 ;
        RECT 145.310 96.945 145.570 98.095 ;
        RECT 145.745 97.005 146.955 98.095 ;
        RECT 145.745 96.465 146.265 97.005 ;
        RECT 143.995 96.095 144.710 96.265 ;
        RECT 143.995 95.715 144.165 96.095 ;
        RECT 144.380 95.545 144.710 95.925 ;
        RECT 144.880 95.715 145.135 96.290 ;
        RECT 145.310 95.545 145.570 96.385 ;
        RECT 146.435 96.295 146.955 96.835 ;
        RECT 145.745 95.545 146.955 96.295 ;
        RECT 17.320 95.375 147.040 95.545 ;
        RECT 17.405 94.625 18.615 95.375 ;
        RECT 17.405 94.085 17.925 94.625 ;
        RECT 18.790 94.535 19.050 95.375 ;
        RECT 19.225 94.630 19.480 95.205 ;
        RECT 19.650 94.995 19.980 95.375 ;
        RECT 20.195 94.825 20.365 95.205 ;
        RECT 19.650 94.655 20.365 94.825 ;
        RECT 18.095 93.915 18.615 94.455 ;
        RECT 17.405 92.825 18.615 93.915 ;
        RECT 18.790 92.825 19.050 93.975 ;
        RECT 19.225 93.900 19.395 94.630 ;
        RECT 19.650 94.465 19.820 94.655 ;
        RECT 20.630 94.535 20.890 95.375 ;
        RECT 21.065 94.630 21.320 95.205 ;
        RECT 21.490 94.995 21.820 95.375 ;
        RECT 22.035 94.825 22.205 95.205 ;
        RECT 21.490 94.655 22.205 94.825 ;
        RECT 19.565 94.135 19.820 94.465 ;
        RECT 19.650 93.925 19.820 94.135 ;
        RECT 20.100 94.105 20.455 94.475 ;
        RECT 19.225 92.995 19.480 93.900 ;
        RECT 19.650 93.755 20.365 93.925 ;
        RECT 19.650 92.825 19.980 93.585 ;
        RECT 20.195 92.995 20.365 93.755 ;
        RECT 20.630 92.825 20.890 93.975 ;
        RECT 21.065 93.900 21.235 94.630 ;
        RECT 21.490 94.465 21.660 94.655 ;
        RECT 22.740 94.565 22.985 95.170 ;
        RECT 23.205 94.840 23.715 95.375 ;
        RECT 21.405 94.135 21.660 94.465 ;
        RECT 21.490 93.925 21.660 94.135 ;
        RECT 21.940 94.105 22.295 94.475 ;
        RECT 22.465 94.395 23.695 94.565 ;
        RECT 21.065 92.995 21.320 93.900 ;
        RECT 21.490 93.755 22.205 93.925 ;
        RECT 21.490 92.825 21.820 93.585 ;
        RECT 22.035 92.995 22.205 93.755 ;
        RECT 22.465 93.585 22.805 94.395 ;
        RECT 22.975 93.830 23.725 94.020 ;
        RECT 22.465 93.175 22.980 93.585 ;
        RECT 23.215 92.825 23.385 93.585 ;
        RECT 23.555 93.165 23.725 93.830 ;
        RECT 23.895 93.845 24.085 95.205 ;
        RECT 24.255 94.695 24.530 95.205 ;
        RECT 24.720 94.840 25.250 95.205 ;
        RECT 25.675 94.975 26.005 95.375 ;
        RECT 25.075 94.805 25.250 94.840 ;
        RECT 24.255 94.525 24.535 94.695 ;
        RECT 24.255 94.045 24.530 94.525 ;
        RECT 24.735 93.845 24.905 94.645 ;
        RECT 23.895 93.675 24.905 93.845 ;
        RECT 25.075 94.635 26.005 94.805 ;
        RECT 26.175 94.635 26.430 95.205 ;
        RECT 25.075 93.505 25.245 94.635 ;
        RECT 25.835 94.465 26.005 94.635 ;
        RECT 24.120 93.335 25.245 93.505 ;
        RECT 25.415 94.135 25.610 94.465 ;
        RECT 25.835 94.135 26.090 94.465 ;
        RECT 25.415 93.165 25.585 94.135 ;
        RECT 26.260 93.965 26.430 94.635 ;
        RECT 23.555 92.995 25.585 93.165 ;
        RECT 25.755 92.825 25.925 93.965 ;
        RECT 26.095 92.995 26.430 93.965 ;
        RECT 26.610 94.635 26.865 95.205 ;
        RECT 27.035 94.975 27.365 95.375 ;
        RECT 27.790 94.840 28.320 95.205 ;
        RECT 27.790 94.805 27.965 94.840 ;
        RECT 27.035 94.635 27.965 94.805 ;
        RECT 26.610 93.965 26.780 94.635 ;
        RECT 27.035 94.465 27.205 94.635 ;
        RECT 26.950 94.135 27.205 94.465 ;
        RECT 27.430 94.135 27.625 94.465 ;
        RECT 26.610 92.995 26.945 93.965 ;
        RECT 27.115 92.825 27.285 93.965 ;
        RECT 27.455 93.165 27.625 94.135 ;
        RECT 27.795 93.505 27.965 94.635 ;
        RECT 28.135 93.845 28.305 94.645 ;
        RECT 28.510 94.355 28.785 95.205 ;
        RECT 28.505 94.185 28.785 94.355 ;
        RECT 28.510 94.045 28.785 94.185 ;
        RECT 28.955 93.845 29.145 95.205 ;
        RECT 29.325 94.840 29.835 95.375 ;
        RECT 30.055 94.565 30.300 95.170 ;
        RECT 31.225 94.565 31.465 95.375 ;
        RECT 31.635 94.565 31.965 95.205 ;
        RECT 32.135 94.565 32.405 95.375 ;
        RECT 32.585 94.700 32.860 95.045 ;
        RECT 33.050 94.975 33.430 95.375 ;
        RECT 33.600 94.805 33.770 95.155 ;
        RECT 33.940 94.975 34.270 95.375 ;
        RECT 34.445 94.805 34.615 95.155 ;
        RECT 34.815 94.875 35.145 95.375 ;
        RECT 29.345 94.395 30.575 94.565 ;
        RECT 28.135 93.675 29.145 93.845 ;
        RECT 29.315 93.830 30.065 94.020 ;
        RECT 27.795 93.335 28.920 93.505 ;
        RECT 29.315 93.165 29.485 93.830 ;
        RECT 30.235 93.585 30.575 94.395 ;
        RECT 31.205 94.135 31.555 94.385 ;
        RECT 31.725 93.965 31.895 94.565 ;
        RECT 32.065 94.135 32.415 94.385 ;
        RECT 32.585 93.965 32.755 94.700 ;
        RECT 33.030 94.635 34.615 94.805 ;
        RECT 33.030 94.465 33.200 94.635 ;
        RECT 35.340 94.465 35.585 95.155 ;
        RECT 35.755 94.875 36.095 95.375 ;
        RECT 32.925 94.135 33.200 94.465 ;
        RECT 33.370 94.135 33.750 94.465 ;
        RECT 33.030 93.965 33.200 94.135 ;
        RECT 27.455 92.995 29.485 93.165 ;
        RECT 29.655 92.825 29.825 93.585 ;
        RECT 30.060 93.175 30.575 93.585 ;
        RECT 31.215 93.795 31.895 93.965 ;
        RECT 31.215 93.010 31.545 93.795 ;
        RECT 32.075 92.825 32.405 93.965 ;
        RECT 32.585 92.995 32.860 93.965 ;
        RECT 33.030 93.795 33.690 93.965 ;
        RECT 33.920 93.845 34.660 94.465 ;
        RECT 34.930 94.135 35.585 94.465 ;
        RECT 35.755 94.135 36.095 94.705 ;
        RECT 36.725 94.635 37.165 95.195 ;
        RECT 37.335 94.635 37.785 95.375 ;
        RECT 37.955 94.805 38.125 95.205 ;
        RECT 38.295 94.975 38.715 95.375 ;
        RECT 38.885 94.805 39.115 95.205 ;
        RECT 37.955 94.635 39.115 94.805 ;
        RECT 39.285 94.635 39.775 95.205 ;
        RECT 33.520 93.675 33.690 93.795 ;
        RECT 34.830 93.675 35.150 93.965 ;
        RECT 33.070 92.825 33.350 93.625 ;
        RECT 33.520 93.505 35.150 93.675 ;
        RECT 35.345 93.540 35.585 94.135 ;
        RECT 33.520 93.045 35.570 93.335 ;
        RECT 35.755 92.825 36.095 93.900 ;
        RECT 36.725 93.625 37.035 94.635 ;
        RECT 37.205 94.015 37.375 94.465 ;
        RECT 37.545 94.185 37.935 94.465 ;
        RECT 38.120 94.135 38.365 94.465 ;
        RECT 37.205 93.845 37.995 94.015 ;
        RECT 36.725 92.995 37.165 93.625 ;
        RECT 37.340 92.825 37.655 93.675 ;
        RECT 37.825 93.165 37.995 93.845 ;
        RECT 38.165 93.335 38.365 94.135 ;
        RECT 38.565 93.335 38.815 94.465 ;
        RECT 39.030 94.135 39.435 94.465 ;
        RECT 39.605 93.965 39.775 94.635 ;
        RECT 40.415 94.565 40.685 95.375 ;
        RECT 40.855 94.565 41.185 95.205 ;
        RECT 41.355 94.565 41.595 95.375 ;
        RECT 41.785 94.625 42.995 95.375 ;
        RECT 43.165 94.650 43.455 95.375 ;
        RECT 43.625 94.830 48.970 95.375 ;
        RECT 49.145 94.830 54.490 95.375 ;
        RECT 40.405 94.135 40.755 94.385 ;
        RECT 40.925 93.965 41.095 94.565 ;
        RECT 41.265 94.135 41.615 94.385 ;
        RECT 41.785 94.085 42.305 94.625 ;
        RECT 39.005 93.795 39.775 93.965 ;
        RECT 39.005 93.165 39.255 93.795 ;
        RECT 37.825 92.995 39.255 93.165 ;
        RECT 39.435 92.825 39.765 93.625 ;
        RECT 40.415 92.825 40.745 93.965 ;
        RECT 40.925 93.795 41.605 93.965 ;
        RECT 42.475 93.915 42.995 94.455 ;
        RECT 45.210 94.000 45.550 94.830 ;
        RECT 41.275 93.010 41.605 93.795 ;
        RECT 41.785 92.825 42.995 93.915 ;
        RECT 43.165 92.825 43.455 93.990 ;
        RECT 47.030 93.260 47.380 94.510 ;
        RECT 50.730 94.000 51.070 94.830 ;
        RECT 54.665 94.605 58.175 95.375 ;
        RECT 58.825 94.685 59.065 95.205 ;
        RECT 59.235 94.880 59.630 95.375 ;
        RECT 60.195 95.045 60.365 95.190 ;
        RECT 59.990 94.850 60.365 95.045 ;
        RECT 52.550 93.260 52.900 94.510 ;
        RECT 54.665 94.085 56.315 94.605 ;
        RECT 56.485 93.915 58.175 94.435 ;
        RECT 43.625 92.825 48.970 93.260 ;
        RECT 49.145 92.825 54.490 93.260 ;
        RECT 54.665 92.825 58.175 93.915 ;
        RECT 58.825 93.880 59.000 94.685 ;
        RECT 59.990 94.515 60.160 94.850 ;
        RECT 60.645 94.805 60.885 95.180 ;
        RECT 61.055 94.870 61.390 95.375 ;
        RECT 61.655 94.825 61.825 95.115 ;
        RECT 61.995 94.995 62.325 95.375 ;
        RECT 60.645 94.655 60.865 94.805 ;
        RECT 59.175 94.155 60.160 94.515 ;
        RECT 60.330 94.325 60.865 94.655 ;
        RECT 59.175 94.135 60.460 94.155 ;
        RECT 59.600 93.985 60.460 94.135 ;
        RECT 58.825 93.095 59.130 93.880 ;
        RECT 59.305 93.505 60.000 93.815 ;
        RECT 59.310 92.825 59.995 93.295 ;
        RECT 60.175 93.040 60.460 93.985 ;
        RECT 60.630 93.675 60.865 94.325 ;
        RECT 61.035 93.845 61.335 94.695 ;
        RECT 61.655 94.655 62.320 94.825 ;
        RECT 61.570 93.835 61.920 94.485 ;
        RECT 60.630 93.445 61.305 93.675 ;
        RECT 62.090 93.665 62.320 94.655 ;
        RECT 60.635 92.825 60.965 93.275 ;
        RECT 61.135 93.015 61.305 93.445 ;
        RECT 61.655 93.495 62.320 93.665 ;
        RECT 61.655 92.995 61.825 93.495 ;
        RECT 61.995 92.825 62.325 93.325 ;
        RECT 62.495 92.995 62.680 95.115 ;
        RECT 62.935 94.915 63.185 95.375 ;
        RECT 63.355 94.925 63.690 95.095 ;
        RECT 63.885 94.925 64.560 95.095 ;
        RECT 63.355 94.785 63.525 94.925 ;
        RECT 62.850 93.795 63.130 94.745 ;
        RECT 63.300 94.655 63.525 94.785 ;
        RECT 63.300 93.550 63.470 94.655 ;
        RECT 63.695 94.505 64.220 94.725 ;
        RECT 63.640 93.740 63.880 94.335 ;
        RECT 64.050 93.805 64.220 94.505 ;
        RECT 64.390 94.145 64.560 94.925 ;
        RECT 64.880 94.875 65.250 95.375 ;
        RECT 65.430 94.925 65.835 95.095 ;
        RECT 66.005 94.925 66.790 95.095 ;
        RECT 65.430 94.695 65.600 94.925 ;
        RECT 64.770 94.395 65.600 94.695 ;
        RECT 65.985 94.425 66.450 94.755 ;
        RECT 64.770 94.365 64.970 94.395 ;
        RECT 65.090 94.145 65.260 94.215 ;
        RECT 64.390 93.975 65.260 94.145 ;
        RECT 64.750 93.885 65.260 93.975 ;
        RECT 63.300 93.420 63.605 93.550 ;
        RECT 64.050 93.440 64.580 93.805 ;
        RECT 62.920 92.825 63.185 93.285 ;
        RECT 63.355 92.995 63.605 93.420 ;
        RECT 64.750 93.270 64.920 93.885 ;
        RECT 63.815 93.100 64.920 93.270 ;
        RECT 65.090 92.825 65.260 93.625 ;
        RECT 65.430 93.325 65.600 94.395 ;
        RECT 65.770 93.495 65.960 94.215 ;
        RECT 66.130 93.465 66.450 94.425 ;
        RECT 66.620 94.465 66.790 94.925 ;
        RECT 67.065 94.845 67.275 95.375 ;
        RECT 67.535 94.635 67.865 95.160 ;
        RECT 68.035 94.765 68.205 95.375 ;
        RECT 68.375 94.720 68.705 95.155 ;
        RECT 68.375 94.635 68.755 94.720 ;
        RECT 68.925 94.650 69.215 95.375 ;
        RECT 67.665 94.465 67.865 94.635 ;
        RECT 68.530 94.595 68.755 94.635 ;
        RECT 66.620 94.135 67.495 94.465 ;
        RECT 67.665 94.135 68.415 94.465 ;
        RECT 65.430 92.995 65.680 93.325 ;
        RECT 66.620 93.295 66.790 94.135 ;
        RECT 67.665 93.930 67.855 94.135 ;
        RECT 68.585 94.015 68.755 94.595 ;
        RECT 68.540 93.965 68.755 94.015 ;
        RECT 69.390 94.635 69.645 95.205 ;
        RECT 69.815 94.975 70.145 95.375 ;
        RECT 70.570 94.840 71.100 95.205 ;
        RECT 71.290 95.035 71.565 95.205 ;
        RECT 71.285 94.865 71.565 95.035 ;
        RECT 70.570 94.805 70.745 94.840 ;
        RECT 69.815 94.635 70.745 94.805 ;
        RECT 66.960 93.555 67.855 93.930 ;
        RECT 68.365 93.885 68.755 93.965 ;
        RECT 65.905 93.125 66.790 93.295 ;
        RECT 66.970 92.825 67.285 93.325 ;
        RECT 67.515 92.995 67.855 93.555 ;
        RECT 68.025 92.825 68.195 93.835 ;
        RECT 68.365 93.040 68.695 93.885 ;
        RECT 68.925 92.825 69.215 93.990 ;
        RECT 69.390 93.965 69.560 94.635 ;
        RECT 69.815 94.465 69.985 94.635 ;
        RECT 69.730 94.135 69.985 94.465 ;
        RECT 70.210 94.135 70.405 94.465 ;
        RECT 69.390 92.995 69.725 93.965 ;
        RECT 69.895 92.825 70.065 93.965 ;
        RECT 70.235 93.165 70.405 94.135 ;
        RECT 70.575 93.505 70.745 94.635 ;
        RECT 70.915 93.845 71.085 94.645 ;
        RECT 71.290 94.045 71.565 94.865 ;
        RECT 71.735 93.845 71.925 95.205 ;
        RECT 72.105 94.840 72.615 95.375 ;
        RECT 72.835 94.565 73.080 95.170 ;
        RECT 73.530 94.870 73.865 95.375 ;
        RECT 74.035 94.805 74.275 95.180 ;
        RECT 74.555 95.045 74.725 95.190 ;
        RECT 74.555 94.850 74.930 95.045 ;
        RECT 75.290 94.880 75.685 95.375 ;
        RECT 72.125 94.395 73.355 94.565 ;
        RECT 70.915 93.675 71.925 93.845 ;
        RECT 72.095 93.830 72.845 94.020 ;
        RECT 70.575 93.335 71.700 93.505 ;
        RECT 72.095 93.165 72.265 93.830 ;
        RECT 73.015 93.585 73.355 94.395 ;
        RECT 73.585 93.845 73.885 94.695 ;
        RECT 74.055 94.655 74.275 94.805 ;
        RECT 74.055 94.325 74.590 94.655 ;
        RECT 74.760 94.515 74.930 94.850 ;
        RECT 75.855 94.685 76.095 95.205 ;
        RECT 74.055 93.675 74.290 94.325 ;
        RECT 74.760 94.155 75.745 94.515 ;
        RECT 70.235 92.995 72.265 93.165 ;
        RECT 72.435 92.825 72.605 93.585 ;
        RECT 72.840 93.175 73.355 93.585 ;
        RECT 73.615 93.445 74.290 93.675 ;
        RECT 74.460 94.135 75.745 94.155 ;
        RECT 74.460 93.985 75.320 94.135 ;
        RECT 73.615 93.015 73.785 93.445 ;
        RECT 73.955 92.825 74.285 93.275 ;
        RECT 74.460 93.040 74.745 93.985 ;
        RECT 75.920 93.880 76.095 94.685 ;
        RECT 74.920 93.505 75.615 93.815 ;
        RECT 74.925 92.825 75.610 93.295 ;
        RECT 75.790 93.095 76.095 93.880 ;
        RECT 76.290 94.635 76.545 95.205 ;
        RECT 76.715 94.975 77.045 95.375 ;
        RECT 77.470 94.840 78.000 95.205 ;
        RECT 77.470 94.805 77.645 94.840 ;
        RECT 76.715 94.635 77.645 94.805 ;
        RECT 76.290 93.965 76.460 94.635 ;
        RECT 76.715 94.465 76.885 94.635 ;
        RECT 76.630 94.135 76.885 94.465 ;
        RECT 77.110 94.135 77.305 94.465 ;
        RECT 76.290 92.995 76.625 93.965 ;
        RECT 76.795 92.825 76.965 93.965 ;
        RECT 77.135 93.165 77.305 94.135 ;
        RECT 77.475 93.505 77.645 94.635 ;
        RECT 77.815 93.845 77.985 94.645 ;
        RECT 78.190 94.355 78.465 95.205 ;
        RECT 78.185 94.185 78.465 94.355 ;
        RECT 78.190 94.045 78.465 94.185 ;
        RECT 78.635 93.845 78.825 95.205 ;
        RECT 79.005 94.840 79.515 95.375 ;
        RECT 79.735 94.565 79.980 95.170 ;
        RECT 80.515 94.825 80.685 95.115 ;
        RECT 80.855 94.995 81.185 95.375 ;
        RECT 80.515 94.655 81.180 94.825 ;
        RECT 79.025 94.395 80.255 94.565 ;
        RECT 77.815 93.675 78.825 93.845 ;
        RECT 78.995 93.830 79.745 94.020 ;
        RECT 77.475 93.335 78.600 93.505 ;
        RECT 78.995 93.165 79.165 93.830 ;
        RECT 79.915 93.585 80.255 94.395 ;
        RECT 80.430 93.835 80.780 94.485 ;
        RECT 80.950 93.665 81.180 94.655 ;
        RECT 77.135 92.995 79.165 93.165 ;
        RECT 79.335 92.825 79.505 93.585 ;
        RECT 79.740 93.175 80.255 93.585 ;
        RECT 80.515 93.495 81.180 93.665 ;
        RECT 80.515 92.995 80.685 93.495 ;
        RECT 80.855 92.825 81.185 93.325 ;
        RECT 81.355 92.995 81.540 95.115 ;
        RECT 81.795 94.915 82.045 95.375 ;
        RECT 82.215 94.925 82.550 95.095 ;
        RECT 82.745 94.925 83.420 95.095 ;
        RECT 82.215 94.785 82.385 94.925 ;
        RECT 81.710 93.795 81.990 94.745 ;
        RECT 82.160 94.655 82.385 94.785 ;
        RECT 82.160 93.550 82.330 94.655 ;
        RECT 82.555 94.505 83.080 94.725 ;
        RECT 82.500 93.740 82.740 94.335 ;
        RECT 82.910 93.805 83.080 94.505 ;
        RECT 83.250 94.145 83.420 94.925 ;
        RECT 83.740 94.875 84.110 95.375 ;
        RECT 84.290 94.925 84.695 95.095 ;
        RECT 84.865 94.925 85.650 95.095 ;
        RECT 84.290 94.695 84.460 94.925 ;
        RECT 83.630 94.395 84.460 94.695 ;
        RECT 84.845 94.425 85.310 94.755 ;
        RECT 83.630 94.365 83.830 94.395 ;
        RECT 83.950 94.145 84.120 94.215 ;
        RECT 83.250 93.975 84.120 94.145 ;
        RECT 83.610 93.885 84.120 93.975 ;
        RECT 82.160 93.420 82.465 93.550 ;
        RECT 82.910 93.440 83.440 93.805 ;
        RECT 81.780 92.825 82.045 93.285 ;
        RECT 82.215 92.995 82.465 93.420 ;
        RECT 83.610 93.270 83.780 93.885 ;
        RECT 82.675 93.100 83.780 93.270 ;
        RECT 83.950 92.825 84.120 93.625 ;
        RECT 84.290 93.325 84.460 94.395 ;
        RECT 84.630 93.495 84.820 94.215 ;
        RECT 84.990 93.465 85.310 94.425 ;
        RECT 85.480 94.465 85.650 94.925 ;
        RECT 85.925 94.845 86.135 95.375 ;
        RECT 86.395 94.635 86.725 95.160 ;
        RECT 86.895 94.765 87.065 95.375 ;
        RECT 87.235 94.720 87.565 95.155 ;
        RECT 87.235 94.635 87.615 94.720 ;
        RECT 86.525 94.465 86.725 94.635 ;
        RECT 87.390 94.595 87.615 94.635 ;
        RECT 85.480 94.135 86.355 94.465 ;
        RECT 86.525 94.135 87.275 94.465 ;
        RECT 84.290 92.995 84.540 93.325 ;
        RECT 85.480 93.295 85.650 94.135 ;
        RECT 86.525 93.930 86.715 94.135 ;
        RECT 87.445 94.015 87.615 94.595 ;
        RECT 87.400 93.965 87.615 94.015 ;
        RECT 85.820 93.555 86.715 93.930 ;
        RECT 87.225 93.885 87.615 93.965 ;
        RECT 87.790 94.635 88.045 95.205 ;
        RECT 88.215 94.975 88.545 95.375 ;
        RECT 88.970 94.840 89.500 95.205 ;
        RECT 89.690 95.035 89.965 95.205 ;
        RECT 89.685 94.865 89.965 95.035 ;
        RECT 88.970 94.805 89.145 94.840 ;
        RECT 88.215 94.635 89.145 94.805 ;
        RECT 87.790 93.965 87.960 94.635 ;
        RECT 88.215 94.465 88.385 94.635 ;
        RECT 88.130 94.135 88.385 94.465 ;
        RECT 88.610 94.135 88.805 94.465 ;
        RECT 84.765 93.125 85.650 93.295 ;
        RECT 85.830 92.825 86.145 93.325 ;
        RECT 86.375 92.995 86.715 93.555 ;
        RECT 86.885 92.825 87.055 93.835 ;
        RECT 87.225 93.040 87.555 93.885 ;
        RECT 87.790 92.995 88.125 93.965 ;
        RECT 88.295 92.825 88.465 93.965 ;
        RECT 88.635 93.165 88.805 94.135 ;
        RECT 88.975 93.505 89.145 94.635 ;
        RECT 89.315 93.845 89.485 94.645 ;
        RECT 89.690 94.045 89.965 94.865 ;
        RECT 90.135 93.845 90.325 95.205 ;
        RECT 90.505 94.840 91.015 95.375 ;
        RECT 91.235 94.565 91.480 95.170 ;
        RECT 91.930 94.870 92.265 95.375 ;
        RECT 92.435 94.805 92.675 95.180 ;
        RECT 92.955 95.045 93.125 95.190 ;
        RECT 92.955 94.850 93.330 95.045 ;
        RECT 93.690 94.880 94.085 95.375 ;
        RECT 90.525 94.395 91.755 94.565 ;
        RECT 89.315 93.675 90.325 93.845 ;
        RECT 90.495 93.830 91.245 94.020 ;
        RECT 88.975 93.335 90.100 93.505 ;
        RECT 90.495 93.165 90.665 93.830 ;
        RECT 91.415 93.585 91.755 94.395 ;
        RECT 91.985 93.845 92.285 94.695 ;
        RECT 92.455 94.655 92.675 94.805 ;
        RECT 92.455 94.325 92.990 94.655 ;
        RECT 93.160 94.515 93.330 94.850 ;
        RECT 94.255 94.685 94.495 95.205 ;
        RECT 92.455 93.675 92.690 94.325 ;
        RECT 93.160 94.155 94.145 94.515 ;
        RECT 88.635 92.995 90.665 93.165 ;
        RECT 90.835 92.825 91.005 93.585 ;
        RECT 91.240 93.175 91.755 93.585 ;
        RECT 92.015 93.445 92.690 93.675 ;
        RECT 92.860 94.135 94.145 94.155 ;
        RECT 92.860 93.985 93.720 94.135 ;
        RECT 94.320 94.015 94.495 94.685 ;
        RECT 94.685 94.650 94.975 95.375 ;
        RECT 95.235 94.825 95.405 95.115 ;
        RECT 95.575 94.995 95.905 95.375 ;
        RECT 95.235 94.655 95.900 94.825 ;
        RECT 92.015 93.015 92.185 93.445 ;
        RECT 92.355 92.825 92.685 93.275 ;
        RECT 92.860 93.040 93.145 93.985 ;
        RECT 94.285 93.880 94.495 94.015 ;
        RECT 93.320 93.505 94.015 93.815 ;
        RECT 93.325 92.825 94.010 93.295 ;
        RECT 94.190 93.095 94.495 93.880 ;
        RECT 94.685 92.825 94.975 93.990 ;
        RECT 95.150 93.835 95.500 94.485 ;
        RECT 95.670 93.665 95.900 94.655 ;
        RECT 95.235 93.495 95.900 93.665 ;
        RECT 95.235 92.995 95.405 93.495 ;
        RECT 95.575 92.825 95.905 93.325 ;
        RECT 96.075 92.995 96.260 95.115 ;
        RECT 96.515 94.915 96.765 95.375 ;
        RECT 96.935 94.925 97.270 95.095 ;
        RECT 97.465 94.925 98.140 95.095 ;
        RECT 96.935 94.785 97.105 94.925 ;
        RECT 96.430 93.795 96.710 94.745 ;
        RECT 96.880 94.655 97.105 94.785 ;
        RECT 96.880 93.550 97.050 94.655 ;
        RECT 97.275 94.505 97.800 94.725 ;
        RECT 97.220 93.740 97.460 94.335 ;
        RECT 97.630 93.805 97.800 94.505 ;
        RECT 97.970 94.145 98.140 94.925 ;
        RECT 98.460 94.875 98.830 95.375 ;
        RECT 99.010 94.925 99.415 95.095 ;
        RECT 99.585 94.925 100.370 95.095 ;
        RECT 99.010 94.695 99.180 94.925 ;
        RECT 98.350 94.395 99.180 94.695 ;
        RECT 99.565 94.425 100.030 94.755 ;
        RECT 98.350 94.365 98.550 94.395 ;
        RECT 98.670 94.145 98.840 94.215 ;
        RECT 97.970 93.975 98.840 94.145 ;
        RECT 98.330 93.885 98.840 93.975 ;
        RECT 96.880 93.420 97.185 93.550 ;
        RECT 97.630 93.440 98.160 93.805 ;
        RECT 96.500 92.825 96.765 93.285 ;
        RECT 96.935 92.995 97.185 93.420 ;
        RECT 98.330 93.270 98.500 93.885 ;
        RECT 97.395 93.100 98.500 93.270 ;
        RECT 98.670 92.825 98.840 93.625 ;
        RECT 99.010 93.325 99.180 94.395 ;
        RECT 99.350 93.495 99.540 94.215 ;
        RECT 99.710 93.465 100.030 94.425 ;
        RECT 100.200 94.465 100.370 94.925 ;
        RECT 100.645 94.845 100.855 95.375 ;
        RECT 101.115 94.635 101.445 95.160 ;
        RECT 101.615 94.765 101.785 95.375 ;
        RECT 101.955 94.720 102.285 95.155 ;
        RECT 101.955 94.635 102.335 94.720 ;
        RECT 101.245 94.465 101.445 94.635 ;
        RECT 102.110 94.595 102.335 94.635 ;
        RECT 100.200 94.135 101.075 94.465 ;
        RECT 101.245 94.135 101.995 94.465 ;
        RECT 99.010 92.995 99.260 93.325 ;
        RECT 100.200 93.295 100.370 94.135 ;
        RECT 101.245 93.930 101.435 94.135 ;
        RECT 102.165 94.015 102.335 94.595 ;
        RECT 102.120 93.965 102.335 94.015 ;
        RECT 100.540 93.555 101.435 93.930 ;
        RECT 101.945 93.885 102.335 93.965 ;
        RECT 102.510 94.635 102.765 95.205 ;
        RECT 102.935 94.975 103.265 95.375 ;
        RECT 103.690 94.840 104.220 95.205 ;
        RECT 104.410 95.035 104.685 95.205 ;
        RECT 104.405 94.865 104.685 95.035 ;
        RECT 103.690 94.805 103.865 94.840 ;
        RECT 102.935 94.635 103.865 94.805 ;
        RECT 102.510 93.965 102.680 94.635 ;
        RECT 102.935 94.465 103.105 94.635 ;
        RECT 102.850 94.135 103.105 94.465 ;
        RECT 103.330 94.135 103.525 94.465 ;
        RECT 99.485 93.125 100.370 93.295 ;
        RECT 100.550 92.825 100.865 93.325 ;
        RECT 101.095 92.995 101.435 93.555 ;
        RECT 101.605 92.825 101.775 93.835 ;
        RECT 101.945 93.040 102.275 93.885 ;
        RECT 102.510 92.995 102.845 93.965 ;
        RECT 103.015 92.825 103.185 93.965 ;
        RECT 103.355 93.165 103.525 94.135 ;
        RECT 103.695 93.505 103.865 94.635 ;
        RECT 104.035 93.845 104.205 94.645 ;
        RECT 104.410 94.045 104.685 94.865 ;
        RECT 104.855 93.845 105.045 95.205 ;
        RECT 105.225 94.840 105.735 95.375 ;
        RECT 105.955 94.565 106.200 95.170 ;
        RECT 107.195 94.825 107.365 95.115 ;
        RECT 107.535 94.995 107.865 95.375 ;
        RECT 107.195 94.655 107.860 94.825 ;
        RECT 105.245 94.395 106.475 94.565 ;
        RECT 104.035 93.675 105.045 93.845 ;
        RECT 105.215 93.830 105.965 94.020 ;
        RECT 103.695 93.335 104.820 93.505 ;
        RECT 105.215 93.165 105.385 93.830 ;
        RECT 106.135 93.585 106.475 94.395 ;
        RECT 107.110 93.835 107.460 94.485 ;
        RECT 107.630 93.665 107.860 94.655 ;
        RECT 103.355 92.995 105.385 93.165 ;
        RECT 105.555 92.825 105.725 93.585 ;
        RECT 105.960 93.175 106.475 93.585 ;
        RECT 107.195 93.495 107.860 93.665 ;
        RECT 107.195 92.995 107.365 93.495 ;
        RECT 107.535 92.825 107.865 93.325 ;
        RECT 108.035 92.995 108.220 95.115 ;
        RECT 108.475 94.915 108.725 95.375 ;
        RECT 108.895 94.925 109.230 95.095 ;
        RECT 109.425 94.925 110.100 95.095 ;
        RECT 108.895 94.785 109.065 94.925 ;
        RECT 108.390 93.795 108.670 94.745 ;
        RECT 108.840 94.655 109.065 94.785 ;
        RECT 108.840 93.550 109.010 94.655 ;
        RECT 109.235 94.505 109.760 94.725 ;
        RECT 109.180 93.740 109.420 94.335 ;
        RECT 109.590 93.805 109.760 94.505 ;
        RECT 109.930 94.145 110.100 94.925 ;
        RECT 110.420 94.875 110.790 95.375 ;
        RECT 110.970 94.925 111.375 95.095 ;
        RECT 111.545 94.925 112.330 95.095 ;
        RECT 110.970 94.695 111.140 94.925 ;
        RECT 110.310 94.395 111.140 94.695 ;
        RECT 111.525 94.425 111.990 94.755 ;
        RECT 110.310 94.365 110.510 94.395 ;
        RECT 110.630 94.145 110.800 94.215 ;
        RECT 109.930 93.975 110.800 94.145 ;
        RECT 110.290 93.885 110.800 93.975 ;
        RECT 108.840 93.420 109.145 93.550 ;
        RECT 109.590 93.440 110.120 93.805 ;
        RECT 108.460 92.825 108.725 93.285 ;
        RECT 108.895 92.995 109.145 93.420 ;
        RECT 110.290 93.270 110.460 93.885 ;
        RECT 109.355 93.100 110.460 93.270 ;
        RECT 110.630 92.825 110.800 93.625 ;
        RECT 110.970 93.325 111.140 94.395 ;
        RECT 111.310 93.495 111.500 94.215 ;
        RECT 111.670 93.465 111.990 94.425 ;
        RECT 112.160 94.465 112.330 94.925 ;
        RECT 112.605 94.845 112.815 95.375 ;
        RECT 113.075 94.635 113.405 95.160 ;
        RECT 113.575 94.765 113.745 95.375 ;
        RECT 113.915 94.720 114.245 95.155 ;
        RECT 113.915 94.635 114.295 94.720 ;
        RECT 113.205 94.465 113.405 94.635 ;
        RECT 114.070 94.595 114.295 94.635 ;
        RECT 112.160 94.135 113.035 94.465 ;
        RECT 113.205 94.135 113.955 94.465 ;
        RECT 110.970 92.995 111.220 93.325 ;
        RECT 112.160 93.295 112.330 94.135 ;
        RECT 113.205 93.930 113.395 94.135 ;
        RECT 114.125 94.015 114.295 94.595 ;
        RECT 114.080 93.965 114.295 94.015 ;
        RECT 112.500 93.555 113.395 93.930 ;
        RECT 113.905 93.885 114.295 93.965 ;
        RECT 114.470 94.635 114.725 95.205 ;
        RECT 114.895 94.975 115.225 95.375 ;
        RECT 115.650 94.840 116.180 95.205 ;
        RECT 115.650 94.805 115.825 94.840 ;
        RECT 114.895 94.635 115.825 94.805 ;
        RECT 116.370 94.695 116.645 95.205 ;
        RECT 114.470 93.965 114.640 94.635 ;
        RECT 114.895 94.465 115.065 94.635 ;
        RECT 114.810 94.135 115.065 94.465 ;
        RECT 115.290 94.135 115.485 94.465 ;
        RECT 111.445 93.125 112.330 93.295 ;
        RECT 112.510 92.825 112.825 93.325 ;
        RECT 113.055 92.995 113.395 93.555 ;
        RECT 113.565 92.825 113.735 93.835 ;
        RECT 113.905 93.040 114.235 93.885 ;
        RECT 114.470 92.995 114.805 93.965 ;
        RECT 114.975 92.825 115.145 93.965 ;
        RECT 115.315 93.165 115.485 94.135 ;
        RECT 115.655 93.505 115.825 94.635 ;
        RECT 115.995 93.845 116.165 94.645 ;
        RECT 116.365 94.525 116.645 94.695 ;
        RECT 116.370 94.045 116.645 94.525 ;
        RECT 116.815 93.845 117.005 95.205 ;
        RECT 117.185 94.840 117.695 95.375 ;
        RECT 117.915 94.565 118.160 95.170 ;
        RECT 118.605 94.605 120.275 95.375 ;
        RECT 120.445 94.650 120.735 95.375 ;
        RECT 120.910 94.635 121.165 95.205 ;
        RECT 121.335 94.975 121.665 95.375 ;
        RECT 122.090 94.840 122.620 95.205 ;
        RECT 122.810 95.035 123.085 95.205 ;
        RECT 122.805 94.865 123.085 95.035 ;
        RECT 122.090 94.805 122.265 94.840 ;
        RECT 121.335 94.635 122.265 94.805 ;
        RECT 117.205 94.395 118.435 94.565 ;
        RECT 115.995 93.675 117.005 93.845 ;
        RECT 117.175 93.830 117.925 94.020 ;
        RECT 115.655 93.335 116.780 93.505 ;
        RECT 117.175 93.165 117.345 93.830 ;
        RECT 118.095 93.585 118.435 94.395 ;
        RECT 118.605 94.085 119.355 94.605 ;
        RECT 119.525 93.915 120.275 94.435 ;
        RECT 115.315 92.995 117.345 93.165 ;
        RECT 117.515 92.825 117.685 93.585 ;
        RECT 117.920 93.175 118.435 93.585 ;
        RECT 118.605 92.825 120.275 93.915 ;
        RECT 120.445 92.825 120.735 93.990 ;
        RECT 120.910 93.965 121.080 94.635 ;
        RECT 121.335 94.465 121.505 94.635 ;
        RECT 121.250 94.135 121.505 94.465 ;
        RECT 121.730 94.135 121.925 94.465 ;
        RECT 120.910 92.995 121.245 93.965 ;
        RECT 121.415 92.825 121.585 93.965 ;
        RECT 121.755 93.165 121.925 94.135 ;
        RECT 122.095 93.505 122.265 94.635 ;
        RECT 122.435 93.845 122.605 94.645 ;
        RECT 122.810 94.045 123.085 94.865 ;
        RECT 123.255 93.845 123.445 95.205 ;
        RECT 123.625 94.840 124.135 95.375 ;
        RECT 124.355 94.565 124.600 95.170 ;
        RECT 125.045 94.625 126.255 95.375 ;
        RECT 126.515 94.825 126.685 95.115 ;
        RECT 126.855 94.995 127.185 95.375 ;
        RECT 126.515 94.655 127.180 94.825 ;
        RECT 123.645 94.395 124.875 94.565 ;
        RECT 122.435 93.675 123.445 93.845 ;
        RECT 123.615 93.830 124.365 94.020 ;
        RECT 122.095 93.335 123.220 93.505 ;
        RECT 123.615 93.165 123.785 93.830 ;
        RECT 124.535 93.585 124.875 94.395 ;
        RECT 125.045 94.085 125.565 94.625 ;
        RECT 125.735 93.915 126.255 94.455 ;
        RECT 121.755 92.995 123.785 93.165 ;
        RECT 123.955 92.825 124.125 93.585 ;
        RECT 124.360 93.175 124.875 93.585 ;
        RECT 125.045 92.825 126.255 93.915 ;
        RECT 126.430 93.835 126.780 94.485 ;
        RECT 126.950 93.665 127.180 94.655 ;
        RECT 126.515 93.495 127.180 93.665 ;
        RECT 126.515 92.995 126.685 93.495 ;
        RECT 126.855 92.825 127.185 93.325 ;
        RECT 127.355 92.995 127.540 95.115 ;
        RECT 127.795 94.915 128.045 95.375 ;
        RECT 128.215 94.925 128.550 95.095 ;
        RECT 128.745 94.925 129.420 95.095 ;
        RECT 128.215 94.785 128.385 94.925 ;
        RECT 127.710 93.795 127.990 94.745 ;
        RECT 128.160 94.655 128.385 94.785 ;
        RECT 128.160 93.550 128.330 94.655 ;
        RECT 128.555 94.505 129.080 94.725 ;
        RECT 128.500 93.740 128.740 94.335 ;
        RECT 128.910 93.805 129.080 94.505 ;
        RECT 129.250 94.145 129.420 94.925 ;
        RECT 129.740 94.875 130.110 95.375 ;
        RECT 130.290 94.925 130.695 95.095 ;
        RECT 130.865 94.925 131.650 95.095 ;
        RECT 130.290 94.695 130.460 94.925 ;
        RECT 129.630 94.395 130.460 94.695 ;
        RECT 130.845 94.425 131.310 94.755 ;
        RECT 129.630 94.365 129.830 94.395 ;
        RECT 129.950 94.145 130.120 94.215 ;
        RECT 129.250 93.975 130.120 94.145 ;
        RECT 129.610 93.885 130.120 93.975 ;
        RECT 128.160 93.420 128.465 93.550 ;
        RECT 128.910 93.440 129.440 93.805 ;
        RECT 127.780 92.825 128.045 93.285 ;
        RECT 128.215 92.995 128.465 93.420 ;
        RECT 129.610 93.270 129.780 93.885 ;
        RECT 128.675 93.100 129.780 93.270 ;
        RECT 129.950 92.825 130.120 93.625 ;
        RECT 130.290 93.325 130.460 94.395 ;
        RECT 130.630 93.495 130.820 94.215 ;
        RECT 130.990 93.465 131.310 94.425 ;
        RECT 131.480 94.465 131.650 94.925 ;
        RECT 131.925 94.845 132.135 95.375 ;
        RECT 132.395 94.635 132.725 95.160 ;
        RECT 132.895 94.765 133.065 95.375 ;
        RECT 133.235 94.720 133.565 95.155 ;
        RECT 133.785 94.875 134.045 95.205 ;
        RECT 134.255 94.895 134.530 95.375 ;
        RECT 133.235 94.635 133.615 94.720 ;
        RECT 132.525 94.465 132.725 94.635 ;
        RECT 133.390 94.595 133.615 94.635 ;
        RECT 131.480 94.135 132.355 94.465 ;
        RECT 132.525 94.135 133.275 94.465 ;
        RECT 130.290 92.995 130.540 93.325 ;
        RECT 131.480 93.295 131.650 94.135 ;
        RECT 132.525 93.930 132.715 94.135 ;
        RECT 133.445 94.015 133.615 94.595 ;
        RECT 133.400 93.965 133.615 94.015 ;
        RECT 131.820 93.555 132.715 93.930 ;
        RECT 133.225 93.885 133.615 93.965 ;
        RECT 133.785 93.965 133.955 94.875 ;
        RECT 134.740 94.805 134.945 95.205 ;
        RECT 135.115 94.975 135.450 95.375 ;
        RECT 134.125 94.135 134.485 94.715 ;
        RECT 134.740 94.635 135.425 94.805 ;
        RECT 134.665 93.965 134.915 94.465 ;
        RECT 130.765 93.125 131.650 93.295 ;
        RECT 131.830 92.825 132.145 93.325 ;
        RECT 132.375 92.995 132.715 93.555 ;
        RECT 132.885 92.825 133.055 93.835 ;
        RECT 133.225 93.040 133.555 93.885 ;
        RECT 133.785 93.795 134.915 93.965 ;
        RECT 133.785 93.025 134.055 93.795 ;
        RECT 135.085 93.605 135.425 94.635 ;
        RECT 134.225 92.825 134.555 93.605 ;
        RECT 134.760 93.430 135.425 93.605 ;
        RECT 136.090 94.635 136.345 95.205 ;
        RECT 136.515 94.975 136.845 95.375 ;
        RECT 137.270 94.840 137.800 95.205 ;
        RECT 137.990 95.035 138.265 95.205 ;
        RECT 137.985 94.865 138.265 95.035 ;
        RECT 137.270 94.805 137.445 94.840 ;
        RECT 136.515 94.635 137.445 94.805 ;
        RECT 136.090 93.965 136.260 94.635 ;
        RECT 136.515 94.465 136.685 94.635 ;
        RECT 136.430 94.135 136.685 94.465 ;
        RECT 136.910 94.135 137.105 94.465 ;
        RECT 134.760 93.025 134.945 93.430 ;
        RECT 135.115 92.825 135.450 93.250 ;
        RECT 136.090 92.995 136.425 93.965 ;
        RECT 136.595 92.825 136.765 93.965 ;
        RECT 136.935 93.165 137.105 94.135 ;
        RECT 137.275 93.505 137.445 94.635 ;
        RECT 137.615 93.845 137.785 94.645 ;
        RECT 137.990 94.045 138.265 94.865 ;
        RECT 138.435 93.845 138.625 95.205 ;
        RECT 138.805 94.840 139.315 95.375 ;
        RECT 139.535 94.565 139.780 95.170 ;
        RECT 140.225 94.875 140.485 95.205 ;
        RECT 140.655 95.015 140.985 95.375 ;
        RECT 141.240 94.995 142.540 95.205 ;
        RECT 138.825 94.395 140.055 94.565 ;
        RECT 137.615 93.675 138.625 93.845 ;
        RECT 138.795 93.830 139.545 94.020 ;
        RECT 137.275 93.335 138.400 93.505 ;
        RECT 138.795 93.165 138.965 93.830 ;
        RECT 139.715 93.585 140.055 94.395 ;
        RECT 136.935 92.995 138.965 93.165 ;
        RECT 139.135 92.825 139.305 93.585 ;
        RECT 139.540 93.175 140.055 93.585 ;
        RECT 140.225 93.675 140.395 94.875 ;
        RECT 141.240 94.845 141.410 94.995 ;
        RECT 140.655 94.720 141.410 94.845 ;
        RECT 140.565 94.675 141.410 94.720 ;
        RECT 140.565 94.555 140.835 94.675 ;
        RECT 140.565 93.980 140.735 94.555 ;
        RECT 140.965 94.115 141.375 94.420 ;
        RECT 141.665 94.385 141.875 94.785 ;
        RECT 141.545 94.175 141.875 94.385 ;
        RECT 142.120 94.385 142.340 94.785 ;
        RECT 142.815 94.610 143.270 95.375 ;
        RECT 143.995 94.825 144.165 95.205 ;
        RECT 144.380 94.995 144.710 95.375 ;
        RECT 143.995 94.655 144.710 94.825 ;
        RECT 142.120 94.175 142.595 94.385 ;
        RECT 142.785 94.185 143.275 94.385 ;
        RECT 143.905 94.105 144.260 94.475 ;
        RECT 144.540 94.465 144.710 94.655 ;
        RECT 144.880 94.630 145.135 95.205 ;
        RECT 144.540 94.135 144.795 94.465 ;
        RECT 140.565 93.945 140.765 93.980 ;
        RECT 142.095 93.945 143.270 94.005 ;
        RECT 140.565 93.835 143.270 93.945 ;
        RECT 144.540 93.925 144.710 94.135 ;
        RECT 140.625 93.775 142.425 93.835 ;
        RECT 142.095 93.745 142.425 93.775 ;
        RECT 140.225 92.995 140.485 93.675 ;
        RECT 140.655 92.825 140.905 93.605 ;
        RECT 141.155 93.575 141.990 93.585 ;
        RECT 142.580 93.575 142.765 93.665 ;
        RECT 141.155 93.375 142.765 93.575 ;
        RECT 141.155 92.995 141.405 93.375 ;
        RECT 142.535 93.335 142.765 93.375 ;
        RECT 143.015 93.215 143.270 93.835 ;
        RECT 141.575 92.825 141.930 93.205 ;
        RECT 142.935 92.995 143.270 93.215 ;
        RECT 143.995 93.755 144.710 93.925 ;
        RECT 144.965 93.900 145.135 94.630 ;
        RECT 145.310 94.535 145.570 95.375 ;
        RECT 145.745 94.625 146.955 95.375 ;
        RECT 143.995 92.995 144.165 93.755 ;
        RECT 144.380 92.825 144.710 93.585 ;
        RECT 144.880 92.995 145.135 93.900 ;
        RECT 145.310 92.825 145.570 93.975 ;
        RECT 145.745 93.915 146.265 94.455 ;
        RECT 146.435 94.085 146.955 94.625 ;
        RECT 145.745 92.825 146.955 93.915 ;
        RECT 17.320 92.655 147.040 92.825 ;
        RECT 17.405 91.565 18.615 92.655 ;
        RECT 18.785 91.565 21.375 92.655 ;
        RECT 21.635 91.985 21.805 92.485 ;
        RECT 21.975 92.155 22.305 92.655 ;
        RECT 21.635 91.815 22.300 91.985 ;
        RECT 17.405 90.855 17.925 91.395 ;
        RECT 18.095 91.025 18.615 91.565 ;
        RECT 18.785 90.875 19.995 91.395 ;
        RECT 20.165 91.045 21.375 91.565 ;
        RECT 21.550 90.995 21.900 91.645 ;
        RECT 17.405 90.105 18.615 90.855 ;
        RECT 18.785 90.105 21.375 90.875 ;
        RECT 22.070 90.825 22.300 91.815 ;
        RECT 21.635 90.655 22.300 90.825 ;
        RECT 21.635 90.365 21.805 90.655 ;
        RECT 21.975 90.105 22.305 90.485 ;
        RECT 22.475 90.365 22.660 92.485 ;
        RECT 22.900 92.195 23.165 92.655 ;
        RECT 23.335 92.060 23.585 92.485 ;
        RECT 23.795 92.210 24.900 92.380 ;
        RECT 23.280 91.930 23.585 92.060 ;
        RECT 22.830 90.735 23.110 91.685 ;
        RECT 23.280 90.825 23.450 91.930 ;
        RECT 23.620 91.145 23.860 91.740 ;
        RECT 24.030 91.675 24.560 92.040 ;
        RECT 24.030 90.975 24.200 91.675 ;
        RECT 24.730 91.595 24.900 92.210 ;
        RECT 25.070 91.855 25.240 92.655 ;
        RECT 25.410 92.155 25.660 92.485 ;
        RECT 25.885 92.185 26.770 92.355 ;
        RECT 24.730 91.505 25.240 91.595 ;
        RECT 23.280 90.695 23.505 90.825 ;
        RECT 23.675 90.755 24.200 90.975 ;
        RECT 24.370 91.335 25.240 91.505 ;
        RECT 22.915 90.105 23.165 90.565 ;
        RECT 23.335 90.555 23.505 90.695 ;
        RECT 24.370 90.555 24.540 91.335 ;
        RECT 25.070 91.265 25.240 91.335 ;
        RECT 24.750 91.085 24.950 91.115 ;
        RECT 25.410 91.085 25.580 92.155 ;
        RECT 25.750 91.265 25.940 91.985 ;
        RECT 24.750 90.785 25.580 91.085 ;
        RECT 26.110 91.055 26.430 92.015 ;
        RECT 23.335 90.385 23.670 90.555 ;
        RECT 23.865 90.385 24.540 90.555 ;
        RECT 24.860 90.105 25.230 90.605 ;
        RECT 25.410 90.555 25.580 90.785 ;
        RECT 25.965 90.725 26.430 91.055 ;
        RECT 26.600 91.345 26.770 92.185 ;
        RECT 26.950 92.155 27.265 92.655 ;
        RECT 27.495 91.925 27.835 92.485 ;
        RECT 26.940 91.550 27.835 91.925 ;
        RECT 28.005 91.645 28.175 92.655 ;
        RECT 27.645 91.345 27.835 91.550 ;
        RECT 28.345 91.595 28.675 92.440 ;
        RECT 28.345 91.515 28.735 91.595 ;
        RECT 28.915 91.515 29.245 92.655 ;
        RECT 29.775 91.685 30.105 92.470 ;
        RECT 29.425 91.515 30.105 91.685 ;
        RECT 28.520 91.465 28.735 91.515 ;
        RECT 26.600 91.015 27.475 91.345 ;
        RECT 27.645 91.015 28.395 91.345 ;
        RECT 26.600 90.555 26.770 91.015 ;
        RECT 27.645 90.845 27.845 91.015 ;
        RECT 28.565 90.885 28.735 91.465 ;
        RECT 28.905 91.095 29.255 91.345 ;
        RECT 29.425 90.915 29.595 91.515 ;
        RECT 30.285 91.490 30.575 92.655 ;
        RECT 31.665 91.500 32.005 92.485 ;
        RECT 32.175 92.225 32.585 92.655 ;
        RECT 33.330 92.235 33.660 92.655 ;
        RECT 33.830 92.055 34.155 92.485 ;
        RECT 32.175 91.885 34.155 92.055 ;
        RECT 29.765 91.095 30.115 91.345 ;
        RECT 28.510 90.845 28.735 90.885 ;
        RECT 25.410 90.385 25.815 90.555 ;
        RECT 25.985 90.385 26.770 90.555 ;
        RECT 27.045 90.105 27.255 90.635 ;
        RECT 27.515 90.320 27.845 90.845 ;
        RECT 28.355 90.760 28.735 90.845 ;
        RECT 28.015 90.105 28.185 90.715 ;
        RECT 28.355 90.325 28.685 90.760 ;
        RECT 28.915 90.105 29.185 90.915 ;
        RECT 29.355 90.275 29.685 90.915 ;
        RECT 29.855 90.105 30.095 90.915 ;
        RECT 31.665 90.845 31.920 91.500 ;
        RECT 32.175 91.345 32.440 91.885 ;
        RECT 32.655 91.545 33.280 91.715 ;
        RECT 32.090 91.015 32.440 91.345 ;
        RECT 32.610 91.015 32.940 91.345 ;
        RECT 33.110 90.845 33.280 91.545 ;
        RECT 30.285 90.105 30.575 90.830 ;
        RECT 31.665 90.470 32.025 90.845 ;
        RECT 32.290 90.105 32.460 90.845 ;
        RECT 32.740 90.675 33.280 90.845 ;
        RECT 33.450 91.475 34.155 91.885 ;
        RECT 34.630 91.555 34.960 92.655 ;
        RECT 35.345 91.500 35.685 92.485 ;
        RECT 35.855 92.225 36.265 92.655 ;
        RECT 37.010 92.235 37.340 92.655 ;
        RECT 37.510 92.055 37.835 92.485 ;
        RECT 35.855 91.885 37.835 92.055 ;
        RECT 32.740 90.470 32.910 90.675 ;
        RECT 33.450 90.275 33.620 91.475 ;
        RECT 33.790 91.095 34.360 91.305 ;
        RECT 34.530 91.095 35.175 91.305 ;
        RECT 33.850 90.755 35.020 90.925 ;
        RECT 33.850 90.275 34.180 90.755 ;
        RECT 34.350 90.105 34.520 90.575 ;
        RECT 34.690 90.290 35.020 90.755 ;
        RECT 35.345 90.845 35.600 91.500 ;
        RECT 35.855 91.345 36.120 91.885 ;
        RECT 36.335 91.545 36.960 91.715 ;
        RECT 35.770 91.015 36.120 91.345 ;
        RECT 36.290 91.015 36.620 91.345 ;
        RECT 36.790 90.845 36.960 91.545 ;
        RECT 35.345 90.470 35.705 90.845 ;
        RECT 35.405 90.445 35.575 90.470 ;
        RECT 35.970 90.105 36.140 90.845 ;
        RECT 36.420 90.675 36.960 90.845 ;
        RECT 37.130 91.475 37.835 91.885 ;
        RECT 38.310 91.555 38.640 92.655 ;
        RECT 39.025 91.500 39.365 92.485 ;
        RECT 39.535 92.225 39.945 92.655 ;
        RECT 40.690 92.235 41.020 92.655 ;
        RECT 41.190 92.055 41.515 92.485 ;
        RECT 39.535 91.885 41.515 92.055 ;
        RECT 36.420 90.470 36.590 90.675 ;
        RECT 37.130 90.275 37.300 91.475 ;
        RECT 37.470 91.095 38.040 91.305 ;
        RECT 38.210 91.095 38.855 91.305 ;
        RECT 37.530 90.755 38.700 90.925 ;
        RECT 37.530 90.275 37.860 90.755 ;
        RECT 38.030 90.105 38.200 90.575 ;
        RECT 38.370 90.290 38.700 90.755 ;
        RECT 39.025 90.845 39.280 91.500 ;
        RECT 39.535 91.345 39.800 91.885 ;
        RECT 40.015 91.545 40.640 91.715 ;
        RECT 39.450 91.015 39.800 91.345 ;
        RECT 39.970 91.015 40.300 91.345 ;
        RECT 40.470 90.845 40.640 91.545 ;
        RECT 39.025 90.470 39.385 90.845 ;
        RECT 39.650 90.105 39.820 90.845 ;
        RECT 40.100 90.675 40.640 90.845 ;
        RECT 40.810 91.475 41.515 91.885 ;
        RECT 41.990 91.555 42.320 92.655 ;
        RECT 42.705 91.500 43.045 92.485 ;
        RECT 43.215 92.225 43.625 92.655 ;
        RECT 44.370 92.235 44.700 92.655 ;
        RECT 44.870 92.055 45.195 92.485 ;
        RECT 43.215 91.885 45.195 92.055 ;
        RECT 40.100 90.470 40.270 90.675 ;
        RECT 40.810 90.275 40.980 91.475 ;
        RECT 41.150 91.095 41.720 91.305 ;
        RECT 41.890 91.095 42.535 91.305 ;
        RECT 41.210 90.755 42.380 90.925 ;
        RECT 41.210 90.275 41.540 90.755 ;
        RECT 41.710 90.105 41.880 90.575 ;
        RECT 42.050 90.290 42.380 90.755 ;
        RECT 42.705 90.845 42.960 91.500 ;
        RECT 43.215 91.345 43.480 91.885 ;
        RECT 43.695 91.545 44.320 91.715 ;
        RECT 43.130 91.015 43.480 91.345 ;
        RECT 43.650 91.015 43.980 91.345 ;
        RECT 44.150 90.845 44.320 91.545 ;
        RECT 42.705 90.470 43.065 90.845 ;
        RECT 43.330 90.105 43.500 90.845 ;
        RECT 43.780 90.675 44.320 90.845 ;
        RECT 44.490 91.475 45.195 91.885 ;
        RECT 45.670 91.555 46.000 92.655 ;
        RECT 46.475 92.035 46.645 92.465 ;
        RECT 46.815 92.205 47.145 92.655 ;
        RECT 46.475 91.805 47.150 92.035 ;
        RECT 43.780 90.470 43.950 90.675 ;
        RECT 44.490 90.275 44.660 91.475 ;
        RECT 44.830 91.095 45.400 91.305 ;
        RECT 45.570 91.095 46.215 91.305 ;
        RECT 44.890 90.755 46.060 90.925 ;
        RECT 46.445 90.785 46.745 91.635 ;
        RECT 46.915 91.155 47.150 91.805 ;
        RECT 47.320 91.495 47.605 92.440 ;
        RECT 47.785 92.185 48.470 92.655 ;
        RECT 47.780 91.665 48.475 91.975 ;
        RECT 48.650 91.600 48.955 92.385 ;
        RECT 49.145 92.220 54.490 92.655 ;
        RECT 47.320 91.345 48.180 91.495 ;
        RECT 48.745 91.465 48.955 91.600 ;
        RECT 47.320 91.325 48.605 91.345 ;
        RECT 46.915 90.825 47.450 91.155 ;
        RECT 47.620 90.965 48.605 91.325 ;
        RECT 44.890 90.275 45.220 90.755 ;
        RECT 45.390 90.105 45.560 90.575 ;
        RECT 45.730 90.290 46.060 90.755 ;
        RECT 46.915 90.675 47.135 90.825 ;
        RECT 46.390 90.105 46.725 90.610 ;
        RECT 46.895 90.300 47.135 90.675 ;
        RECT 47.620 90.630 47.790 90.965 ;
        RECT 48.780 90.795 48.955 91.465 ;
        RECT 47.415 90.435 47.790 90.630 ;
        RECT 47.415 90.290 47.585 90.435 ;
        RECT 48.150 90.105 48.545 90.600 ;
        RECT 48.715 90.275 48.955 90.795 ;
        RECT 50.730 90.650 51.070 91.480 ;
        RECT 52.550 90.970 52.900 92.220 ;
        RECT 54.665 91.565 55.875 92.655 ;
        RECT 54.665 90.855 55.185 91.395 ;
        RECT 55.355 91.025 55.875 91.565 ;
        RECT 56.045 91.490 56.335 92.655 ;
        RECT 56.505 91.565 57.715 92.655 ;
        RECT 57.975 91.985 58.145 92.485 ;
        RECT 58.315 92.155 58.645 92.655 ;
        RECT 57.975 91.815 58.640 91.985 ;
        RECT 56.505 90.855 57.025 91.395 ;
        RECT 57.195 91.025 57.715 91.565 ;
        RECT 57.890 90.995 58.240 91.645 ;
        RECT 49.145 90.105 54.490 90.650 ;
        RECT 54.665 90.105 55.875 90.855 ;
        RECT 56.045 90.105 56.335 90.830 ;
        RECT 56.505 90.105 57.715 90.855 ;
        RECT 58.410 90.825 58.640 91.815 ;
        RECT 57.975 90.655 58.640 90.825 ;
        RECT 57.975 90.365 58.145 90.655 ;
        RECT 58.315 90.105 58.645 90.485 ;
        RECT 58.815 90.365 59.000 92.485 ;
        RECT 59.240 92.195 59.505 92.655 ;
        RECT 59.675 92.060 59.925 92.485 ;
        RECT 60.135 92.210 61.240 92.380 ;
        RECT 59.620 91.930 59.925 92.060 ;
        RECT 59.170 90.735 59.450 91.685 ;
        RECT 59.620 90.825 59.790 91.930 ;
        RECT 59.960 91.145 60.200 91.740 ;
        RECT 60.370 91.675 60.900 92.040 ;
        RECT 60.370 90.975 60.540 91.675 ;
        RECT 61.070 91.595 61.240 92.210 ;
        RECT 61.410 91.855 61.580 92.655 ;
        RECT 61.750 92.155 62.000 92.485 ;
        RECT 62.225 92.185 63.110 92.355 ;
        RECT 61.070 91.505 61.580 91.595 ;
        RECT 59.620 90.695 59.845 90.825 ;
        RECT 60.015 90.755 60.540 90.975 ;
        RECT 60.710 91.335 61.580 91.505 ;
        RECT 59.255 90.105 59.505 90.565 ;
        RECT 59.675 90.555 59.845 90.695 ;
        RECT 60.710 90.555 60.880 91.335 ;
        RECT 61.410 91.265 61.580 91.335 ;
        RECT 61.090 91.085 61.290 91.115 ;
        RECT 61.750 91.085 61.920 92.155 ;
        RECT 62.090 91.265 62.280 91.985 ;
        RECT 61.090 90.785 61.920 91.085 ;
        RECT 62.450 91.055 62.770 92.015 ;
        RECT 59.675 90.385 60.010 90.555 ;
        RECT 60.205 90.385 60.880 90.555 ;
        RECT 61.200 90.105 61.570 90.605 ;
        RECT 61.750 90.555 61.920 90.785 ;
        RECT 62.305 90.725 62.770 91.055 ;
        RECT 62.940 91.345 63.110 92.185 ;
        RECT 63.290 92.155 63.605 92.655 ;
        RECT 63.835 91.925 64.175 92.485 ;
        RECT 63.280 91.550 64.175 91.925 ;
        RECT 64.345 91.645 64.515 92.655 ;
        RECT 63.985 91.345 64.175 91.550 ;
        RECT 64.685 91.595 65.015 92.440 ;
        RECT 65.335 91.985 65.505 92.485 ;
        RECT 65.675 92.155 66.005 92.655 ;
        RECT 65.335 91.815 66.000 91.985 ;
        RECT 64.685 91.515 65.075 91.595 ;
        RECT 64.860 91.465 65.075 91.515 ;
        RECT 62.940 91.015 63.815 91.345 ;
        RECT 63.985 91.015 64.735 91.345 ;
        RECT 62.940 90.555 63.110 91.015 ;
        RECT 63.985 90.845 64.185 91.015 ;
        RECT 64.905 90.885 65.075 91.465 ;
        RECT 65.250 90.995 65.600 91.645 ;
        RECT 64.850 90.845 65.075 90.885 ;
        RECT 61.750 90.385 62.155 90.555 ;
        RECT 62.325 90.385 63.110 90.555 ;
        RECT 63.385 90.105 63.595 90.635 ;
        RECT 63.855 90.320 64.185 90.845 ;
        RECT 64.695 90.760 65.075 90.845 ;
        RECT 65.770 90.825 66.000 91.815 ;
        RECT 64.355 90.105 64.525 90.715 ;
        RECT 64.695 90.325 65.025 90.760 ;
        RECT 65.335 90.655 66.000 90.825 ;
        RECT 65.335 90.365 65.505 90.655 ;
        RECT 65.675 90.105 66.005 90.485 ;
        RECT 66.175 90.365 66.360 92.485 ;
        RECT 66.600 92.195 66.865 92.655 ;
        RECT 67.035 92.060 67.285 92.485 ;
        RECT 67.495 92.210 68.600 92.380 ;
        RECT 66.980 91.930 67.285 92.060 ;
        RECT 66.530 90.735 66.810 91.685 ;
        RECT 66.980 90.825 67.150 91.930 ;
        RECT 67.320 91.145 67.560 91.740 ;
        RECT 67.730 91.675 68.260 92.040 ;
        RECT 67.730 90.975 67.900 91.675 ;
        RECT 68.430 91.595 68.600 92.210 ;
        RECT 68.770 91.855 68.940 92.655 ;
        RECT 69.110 92.155 69.360 92.485 ;
        RECT 69.585 92.185 70.470 92.355 ;
        RECT 68.430 91.505 68.940 91.595 ;
        RECT 66.980 90.695 67.205 90.825 ;
        RECT 67.375 90.755 67.900 90.975 ;
        RECT 68.070 91.335 68.940 91.505 ;
        RECT 66.615 90.105 66.865 90.565 ;
        RECT 67.035 90.555 67.205 90.695 ;
        RECT 68.070 90.555 68.240 91.335 ;
        RECT 68.770 91.265 68.940 91.335 ;
        RECT 68.450 91.085 68.650 91.115 ;
        RECT 69.110 91.085 69.280 92.155 ;
        RECT 69.450 91.265 69.640 91.985 ;
        RECT 68.450 90.785 69.280 91.085 ;
        RECT 69.810 91.055 70.130 92.015 ;
        RECT 67.035 90.385 67.370 90.555 ;
        RECT 67.565 90.385 68.240 90.555 ;
        RECT 68.560 90.105 68.930 90.605 ;
        RECT 69.110 90.555 69.280 90.785 ;
        RECT 69.665 90.725 70.130 91.055 ;
        RECT 70.300 91.345 70.470 92.185 ;
        RECT 70.650 92.155 70.965 92.655 ;
        RECT 71.195 91.925 71.535 92.485 ;
        RECT 70.640 91.550 71.535 91.925 ;
        RECT 71.705 91.645 71.875 92.655 ;
        RECT 71.345 91.345 71.535 91.550 ;
        RECT 72.045 91.595 72.375 92.440 ;
        RECT 72.695 91.725 72.865 92.485 ;
        RECT 73.080 91.895 73.410 92.655 ;
        RECT 72.045 91.515 72.435 91.595 ;
        RECT 72.695 91.555 73.410 91.725 ;
        RECT 73.580 91.580 73.835 92.485 ;
        RECT 72.220 91.465 72.435 91.515 ;
        RECT 70.300 91.015 71.175 91.345 ;
        RECT 71.345 91.015 72.095 91.345 ;
        RECT 70.300 90.555 70.470 91.015 ;
        RECT 71.345 90.845 71.545 91.015 ;
        RECT 72.265 90.885 72.435 91.465 ;
        RECT 72.605 91.005 72.960 91.375 ;
        RECT 73.240 91.345 73.410 91.555 ;
        RECT 73.240 91.015 73.495 91.345 ;
        RECT 72.210 90.845 72.435 90.885 ;
        RECT 69.110 90.385 69.515 90.555 ;
        RECT 69.685 90.385 70.470 90.555 ;
        RECT 70.745 90.105 70.955 90.635 ;
        RECT 71.215 90.320 71.545 90.845 ;
        RECT 72.055 90.760 72.435 90.845 ;
        RECT 73.240 90.825 73.410 91.015 ;
        RECT 73.665 90.850 73.835 91.580 ;
        RECT 74.010 91.505 74.270 92.655 ;
        RECT 74.535 91.985 74.705 92.485 ;
        RECT 74.875 92.155 75.205 92.655 ;
        RECT 74.535 91.815 75.200 91.985 ;
        RECT 74.450 90.995 74.800 91.645 ;
        RECT 71.715 90.105 71.885 90.715 ;
        RECT 72.055 90.325 72.385 90.760 ;
        RECT 72.695 90.655 73.410 90.825 ;
        RECT 72.695 90.275 72.865 90.655 ;
        RECT 73.080 90.105 73.410 90.485 ;
        RECT 73.580 90.275 73.835 90.850 ;
        RECT 74.010 90.105 74.270 90.945 ;
        RECT 74.970 90.825 75.200 91.815 ;
        RECT 74.535 90.655 75.200 90.825 ;
        RECT 74.535 90.365 74.705 90.655 ;
        RECT 74.875 90.105 75.205 90.485 ;
        RECT 75.375 90.365 75.560 92.485 ;
        RECT 75.800 92.195 76.065 92.655 ;
        RECT 76.235 92.060 76.485 92.485 ;
        RECT 76.695 92.210 77.800 92.380 ;
        RECT 76.180 91.930 76.485 92.060 ;
        RECT 75.730 90.735 76.010 91.685 ;
        RECT 76.180 90.825 76.350 91.930 ;
        RECT 76.520 91.145 76.760 91.740 ;
        RECT 76.930 91.675 77.460 92.040 ;
        RECT 76.930 90.975 77.100 91.675 ;
        RECT 77.630 91.595 77.800 92.210 ;
        RECT 77.970 91.855 78.140 92.655 ;
        RECT 78.310 92.155 78.560 92.485 ;
        RECT 78.785 92.185 79.670 92.355 ;
        RECT 77.630 91.505 78.140 91.595 ;
        RECT 76.180 90.695 76.405 90.825 ;
        RECT 76.575 90.755 77.100 90.975 ;
        RECT 77.270 91.335 78.140 91.505 ;
        RECT 75.815 90.105 76.065 90.565 ;
        RECT 76.235 90.555 76.405 90.695 ;
        RECT 77.270 90.555 77.440 91.335 ;
        RECT 77.970 91.265 78.140 91.335 ;
        RECT 77.650 91.085 77.850 91.115 ;
        RECT 78.310 91.085 78.480 92.155 ;
        RECT 78.650 91.265 78.840 91.985 ;
        RECT 77.650 90.785 78.480 91.085 ;
        RECT 79.010 91.055 79.330 92.015 ;
        RECT 76.235 90.385 76.570 90.555 ;
        RECT 76.765 90.385 77.440 90.555 ;
        RECT 77.760 90.105 78.130 90.605 ;
        RECT 78.310 90.555 78.480 90.785 ;
        RECT 78.865 90.725 79.330 91.055 ;
        RECT 79.500 91.345 79.670 92.185 ;
        RECT 79.850 92.155 80.165 92.655 ;
        RECT 80.395 91.925 80.735 92.485 ;
        RECT 79.840 91.550 80.735 91.925 ;
        RECT 80.905 91.645 81.075 92.655 ;
        RECT 80.545 91.345 80.735 91.550 ;
        RECT 81.245 91.595 81.575 92.440 ;
        RECT 81.245 91.515 81.635 91.595 ;
        RECT 81.420 91.465 81.635 91.515 ;
        RECT 81.805 91.490 82.095 92.655 ;
        RECT 82.270 92.265 82.605 92.485 ;
        RECT 83.610 92.275 83.965 92.655 ;
        RECT 82.270 91.645 82.525 92.265 ;
        RECT 82.775 92.105 83.005 92.145 ;
        RECT 84.135 92.105 84.385 92.485 ;
        RECT 82.775 91.905 84.385 92.105 ;
        RECT 82.775 91.815 82.960 91.905 ;
        RECT 83.550 91.895 84.385 91.905 ;
        RECT 84.635 91.875 84.885 92.655 ;
        RECT 85.055 91.805 85.315 92.485 ;
        RECT 83.115 91.705 83.445 91.735 ;
        RECT 83.115 91.645 84.915 91.705 ;
        RECT 82.270 91.535 84.975 91.645 ;
        RECT 82.270 91.475 83.445 91.535 ;
        RECT 84.775 91.500 84.975 91.535 ;
        RECT 79.500 91.015 80.375 91.345 ;
        RECT 80.545 91.015 81.295 91.345 ;
        RECT 79.500 90.555 79.670 91.015 ;
        RECT 80.545 90.845 80.745 91.015 ;
        RECT 81.465 90.885 81.635 91.465 ;
        RECT 82.265 91.095 82.755 91.295 ;
        RECT 82.945 91.095 83.420 91.305 ;
        RECT 81.410 90.845 81.635 90.885 ;
        RECT 78.310 90.385 78.715 90.555 ;
        RECT 78.885 90.385 79.670 90.555 ;
        RECT 79.945 90.105 80.155 90.635 ;
        RECT 80.415 90.320 80.745 90.845 ;
        RECT 81.255 90.760 81.635 90.845 ;
        RECT 80.915 90.105 81.085 90.715 ;
        RECT 81.255 90.325 81.585 90.760 ;
        RECT 81.805 90.105 82.095 90.830 ;
        RECT 82.270 90.105 82.725 90.870 ;
        RECT 83.200 90.695 83.420 91.095 ;
        RECT 83.665 91.095 83.995 91.305 ;
        RECT 83.665 90.695 83.875 91.095 ;
        RECT 84.165 91.060 84.575 91.365 ;
        RECT 84.805 90.925 84.975 91.500 ;
        RECT 84.705 90.805 84.975 90.925 ;
        RECT 84.130 90.760 84.975 90.805 ;
        RECT 84.130 90.635 84.885 90.760 ;
        RECT 84.130 90.485 84.300 90.635 ;
        RECT 85.145 90.605 85.315 91.805 ;
        RECT 85.485 91.565 87.155 92.655 ;
        RECT 87.415 91.985 87.585 92.485 ;
        RECT 87.755 92.155 88.085 92.655 ;
        RECT 87.415 91.815 88.080 91.985 ;
        RECT 83.000 90.275 84.300 90.485 ;
        RECT 84.555 90.105 84.885 90.465 ;
        RECT 85.055 90.275 85.315 90.605 ;
        RECT 85.485 90.875 86.235 91.395 ;
        RECT 86.405 91.045 87.155 91.565 ;
        RECT 87.330 90.995 87.680 91.645 ;
        RECT 85.485 90.105 87.155 90.875 ;
        RECT 87.850 90.825 88.080 91.815 ;
        RECT 87.415 90.655 88.080 90.825 ;
        RECT 87.415 90.365 87.585 90.655 ;
        RECT 87.755 90.105 88.085 90.485 ;
        RECT 88.255 90.365 88.440 92.485 ;
        RECT 88.680 92.195 88.945 92.655 ;
        RECT 89.115 92.060 89.365 92.485 ;
        RECT 89.575 92.210 90.680 92.380 ;
        RECT 89.060 91.930 89.365 92.060 ;
        RECT 88.610 90.735 88.890 91.685 ;
        RECT 89.060 90.825 89.230 91.930 ;
        RECT 89.400 91.145 89.640 91.740 ;
        RECT 89.810 91.675 90.340 92.040 ;
        RECT 89.810 90.975 89.980 91.675 ;
        RECT 90.510 91.595 90.680 92.210 ;
        RECT 90.850 91.855 91.020 92.655 ;
        RECT 91.190 92.155 91.440 92.485 ;
        RECT 91.665 92.185 92.550 92.355 ;
        RECT 90.510 91.505 91.020 91.595 ;
        RECT 89.060 90.695 89.285 90.825 ;
        RECT 89.455 90.755 89.980 90.975 ;
        RECT 90.150 91.335 91.020 91.505 ;
        RECT 88.695 90.105 88.945 90.565 ;
        RECT 89.115 90.555 89.285 90.695 ;
        RECT 90.150 90.555 90.320 91.335 ;
        RECT 90.850 91.265 91.020 91.335 ;
        RECT 90.530 91.085 90.730 91.115 ;
        RECT 91.190 91.085 91.360 92.155 ;
        RECT 91.530 91.265 91.720 91.985 ;
        RECT 90.530 90.785 91.360 91.085 ;
        RECT 91.890 91.055 92.210 92.015 ;
        RECT 89.115 90.385 89.450 90.555 ;
        RECT 89.645 90.385 90.320 90.555 ;
        RECT 90.640 90.105 91.010 90.605 ;
        RECT 91.190 90.555 91.360 90.785 ;
        RECT 91.745 90.725 92.210 91.055 ;
        RECT 92.380 91.345 92.550 92.185 ;
        RECT 92.730 92.155 93.045 92.655 ;
        RECT 93.275 91.925 93.615 92.485 ;
        RECT 92.720 91.550 93.615 91.925 ;
        RECT 93.785 91.645 93.955 92.655 ;
        RECT 93.425 91.345 93.615 91.550 ;
        RECT 94.125 91.595 94.455 92.440 ;
        RECT 94.125 91.515 94.515 91.595 ;
        RECT 94.300 91.465 94.515 91.515 ;
        RECT 92.380 91.015 93.255 91.345 ;
        RECT 93.425 91.015 94.175 91.345 ;
        RECT 92.380 90.555 92.550 91.015 ;
        RECT 93.425 90.845 93.625 91.015 ;
        RECT 94.345 90.885 94.515 91.465 ;
        RECT 94.290 90.845 94.515 90.885 ;
        RECT 91.190 90.385 91.595 90.555 ;
        RECT 91.765 90.385 92.550 90.555 ;
        RECT 92.825 90.105 93.035 90.635 ;
        RECT 93.295 90.320 93.625 90.845 ;
        RECT 94.135 90.760 94.515 90.845 ;
        RECT 94.685 91.580 94.955 92.485 ;
        RECT 95.125 91.895 95.455 92.655 ;
        RECT 95.635 91.725 95.815 92.485 ;
        RECT 96.155 91.985 96.325 92.485 ;
        RECT 96.495 92.155 96.825 92.655 ;
        RECT 96.155 91.815 96.820 91.985 ;
        RECT 94.685 90.780 94.865 91.580 ;
        RECT 95.140 91.555 95.815 91.725 ;
        RECT 95.140 91.410 95.310 91.555 ;
        RECT 95.035 91.080 95.310 91.410 ;
        RECT 95.140 90.825 95.310 91.080 ;
        RECT 95.535 91.005 95.875 91.375 ;
        RECT 96.070 90.995 96.420 91.645 ;
        RECT 96.590 90.825 96.820 91.815 ;
        RECT 93.795 90.105 93.965 90.715 ;
        RECT 94.135 90.325 94.465 90.760 ;
        RECT 94.685 90.275 94.945 90.780 ;
        RECT 95.140 90.655 95.805 90.825 ;
        RECT 95.125 90.105 95.455 90.485 ;
        RECT 95.635 90.275 95.805 90.655 ;
        RECT 96.155 90.655 96.820 90.825 ;
        RECT 96.155 90.365 96.325 90.655 ;
        RECT 96.495 90.105 96.825 90.485 ;
        RECT 96.995 90.365 97.180 92.485 ;
        RECT 97.420 92.195 97.685 92.655 ;
        RECT 97.855 92.060 98.105 92.485 ;
        RECT 98.315 92.210 99.420 92.380 ;
        RECT 97.800 91.930 98.105 92.060 ;
        RECT 97.350 90.735 97.630 91.685 ;
        RECT 97.800 90.825 97.970 91.930 ;
        RECT 98.140 91.145 98.380 91.740 ;
        RECT 98.550 91.675 99.080 92.040 ;
        RECT 98.550 90.975 98.720 91.675 ;
        RECT 99.250 91.595 99.420 92.210 ;
        RECT 99.590 91.855 99.760 92.655 ;
        RECT 99.930 92.155 100.180 92.485 ;
        RECT 100.405 92.185 101.290 92.355 ;
        RECT 99.250 91.505 99.760 91.595 ;
        RECT 97.800 90.695 98.025 90.825 ;
        RECT 98.195 90.755 98.720 90.975 ;
        RECT 98.890 91.335 99.760 91.505 ;
        RECT 97.435 90.105 97.685 90.565 ;
        RECT 97.855 90.555 98.025 90.695 ;
        RECT 98.890 90.555 99.060 91.335 ;
        RECT 99.590 91.265 99.760 91.335 ;
        RECT 99.270 91.085 99.470 91.115 ;
        RECT 99.930 91.085 100.100 92.155 ;
        RECT 100.270 91.265 100.460 91.985 ;
        RECT 99.270 90.785 100.100 91.085 ;
        RECT 100.630 91.055 100.950 92.015 ;
        RECT 97.855 90.385 98.190 90.555 ;
        RECT 98.385 90.385 99.060 90.555 ;
        RECT 99.380 90.105 99.750 90.605 ;
        RECT 99.930 90.555 100.100 90.785 ;
        RECT 100.485 90.725 100.950 91.055 ;
        RECT 101.120 91.345 101.290 92.185 ;
        RECT 101.470 92.155 101.785 92.655 ;
        RECT 102.015 91.925 102.355 92.485 ;
        RECT 101.460 91.550 102.355 91.925 ;
        RECT 102.525 91.645 102.695 92.655 ;
        RECT 102.165 91.345 102.355 91.550 ;
        RECT 102.865 91.595 103.195 92.440 ;
        RECT 103.515 91.645 103.685 92.485 ;
        RECT 103.855 92.315 105.025 92.485 ;
        RECT 103.855 91.815 104.185 92.315 ;
        RECT 104.695 92.275 105.025 92.315 ;
        RECT 105.215 92.235 105.570 92.655 ;
        RECT 104.355 92.055 104.585 92.145 ;
        RECT 105.740 92.055 105.990 92.485 ;
        RECT 104.355 91.815 105.990 92.055 ;
        RECT 106.160 91.895 106.490 92.655 ;
        RECT 106.660 91.815 106.915 92.485 ;
        RECT 102.865 91.515 103.255 91.595 ;
        RECT 103.040 91.465 103.255 91.515 ;
        RECT 103.515 91.475 106.575 91.645 ;
        RECT 101.120 91.015 101.995 91.345 ;
        RECT 102.165 91.015 102.915 91.345 ;
        RECT 101.120 90.555 101.290 91.015 ;
        RECT 102.165 90.845 102.365 91.015 ;
        RECT 103.085 90.885 103.255 91.465 ;
        RECT 103.430 91.095 103.780 91.305 ;
        RECT 103.950 91.095 104.395 91.295 ;
        RECT 104.565 91.095 105.040 91.295 ;
        RECT 103.030 90.845 103.255 90.885 ;
        RECT 99.930 90.385 100.335 90.555 ;
        RECT 100.505 90.385 101.290 90.555 ;
        RECT 101.565 90.105 101.775 90.635 ;
        RECT 102.035 90.320 102.365 90.845 ;
        RECT 102.875 90.760 103.255 90.845 ;
        RECT 102.535 90.105 102.705 90.715 ;
        RECT 102.875 90.325 103.205 90.760 ;
        RECT 103.515 90.755 104.580 90.925 ;
        RECT 103.515 90.275 103.685 90.755 ;
        RECT 103.855 90.105 104.185 90.585 ;
        RECT 104.410 90.525 104.580 90.755 ;
        RECT 104.760 90.695 105.040 91.095 ;
        RECT 105.310 91.095 105.640 91.295 ;
        RECT 105.810 91.095 106.175 91.295 ;
        RECT 105.310 90.695 105.595 91.095 ;
        RECT 106.405 90.925 106.575 91.475 ;
        RECT 105.775 90.755 106.575 90.925 ;
        RECT 105.775 90.525 105.945 90.755 ;
        RECT 106.745 90.685 106.915 91.815 ;
        RECT 107.565 91.490 107.855 92.655 ;
        RECT 108.115 91.985 108.285 92.485 ;
        RECT 108.455 92.155 108.785 92.655 ;
        RECT 108.115 91.815 108.780 91.985 ;
        RECT 108.030 90.995 108.380 91.645 ;
        RECT 106.730 90.605 106.915 90.685 ;
        RECT 104.410 90.275 105.945 90.525 ;
        RECT 106.115 90.105 106.445 90.585 ;
        RECT 106.660 90.275 106.915 90.605 ;
        RECT 107.565 90.105 107.855 90.830 ;
        RECT 108.550 90.825 108.780 91.815 ;
        RECT 108.115 90.655 108.780 90.825 ;
        RECT 108.115 90.365 108.285 90.655 ;
        RECT 108.455 90.105 108.785 90.485 ;
        RECT 108.955 90.365 109.140 92.485 ;
        RECT 109.380 92.195 109.645 92.655 ;
        RECT 109.815 92.060 110.065 92.485 ;
        RECT 110.275 92.210 111.380 92.380 ;
        RECT 109.760 91.930 110.065 92.060 ;
        RECT 109.310 90.735 109.590 91.685 ;
        RECT 109.760 90.825 109.930 91.930 ;
        RECT 110.100 91.145 110.340 91.740 ;
        RECT 110.510 91.675 111.040 92.040 ;
        RECT 110.510 90.975 110.680 91.675 ;
        RECT 111.210 91.595 111.380 92.210 ;
        RECT 111.550 91.855 111.720 92.655 ;
        RECT 111.890 92.155 112.140 92.485 ;
        RECT 112.365 92.185 113.250 92.355 ;
        RECT 111.210 91.505 111.720 91.595 ;
        RECT 109.760 90.695 109.985 90.825 ;
        RECT 110.155 90.755 110.680 90.975 ;
        RECT 110.850 91.335 111.720 91.505 ;
        RECT 109.395 90.105 109.645 90.565 ;
        RECT 109.815 90.555 109.985 90.695 ;
        RECT 110.850 90.555 111.020 91.335 ;
        RECT 111.550 91.265 111.720 91.335 ;
        RECT 111.230 91.085 111.430 91.115 ;
        RECT 111.890 91.085 112.060 92.155 ;
        RECT 112.230 91.265 112.420 91.985 ;
        RECT 111.230 90.785 112.060 91.085 ;
        RECT 112.590 91.055 112.910 92.015 ;
        RECT 109.815 90.385 110.150 90.555 ;
        RECT 110.345 90.385 111.020 90.555 ;
        RECT 111.340 90.105 111.710 90.605 ;
        RECT 111.890 90.555 112.060 90.785 ;
        RECT 112.445 90.725 112.910 91.055 ;
        RECT 113.080 91.345 113.250 92.185 ;
        RECT 113.430 92.155 113.745 92.655 ;
        RECT 113.975 91.925 114.315 92.485 ;
        RECT 113.420 91.550 114.315 91.925 ;
        RECT 114.485 91.645 114.655 92.655 ;
        RECT 114.125 91.345 114.315 91.550 ;
        RECT 114.825 91.595 115.155 92.440 ;
        RECT 115.475 91.985 115.645 92.485 ;
        RECT 115.815 92.155 116.145 92.655 ;
        RECT 115.475 91.815 116.140 91.985 ;
        RECT 114.825 91.515 115.215 91.595 ;
        RECT 115.000 91.465 115.215 91.515 ;
        RECT 113.080 91.015 113.955 91.345 ;
        RECT 114.125 91.015 114.875 91.345 ;
        RECT 113.080 90.555 113.250 91.015 ;
        RECT 114.125 90.845 114.325 91.015 ;
        RECT 115.045 90.885 115.215 91.465 ;
        RECT 115.390 90.995 115.740 91.645 ;
        RECT 114.990 90.845 115.215 90.885 ;
        RECT 111.890 90.385 112.295 90.555 ;
        RECT 112.465 90.385 113.250 90.555 ;
        RECT 113.525 90.105 113.735 90.635 ;
        RECT 113.995 90.320 114.325 90.845 ;
        RECT 114.835 90.760 115.215 90.845 ;
        RECT 115.910 90.825 116.140 91.815 ;
        RECT 114.495 90.105 114.665 90.715 ;
        RECT 114.835 90.325 115.165 90.760 ;
        RECT 115.475 90.655 116.140 90.825 ;
        RECT 115.475 90.365 115.645 90.655 ;
        RECT 115.815 90.105 116.145 90.485 ;
        RECT 116.315 90.365 116.500 92.485 ;
        RECT 116.740 92.195 117.005 92.655 ;
        RECT 117.175 92.060 117.425 92.485 ;
        RECT 117.635 92.210 118.740 92.380 ;
        RECT 117.120 91.930 117.425 92.060 ;
        RECT 116.670 90.735 116.950 91.685 ;
        RECT 117.120 90.825 117.290 91.930 ;
        RECT 117.460 91.145 117.700 91.740 ;
        RECT 117.870 91.675 118.400 92.040 ;
        RECT 117.870 90.975 118.040 91.675 ;
        RECT 118.570 91.595 118.740 92.210 ;
        RECT 118.910 91.855 119.080 92.655 ;
        RECT 119.250 92.155 119.500 92.485 ;
        RECT 119.725 92.185 120.610 92.355 ;
        RECT 118.570 91.505 119.080 91.595 ;
        RECT 117.120 90.695 117.345 90.825 ;
        RECT 117.515 90.755 118.040 90.975 ;
        RECT 118.210 91.335 119.080 91.505 ;
        RECT 116.755 90.105 117.005 90.565 ;
        RECT 117.175 90.555 117.345 90.695 ;
        RECT 118.210 90.555 118.380 91.335 ;
        RECT 118.910 91.265 119.080 91.335 ;
        RECT 118.590 91.085 118.790 91.115 ;
        RECT 119.250 91.085 119.420 92.155 ;
        RECT 119.590 91.265 119.780 91.985 ;
        RECT 118.590 90.785 119.420 91.085 ;
        RECT 119.950 91.055 120.270 92.015 ;
        RECT 117.175 90.385 117.510 90.555 ;
        RECT 117.705 90.385 118.380 90.555 ;
        RECT 118.700 90.105 119.070 90.605 ;
        RECT 119.250 90.555 119.420 90.785 ;
        RECT 119.805 90.725 120.270 91.055 ;
        RECT 120.440 91.345 120.610 92.185 ;
        RECT 120.790 92.155 121.105 92.655 ;
        RECT 121.335 91.925 121.675 92.485 ;
        RECT 120.780 91.550 121.675 91.925 ;
        RECT 121.845 91.645 122.015 92.655 ;
        RECT 121.485 91.345 121.675 91.550 ;
        RECT 122.185 91.595 122.515 92.440 ;
        RECT 122.835 91.985 123.005 92.485 ;
        RECT 123.175 92.155 123.505 92.655 ;
        RECT 122.835 91.815 123.500 91.985 ;
        RECT 122.185 91.515 122.575 91.595 ;
        RECT 122.360 91.465 122.575 91.515 ;
        RECT 120.440 91.015 121.315 91.345 ;
        RECT 121.485 91.015 122.235 91.345 ;
        RECT 120.440 90.555 120.610 91.015 ;
        RECT 121.485 90.845 121.685 91.015 ;
        RECT 122.405 90.885 122.575 91.465 ;
        RECT 122.750 90.995 123.100 91.645 ;
        RECT 122.350 90.845 122.575 90.885 ;
        RECT 119.250 90.385 119.655 90.555 ;
        RECT 119.825 90.385 120.610 90.555 ;
        RECT 120.885 90.105 121.095 90.635 ;
        RECT 121.355 90.320 121.685 90.845 ;
        RECT 122.195 90.760 122.575 90.845 ;
        RECT 123.270 90.825 123.500 91.815 ;
        RECT 121.855 90.105 122.025 90.715 ;
        RECT 122.195 90.325 122.525 90.760 ;
        RECT 122.835 90.655 123.500 90.825 ;
        RECT 122.835 90.365 123.005 90.655 ;
        RECT 123.175 90.105 123.505 90.485 ;
        RECT 123.675 90.365 123.860 92.485 ;
        RECT 124.100 92.195 124.365 92.655 ;
        RECT 124.535 92.060 124.785 92.485 ;
        RECT 124.995 92.210 126.100 92.380 ;
        RECT 124.480 91.930 124.785 92.060 ;
        RECT 124.030 90.735 124.310 91.685 ;
        RECT 124.480 90.825 124.650 91.930 ;
        RECT 124.820 91.145 125.060 91.740 ;
        RECT 125.230 91.675 125.760 92.040 ;
        RECT 125.230 90.975 125.400 91.675 ;
        RECT 125.930 91.595 126.100 92.210 ;
        RECT 126.270 91.855 126.440 92.655 ;
        RECT 126.610 92.155 126.860 92.485 ;
        RECT 127.085 92.185 127.970 92.355 ;
        RECT 125.930 91.505 126.440 91.595 ;
        RECT 124.480 90.695 124.705 90.825 ;
        RECT 124.875 90.755 125.400 90.975 ;
        RECT 125.570 91.335 126.440 91.505 ;
        RECT 124.115 90.105 124.365 90.565 ;
        RECT 124.535 90.555 124.705 90.695 ;
        RECT 125.570 90.555 125.740 91.335 ;
        RECT 126.270 91.265 126.440 91.335 ;
        RECT 125.950 91.085 126.150 91.115 ;
        RECT 126.610 91.085 126.780 92.155 ;
        RECT 126.950 91.265 127.140 91.985 ;
        RECT 125.950 90.785 126.780 91.085 ;
        RECT 127.310 91.055 127.630 92.015 ;
        RECT 124.535 90.385 124.870 90.555 ;
        RECT 125.065 90.385 125.740 90.555 ;
        RECT 126.060 90.105 126.430 90.605 ;
        RECT 126.610 90.555 126.780 90.785 ;
        RECT 127.165 90.725 127.630 91.055 ;
        RECT 127.800 91.345 127.970 92.185 ;
        RECT 128.150 92.155 128.465 92.655 ;
        RECT 128.695 91.925 129.035 92.485 ;
        RECT 128.140 91.550 129.035 91.925 ;
        RECT 129.205 91.645 129.375 92.655 ;
        RECT 128.845 91.345 129.035 91.550 ;
        RECT 129.545 91.595 129.875 92.440 ;
        RECT 130.125 91.600 130.430 92.385 ;
        RECT 130.610 92.185 131.295 92.655 ;
        RECT 130.605 91.665 131.300 91.975 ;
        RECT 129.545 91.515 129.935 91.595 ;
        RECT 129.720 91.465 129.935 91.515 ;
        RECT 127.800 91.015 128.675 91.345 ;
        RECT 128.845 91.015 129.595 91.345 ;
        RECT 127.800 90.555 127.970 91.015 ;
        RECT 128.845 90.845 129.045 91.015 ;
        RECT 129.765 90.885 129.935 91.465 ;
        RECT 129.710 90.845 129.935 90.885 ;
        RECT 126.610 90.385 127.015 90.555 ;
        RECT 127.185 90.385 127.970 90.555 ;
        RECT 128.245 90.105 128.455 90.635 ;
        RECT 128.715 90.320 129.045 90.845 ;
        RECT 129.555 90.760 129.935 90.845 ;
        RECT 130.125 90.795 130.300 91.600 ;
        RECT 131.475 91.495 131.760 92.440 ;
        RECT 131.935 92.205 132.265 92.655 ;
        RECT 132.435 92.035 132.605 92.465 ;
        RECT 130.900 91.345 131.760 91.495 ;
        RECT 130.475 91.325 131.760 91.345 ;
        RECT 131.930 91.805 132.605 92.035 ;
        RECT 130.475 90.965 131.460 91.325 ;
        RECT 131.930 91.155 132.165 91.805 ;
        RECT 129.215 90.105 129.385 90.715 ;
        RECT 129.555 90.325 129.885 90.760 ;
        RECT 130.125 90.275 130.365 90.795 ;
        RECT 131.290 90.630 131.460 90.965 ;
        RECT 131.630 90.825 132.165 91.155 ;
        RECT 131.945 90.675 132.165 90.825 ;
        RECT 132.335 90.785 132.635 91.635 ;
        RECT 133.325 91.490 133.615 92.655 ;
        RECT 134.335 91.985 134.505 92.485 ;
        RECT 134.675 92.155 135.005 92.655 ;
        RECT 134.335 91.815 135.000 91.985 ;
        RECT 134.250 90.995 134.600 91.645 ;
        RECT 130.535 90.105 130.930 90.600 ;
        RECT 131.290 90.435 131.665 90.630 ;
        RECT 131.495 90.290 131.665 90.435 ;
        RECT 131.945 90.300 132.185 90.675 ;
        RECT 132.355 90.105 132.690 90.610 ;
        RECT 133.325 90.105 133.615 90.830 ;
        RECT 134.770 90.825 135.000 91.815 ;
        RECT 134.335 90.655 135.000 90.825 ;
        RECT 134.335 90.365 134.505 90.655 ;
        RECT 134.675 90.105 135.005 90.485 ;
        RECT 135.175 90.365 135.360 92.485 ;
        RECT 135.600 92.195 135.865 92.655 ;
        RECT 136.035 92.060 136.285 92.485 ;
        RECT 136.495 92.210 137.600 92.380 ;
        RECT 135.980 91.930 136.285 92.060 ;
        RECT 135.530 90.735 135.810 91.685 ;
        RECT 135.980 90.825 136.150 91.930 ;
        RECT 136.320 91.145 136.560 91.740 ;
        RECT 136.730 91.675 137.260 92.040 ;
        RECT 136.730 90.975 136.900 91.675 ;
        RECT 137.430 91.595 137.600 92.210 ;
        RECT 137.770 91.855 137.940 92.655 ;
        RECT 138.110 92.155 138.360 92.485 ;
        RECT 138.585 92.185 139.470 92.355 ;
        RECT 137.430 91.505 137.940 91.595 ;
        RECT 135.980 90.695 136.205 90.825 ;
        RECT 136.375 90.755 136.900 90.975 ;
        RECT 137.070 91.335 137.940 91.505 ;
        RECT 135.615 90.105 135.865 90.565 ;
        RECT 136.035 90.555 136.205 90.695 ;
        RECT 137.070 90.555 137.240 91.335 ;
        RECT 137.770 91.265 137.940 91.335 ;
        RECT 137.450 91.085 137.650 91.115 ;
        RECT 138.110 91.085 138.280 92.155 ;
        RECT 138.450 91.265 138.640 91.985 ;
        RECT 137.450 90.785 138.280 91.085 ;
        RECT 138.810 91.055 139.130 92.015 ;
        RECT 136.035 90.385 136.370 90.555 ;
        RECT 136.565 90.385 137.240 90.555 ;
        RECT 137.560 90.105 137.930 90.605 ;
        RECT 138.110 90.555 138.280 90.785 ;
        RECT 138.665 90.725 139.130 91.055 ;
        RECT 139.300 91.345 139.470 92.185 ;
        RECT 139.650 92.155 139.965 92.655 ;
        RECT 140.195 91.925 140.535 92.485 ;
        RECT 139.640 91.550 140.535 91.925 ;
        RECT 140.705 91.645 140.875 92.655 ;
        RECT 140.345 91.345 140.535 91.550 ;
        RECT 141.045 91.595 141.375 92.440 ;
        RECT 141.045 91.515 141.435 91.595 ;
        RECT 141.220 91.465 141.435 91.515 ;
        RECT 139.300 91.015 140.175 91.345 ;
        RECT 140.345 91.015 141.095 91.345 ;
        RECT 139.300 90.555 139.470 91.015 ;
        RECT 140.345 90.845 140.545 91.015 ;
        RECT 141.265 90.885 141.435 91.465 ;
        RECT 141.210 90.845 141.435 90.885 ;
        RECT 138.110 90.385 138.515 90.555 ;
        RECT 138.685 90.385 139.470 90.555 ;
        RECT 139.745 90.105 139.955 90.635 ;
        RECT 140.215 90.320 140.545 90.845 ;
        RECT 141.055 90.760 141.435 90.845 ;
        RECT 141.610 91.515 141.945 92.485 ;
        RECT 142.115 91.515 142.285 92.655 ;
        RECT 142.455 92.315 144.485 92.485 ;
        RECT 141.610 90.845 141.780 91.515 ;
        RECT 142.455 91.345 142.625 92.315 ;
        RECT 141.950 91.015 142.205 91.345 ;
        RECT 142.430 91.015 142.625 91.345 ;
        RECT 142.795 91.975 143.920 92.145 ;
        RECT 142.035 90.845 142.205 91.015 ;
        RECT 142.795 90.845 142.965 91.975 ;
        RECT 140.715 90.105 140.885 90.715 ;
        RECT 141.055 90.325 141.385 90.760 ;
        RECT 141.610 90.275 141.865 90.845 ;
        RECT 142.035 90.675 142.965 90.845 ;
        RECT 143.135 91.635 144.145 91.805 ;
        RECT 143.135 90.835 143.305 91.635 ;
        RECT 143.510 90.955 143.785 91.435 ;
        RECT 143.505 90.785 143.785 90.955 ;
        RECT 142.790 90.640 142.965 90.675 ;
        RECT 142.035 90.105 142.365 90.505 ;
        RECT 142.790 90.275 143.320 90.640 ;
        RECT 143.510 90.275 143.785 90.785 ;
        RECT 143.955 90.275 144.145 91.635 ;
        RECT 144.315 91.650 144.485 92.315 ;
        RECT 144.655 91.895 144.825 92.655 ;
        RECT 145.060 91.895 145.575 92.305 ;
        RECT 144.315 91.460 145.065 91.650 ;
        RECT 145.235 91.085 145.575 91.895 ;
        RECT 144.345 90.915 145.575 91.085 ;
        RECT 145.745 91.565 146.955 92.655 ;
        RECT 145.745 91.025 146.265 91.565 ;
        RECT 144.325 90.105 144.835 90.640 ;
        RECT 145.055 90.310 145.300 90.915 ;
        RECT 146.435 90.855 146.955 91.395 ;
        RECT 145.745 90.105 146.955 90.855 ;
        RECT 17.320 89.935 147.040 90.105 ;
        RECT 17.405 89.185 18.615 89.935 ;
        RECT 19.295 89.280 19.625 89.715 ;
        RECT 19.795 89.325 19.965 89.935 ;
        RECT 19.245 89.195 19.625 89.280 ;
        RECT 20.135 89.195 20.465 89.720 ;
        RECT 20.725 89.405 20.935 89.935 ;
        RECT 21.210 89.485 21.995 89.655 ;
        RECT 22.165 89.485 22.570 89.655 ;
        RECT 17.405 88.645 17.925 89.185 ;
        RECT 19.245 89.155 19.470 89.195 ;
        RECT 18.095 88.475 18.615 89.015 ;
        RECT 17.405 87.385 18.615 88.475 ;
        RECT 19.245 88.575 19.415 89.155 ;
        RECT 20.135 89.025 20.335 89.195 ;
        RECT 21.210 89.025 21.380 89.485 ;
        RECT 19.585 88.695 20.335 89.025 ;
        RECT 20.505 88.695 21.380 89.025 ;
        RECT 19.245 88.525 19.460 88.575 ;
        RECT 19.245 88.445 19.635 88.525 ;
        RECT 19.305 87.600 19.635 88.445 ;
        RECT 20.145 88.490 20.335 88.695 ;
        RECT 19.805 87.385 19.975 88.395 ;
        RECT 20.145 88.115 21.040 88.490 ;
        RECT 20.145 87.555 20.485 88.115 ;
        RECT 20.715 87.385 21.030 87.885 ;
        RECT 21.210 87.855 21.380 88.695 ;
        RECT 21.550 88.985 22.015 89.315 ;
        RECT 22.400 89.255 22.570 89.485 ;
        RECT 22.750 89.435 23.120 89.935 ;
        RECT 23.440 89.485 24.115 89.655 ;
        RECT 24.310 89.485 24.645 89.655 ;
        RECT 21.550 88.025 21.870 88.985 ;
        RECT 22.400 88.955 23.230 89.255 ;
        RECT 22.040 88.055 22.230 88.775 ;
        RECT 22.400 87.885 22.570 88.955 ;
        RECT 23.030 88.925 23.230 88.955 ;
        RECT 22.740 88.705 22.910 88.775 ;
        RECT 23.440 88.705 23.610 89.485 ;
        RECT 24.475 89.345 24.645 89.485 ;
        RECT 24.815 89.475 25.065 89.935 ;
        RECT 22.740 88.535 23.610 88.705 ;
        RECT 23.780 89.065 24.305 89.285 ;
        RECT 24.475 89.215 24.700 89.345 ;
        RECT 22.740 88.445 23.250 88.535 ;
        RECT 21.210 87.685 22.095 87.855 ;
        RECT 22.320 87.555 22.570 87.885 ;
        RECT 22.740 87.385 22.910 88.185 ;
        RECT 23.080 87.830 23.250 88.445 ;
        RECT 23.780 88.365 23.950 89.065 ;
        RECT 23.420 88.000 23.950 88.365 ;
        RECT 24.120 88.300 24.360 88.895 ;
        RECT 24.530 88.110 24.700 89.215 ;
        RECT 24.870 88.355 25.150 89.305 ;
        RECT 24.395 87.980 24.700 88.110 ;
        RECT 23.080 87.660 24.185 87.830 ;
        RECT 24.395 87.555 24.645 87.980 ;
        RECT 24.815 87.385 25.080 87.845 ;
        RECT 25.320 87.555 25.505 89.675 ;
        RECT 25.675 89.555 26.005 89.935 ;
        RECT 26.175 89.385 26.345 89.675 ;
        RECT 25.680 89.215 26.345 89.385 ;
        RECT 25.680 88.225 25.910 89.215 ;
        RECT 26.610 89.195 26.865 89.765 ;
        RECT 27.035 89.535 27.365 89.935 ;
        RECT 27.790 89.400 28.320 89.765 ;
        RECT 28.510 89.595 28.785 89.765 ;
        RECT 28.505 89.425 28.785 89.595 ;
        RECT 27.790 89.365 27.965 89.400 ;
        RECT 27.035 89.195 27.965 89.365 ;
        RECT 26.080 88.395 26.430 89.045 ;
        RECT 26.610 88.525 26.780 89.195 ;
        RECT 27.035 89.025 27.205 89.195 ;
        RECT 26.950 88.695 27.205 89.025 ;
        RECT 27.430 88.695 27.625 89.025 ;
        RECT 25.680 88.055 26.345 88.225 ;
        RECT 25.675 87.385 26.005 87.885 ;
        RECT 26.175 87.555 26.345 88.055 ;
        RECT 26.610 87.555 26.945 88.525 ;
        RECT 27.115 87.385 27.285 88.525 ;
        RECT 27.455 87.725 27.625 88.695 ;
        RECT 27.795 88.065 27.965 89.195 ;
        RECT 28.135 88.405 28.305 89.205 ;
        RECT 28.510 88.605 28.785 89.425 ;
        RECT 28.955 88.405 29.145 89.765 ;
        RECT 29.325 89.400 29.835 89.935 ;
        RECT 30.055 89.125 30.300 89.730 ;
        RECT 31.675 89.210 32.005 89.720 ;
        RECT 32.175 89.535 32.505 89.935 ;
        RECT 33.555 89.365 33.885 89.705 ;
        RECT 34.055 89.535 34.385 89.935 ;
        RECT 29.345 88.955 30.575 89.125 ;
        RECT 28.135 88.235 29.145 88.405 ;
        RECT 29.315 88.390 30.065 88.580 ;
        RECT 27.795 87.895 28.920 88.065 ;
        RECT 29.315 87.725 29.485 88.390 ;
        RECT 30.235 88.145 30.575 88.955 ;
        RECT 27.455 87.555 29.485 87.725 ;
        RECT 29.655 87.385 29.825 88.145 ;
        RECT 30.060 87.735 30.575 88.145 ;
        RECT 31.675 88.445 31.865 89.210 ;
        RECT 32.175 89.195 34.540 89.365 ;
        RECT 32.175 89.025 32.345 89.195 ;
        RECT 32.035 88.695 32.345 89.025 ;
        RECT 32.515 88.695 32.820 89.025 ;
        RECT 31.675 87.595 32.005 88.445 ;
        RECT 32.175 87.385 32.425 88.525 ;
        RECT 32.605 88.365 32.820 88.695 ;
        RECT 32.995 88.365 33.280 89.025 ;
        RECT 33.475 88.365 33.740 89.025 ;
        RECT 33.955 88.365 34.200 89.025 ;
        RECT 34.370 88.195 34.540 89.195 ;
        RECT 32.615 88.025 33.905 88.195 ;
        RECT 32.615 87.605 32.865 88.025 ;
        RECT 33.095 87.385 33.425 87.855 ;
        RECT 33.655 87.605 33.905 88.025 ;
        RECT 34.085 88.025 34.540 88.195 ;
        RECT 34.885 89.195 35.245 89.570 ;
        RECT 35.510 89.195 35.680 89.935 ;
        RECT 35.960 89.365 36.130 89.570 ;
        RECT 35.960 89.195 36.500 89.365 ;
        RECT 34.885 88.540 35.140 89.195 ;
        RECT 35.310 88.695 35.660 89.025 ;
        RECT 35.830 88.695 36.160 89.025 ;
        RECT 34.085 87.595 34.415 88.025 ;
        RECT 34.885 87.555 35.225 88.540 ;
        RECT 35.395 88.155 35.660 88.695 ;
        RECT 36.330 88.495 36.500 89.195 ;
        RECT 35.875 88.325 36.500 88.495 ;
        RECT 36.670 88.565 36.840 89.765 ;
        RECT 37.070 89.285 37.400 89.765 ;
        RECT 37.570 89.465 37.740 89.935 ;
        RECT 37.910 89.285 38.240 89.750 ;
        RECT 37.070 89.115 38.240 89.285 ;
        RECT 38.565 89.260 38.835 89.605 ;
        RECT 39.025 89.535 39.405 89.935 ;
        RECT 39.575 89.365 39.745 89.715 ;
        RECT 39.915 89.535 40.245 89.935 ;
        RECT 40.445 89.365 40.615 89.715 ;
        RECT 40.815 89.435 41.145 89.935 ;
        RECT 37.010 88.735 37.580 88.945 ;
        RECT 37.750 88.735 38.395 88.945 ;
        RECT 36.670 88.155 37.375 88.565 ;
        RECT 38.565 88.525 38.735 89.260 ;
        RECT 39.005 89.195 40.615 89.365 ;
        RECT 39.005 89.025 39.175 89.195 ;
        RECT 38.905 88.695 39.175 89.025 ;
        RECT 39.345 88.695 39.750 89.025 ;
        RECT 39.005 88.525 39.175 88.695 ;
        RECT 35.395 87.985 37.375 88.155 ;
        RECT 35.395 87.385 35.805 87.815 ;
        RECT 36.550 87.385 36.880 87.805 ;
        RECT 37.050 87.555 37.375 87.985 ;
        RECT 37.850 87.385 38.180 88.485 ;
        RECT 38.565 87.555 38.835 88.525 ;
        RECT 39.005 88.355 39.730 88.525 ;
        RECT 39.920 88.405 40.630 89.025 ;
        RECT 40.800 88.695 41.150 89.265 ;
        RECT 41.345 89.125 41.585 89.935 ;
        RECT 41.755 89.125 42.085 89.765 ;
        RECT 42.255 89.125 42.525 89.935 ;
        RECT 43.165 89.210 43.455 89.935 ;
        RECT 41.325 88.695 41.675 88.945 ;
        RECT 41.845 88.525 42.015 89.125 ;
        RECT 43.625 88.990 43.965 89.765 ;
        RECT 44.135 89.475 44.305 89.935 ;
        RECT 44.545 89.500 44.905 89.765 ;
        RECT 44.545 89.495 44.900 89.500 ;
        RECT 44.545 89.485 44.895 89.495 ;
        RECT 44.545 89.480 44.890 89.485 ;
        RECT 44.545 89.470 44.885 89.480 ;
        RECT 45.535 89.475 45.705 89.935 ;
        RECT 44.545 89.465 44.880 89.470 ;
        RECT 44.545 89.455 44.870 89.465 ;
        RECT 44.545 89.445 44.860 89.455 ;
        RECT 44.545 89.305 44.845 89.445 ;
        RECT 44.135 89.115 44.845 89.305 ;
        RECT 45.035 89.305 45.365 89.385 ;
        RECT 45.875 89.305 46.215 89.765 ;
        RECT 46.385 89.390 51.730 89.935 ;
        RECT 51.905 89.390 57.250 89.935 ;
        RECT 45.035 89.115 46.215 89.305 ;
        RECT 42.185 88.695 42.535 88.945 ;
        RECT 39.560 88.235 39.730 88.355 ;
        RECT 40.830 88.235 41.150 88.525 ;
        RECT 39.045 87.385 39.325 88.185 ;
        RECT 39.560 88.065 41.150 88.235 ;
        RECT 41.335 88.355 42.015 88.525 ;
        RECT 39.495 87.605 41.150 87.895 ;
        RECT 41.335 87.570 41.665 88.355 ;
        RECT 42.195 87.385 42.525 88.525 ;
        RECT 43.165 87.385 43.455 88.550 ;
        RECT 43.625 87.555 43.905 88.990 ;
        RECT 44.135 88.545 44.420 89.115 ;
        RECT 44.605 88.715 45.075 88.945 ;
        RECT 45.245 88.925 45.575 88.945 ;
        RECT 45.245 88.745 45.695 88.925 ;
        RECT 45.885 88.745 46.215 88.945 ;
        RECT 44.135 88.330 45.285 88.545 ;
        RECT 44.075 87.385 44.785 88.160 ;
        RECT 44.955 87.555 45.285 88.330 ;
        RECT 45.480 87.630 45.695 88.745 ;
        RECT 45.985 88.405 46.215 88.745 ;
        RECT 47.970 88.560 48.310 89.390 ;
        RECT 45.875 87.385 46.205 88.105 ;
        RECT 49.790 87.820 50.140 89.070 ;
        RECT 53.490 88.560 53.830 89.390 ;
        RECT 57.425 89.260 57.685 89.765 ;
        RECT 57.865 89.555 58.195 89.935 ;
        RECT 58.375 89.385 58.545 89.765 ;
        RECT 55.310 87.820 55.660 89.070 ;
        RECT 57.425 88.460 57.595 89.260 ;
        RECT 57.880 89.215 58.545 89.385 ;
        RECT 57.880 88.960 58.050 89.215 ;
        RECT 58.805 89.165 60.475 89.935 ;
        RECT 60.735 89.385 60.905 89.675 ;
        RECT 61.075 89.555 61.405 89.935 ;
        RECT 60.735 89.215 61.400 89.385 ;
        RECT 57.765 88.630 58.050 88.960 ;
        RECT 58.285 88.665 58.615 89.035 ;
        RECT 58.805 88.645 59.555 89.165 ;
        RECT 57.880 88.485 58.050 88.630 ;
        RECT 46.385 87.385 51.730 87.820 ;
        RECT 51.905 87.385 57.250 87.820 ;
        RECT 57.425 87.555 57.695 88.460 ;
        RECT 57.880 88.315 58.545 88.485 ;
        RECT 59.725 88.475 60.475 88.995 ;
        RECT 57.865 87.385 58.195 88.145 ;
        RECT 58.375 87.555 58.545 88.315 ;
        RECT 58.805 87.385 60.475 88.475 ;
        RECT 60.650 88.395 61.000 89.045 ;
        RECT 61.170 88.225 61.400 89.215 ;
        RECT 60.735 88.055 61.400 88.225 ;
        RECT 60.735 87.555 60.905 88.055 ;
        RECT 61.075 87.385 61.405 87.885 ;
        RECT 61.575 87.555 61.760 89.675 ;
        RECT 62.015 89.475 62.265 89.935 ;
        RECT 62.435 89.485 62.770 89.655 ;
        RECT 62.965 89.485 63.640 89.655 ;
        RECT 62.435 89.345 62.605 89.485 ;
        RECT 61.930 88.355 62.210 89.305 ;
        RECT 62.380 89.215 62.605 89.345 ;
        RECT 62.380 88.110 62.550 89.215 ;
        RECT 62.775 89.065 63.300 89.285 ;
        RECT 62.720 88.300 62.960 88.895 ;
        RECT 63.130 88.365 63.300 89.065 ;
        RECT 63.470 88.705 63.640 89.485 ;
        RECT 63.960 89.435 64.330 89.935 ;
        RECT 64.510 89.485 64.915 89.655 ;
        RECT 65.085 89.485 65.870 89.655 ;
        RECT 64.510 89.255 64.680 89.485 ;
        RECT 63.850 88.955 64.680 89.255 ;
        RECT 65.065 88.985 65.530 89.315 ;
        RECT 63.850 88.925 64.050 88.955 ;
        RECT 64.170 88.705 64.340 88.775 ;
        RECT 63.470 88.535 64.340 88.705 ;
        RECT 63.830 88.445 64.340 88.535 ;
        RECT 62.380 87.980 62.685 88.110 ;
        RECT 63.130 88.000 63.660 88.365 ;
        RECT 62.000 87.385 62.265 87.845 ;
        RECT 62.435 87.555 62.685 87.980 ;
        RECT 63.830 87.830 64.000 88.445 ;
        RECT 62.895 87.660 64.000 87.830 ;
        RECT 64.170 87.385 64.340 88.185 ;
        RECT 64.510 87.885 64.680 88.955 ;
        RECT 64.850 88.055 65.040 88.775 ;
        RECT 65.210 88.025 65.530 88.985 ;
        RECT 65.700 89.025 65.870 89.485 ;
        RECT 66.145 89.405 66.355 89.935 ;
        RECT 66.615 89.195 66.945 89.720 ;
        RECT 67.115 89.325 67.285 89.935 ;
        RECT 67.455 89.280 67.785 89.715 ;
        RECT 67.455 89.195 67.835 89.280 ;
        RECT 68.925 89.210 69.215 89.935 ;
        RECT 66.745 89.025 66.945 89.195 ;
        RECT 67.610 89.155 67.835 89.195 ;
        RECT 65.700 88.695 66.575 89.025 ;
        RECT 66.745 88.695 67.495 89.025 ;
        RECT 64.510 87.555 64.760 87.885 ;
        RECT 65.700 87.855 65.870 88.695 ;
        RECT 66.745 88.490 66.935 88.695 ;
        RECT 67.665 88.575 67.835 89.155 ;
        RECT 67.620 88.525 67.835 88.575 ;
        RECT 69.390 89.195 69.645 89.765 ;
        RECT 69.815 89.535 70.145 89.935 ;
        RECT 70.570 89.400 71.100 89.765 ;
        RECT 70.570 89.365 70.745 89.400 ;
        RECT 69.815 89.195 70.745 89.365 ;
        RECT 66.040 88.115 66.935 88.490 ;
        RECT 67.445 88.445 67.835 88.525 ;
        RECT 64.985 87.685 65.870 87.855 ;
        RECT 66.050 87.385 66.365 87.885 ;
        RECT 66.595 87.555 66.935 88.115 ;
        RECT 67.105 87.385 67.275 88.395 ;
        RECT 67.445 87.600 67.775 88.445 ;
        RECT 68.925 87.385 69.215 88.550 ;
        RECT 69.390 88.525 69.560 89.195 ;
        RECT 69.815 89.025 69.985 89.195 ;
        RECT 69.730 88.695 69.985 89.025 ;
        RECT 70.210 88.695 70.405 89.025 ;
        RECT 69.390 87.555 69.725 88.525 ;
        RECT 69.895 87.385 70.065 88.525 ;
        RECT 70.235 87.725 70.405 88.695 ;
        RECT 70.575 88.065 70.745 89.195 ;
        RECT 70.915 88.405 71.085 89.205 ;
        RECT 71.290 88.915 71.565 89.765 ;
        RECT 71.285 88.745 71.565 88.915 ;
        RECT 71.290 88.605 71.565 88.745 ;
        RECT 71.735 88.405 71.925 89.765 ;
        RECT 72.105 89.400 72.615 89.935 ;
        RECT 72.835 89.125 73.080 89.730 ;
        RECT 73.530 89.170 73.985 89.935 ;
        RECT 74.260 89.555 75.560 89.765 ;
        RECT 75.815 89.575 76.145 89.935 ;
        RECT 75.390 89.405 75.560 89.555 ;
        RECT 76.315 89.435 76.575 89.765 ;
        RECT 76.345 89.425 76.575 89.435 ;
        RECT 72.125 88.955 73.355 89.125 ;
        RECT 70.915 88.235 71.925 88.405 ;
        RECT 72.095 88.390 72.845 88.580 ;
        RECT 70.575 87.895 71.700 88.065 ;
        RECT 72.095 87.725 72.265 88.390 ;
        RECT 73.015 88.145 73.355 88.955 ;
        RECT 74.460 88.945 74.680 89.345 ;
        RECT 73.525 88.745 74.015 88.945 ;
        RECT 74.205 88.735 74.680 88.945 ;
        RECT 74.925 88.945 75.135 89.345 ;
        RECT 75.390 89.280 76.145 89.405 ;
        RECT 75.390 89.235 76.235 89.280 ;
        RECT 75.965 89.115 76.235 89.235 ;
        RECT 74.925 88.735 75.255 88.945 ;
        RECT 75.425 88.675 75.835 88.980 ;
        RECT 70.235 87.555 72.265 87.725 ;
        RECT 72.435 87.385 72.605 88.145 ;
        RECT 72.840 87.735 73.355 88.145 ;
        RECT 73.530 88.505 74.705 88.565 ;
        RECT 76.065 88.540 76.235 89.115 ;
        RECT 76.035 88.505 76.235 88.540 ;
        RECT 73.530 88.395 76.235 88.505 ;
        RECT 73.530 87.775 73.785 88.395 ;
        RECT 74.375 88.335 76.175 88.395 ;
        RECT 74.375 88.305 74.705 88.335 ;
        RECT 76.405 88.235 76.575 89.425 ;
        RECT 76.745 89.390 82.090 89.935 ;
        RECT 78.330 88.560 78.670 89.390 ;
        RECT 82.265 89.185 83.475 89.935 ;
        RECT 83.735 89.385 83.905 89.675 ;
        RECT 84.075 89.555 84.405 89.935 ;
        RECT 83.735 89.215 84.400 89.385 ;
        RECT 74.035 88.135 74.220 88.225 ;
        RECT 74.810 88.135 75.645 88.145 ;
        RECT 74.035 87.935 75.645 88.135 ;
        RECT 74.035 87.895 74.265 87.935 ;
        RECT 73.530 87.555 73.865 87.775 ;
        RECT 74.870 87.385 75.225 87.765 ;
        RECT 75.395 87.555 75.645 87.935 ;
        RECT 75.895 87.385 76.145 88.165 ;
        RECT 76.315 87.555 76.575 88.235 ;
        RECT 80.150 87.820 80.500 89.070 ;
        RECT 82.265 88.645 82.785 89.185 ;
        RECT 82.955 88.475 83.475 89.015 ;
        RECT 76.745 87.385 82.090 87.820 ;
        RECT 82.265 87.385 83.475 88.475 ;
        RECT 83.650 88.395 84.000 89.045 ;
        RECT 84.170 88.225 84.400 89.215 ;
        RECT 83.735 88.055 84.400 88.225 ;
        RECT 83.735 87.555 83.905 88.055 ;
        RECT 84.075 87.385 84.405 87.885 ;
        RECT 84.575 87.555 84.760 89.675 ;
        RECT 85.015 89.475 85.265 89.935 ;
        RECT 85.435 89.485 85.770 89.655 ;
        RECT 85.965 89.485 86.640 89.655 ;
        RECT 85.435 89.345 85.605 89.485 ;
        RECT 84.930 88.355 85.210 89.305 ;
        RECT 85.380 89.215 85.605 89.345 ;
        RECT 85.380 88.110 85.550 89.215 ;
        RECT 85.775 89.065 86.300 89.285 ;
        RECT 85.720 88.300 85.960 88.895 ;
        RECT 86.130 88.365 86.300 89.065 ;
        RECT 86.470 88.705 86.640 89.485 ;
        RECT 86.960 89.435 87.330 89.935 ;
        RECT 87.510 89.485 87.915 89.655 ;
        RECT 88.085 89.485 88.870 89.655 ;
        RECT 87.510 89.255 87.680 89.485 ;
        RECT 86.850 88.955 87.680 89.255 ;
        RECT 88.065 88.985 88.530 89.315 ;
        RECT 86.850 88.925 87.050 88.955 ;
        RECT 87.170 88.705 87.340 88.775 ;
        RECT 86.470 88.535 87.340 88.705 ;
        RECT 86.830 88.445 87.340 88.535 ;
        RECT 85.380 87.980 85.685 88.110 ;
        RECT 86.130 88.000 86.660 88.365 ;
        RECT 85.000 87.385 85.265 87.845 ;
        RECT 85.435 87.555 85.685 87.980 ;
        RECT 86.830 87.830 87.000 88.445 ;
        RECT 85.895 87.660 87.000 87.830 ;
        RECT 87.170 87.385 87.340 88.185 ;
        RECT 87.510 87.885 87.680 88.955 ;
        RECT 87.850 88.055 88.040 88.775 ;
        RECT 88.210 88.025 88.530 88.985 ;
        RECT 88.700 89.025 88.870 89.485 ;
        RECT 89.145 89.405 89.355 89.935 ;
        RECT 89.615 89.195 89.945 89.720 ;
        RECT 90.115 89.325 90.285 89.935 ;
        RECT 90.455 89.280 90.785 89.715 ;
        RECT 91.095 89.285 91.265 89.765 ;
        RECT 91.435 89.455 91.765 89.935 ;
        RECT 91.990 89.515 93.525 89.765 ;
        RECT 91.990 89.285 92.160 89.515 ;
        RECT 90.455 89.195 90.835 89.280 ;
        RECT 89.745 89.025 89.945 89.195 ;
        RECT 90.610 89.155 90.835 89.195 ;
        RECT 88.700 88.695 89.575 89.025 ;
        RECT 89.745 88.695 90.495 89.025 ;
        RECT 87.510 87.555 87.760 87.885 ;
        RECT 88.700 87.855 88.870 88.695 ;
        RECT 89.745 88.490 89.935 88.695 ;
        RECT 90.665 88.575 90.835 89.155 ;
        RECT 91.095 89.115 92.160 89.285 ;
        RECT 92.340 88.945 92.620 89.345 ;
        RECT 91.010 88.735 91.360 88.945 ;
        RECT 91.530 88.745 91.975 88.945 ;
        RECT 92.145 88.745 92.620 88.945 ;
        RECT 92.890 88.945 93.175 89.345 ;
        RECT 93.355 89.285 93.525 89.515 ;
        RECT 93.695 89.455 94.025 89.935 ;
        RECT 94.240 89.435 94.495 89.765 ;
        RECT 94.285 89.425 94.495 89.435 ;
        RECT 94.310 89.355 94.495 89.425 ;
        RECT 93.355 89.115 94.155 89.285 ;
        RECT 92.890 88.745 93.220 88.945 ;
        RECT 93.390 88.745 93.755 88.945 ;
        RECT 90.620 88.525 90.835 88.575 ;
        RECT 93.985 88.565 94.155 89.115 ;
        RECT 89.040 88.115 89.935 88.490 ;
        RECT 90.445 88.445 90.835 88.525 ;
        RECT 87.985 87.685 88.870 87.855 ;
        RECT 89.050 87.385 89.365 87.885 ;
        RECT 89.595 87.555 89.935 88.115 ;
        RECT 90.105 87.385 90.275 88.395 ;
        RECT 90.445 87.600 90.775 88.445 ;
        RECT 91.095 88.395 94.155 88.565 ;
        RECT 91.095 87.555 91.265 88.395 ;
        RECT 94.325 88.225 94.495 89.355 ;
        RECT 94.685 89.210 94.975 89.935 ;
        RECT 95.150 89.195 95.405 89.765 ;
        RECT 95.575 89.535 95.905 89.935 ;
        RECT 96.330 89.400 96.860 89.765 ;
        RECT 96.330 89.365 96.505 89.400 ;
        RECT 95.575 89.195 96.505 89.365 ;
        RECT 91.435 87.725 91.765 88.225 ;
        RECT 91.935 87.985 93.570 88.225 ;
        RECT 91.935 87.895 92.165 87.985 ;
        RECT 92.275 87.725 92.605 87.765 ;
        RECT 91.435 87.555 92.605 87.725 ;
        RECT 92.795 87.385 93.150 87.805 ;
        RECT 93.320 87.555 93.570 87.985 ;
        RECT 93.740 87.385 94.070 88.145 ;
        RECT 94.240 87.555 94.495 88.225 ;
        RECT 94.685 87.385 94.975 88.550 ;
        RECT 95.150 88.525 95.320 89.195 ;
        RECT 95.575 89.025 95.745 89.195 ;
        RECT 95.490 88.695 95.745 89.025 ;
        RECT 95.970 88.695 96.165 89.025 ;
        RECT 95.150 87.555 95.485 88.525 ;
        RECT 95.655 87.385 95.825 88.525 ;
        RECT 95.995 87.725 96.165 88.695 ;
        RECT 96.335 88.065 96.505 89.195 ;
        RECT 96.675 88.405 96.845 89.205 ;
        RECT 97.050 88.915 97.325 89.765 ;
        RECT 97.045 88.745 97.325 88.915 ;
        RECT 97.050 88.605 97.325 88.745 ;
        RECT 97.495 88.405 97.685 89.765 ;
        RECT 97.865 89.400 98.375 89.935 ;
        RECT 98.595 89.125 98.840 89.730 ;
        RECT 99.290 89.430 99.625 89.935 ;
        RECT 99.795 89.365 100.035 89.740 ;
        RECT 100.315 89.605 100.485 89.750 ;
        RECT 100.315 89.410 100.690 89.605 ;
        RECT 101.050 89.440 101.445 89.935 ;
        RECT 97.885 88.955 99.115 89.125 ;
        RECT 96.675 88.235 97.685 88.405 ;
        RECT 97.855 88.390 98.605 88.580 ;
        RECT 96.335 87.895 97.460 88.065 ;
        RECT 97.855 87.725 98.025 88.390 ;
        RECT 98.775 88.145 99.115 88.955 ;
        RECT 99.345 88.405 99.645 89.255 ;
        RECT 99.815 89.215 100.035 89.365 ;
        RECT 99.815 88.885 100.350 89.215 ;
        RECT 100.520 89.075 100.690 89.410 ;
        RECT 101.615 89.245 101.855 89.765 ;
        RECT 99.815 88.235 100.050 88.885 ;
        RECT 100.520 88.715 101.505 89.075 ;
        RECT 95.995 87.555 98.025 87.725 ;
        RECT 98.195 87.385 98.365 88.145 ;
        RECT 98.600 87.735 99.115 88.145 ;
        RECT 99.375 88.005 100.050 88.235 ;
        RECT 100.220 88.695 101.505 88.715 ;
        RECT 100.220 88.545 101.080 88.695 ;
        RECT 99.375 87.575 99.545 88.005 ;
        RECT 99.715 87.385 100.045 87.835 ;
        RECT 100.220 87.600 100.505 88.545 ;
        RECT 101.680 88.440 101.855 89.245 ;
        RECT 102.045 89.165 104.635 89.935 ;
        RECT 104.810 89.430 105.145 89.935 ;
        RECT 105.315 89.365 105.555 89.740 ;
        RECT 105.835 89.605 106.005 89.750 ;
        RECT 105.835 89.410 106.210 89.605 ;
        RECT 106.570 89.440 106.965 89.935 ;
        RECT 102.045 88.645 103.255 89.165 ;
        RECT 103.425 88.475 104.635 88.995 ;
        RECT 100.680 88.065 101.375 88.375 ;
        RECT 100.685 87.385 101.370 87.855 ;
        RECT 101.550 87.655 101.855 88.440 ;
        RECT 102.045 87.385 104.635 88.475 ;
        RECT 104.865 88.405 105.165 89.255 ;
        RECT 105.335 89.215 105.555 89.365 ;
        RECT 105.335 88.885 105.870 89.215 ;
        RECT 106.040 89.075 106.210 89.410 ;
        RECT 107.135 89.245 107.375 89.765 ;
        RECT 105.335 88.235 105.570 88.885 ;
        RECT 106.040 88.715 107.025 89.075 ;
        RECT 104.895 88.005 105.570 88.235 ;
        RECT 105.740 88.695 107.025 88.715 ;
        RECT 105.740 88.545 106.600 88.695 ;
        RECT 104.895 87.575 105.065 88.005 ;
        RECT 105.235 87.385 105.565 87.835 ;
        RECT 105.740 87.600 106.025 88.545 ;
        RECT 107.200 88.440 107.375 89.245 ;
        RECT 107.565 89.165 111.075 89.935 ;
        RECT 111.245 89.185 112.455 89.935 ;
        RECT 112.630 89.430 112.965 89.935 ;
        RECT 113.135 89.365 113.375 89.740 ;
        RECT 113.655 89.605 113.825 89.750 ;
        RECT 113.655 89.410 114.030 89.605 ;
        RECT 114.390 89.440 114.785 89.935 ;
        RECT 107.565 88.645 109.215 89.165 ;
        RECT 109.385 88.475 111.075 88.995 ;
        RECT 111.245 88.645 111.765 89.185 ;
        RECT 111.935 88.475 112.455 89.015 ;
        RECT 106.200 88.065 106.895 88.375 ;
        RECT 106.205 87.385 106.890 87.855 ;
        RECT 107.070 87.655 107.375 88.440 ;
        RECT 107.565 87.385 111.075 88.475 ;
        RECT 111.245 87.385 112.455 88.475 ;
        RECT 112.685 88.405 112.985 89.255 ;
        RECT 113.155 89.215 113.375 89.365 ;
        RECT 113.155 88.885 113.690 89.215 ;
        RECT 113.860 89.075 114.030 89.410 ;
        RECT 114.955 89.245 115.195 89.765 ;
        RECT 113.155 88.235 113.390 88.885 ;
        RECT 113.860 88.715 114.845 89.075 ;
        RECT 112.715 88.005 113.390 88.235 ;
        RECT 113.560 88.695 114.845 88.715 ;
        RECT 113.560 88.545 114.420 88.695 ;
        RECT 112.715 87.575 112.885 88.005 ;
        RECT 113.055 87.385 113.385 87.835 ;
        RECT 113.560 87.600 113.845 88.545 ;
        RECT 115.020 88.440 115.195 89.245 ;
        RECT 114.020 88.065 114.715 88.375 ;
        RECT 114.025 87.385 114.710 87.855 ;
        RECT 114.890 87.655 115.195 88.440 ;
        RECT 115.850 89.195 116.105 89.765 ;
        RECT 116.275 89.535 116.605 89.935 ;
        RECT 117.030 89.400 117.560 89.765 ;
        RECT 117.750 89.595 118.025 89.765 ;
        RECT 117.745 89.425 118.025 89.595 ;
        RECT 117.030 89.365 117.205 89.400 ;
        RECT 116.275 89.195 117.205 89.365 ;
        RECT 115.850 88.525 116.020 89.195 ;
        RECT 116.275 89.025 116.445 89.195 ;
        RECT 116.190 88.695 116.445 89.025 ;
        RECT 116.670 88.695 116.865 89.025 ;
        RECT 115.850 87.555 116.185 88.525 ;
        RECT 116.355 87.385 116.525 88.525 ;
        RECT 116.695 87.725 116.865 88.695 ;
        RECT 117.035 88.065 117.205 89.195 ;
        RECT 117.375 88.405 117.545 89.205 ;
        RECT 117.750 88.605 118.025 89.425 ;
        RECT 118.195 88.405 118.385 89.765 ;
        RECT 118.565 89.400 119.075 89.935 ;
        RECT 119.295 89.125 119.540 89.730 ;
        RECT 120.445 89.210 120.735 89.935 ;
        RECT 120.905 89.165 123.495 89.935 ;
        RECT 123.755 89.385 123.925 89.675 ;
        RECT 124.095 89.555 124.425 89.935 ;
        RECT 123.755 89.215 124.420 89.385 ;
        RECT 118.585 88.955 119.815 89.125 ;
        RECT 117.375 88.235 118.385 88.405 ;
        RECT 118.555 88.390 119.305 88.580 ;
        RECT 117.035 87.895 118.160 88.065 ;
        RECT 118.555 87.725 118.725 88.390 ;
        RECT 119.475 88.145 119.815 88.955 ;
        RECT 120.905 88.645 122.115 89.165 ;
        RECT 116.695 87.555 118.725 87.725 ;
        RECT 118.895 87.385 119.065 88.145 ;
        RECT 119.300 87.735 119.815 88.145 ;
        RECT 120.445 87.385 120.735 88.550 ;
        RECT 122.285 88.475 123.495 88.995 ;
        RECT 120.905 87.385 123.495 88.475 ;
        RECT 123.670 88.395 124.020 89.045 ;
        RECT 124.190 88.225 124.420 89.215 ;
        RECT 123.755 88.055 124.420 88.225 ;
        RECT 123.755 87.555 123.925 88.055 ;
        RECT 124.095 87.385 124.425 87.885 ;
        RECT 124.595 87.555 124.780 89.675 ;
        RECT 125.035 89.475 125.285 89.935 ;
        RECT 125.455 89.485 125.790 89.655 ;
        RECT 125.985 89.485 126.660 89.655 ;
        RECT 125.455 89.345 125.625 89.485 ;
        RECT 124.950 88.355 125.230 89.305 ;
        RECT 125.400 89.215 125.625 89.345 ;
        RECT 125.400 88.110 125.570 89.215 ;
        RECT 125.795 89.065 126.320 89.285 ;
        RECT 125.740 88.300 125.980 88.895 ;
        RECT 126.150 88.365 126.320 89.065 ;
        RECT 126.490 88.705 126.660 89.485 ;
        RECT 126.980 89.435 127.350 89.935 ;
        RECT 127.530 89.485 127.935 89.655 ;
        RECT 128.105 89.485 128.890 89.655 ;
        RECT 127.530 89.255 127.700 89.485 ;
        RECT 126.870 88.955 127.700 89.255 ;
        RECT 128.085 88.985 128.550 89.315 ;
        RECT 126.870 88.925 127.070 88.955 ;
        RECT 127.190 88.705 127.360 88.775 ;
        RECT 126.490 88.535 127.360 88.705 ;
        RECT 126.850 88.445 127.360 88.535 ;
        RECT 125.400 87.980 125.705 88.110 ;
        RECT 126.150 88.000 126.680 88.365 ;
        RECT 125.020 87.385 125.285 87.845 ;
        RECT 125.455 87.555 125.705 87.980 ;
        RECT 126.850 87.830 127.020 88.445 ;
        RECT 125.915 87.660 127.020 87.830 ;
        RECT 127.190 87.385 127.360 88.185 ;
        RECT 127.530 87.885 127.700 88.955 ;
        RECT 127.870 88.055 128.060 88.775 ;
        RECT 128.230 88.025 128.550 88.985 ;
        RECT 128.720 89.025 128.890 89.485 ;
        RECT 129.165 89.405 129.375 89.935 ;
        RECT 129.635 89.195 129.965 89.720 ;
        RECT 130.135 89.325 130.305 89.935 ;
        RECT 130.475 89.280 130.805 89.715 ;
        RECT 130.475 89.195 130.855 89.280 ;
        RECT 129.765 89.025 129.965 89.195 ;
        RECT 130.630 89.155 130.855 89.195 ;
        RECT 128.720 88.695 129.595 89.025 ;
        RECT 129.765 88.695 130.515 89.025 ;
        RECT 127.530 87.555 127.780 87.885 ;
        RECT 128.720 87.855 128.890 88.695 ;
        RECT 129.765 88.490 129.955 88.695 ;
        RECT 130.685 88.575 130.855 89.155 ;
        RECT 130.640 88.525 130.855 88.575 ;
        RECT 129.060 88.115 129.955 88.490 ;
        RECT 130.465 88.445 130.855 88.525 ;
        RECT 131.030 89.195 131.285 89.765 ;
        RECT 131.455 89.535 131.785 89.935 ;
        RECT 132.210 89.400 132.740 89.765 ;
        RECT 132.930 89.595 133.205 89.765 ;
        RECT 132.925 89.425 133.205 89.595 ;
        RECT 132.210 89.365 132.385 89.400 ;
        RECT 131.455 89.195 132.385 89.365 ;
        RECT 131.030 88.525 131.200 89.195 ;
        RECT 131.455 89.025 131.625 89.195 ;
        RECT 131.370 88.695 131.625 89.025 ;
        RECT 131.850 88.695 132.045 89.025 ;
        RECT 128.005 87.685 128.890 87.855 ;
        RECT 129.070 87.385 129.385 87.885 ;
        RECT 129.615 87.555 129.955 88.115 ;
        RECT 130.125 87.385 130.295 88.395 ;
        RECT 130.465 87.600 130.795 88.445 ;
        RECT 131.030 87.555 131.365 88.525 ;
        RECT 131.535 87.385 131.705 88.525 ;
        RECT 131.875 87.725 132.045 88.695 ;
        RECT 132.215 88.065 132.385 89.195 ;
        RECT 132.555 88.405 132.725 89.205 ;
        RECT 132.930 88.605 133.205 89.425 ;
        RECT 133.375 88.405 133.565 89.765 ;
        RECT 133.745 89.400 134.255 89.935 ;
        RECT 134.475 89.125 134.720 89.730 ;
        RECT 135.165 89.260 135.425 89.765 ;
        RECT 135.605 89.555 135.935 89.935 ;
        RECT 136.115 89.385 136.285 89.765 ;
        RECT 133.765 88.955 134.995 89.125 ;
        RECT 132.555 88.235 133.565 88.405 ;
        RECT 133.735 88.390 134.485 88.580 ;
        RECT 132.215 87.895 133.340 88.065 ;
        RECT 133.735 87.725 133.905 88.390 ;
        RECT 134.655 88.145 134.995 88.955 ;
        RECT 131.875 87.555 133.905 87.725 ;
        RECT 134.075 87.385 134.245 88.145 ;
        RECT 134.480 87.735 134.995 88.145 ;
        RECT 135.165 88.460 135.345 89.260 ;
        RECT 135.620 89.215 136.285 89.385 ;
        RECT 136.635 89.385 136.805 89.675 ;
        RECT 136.975 89.555 137.305 89.935 ;
        RECT 136.635 89.215 137.300 89.385 ;
        RECT 135.620 88.960 135.790 89.215 ;
        RECT 135.515 88.630 135.790 88.960 ;
        RECT 136.015 88.665 136.355 89.035 ;
        RECT 135.620 88.485 135.790 88.630 ;
        RECT 135.165 87.555 135.435 88.460 ;
        RECT 135.620 88.315 136.295 88.485 ;
        RECT 136.550 88.395 136.900 89.045 ;
        RECT 135.605 87.385 135.935 88.145 ;
        RECT 136.115 87.555 136.295 88.315 ;
        RECT 137.070 88.225 137.300 89.215 ;
        RECT 136.635 88.055 137.300 88.225 ;
        RECT 136.635 87.555 136.805 88.055 ;
        RECT 136.975 87.385 137.305 87.885 ;
        RECT 137.475 87.555 137.660 89.675 ;
        RECT 137.915 89.475 138.165 89.935 ;
        RECT 138.335 89.485 138.670 89.655 ;
        RECT 138.865 89.485 139.540 89.655 ;
        RECT 138.335 89.345 138.505 89.485 ;
        RECT 137.830 88.355 138.110 89.305 ;
        RECT 138.280 89.215 138.505 89.345 ;
        RECT 138.280 88.110 138.450 89.215 ;
        RECT 138.675 89.065 139.200 89.285 ;
        RECT 138.620 88.300 138.860 88.895 ;
        RECT 139.030 88.365 139.200 89.065 ;
        RECT 139.370 88.705 139.540 89.485 ;
        RECT 139.860 89.435 140.230 89.935 ;
        RECT 140.410 89.485 140.815 89.655 ;
        RECT 140.985 89.485 141.770 89.655 ;
        RECT 140.410 89.255 140.580 89.485 ;
        RECT 139.750 88.955 140.580 89.255 ;
        RECT 140.965 88.985 141.430 89.315 ;
        RECT 139.750 88.925 139.950 88.955 ;
        RECT 140.070 88.705 140.240 88.775 ;
        RECT 139.370 88.535 140.240 88.705 ;
        RECT 139.730 88.445 140.240 88.535 ;
        RECT 138.280 87.980 138.585 88.110 ;
        RECT 139.030 88.000 139.560 88.365 ;
        RECT 137.900 87.385 138.165 87.845 ;
        RECT 138.335 87.555 138.585 87.980 ;
        RECT 139.730 87.830 139.900 88.445 ;
        RECT 138.795 87.660 139.900 87.830 ;
        RECT 140.070 87.385 140.240 88.185 ;
        RECT 140.410 87.885 140.580 88.955 ;
        RECT 140.750 88.055 140.940 88.775 ;
        RECT 141.110 88.025 141.430 88.985 ;
        RECT 141.600 89.025 141.770 89.485 ;
        RECT 142.045 89.405 142.255 89.935 ;
        RECT 142.515 89.195 142.845 89.720 ;
        RECT 143.015 89.325 143.185 89.935 ;
        RECT 143.355 89.280 143.685 89.715 ;
        RECT 143.995 89.385 144.165 89.765 ;
        RECT 144.380 89.555 144.710 89.935 ;
        RECT 143.355 89.195 143.735 89.280 ;
        RECT 143.995 89.215 144.710 89.385 ;
        RECT 142.645 89.025 142.845 89.195 ;
        RECT 143.510 89.155 143.735 89.195 ;
        RECT 141.600 88.695 142.475 89.025 ;
        RECT 142.645 88.695 143.395 89.025 ;
        RECT 140.410 87.555 140.660 87.885 ;
        RECT 141.600 87.855 141.770 88.695 ;
        RECT 142.645 88.490 142.835 88.695 ;
        RECT 143.565 88.575 143.735 89.155 ;
        RECT 143.905 88.665 144.260 89.035 ;
        RECT 144.540 89.025 144.710 89.215 ;
        RECT 144.880 89.190 145.135 89.765 ;
        RECT 144.540 88.695 144.795 89.025 ;
        RECT 143.520 88.525 143.735 88.575 ;
        RECT 141.940 88.115 142.835 88.490 ;
        RECT 143.345 88.445 143.735 88.525 ;
        RECT 144.540 88.485 144.710 88.695 ;
        RECT 140.885 87.685 141.770 87.855 ;
        RECT 141.950 87.385 142.265 87.885 ;
        RECT 142.495 87.555 142.835 88.115 ;
        RECT 143.005 87.385 143.175 88.395 ;
        RECT 143.345 87.600 143.675 88.445 ;
        RECT 143.995 88.315 144.710 88.485 ;
        RECT 144.965 88.460 145.135 89.190 ;
        RECT 145.310 89.095 145.570 89.935 ;
        RECT 145.745 89.185 146.955 89.935 ;
        RECT 143.995 87.555 144.165 88.315 ;
        RECT 144.380 87.385 144.710 88.145 ;
        RECT 144.880 87.555 145.135 88.460 ;
        RECT 145.310 87.385 145.570 88.535 ;
        RECT 145.745 88.475 146.265 89.015 ;
        RECT 146.435 88.645 146.955 89.185 ;
        RECT 145.745 87.385 146.955 88.475 ;
        RECT 17.320 87.215 147.040 87.385 ;
        RECT 17.405 86.125 18.615 87.215 ;
        RECT 17.405 85.415 17.925 85.955 ;
        RECT 18.095 85.585 18.615 86.125 ;
        RECT 18.865 86.285 19.045 87.045 ;
        RECT 19.225 86.455 19.555 87.215 ;
        RECT 18.865 86.115 19.540 86.285 ;
        RECT 19.725 86.140 19.995 87.045 ;
        RECT 19.370 85.970 19.540 86.115 ;
        RECT 18.805 85.565 19.145 85.935 ;
        RECT 19.370 85.640 19.645 85.970 ;
        RECT 17.405 84.665 18.615 85.415 ;
        RECT 19.370 85.385 19.540 85.640 ;
        RECT 18.875 85.215 19.540 85.385 ;
        RECT 19.815 85.340 19.995 86.140 ;
        RECT 20.255 86.285 20.425 87.045 ;
        RECT 20.605 86.455 20.935 87.215 ;
        RECT 20.255 86.115 20.920 86.285 ;
        RECT 21.105 86.140 21.375 87.045 ;
        RECT 20.750 85.970 20.920 86.115 ;
        RECT 20.185 85.565 20.515 85.935 ;
        RECT 20.750 85.640 21.035 85.970 ;
        RECT 20.750 85.385 20.920 85.640 ;
        RECT 18.875 84.835 19.045 85.215 ;
        RECT 19.225 84.665 19.555 85.045 ;
        RECT 19.735 84.835 19.995 85.340 ;
        RECT 20.255 85.215 20.920 85.385 ;
        RECT 21.205 85.340 21.375 86.140 ;
        RECT 22.010 86.065 22.270 87.215 ;
        RECT 22.445 86.140 22.700 87.045 ;
        RECT 22.870 86.455 23.200 87.215 ;
        RECT 23.415 86.285 23.585 87.045 ;
        RECT 20.255 84.835 20.425 85.215 ;
        RECT 20.605 84.665 20.935 85.045 ;
        RECT 21.115 84.835 21.375 85.340 ;
        RECT 22.010 84.665 22.270 85.505 ;
        RECT 22.445 85.410 22.615 86.140 ;
        RECT 22.870 86.115 23.585 86.285 ;
        RECT 23.925 86.285 24.105 87.045 ;
        RECT 24.285 86.455 24.615 87.215 ;
        RECT 23.925 86.115 24.600 86.285 ;
        RECT 24.785 86.140 25.055 87.045 ;
        RECT 22.870 85.905 23.040 86.115 ;
        RECT 24.430 85.970 24.600 86.115 ;
        RECT 22.785 85.575 23.040 85.905 ;
        RECT 22.445 84.835 22.700 85.410 ;
        RECT 22.870 85.385 23.040 85.575 ;
        RECT 23.320 85.565 23.675 85.935 ;
        RECT 23.865 85.565 24.205 85.935 ;
        RECT 24.430 85.640 24.705 85.970 ;
        RECT 24.430 85.385 24.600 85.640 ;
        RECT 22.870 85.215 23.585 85.385 ;
        RECT 22.870 84.665 23.200 85.045 ;
        RECT 23.415 84.835 23.585 85.215 ;
        RECT 23.935 85.215 24.600 85.385 ;
        RECT 24.875 85.340 25.055 86.140 ;
        RECT 25.305 86.285 25.485 87.045 ;
        RECT 25.665 86.455 25.995 87.215 ;
        RECT 25.305 86.115 25.980 86.285 ;
        RECT 26.165 86.140 26.435 87.045 ;
        RECT 25.810 85.970 25.980 86.115 ;
        RECT 25.245 85.565 25.585 85.935 ;
        RECT 25.810 85.640 26.085 85.970 ;
        RECT 25.810 85.385 25.980 85.640 ;
        RECT 23.935 84.835 24.105 85.215 ;
        RECT 24.285 84.665 24.615 85.045 ;
        RECT 24.795 84.835 25.055 85.340 ;
        RECT 25.315 85.215 25.980 85.385 ;
        RECT 26.255 85.340 26.435 86.140 ;
        RECT 26.605 86.125 28.275 87.215 ;
        RECT 25.315 84.835 25.485 85.215 ;
        RECT 25.665 84.665 25.995 85.045 ;
        RECT 26.175 84.835 26.435 85.340 ;
        RECT 26.605 85.435 27.355 85.955 ;
        RECT 27.525 85.605 28.275 86.125 ;
        RECT 28.535 86.285 28.705 87.045 ;
        RECT 28.920 86.455 29.250 87.215 ;
        RECT 28.535 86.115 29.250 86.285 ;
        RECT 29.420 86.140 29.675 87.045 ;
        RECT 28.445 85.565 28.800 85.935 ;
        RECT 29.080 85.905 29.250 86.115 ;
        RECT 29.080 85.575 29.335 85.905 ;
        RECT 26.605 84.665 28.275 85.435 ;
        RECT 29.080 85.385 29.250 85.575 ;
        RECT 29.505 85.410 29.675 86.140 ;
        RECT 29.850 86.065 30.110 87.215 ;
        RECT 30.285 86.050 30.575 87.215 ;
        RECT 30.825 86.285 31.005 87.045 ;
        RECT 31.185 86.455 31.515 87.215 ;
        RECT 30.825 86.115 31.500 86.285 ;
        RECT 31.685 86.140 31.955 87.045 ;
        RECT 31.330 85.970 31.500 86.115 ;
        RECT 30.765 85.565 31.105 85.935 ;
        RECT 31.330 85.640 31.605 85.970 ;
        RECT 28.535 85.215 29.250 85.385 ;
        RECT 28.535 84.835 28.705 85.215 ;
        RECT 28.920 84.665 29.250 85.045 ;
        RECT 29.420 84.835 29.675 85.410 ;
        RECT 29.850 84.665 30.110 85.505 ;
        RECT 30.285 84.665 30.575 85.390 ;
        RECT 31.330 85.385 31.500 85.640 ;
        RECT 30.835 85.215 31.500 85.385 ;
        RECT 31.775 85.340 31.955 86.140 ;
        RECT 30.835 84.835 31.005 85.215 ;
        RECT 31.185 84.665 31.515 85.045 ;
        RECT 31.695 84.835 31.955 85.340 ;
        RECT 32.125 86.415 32.565 87.045 ;
        RECT 32.125 85.405 32.435 86.415 ;
        RECT 32.740 86.365 33.055 87.215 ;
        RECT 33.225 86.875 34.655 87.045 ;
        RECT 33.225 86.195 33.395 86.875 ;
        RECT 32.605 86.025 33.395 86.195 ;
        RECT 32.605 85.575 32.775 86.025 ;
        RECT 33.565 85.905 33.765 86.705 ;
        RECT 32.945 85.575 33.335 85.855 ;
        RECT 33.520 85.575 33.765 85.905 ;
        RECT 33.965 85.575 34.215 86.705 ;
        RECT 34.405 86.245 34.655 86.875 ;
        RECT 34.835 86.415 35.165 87.215 ;
        RECT 35.435 86.285 35.605 87.045 ;
        RECT 35.785 86.455 36.115 87.215 ;
        RECT 34.405 86.075 35.175 86.245 ;
        RECT 35.435 86.115 36.100 86.285 ;
        RECT 36.285 86.140 36.555 87.045 ;
        RECT 34.430 85.575 34.835 85.905 ;
        RECT 35.005 85.405 35.175 86.075 ;
        RECT 35.930 85.970 36.100 86.115 ;
        RECT 35.365 85.565 35.695 85.935 ;
        RECT 35.930 85.640 36.215 85.970 ;
        RECT 32.125 84.845 32.565 85.405 ;
        RECT 32.735 84.665 33.185 85.405 ;
        RECT 33.355 85.235 34.515 85.405 ;
        RECT 33.355 84.835 33.525 85.235 ;
        RECT 33.695 84.665 34.115 85.065 ;
        RECT 34.285 84.835 34.515 85.235 ;
        RECT 34.685 84.835 35.175 85.405 ;
        RECT 35.930 85.385 36.100 85.640 ;
        RECT 35.435 85.215 36.100 85.385 ;
        RECT 36.385 85.340 36.555 86.140 ;
        RECT 36.725 86.125 37.935 87.215 ;
        RECT 35.435 84.835 35.605 85.215 ;
        RECT 35.785 84.665 36.115 85.045 ;
        RECT 36.295 84.835 36.555 85.340 ;
        RECT 36.725 85.415 37.245 85.955 ;
        RECT 37.415 85.585 37.935 86.125 ;
        RECT 38.195 86.285 38.365 87.045 ;
        RECT 38.545 86.455 38.875 87.215 ;
        RECT 38.195 86.115 38.860 86.285 ;
        RECT 39.045 86.140 39.315 87.045 ;
        RECT 38.690 85.970 38.860 86.115 ;
        RECT 38.125 85.565 38.455 85.935 ;
        RECT 38.690 85.640 38.975 85.970 ;
        RECT 36.725 84.665 37.935 85.415 ;
        RECT 38.690 85.385 38.860 85.640 ;
        RECT 38.195 85.215 38.860 85.385 ;
        RECT 39.145 85.340 39.315 86.140 ;
        RECT 39.485 86.125 41.155 87.215 ;
        RECT 38.195 84.835 38.365 85.215 ;
        RECT 38.545 84.665 38.875 85.045 ;
        RECT 39.055 84.835 39.315 85.340 ;
        RECT 39.485 85.435 40.235 85.955 ;
        RECT 40.405 85.605 41.155 86.125 ;
        RECT 41.325 86.140 41.595 87.045 ;
        RECT 41.765 86.455 42.095 87.215 ;
        RECT 42.275 86.285 42.455 87.045 ;
        RECT 39.485 84.665 41.155 85.435 ;
        RECT 41.325 85.340 41.505 86.140 ;
        RECT 41.780 86.115 42.455 86.285 ;
        RECT 41.780 85.970 41.950 86.115 ;
        RECT 43.165 86.050 43.455 87.215 ;
        RECT 44.545 86.140 44.815 87.045 ;
        RECT 44.985 86.455 45.315 87.215 ;
        RECT 45.495 86.285 45.675 87.045 ;
        RECT 41.675 85.640 41.950 85.970 ;
        RECT 41.780 85.385 41.950 85.640 ;
        RECT 42.175 85.565 42.515 85.935 ;
        RECT 41.325 84.835 41.585 85.340 ;
        RECT 41.780 85.215 42.445 85.385 ;
        RECT 41.765 84.665 42.095 85.045 ;
        RECT 42.275 84.835 42.445 85.215 ;
        RECT 43.165 84.665 43.455 85.390 ;
        RECT 44.545 85.340 44.725 86.140 ;
        RECT 45.000 86.115 45.675 86.285 ;
        RECT 45.925 86.125 47.595 87.215 ;
        RECT 45.000 85.970 45.170 86.115 ;
        RECT 44.895 85.640 45.170 85.970 ;
        RECT 45.000 85.385 45.170 85.640 ;
        RECT 45.395 85.565 45.735 85.935 ;
        RECT 45.925 85.435 46.675 85.955 ;
        RECT 46.845 85.605 47.595 86.125 ;
        RECT 47.765 86.140 48.035 87.045 ;
        RECT 48.205 86.455 48.535 87.215 ;
        RECT 48.715 86.285 48.895 87.045 ;
        RECT 44.545 84.835 44.805 85.340 ;
        RECT 45.000 85.215 45.665 85.385 ;
        RECT 44.985 84.665 45.315 85.045 ;
        RECT 45.495 84.835 45.665 85.215 ;
        RECT 45.925 84.665 47.595 85.435 ;
        RECT 47.765 85.340 47.945 86.140 ;
        RECT 48.220 86.115 48.895 86.285 ;
        RECT 49.145 86.125 50.815 87.215 ;
        RECT 48.220 85.970 48.390 86.115 ;
        RECT 48.115 85.640 48.390 85.970 ;
        RECT 48.220 85.385 48.390 85.640 ;
        RECT 48.615 85.565 48.955 85.935 ;
        RECT 49.145 85.435 49.895 85.955 ;
        RECT 50.065 85.605 50.815 86.125 ;
        RECT 50.985 86.140 51.255 87.045 ;
        RECT 51.425 86.455 51.755 87.215 ;
        RECT 51.935 86.285 52.105 87.045 ;
        RECT 47.765 84.835 48.025 85.340 ;
        RECT 48.220 85.215 48.885 85.385 ;
        RECT 48.205 84.665 48.535 85.045 ;
        RECT 48.715 84.835 48.885 85.215 ;
        RECT 49.145 84.665 50.815 85.435 ;
        RECT 50.985 85.340 51.155 86.140 ;
        RECT 51.440 86.115 52.105 86.285 ;
        RECT 52.365 86.125 54.035 87.215 ;
        RECT 51.440 85.970 51.610 86.115 ;
        RECT 51.325 85.640 51.610 85.970 ;
        RECT 51.440 85.385 51.610 85.640 ;
        RECT 51.845 85.565 52.175 85.935 ;
        RECT 52.365 85.435 53.115 85.955 ;
        RECT 53.285 85.605 54.035 86.125 ;
        RECT 54.205 86.140 54.475 87.045 ;
        RECT 54.645 86.455 54.975 87.215 ;
        RECT 55.155 86.285 55.325 87.045 ;
        RECT 50.985 84.835 51.245 85.340 ;
        RECT 51.440 85.215 52.105 85.385 ;
        RECT 51.425 84.665 51.755 85.045 ;
        RECT 51.935 84.835 52.105 85.215 ;
        RECT 52.365 84.665 54.035 85.435 ;
        RECT 54.205 85.340 54.375 86.140 ;
        RECT 54.660 86.115 55.325 86.285 ;
        RECT 54.660 85.970 54.830 86.115 ;
        RECT 56.045 86.050 56.335 87.215 ;
        RECT 56.510 86.065 56.770 87.215 ;
        RECT 56.945 86.140 57.200 87.045 ;
        RECT 57.370 86.455 57.700 87.215 ;
        RECT 57.915 86.285 58.085 87.045 ;
        RECT 54.545 85.640 54.830 85.970 ;
        RECT 54.660 85.385 54.830 85.640 ;
        RECT 55.065 85.565 55.395 85.935 ;
        RECT 54.205 84.835 54.465 85.340 ;
        RECT 54.660 85.215 55.325 85.385 ;
        RECT 54.645 84.665 54.975 85.045 ;
        RECT 55.155 84.835 55.325 85.215 ;
        RECT 56.045 84.665 56.335 85.390 ;
        RECT 56.510 84.665 56.770 85.505 ;
        RECT 56.945 85.410 57.115 86.140 ;
        RECT 57.370 86.115 58.085 86.285 ;
        RECT 57.370 85.905 57.540 86.115 ;
        RECT 58.350 86.065 58.610 87.215 ;
        RECT 58.785 86.140 59.040 87.045 ;
        RECT 59.210 86.455 59.540 87.215 ;
        RECT 59.755 86.285 59.925 87.045 ;
        RECT 57.285 85.575 57.540 85.905 ;
        RECT 56.945 84.835 57.200 85.410 ;
        RECT 57.370 85.385 57.540 85.575 ;
        RECT 57.820 85.565 58.175 85.935 ;
        RECT 57.370 85.215 58.085 85.385 ;
        RECT 57.370 84.665 57.700 85.045 ;
        RECT 57.915 84.835 58.085 85.215 ;
        RECT 58.350 84.665 58.610 85.505 ;
        RECT 58.785 85.410 58.955 86.140 ;
        RECT 59.210 86.115 59.925 86.285 ;
        RECT 59.210 85.905 59.380 86.115 ;
        RECT 60.190 86.065 60.450 87.215 ;
        RECT 60.625 86.140 60.880 87.045 ;
        RECT 61.050 86.455 61.380 87.215 ;
        RECT 61.595 86.285 61.765 87.045 ;
        RECT 59.125 85.575 59.380 85.905 ;
        RECT 58.785 84.835 59.040 85.410 ;
        RECT 59.210 85.385 59.380 85.575 ;
        RECT 59.660 85.565 60.015 85.935 ;
        RECT 59.210 85.215 59.925 85.385 ;
        RECT 59.210 84.665 59.540 85.045 ;
        RECT 59.755 84.835 59.925 85.215 ;
        RECT 60.190 84.665 60.450 85.505 ;
        RECT 60.625 85.410 60.795 86.140 ;
        RECT 61.050 86.115 61.765 86.285 ;
        RECT 62.045 86.160 62.350 86.945 ;
        RECT 62.530 86.745 63.215 87.215 ;
        RECT 62.525 86.225 63.220 86.535 ;
        RECT 61.050 85.905 61.220 86.115 ;
        RECT 60.965 85.575 61.220 85.905 ;
        RECT 60.625 84.835 60.880 85.410 ;
        RECT 61.050 85.385 61.220 85.575 ;
        RECT 61.500 85.565 61.855 85.935 ;
        RECT 61.050 85.215 61.765 85.385 ;
        RECT 61.050 84.665 61.380 85.045 ;
        RECT 61.595 84.835 61.765 85.215 ;
        RECT 62.045 85.355 62.220 86.160 ;
        RECT 63.395 86.055 63.680 87.000 ;
        RECT 63.855 86.765 64.185 87.215 ;
        RECT 64.355 86.595 64.525 87.025 ;
        RECT 62.820 85.905 63.680 86.055 ;
        RECT 62.395 85.885 63.680 85.905 ;
        RECT 63.850 86.365 64.525 86.595 ;
        RECT 65.795 86.595 65.965 87.025 ;
        RECT 66.135 86.765 66.465 87.215 ;
        RECT 65.795 86.365 66.470 86.595 ;
        RECT 62.395 85.525 63.380 85.885 ;
        RECT 63.850 85.715 64.085 86.365 ;
        RECT 62.045 84.835 62.285 85.355 ;
        RECT 63.210 85.190 63.380 85.525 ;
        RECT 63.550 85.385 64.085 85.715 ;
        RECT 63.865 85.235 64.085 85.385 ;
        RECT 64.255 85.345 64.555 86.195 ;
        RECT 65.765 85.345 66.065 86.195 ;
        RECT 66.235 85.715 66.470 86.365 ;
        RECT 66.640 86.055 66.925 87.000 ;
        RECT 67.105 86.745 67.790 87.215 ;
        RECT 67.100 86.225 67.795 86.535 ;
        RECT 67.970 86.160 68.275 86.945 ;
        RECT 66.640 85.905 67.500 86.055 ;
        RECT 66.640 85.885 67.925 85.905 ;
        RECT 66.235 85.385 66.770 85.715 ;
        RECT 66.940 85.525 67.925 85.885 ;
        RECT 66.235 85.235 66.455 85.385 ;
        RECT 62.455 84.665 62.850 85.160 ;
        RECT 63.210 84.995 63.585 85.190 ;
        RECT 63.415 84.850 63.585 84.995 ;
        RECT 63.865 84.860 64.105 85.235 ;
        RECT 64.275 84.665 64.610 85.170 ;
        RECT 65.710 84.665 66.045 85.170 ;
        RECT 66.215 84.860 66.455 85.235 ;
        RECT 66.940 85.190 67.110 85.525 ;
        RECT 68.100 85.355 68.275 86.160 ;
        RECT 68.925 86.050 69.215 87.215 ;
        RECT 69.390 86.075 69.725 87.045 ;
        RECT 69.895 86.075 70.065 87.215 ;
        RECT 70.235 86.875 72.265 87.045 ;
        RECT 69.390 85.405 69.560 86.075 ;
        RECT 70.235 85.905 70.405 86.875 ;
        RECT 69.730 85.575 69.985 85.905 ;
        RECT 70.210 85.575 70.405 85.905 ;
        RECT 70.575 86.535 71.700 86.705 ;
        RECT 69.815 85.405 69.985 85.575 ;
        RECT 70.575 85.405 70.745 86.535 ;
        RECT 66.735 84.995 67.110 85.190 ;
        RECT 66.735 84.850 66.905 84.995 ;
        RECT 67.470 84.665 67.865 85.160 ;
        RECT 68.035 84.835 68.275 85.355 ;
        RECT 68.925 84.665 69.215 85.390 ;
        RECT 69.390 84.835 69.645 85.405 ;
        RECT 69.815 85.235 70.745 85.405 ;
        RECT 70.915 86.195 71.925 86.365 ;
        RECT 70.915 85.395 71.085 86.195 ;
        RECT 71.290 85.855 71.565 85.995 ;
        RECT 71.285 85.685 71.565 85.855 ;
        RECT 70.570 85.200 70.745 85.235 ;
        RECT 69.815 84.665 70.145 85.065 ;
        RECT 70.570 84.835 71.100 85.200 ;
        RECT 71.290 84.835 71.565 85.685 ;
        RECT 71.735 84.835 71.925 86.195 ;
        RECT 72.095 86.210 72.265 86.875 ;
        RECT 72.435 86.455 72.605 87.215 ;
        RECT 72.840 86.455 73.355 86.865 ;
        RECT 72.095 86.020 72.845 86.210 ;
        RECT 73.015 85.645 73.355 86.455 ;
        RECT 73.615 86.285 73.785 87.045 ;
        RECT 74.000 86.455 74.330 87.215 ;
        RECT 73.615 86.115 74.330 86.285 ;
        RECT 74.500 86.140 74.755 87.045 ;
        RECT 72.125 85.475 73.355 85.645 ;
        RECT 73.525 85.565 73.880 85.935 ;
        RECT 74.160 85.905 74.330 86.115 ;
        RECT 74.160 85.575 74.415 85.905 ;
        RECT 72.105 84.665 72.615 85.200 ;
        RECT 72.835 84.870 73.080 85.475 ;
        RECT 74.160 85.385 74.330 85.575 ;
        RECT 74.585 85.410 74.755 86.140 ;
        RECT 74.930 86.065 75.190 87.215 ;
        RECT 76.290 86.065 76.550 87.215 ;
        RECT 76.725 86.140 76.980 87.045 ;
        RECT 77.150 86.455 77.480 87.215 ;
        RECT 77.695 86.285 77.865 87.045 ;
        RECT 73.615 85.215 74.330 85.385 ;
        RECT 73.615 84.835 73.785 85.215 ;
        RECT 74.000 84.665 74.330 85.045 ;
        RECT 74.500 84.835 74.755 85.410 ;
        RECT 74.930 84.665 75.190 85.505 ;
        RECT 76.290 84.665 76.550 85.505 ;
        RECT 76.725 85.410 76.895 86.140 ;
        RECT 77.150 86.115 77.865 86.285 ;
        RECT 78.215 86.285 78.385 87.045 ;
        RECT 78.600 86.455 78.930 87.215 ;
        RECT 78.215 86.115 78.930 86.285 ;
        RECT 79.100 86.140 79.355 87.045 ;
        RECT 77.150 85.905 77.320 86.115 ;
        RECT 77.065 85.575 77.320 85.905 ;
        RECT 76.725 84.835 76.980 85.410 ;
        RECT 77.150 85.385 77.320 85.575 ;
        RECT 77.600 85.565 77.955 85.935 ;
        RECT 78.125 85.565 78.480 85.935 ;
        RECT 78.760 85.905 78.930 86.115 ;
        RECT 78.760 85.575 79.015 85.905 ;
        RECT 78.760 85.385 78.930 85.575 ;
        RECT 79.185 85.410 79.355 86.140 ;
        RECT 79.530 86.065 79.790 87.215 ;
        RECT 80.055 86.285 80.225 87.045 ;
        RECT 80.440 86.455 80.770 87.215 ;
        RECT 80.055 86.115 80.770 86.285 ;
        RECT 80.940 86.140 81.195 87.045 ;
        RECT 79.965 85.565 80.320 85.935 ;
        RECT 80.600 85.905 80.770 86.115 ;
        RECT 80.600 85.575 80.855 85.905 ;
        RECT 77.150 85.215 77.865 85.385 ;
        RECT 77.150 84.665 77.480 85.045 ;
        RECT 77.695 84.835 77.865 85.215 ;
        RECT 78.215 85.215 78.930 85.385 ;
        RECT 78.215 84.835 78.385 85.215 ;
        RECT 78.600 84.665 78.930 85.045 ;
        RECT 79.100 84.835 79.355 85.410 ;
        RECT 79.530 84.665 79.790 85.505 ;
        RECT 80.600 85.385 80.770 85.575 ;
        RECT 81.025 85.410 81.195 86.140 ;
        RECT 81.370 86.065 81.630 87.215 ;
        RECT 81.805 86.050 82.095 87.215 ;
        RECT 82.265 86.125 83.475 87.215 ;
        RECT 83.735 86.595 83.905 87.025 ;
        RECT 84.075 86.765 84.405 87.215 ;
        RECT 83.735 86.365 84.410 86.595 ;
        RECT 80.055 85.215 80.770 85.385 ;
        RECT 80.055 84.835 80.225 85.215 ;
        RECT 80.440 84.665 80.770 85.045 ;
        RECT 80.940 84.835 81.195 85.410 ;
        RECT 81.370 84.665 81.630 85.505 ;
        RECT 82.265 85.415 82.785 85.955 ;
        RECT 82.955 85.585 83.475 86.125 ;
        RECT 81.805 84.665 82.095 85.390 ;
        RECT 82.265 84.665 83.475 85.415 ;
        RECT 83.705 85.345 84.005 86.195 ;
        RECT 84.175 85.715 84.410 86.365 ;
        RECT 84.580 86.055 84.865 87.000 ;
        RECT 85.045 86.745 85.730 87.215 ;
        RECT 85.040 86.225 85.735 86.535 ;
        RECT 85.910 86.160 86.215 86.945 ;
        RECT 87.415 86.595 87.585 87.025 ;
        RECT 87.755 86.765 88.085 87.215 ;
        RECT 87.415 86.365 88.090 86.595 ;
        RECT 84.580 85.905 85.440 86.055 ;
        RECT 84.580 85.885 85.865 85.905 ;
        RECT 84.175 85.385 84.710 85.715 ;
        RECT 84.880 85.525 85.865 85.885 ;
        RECT 84.175 85.235 84.395 85.385 ;
        RECT 83.650 84.665 83.985 85.170 ;
        RECT 84.155 84.860 84.395 85.235 ;
        RECT 84.880 85.190 85.050 85.525 ;
        RECT 86.040 85.355 86.215 86.160 ;
        RECT 84.675 84.995 85.050 85.190 ;
        RECT 84.675 84.850 84.845 84.995 ;
        RECT 85.410 84.665 85.805 85.160 ;
        RECT 85.975 84.835 86.215 85.355 ;
        RECT 87.385 85.345 87.685 86.195 ;
        RECT 87.855 85.715 88.090 86.365 ;
        RECT 88.260 86.055 88.545 87.000 ;
        RECT 88.725 86.745 89.410 87.215 ;
        RECT 88.720 86.225 89.415 86.535 ;
        RECT 89.590 86.160 89.895 86.945 ;
        RECT 88.260 85.905 89.120 86.055 ;
        RECT 88.260 85.885 89.545 85.905 ;
        RECT 87.855 85.385 88.390 85.715 ;
        RECT 88.560 85.525 89.545 85.885 ;
        RECT 87.855 85.235 88.075 85.385 ;
        RECT 87.330 84.665 87.665 85.170 ;
        RECT 87.835 84.860 88.075 85.235 ;
        RECT 88.560 85.190 88.730 85.525 ;
        RECT 89.720 85.355 89.895 86.160 ;
        RECT 90.090 86.065 90.350 87.215 ;
        RECT 90.525 86.140 90.780 87.045 ;
        RECT 90.950 86.455 91.280 87.215 ;
        RECT 91.495 86.285 91.665 87.045 ;
        RECT 88.355 84.995 88.730 85.190 ;
        RECT 88.355 84.850 88.525 84.995 ;
        RECT 89.090 84.665 89.485 85.160 ;
        RECT 89.655 84.835 89.895 85.355 ;
        RECT 90.090 84.665 90.350 85.505 ;
        RECT 90.525 85.410 90.695 86.140 ;
        RECT 90.950 86.115 91.665 86.285 ;
        RECT 92.015 86.285 92.185 87.045 ;
        RECT 92.400 86.455 92.730 87.215 ;
        RECT 92.015 86.115 92.730 86.285 ;
        RECT 92.900 86.140 93.155 87.045 ;
        RECT 90.950 85.905 91.120 86.115 ;
        RECT 90.865 85.575 91.120 85.905 ;
        RECT 90.525 84.835 90.780 85.410 ;
        RECT 90.950 85.385 91.120 85.575 ;
        RECT 91.400 85.565 91.755 85.935 ;
        RECT 91.925 85.565 92.280 85.935 ;
        RECT 92.560 85.905 92.730 86.115 ;
        RECT 92.560 85.575 92.815 85.905 ;
        RECT 92.560 85.385 92.730 85.575 ;
        RECT 92.985 85.410 93.155 86.140 ;
        RECT 93.330 86.065 93.590 87.215 ;
        RECT 94.685 86.050 94.975 87.215 ;
        RECT 95.235 86.285 95.405 87.045 ;
        RECT 95.620 86.455 95.950 87.215 ;
        RECT 95.235 86.115 95.950 86.285 ;
        RECT 96.120 86.140 96.375 87.045 ;
        RECT 95.145 85.565 95.500 85.935 ;
        RECT 95.780 85.905 95.950 86.115 ;
        RECT 95.780 85.575 96.035 85.905 ;
        RECT 90.950 85.215 91.665 85.385 ;
        RECT 90.950 84.665 91.280 85.045 ;
        RECT 91.495 84.835 91.665 85.215 ;
        RECT 92.015 85.215 92.730 85.385 ;
        RECT 92.015 84.835 92.185 85.215 ;
        RECT 92.400 84.665 92.730 85.045 ;
        RECT 92.900 84.835 93.155 85.410 ;
        RECT 93.330 84.665 93.590 85.505 ;
        RECT 94.685 84.665 94.975 85.390 ;
        RECT 95.780 85.385 95.950 85.575 ;
        RECT 96.205 85.410 96.375 86.140 ;
        RECT 96.550 86.065 96.810 87.215 ;
        RECT 97.075 86.285 97.245 87.045 ;
        RECT 97.460 86.455 97.790 87.215 ;
        RECT 97.075 86.115 97.790 86.285 ;
        RECT 97.960 86.140 98.215 87.045 ;
        RECT 96.985 85.565 97.340 85.935 ;
        RECT 97.620 85.905 97.790 86.115 ;
        RECT 97.620 85.575 97.875 85.905 ;
        RECT 95.235 85.215 95.950 85.385 ;
        RECT 95.235 84.835 95.405 85.215 ;
        RECT 95.620 84.665 95.950 85.045 ;
        RECT 96.120 84.835 96.375 85.410 ;
        RECT 96.550 84.665 96.810 85.505 ;
        RECT 97.620 85.385 97.790 85.575 ;
        RECT 98.045 85.410 98.215 86.140 ;
        RECT 98.390 86.065 98.650 87.215 ;
        RECT 99.290 86.065 99.550 87.215 ;
        RECT 99.725 86.140 99.980 87.045 ;
        RECT 100.150 86.455 100.480 87.215 ;
        RECT 100.695 86.285 100.865 87.045 ;
        RECT 97.075 85.215 97.790 85.385 ;
        RECT 97.075 84.835 97.245 85.215 ;
        RECT 97.460 84.665 97.790 85.045 ;
        RECT 97.960 84.835 98.215 85.410 ;
        RECT 98.390 84.665 98.650 85.505 ;
        RECT 99.290 84.665 99.550 85.505 ;
        RECT 99.725 85.410 99.895 86.140 ;
        RECT 100.150 86.115 100.865 86.285 ;
        RECT 101.125 86.125 102.335 87.215 ;
        RECT 100.150 85.905 100.320 86.115 ;
        RECT 100.065 85.575 100.320 85.905 ;
        RECT 99.725 84.835 99.980 85.410 ;
        RECT 100.150 85.385 100.320 85.575 ;
        RECT 100.600 85.565 100.955 85.935 ;
        RECT 101.125 85.415 101.645 85.955 ;
        RECT 101.815 85.585 102.335 86.125 ;
        RECT 102.510 86.065 102.770 87.215 ;
        RECT 102.945 86.140 103.200 87.045 ;
        RECT 103.370 86.455 103.700 87.215 ;
        RECT 103.915 86.285 104.085 87.045 ;
        RECT 100.150 85.215 100.865 85.385 ;
        RECT 100.150 84.665 100.480 85.045 ;
        RECT 100.695 84.835 100.865 85.215 ;
        RECT 101.125 84.665 102.335 85.415 ;
        RECT 102.510 84.665 102.770 85.505 ;
        RECT 102.945 85.410 103.115 86.140 ;
        RECT 103.370 86.115 104.085 86.285 ;
        RECT 104.345 86.125 105.555 87.215 ;
        RECT 103.370 85.905 103.540 86.115 ;
        RECT 103.285 85.575 103.540 85.905 ;
        RECT 102.945 84.835 103.200 85.410 ;
        RECT 103.370 85.385 103.540 85.575 ;
        RECT 103.820 85.565 104.175 85.935 ;
        RECT 104.345 85.415 104.865 85.955 ;
        RECT 105.035 85.585 105.555 86.125 ;
        RECT 105.730 86.065 105.990 87.215 ;
        RECT 106.165 86.140 106.420 87.045 ;
        RECT 106.590 86.455 106.920 87.215 ;
        RECT 107.135 86.285 107.305 87.045 ;
        RECT 103.370 85.215 104.085 85.385 ;
        RECT 103.370 84.665 103.700 85.045 ;
        RECT 103.915 84.835 104.085 85.215 ;
        RECT 104.345 84.665 105.555 85.415 ;
        RECT 105.730 84.665 105.990 85.505 ;
        RECT 106.165 85.410 106.335 86.140 ;
        RECT 106.590 86.115 107.305 86.285 ;
        RECT 106.590 85.905 106.760 86.115 ;
        RECT 107.565 86.050 107.855 87.215 ;
        RECT 108.950 86.065 109.210 87.215 ;
        RECT 109.385 86.140 109.640 87.045 ;
        RECT 109.810 86.455 110.140 87.215 ;
        RECT 110.355 86.285 110.525 87.045 ;
        RECT 106.505 85.575 106.760 85.905 ;
        RECT 106.165 84.835 106.420 85.410 ;
        RECT 106.590 85.385 106.760 85.575 ;
        RECT 107.040 85.565 107.395 85.935 ;
        RECT 106.590 85.215 107.305 85.385 ;
        RECT 106.590 84.665 106.920 85.045 ;
        RECT 107.135 84.835 107.305 85.215 ;
        RECT 107.565 84.665 107.855 85.390 ;
        RECT 108.950 84.665 109.210 85.505 ;
        RECT 109.385 85.410 109.555 86.140 ;
        RECT 109.810 86.115 110.525 86.285 ;
        RECT 110.785 86.125 111.995 87.215 ;
        RECT 109.810 85.905 109.980 86.115 ;
        RECT 109.725 85.575 109.980 85.905 ;
        RECT 109.385 84.835 109.640 85.410 ;
        RECT 109.810 85.385 109.980 85.575 ;
        RECT 110.260 85.565 110.615 85.935 ;
        RECT 110.785 85.415 111.305 85.955 ;
        RECT 111.475 85.585 111.995 86.125 ;
        RECT 112.170 86.065 112.430 87.215 ;
        RECT 112.605 86.140 112.860 87.045 ;
        RECT 113.030 86.455 113.360 87.215 ;
        RECT 113.575 86.285 113.745 87.045 ;
        RECT 114.095 86.595 114.265 87.025 ;
        RECT 114.435 86.765 114.765 87.215 ;
        RECT 114.095 86.365 114.770 86.595 ;
        RECT 109.810 85.215 110.525 85.385 ;
        RECT 109.810 84.665 110.140 85.045 ;
        RECT 110.355 84.835 110.525 85.215 ;
        RECT 110.785 84.665 111.995 85.415 ;
        RECT 112.170 84.665 112.430 85.505 ;
        RECT 112.605 85.410 112.775 86.140 ;
        RECT 113.030 86.115 113.745 86.285 ;
        RECT 113.030 85.905 113.200 86.115 ;
        RECT 112.945 85.575 113.200 85.905 ;
        RECT 112.605 84.835 112.860 85.410 ;
        RECT 113.030 85.385 113.200 85.575 ;
        RECT 113.480 85.565 113.835 85.935 ;
        RECT 113.030 85.215 113.745 85.385 ;
        RECT 114.065 85.345 114.365 86.195 ;
        RECT 114.535 85.715 114.770 86.365 ;
        RECT 114.940 86.055 115.225 87.000 ;
        RECT 115.405 86.745 116.090 87.215 ;
        RECT 115.400 86.225 116.095 86.535 ;
        RECT 116.270 86.160 116.575 86.945 ;
        RECT 114.940 85.905 115.800 86.055 ;
        RECT 114.940 85.885 116.225 85.905 ;
        RECT 114.535 85.385 115.070 85.715 ;
        RECT 115.240 85.525 116.225 85.885 ;
        RECT 114.535 85.235 114.755 85.385 ;
        RECT 113.030 84.665 113.360 85.045 ;
        RECT 113.575 84.835 113.745 85.215 ;
        RECT 114.010 84.665 114.345 85.170 ;
        RECT 114.515 84.860 114.755 85.235 ;
        RECT 115.240 85.190 115.410 85.525 ;
        RECT 116.400 85.355 116.575 86.160 ;
        RECT 115.035 84.995 115.410 85.190 ;
        RECT 115.035 84.850 115.205 84.995 ;
        RECT 115.770 84.665 116.165 85.160 ;
        RECT 116.335 84.835 116.575 85.355 ;
        RECT 117.225 86.365 117.485 87.045 ;
        RECT 117.655 86.435 117.905 87.215 ;
        RECT 118.155 86.665 118.405 87.045 ;
        RECT 118.575 86.835 118.930 87.215 ;
        RECT 119.935 86.825 120.270 87.045 ;
        RECT 119.535 86.665 119.765 86.705 ;
        RECT 118.155 86.465 119.765 86.665 ;
        RECT 118.155 86.455 118.990 86.465 ;
        RECT 119.580 86.375 119.765 86.465 ;
        RECT 117.225 85.165 117.395 86.365 ;
        RECT 119.095 86.265 119.425 86.295 ;
        RECT 117.625 86.205 119.425 86.265 ;
        RECT 120.015 86.205 120.270 86.825 ;
        RECT 117.565 86.095 120.270 86.205 ;
        RECT 117.565 86.060 117.765 86.095 ;
        RECT 117.565 85.485 117.735 86.060 ;
        RECT 119.095 86.035 120.270 86.095 ;
        RECT 120.445 86.050 120.735 87.215 ;
        RECT 120.995 86.285 121.165 87.045 ;
        RECT 121.380 86.455 121.710 87.215 ;
        RECT 120.995 86.115 121.710 86.285 ;
        RECT 121.880 86.140 122.135 87.045 ;
        RECT 117.965 85.620 118.375 85.925 ;
        RECT 118.545 85.655 118.875 85.865 ;
        RECT 117.565 85.365 117.835 85.485 ;
        RECT 117.565 85.320 118.410 85.365 ;
        RECT 117.655 85.195 118.410 85.320 ;
        RECT 118.665 85.255 118.875 85.655 ;
        RECT 119.120 85.655 119.595 85.865 ;
        RECT 119.785 85.655 120.275 85.855 ;
        RECT 119.120 85.255 119.340 85.655 ;
        RECT 120.905 85.565 121.260 85.935 ;
        RECT 121.540 85.905 121.710 86.115 ;
        RECT 121.540 85.575 121.795 85.905 ;
        RECT 117.225 84.835 117.485 85.165 ;
        RECT 118.240 85.045 118.410 85.195 ;
        RECT 117.655 84.665 117.985 85.025 ;
        RECT 118.240 84.835 119.540 85.045 ;
        RECT 119.815 84.665 120.270 85.430 ;
        RECT 120.445 84.665 120.735 85.390 ;
        RECT 121.540 85.385 121.710 85.575 ;
        RECT 121.965 85.410 122.135 86.140 ;
        RECT 122.310 86.065 122.570 87.215 ;
        RECT 122.835 86.285 123.005 87.045 ;
        RECT 123.220 86.455 123.550 87.215 ;
        RECT 122.835 86.115 123.550 86.285 ;
        RECT 123.720 86.140 123.975 87.045 ;
        RECT 122.745 85.565 123.100 85.935 ;
        RECT 123.380 85.905 123.550 86.115 ;
        RECT 123.380 85.575 123.635 85.905 ;
        RECT 120.995 85.215 121.710 85.385 ;
        RECT 120.995 84.835 121.165 85.215 ;
        RECT 121.380 84.665 121.710 85.045 ;
        RECT 121.880 84.835 122.135 85.410 ;
        RECT 122.310 84.665 122.570 85.505 ;
        RECT 123.380 85.385 123.550 85.575 ;
        RECT 123.805 85.410 123.975 86.140 ;
        RECT 124.150 86.065 124.410 87.215 ;
        RECT 124.590 86.065 124.850 87.215 ;
        RECT 125.025 86.140 125.280 87.045 ;
        RECT 125.450 86.455 125.780 87.215 ;
        RECT 125.995 86.285 126.165 87.045 ;
        RECT 122.835 85.215 123.550 85.385 ;
        RECT 122.835 84.835 123.005 85.215 ;
        RECT 123.220 84.665 123.550 85.045 ;
        RECT 123.720 84.835 123.975 85.410 ;
        RECT 124.150 84.665 124.410 85.505 ;
        RECT 124.590 84.665 124.850 85.505 ;
        RECT 125.025 85.410 125.195 86.140 ;
        RECT 125.450 86.115 126.165 86.285 ;
        RECT 126.425 86.455 126.940 86.865 ;
        RECT 127.175 86.455 127.345 87.215 ;
        RECT 127.515 86.875 129.545 87.045 ;
        RECT 125.450 85.905 125.620 86.115 ;
        RECT 125.365 85.575 125.620 85.905 ;
        RECT 125.025 84.835 125.280 85.410 ;
        RECT 125.450 85.385 125.620 85.575 ;
        RECT 125.900 85.565 126.255 85.935 ;
        RECT 126.425 85.645 126.765 86.455 ;
        RECT 127.515 86.210 127.685 86.875 ;
        RECT 128.080 86.535 129.205 86.705 ;
        RECT 126.935 86.020 127.685 86.210 ;
        RECT 127.855 86.195 128.865 86.365 ;
        RECT 126.425 85.475 127.655 85.645 ;
        RECT 125.450 85.215 126.165 85.385 ;
        RECT 125.450 84.665 125.780 85.045 ;
        RECT 125.995 84.835 126.165 85.215 ;
        RECT 126.700 84.870 126.945 85.475 ;
        RECT 127.165 84.665 127.675 85.200 ;
        RECT 127.855 84.835 128.045 86.195 ;
        RECT 128.215 85.175 128.490 85.995 ;
        RECT 128.695 85.395 128.865 86.195 ;
        RECT 129.035 85.405 129.205 86.535 ;
        RECT 129.375 85.905 129.545 86.875 ;
        RECT 129.715 86.075 129.885 87.215 ;
        RECT 130.055 86.075 130.390 87.045 ;
        RECT 130.655 86.285 130.825 87.045 ;
        RECT 131.040 86.455 131.370 87.215 ;
        RECT 130.655 86.115 131.370 86.285 ;
        RECT 131.540 86.140 131.795 87.045 ;
        RECT 129.375 85.575 129.570 85.905 ;
        RECT 129.795 85.575 130.050 85.905 ;
        RECT 129.795 85.405 129.965 85.575 ;
        RECT 130.220 85.405 130.390 86.075 ;
        RECT 130.565 85.565 130.920 85.935 ;
        RECT 131.200 85.905 131.370 86.115 ;
        RECT 131.200 85.575 131.455 85.905 ;
        RECT 129.035 85.235 129.965 85.405 ;
        RECT 129.035 85.200 129.210 85.235 ;
        RECT 128.215 85.005 128.495 85.175 ;
        RECT 128.215 84.835 128.490 85.005 ;
        RECT 128.680 84.835 129.210 85.200 ;
        RECT 129.635 84.665 129.965 85.065 ;
        RECT 130.135 84.835 130.390 85.405 ;
        RECT 131.200 85.385 131.370 85.575 ;
        RECT 131.625 85.410 131.795 86.140 ;
        RECT 131.970 86.065 132.230 87.215 ;
        RECT 133.325 86.050 133.615 87.215 ;
        RECT 133.805 86.375 134.060 87.045 ;
        RECT 134.230 86.455 134.560 87.215 ;
        RECT 134.730 86.615 134.980 87.045 ;
        RECT 135.150 86.795 135.505 87.215 ;
        RECT 135.695 86.875 136.865 87.045 ;
        RECT 135.695 86.835 136.025 86.875 ;
        RECT 136.135 86.615 136.365 86.705 ;
        RECT 134.730 86.375 136.365 86.615 ;
        RECT 136.535 86.375 136.865 86.875 ;
        RECT 130.655 85.215 131.370 85.385 ;
        RECT 130.655 84.835 130.825 85.215 ;
        RECT 131.040 84.665 131.370 85.045 ;
        RECT 131.540 84.835 131.795 85.410 ;
        RECT 131.970 84.665 132.230 85.505 ;
        RECT 133.325 84.665 133.615 85.390 ;
        RECT 133.805 85.245 133.975 86.375 ;
        RECT 137.035 86.205 137.205 87.045 ;
        RECT 137.555 86.595 137.725 87.025 ;
        RECT 137.895 86.765 138.225 87.215 ;
        RECT 137.555 86.365 138.230 86.595 ;
        RECT 134.145 86.035 137.205 86.205 ;
        RECT 134.145 85.485 134.315 86.035 ;
        RECT 134.535 85.685 134.910 85.855 ;
        RECT 134.545 85.655 134.910 85.685 ;
        RECT 135.080 85.655 135.410 85.855 ;
        RECT 134.145 85.315 134.945 85.485 ;
        RECT 133.805 85.165 133.990 85.245 ;
        RECT 133.805 84.835 134.060 85.165 ;
        RECT 134.275 84.665 134.605 85.145 ;
        RECT 134.775 85.085 134.945 85.315 ;
        RECT 135.125 85.255 135.410 85.655 ;
        RECT 135.680 85.655 136.155 85.855 ;
        RECT 136.325 85.655 136.770 85.855 ;
        RECT 136.940 85.655 137.290 85.865 ;
        RECT 135.680 85.255 135.960 85.655 ;
        RECT 136.140 85.315 137.205 85.485 ;
        RECT 137.525 85.345 137.825 86.195 ;
        RECT 137.995 85.715 138.230 86.365 ;
        RECT 138.400 86.055 138.685 87.000 ;
        RECT 138.865 86.745 139.550 87.215 ;
        RECT 138.860 86.225 139.555 86.535 ;
        RECT 139.730 86.160 140.035 86.945 ;
        RECT 138.400 85.905 139.260 86.055 ;
        RECT 138.400 85.885 139.685 85.905 ;
        RECT 137.995 85.385 138.530 85.715 ;
        RECT 138.700 85.525 139.685 85.885 ;
        RECT 136.140 85.085 136.310 85.315 ;
        RECT 134.775 84.835 136.310 85.085 ;
        RECT 136.535 84.665 136.865 85.145 ;
        RECT 137.035 84.835 137.205 85.315 ;
        RECT 137.995 85.235 138.215 85.385 ;
        RECT 137.470 84.665 137.805 85.170 ;
        RECT 137.975 84.860 138.215 85.235 ;
        RECT 138.700 85.190 138.870 85.525 ;
        RECT 139.860 85.355 140.035 86.160 ;
        RECT 140.315 86.285 140.485 87.045 ;
        RECT 140.700 86.455 141.030 87.215 ;
        RECT 140.315 86.115 141.030 86.285 ;
        RECT 141.200 86.140 141.455 87.045 ;
        RECT 140.225 85.565 140.580 85.935 ;
        RECT 140.860 85.905 141.030 86.115 ;
        RECT 140.860 85.575 141.115 85.905 ;
        RECT 140.860 85.385 141.030 85.575 ;
        RECT 141.285 85.410 141.455 86.140 ;
        RECT 141.630 86.065 141.890 87.215 ;
        RECT 142.155 86.285 142.325 87.045 ;
        RECT 142.540 86.455 142.870 87.215 ;
        RECT 142.155 86.115 142.870 86.285 ;
        RECT 143.040 86.140 143.295 87.045 ;
        RECT 142.065 85.565 142.420 85.935 ;
        RECT 142.700 85.905 142.870 86.115 ;
        RECT 142.700 85.575 142.955 85.905 ;
        RECT 138.495 84.995 138.870 85.190 ;
        RECT 138.495 84.850 138.665 84.995 ;
        RECT 139.230 84.665 139.625 85.160 ;
        RECT 139.795 84.835 140.035 85.355 ;
        RECT 140.315 85.215 141.030 85.385 ;
        RECT 140.315 84.835 140.485 85.215 ;
        RECT 140.700 84.665 141.030 85.045 ;
        RECT 141.200 84.835 141.455 85.410 ;
        RECT 141.630 84.665 141.890 85.505 ;
        RECT 142.700 85.385 142.870 85.575 ;
        RECT 143.125 85.410 143.295 86.140 ;
        RECT 143.470 86.065 143.730 87.215 ;
        RECT 143.995 86.285 144.165 87.045 ;
        RECT 144.380 86.455 144.710 87.215 ;
        RECT 143.995 86.115 144.710 86.285 ;
        RECT 144.880 86.140 145.135 87.045 ;
        RECT 143.905 85.565 144.260 85.935 ;
        RECT 144.540 85.905 144.710 86.115 ;
        RECT 144.540 85.575 144.795 85.905 ;
        RECT 142.155 85.215 142.870 85.385 ;
        RECT 142.155 84.835 142.325 85.215 ;
        RECT 142.540 84.665 142.870 85.045 ;
        RECT 143.040 84.835 143.295 85.410 ;
        RECT 143.470 84.665 143.730 85.505 ;
        RECT 144.540 85.385 144.710 85.575 ;
        RECT 144.965 85.410 145.135 86.140 ;
        RECT 145.310 86.065 145.570 87.215 ;
        RECT 145.745 86.125 146.955 87.215 ;
        RECT 145.745 85.585 146.265 86.125 ;
        RECT 143.995 85.215 144.710 85.385 ;
        RECT 143.995 84.835 144.165 85.215 ;
        RECT 144.380 84.665 144.710 85.045 ;
        RECT 144.880 84.835 145.135 85.410 ;
        RECT 145.310 84.665 145.570 85.505 ;
        RECT 146.435 85.415 146.955 85.955 ;
        RECT 145.745 84.665 146.955 85.415 ;
        RECT 17.320 84.495 147.040 84.665 ;
      LAYER met1 ;
        RECT 7.615 222.450 39.790 222.970 ;
        RECT 0.510 219.970 39.790 222.450 ;
        RECT 0.510 7.020 2.990 219.970 ;
        RECT 7.615 219.860 39.790 219.970 ;
        RECT 7.615 7.555 10.725 219.860 ;
        RECT 17.320 212.180 147.040 212.660 ;
        RECT 79.490 211.640 79.810 211.700 ;
        RECT 80.425 211.640 80.715 211.685 ;
        RECT 79.490 211.500 80.715 211.640 ;
        RECT 79.490 211.440 79.810 211.500 ;
        RECT 80.425 211.455 80.715 211.500 ;
        RECT 84.105 211.640 84.395 211.685 ;
        RECT 87.770 211.640 88.090 211.700 ;
        RECT 84.105 211.500 88.090 211.640 ;
        RECT 84.105 211.455 84.395 211.500 ;
        RECT 87.770 211.440 88.090 211.500 ;
        RECT 95.590 211.640 95.910 211.700 ;
        RECT 96.525 211.640 96.815 211.685 ;
        RECT 95.590 211.500 96.815 211.640 ;
        RECT 95.590 211.440 95.910 211.500 ;
        RECT 96.525 211.455 96.815 211.500 ;
        RECT 85.930 211.300 86.250 211.360 ;
        RECT 85.930 211.160 88.000 211.300 ;
        RECT 85.930 211.100 86.250 211.160 ;
        RECT 60.170 210.960 60.490 211.020 ;
        RECT 60.645 210.960 60.935 211.005 ;
        RECT 60.170 210.820 60.935 210.960 ;
        RECT 60.170 210.760 60.490 210.820 ;
        RECT 60.645 210.775 60.935 210.820 ;
        RECT 81.345 210.775 81.635 211.005 ;
        RECT 82.710 210.960 83.030 211.020 ;
        RECT 83.185 210.960 83.475 211.005 ;
        RECT 82.710 210.820 83.475 210.960 ;
        RECT 51.890 210.620 52.210 210.680 ;
        RECT 62.025 210.620 62.315 210.665 ;
        RECT 51.890 210.480 62.315 210.620 ;
        RECT 81.420 210.620 81.560 210.775 ;
        RECT 82.710 210.760 83.030 210.820 ;
        RECT 83.185 210.775 83.475 210.820 ;
        RECT 86.405 210.775 86.695 211.005 ;
        RECT 84.550 210.620 84.870 210.680 ;
        RECT 81.420 210.480 84.870 210.620 ;
        RECT 86.480 210.620 86.620 210.775 ;
        RECT 87.310 210.760 87.630 211.020 ;
        RECT 87.860 211.005 88.000 211.160 ;
        RECT 87.785 210.775 88.075 211.005 ;
        RECT 89.150 210.960 89.470 211.020 ;
        RECT 90.545 210.960 90.835 211.005 ;
        RECT 89.150 210.820 90.835 210.960 ;
        RECT 89.150 210.760 89.470 210.820 ;
        RECT 90.545 210.775 90.835 210.820 ;
        RECT 97.445 210.960 97.735 211.005 ;
        RECT 103.410 210.960 103.730 211.020 ;
        RECT 97.445 210.820 103.730 210.960 ;
        RECT 97.445 210.775 97.735 210.820 ;
        RECT 103.410 210.760 103.730 210.820 ;
        RECT 89.610 210.620 89.930 210.680 ;
        RECT 86.480 210.480 89.930 210.620 ;
        RECT 51.890 210.420 52.210 210.480 ;
        RECT 62.025 210.435 62.315 210.480 ;
        RECT 84.550 210.420 84.870 210.480 ;
        RECT 89.610 210.420 89.930 210.480 ;
        RECT 85.470 210.080 85.790 210.340 ;
        RECT 88.230 210.280 88.550 210.340 ;
        RECT 88.705 210.280 88.995 210.325 ;
        RECT 88.230 210.140 88.995 210.280 ;
        RECT 88.230 210.080 88.550 210.140 ;
        RECT 88.705 210.095 88.995 210.140 ;
        RECT 90.990 210.080 91.310 210.340 ;
        RECT 17.320 209.460 147.040 209.940 ;
        RECT 55.110 209.260 55.430 209.320 ;
        RECT 55.110 209.120 70.520 209.260 ;
        RECT 55.110 209.060 55.430 209.120 ;
        RECT 60.185 208.920 60.475 208.965 ;
        RECT 64.310 208.920 64.630 208.980 ;
        RECT 67.545 208.920 67.835 208.965 ;
        RECT 53.360 208.780 58.560 208.920 ;
        RECT 53.360 208.625 53.500 208.780 ;
        RECT 53.285 208.395 53.575 208.625 ;
        RECT 53.730 208.380 54.050 208.640 ;
        RECT 54.205 208.580 54.495 208.625 ;
        RECT 55.110 208.580 55.430 208.640 ;
        RECT 54.205 208.440 55.430 208.580 ;
        RECT 54.205 208.395 54.495 208.440 ;
        RECT 55.110 208.380 55.430 208.440 ;
        RECT 55.585 208.580 55.875 208.625 ;
        RECT 58.420 208.580 58.560 208.780 ;
        RECT 60.185 208.780 61.780 208.920 ;
        RECT 60.185 208.735 60.475 208.780 ;
        RECT 60.630 208.580 60.950 208.640 ;
        RECT 61.640 208.625 61.780 208.780 ;
        RECT 64.310 208.780 67.835 208.920 ;
        RECT 64.310 208.720 64.630 208.780 ;
        RECT 67.545 208.735 67.835 208.780 ;
        RECT 55.585 208.440 58.100 208.580 ;
        RECT 58.420 208.440 60.950 208.580 ;
        RECT 55.585 208.395 55.875 208.440 ;
        RECT 52.350 208.040 52.670 208.300 ;
        RECT 56.950 208.040 57.270 208.300 ;
        RECT 57.960 208.240 58.100 208.440 ;
        RECT 60.630 208.380 60.950 208.440 ;
        RECT 61.565 208.395 61.855 208.625 ;
        RECT 67.085 208.395 67.375 208.625 ;
        RECT 61.105 208.240 61.395 208.285 ;
        RECT 57.960 208.100 61.395 208.240 ;
        RECT 61.105 208.055 61.395 208.100 ;
        RECT 55.125 207.900 55.415 207.945 ;
        RECT 60.170 207.900 60.490 207.960 ;
        RECT 67.160 207.900 67.300 208.395 ;
        RECT 68.450 208.380 68.770 208.640 ;
        RECT 68.910 208.580 69.230 208.640 ;
        RECT 70.380 208.625 70.520 209.120 ;
        RECT 89.150 209.060 89.470 209.320 ;
        RECT 89.610 209.060 89.930 209.320 ;
        RECT 93.290 209.260 93.610 209.320 ;
        RECT 90.160 209.120 93.610 209.260 ;
        RECT 69.385 208.580 69.675 208.625 ;
        RECT 68.910 208.440 69.675 208.580 ;
        RECT 68.910 208.380 69.230 208.440 ;
        RECT 69.385 208.395 69.675 208.440 ;
        RECT 70.305 208.580 70.595 208.625 ;
        RECT 70.750 208.580 71.070 208.640 ;
        RECT 70.305 208.440 71.070 208.580 ;
        RECT 70.305 208.395 70.595 208.440 ;
        RECT 70.750 208.380 71.070 208.440 ;
        RECT 81.345 208.240 81.635 208.285 ;
        RECT 82.710 208.240 83.030 208.300 ;
        RECT 81.345 208.100 83.030 208.240 ;
        RECT 81.345 208.055 81.635 208.100 ;
        RECT 82.710 208.040 83.030 208.100 ;
        RECT 85.930 208.240 86.250 208.300 ;
        RECT 90.160 208.240 90.300 209.120 ;
        RECT 93.290 209.060 93.610 209.120 ;
        RECT 97.905 209.075 98.195 209.305 ;
        RECT 90.530 208.920 90.850 208.980 ;
        RECT 95.590 208.920 95.910 208.980 ;
        RECT 96.985 208.920 97.275 208.965 ;
        RECT 90.530 208.780 91.245 208.920 ;
        RECT 90.530 208.720 90.850 208.780 ;
        RECT 91.105 208.625 91.245 208.780 ;
        RECT 92.000 208.780 97.275 208.920 ;
        RECT 91.005 208.395 91.295 208.625 ;
        RECT 92.000 208.570 92.140 208.780 ;
        RECT 95.590 208.720 95.910 208.780 ;
        RECT 96.985 208.735 97.275 208.780 ;
        RECT 97.430 208.920 97.750 208.980 ;
        RECT 97.980 208.920 98.120 209.075 ;
        RECT 102.505 208.920 102.795 208.965 ;
        RECT 97.430 208.780 102.795 208.920 ;
        RECT 91.540 208.430 92.140 208.570 ;
        RECT 91.540 208.285 91.680 208.430 ;
        RECT 93.290 208.380 93.610 208.640 ;
        RECT 94.225 208.580 94.515 208.625 ;
        RECT 96.510 208.580 96.830 208.640 ;
        RECT 94.225 208.440 96.830 208.580 ;
        RECT 97.060 208.580 97.200 208.735 ;
        RECT 97.430 208.720 97.750 208.780 ;
        RECT 102.505 208.735 102.795 208.780 ;
        RECT 103.410 208.720 103.730 208.980 ;
        RECT 100.205 208.580 100.495 208.625 ;
        RECT 97.060 208.440 100.495 208.580 ;
        RECT 94.225 208.395 94.515 208.440 ;
        RECT 96.510 208.380 96.830 208.440 ;
        RECT 100.205 208.395 100.495 208.440 ;
        RECT 90.545 208.240 90.835 208.285 ;
        RECT 85.930 208.100 90.835 208.240 ;
        RECT 85.930 208.040 86.250 208.100 ;
        RECT 90.545 208.055 90.835 208.100 ;
        RECT 91.465 208.055 91.755 208.285 ;
        RECT 91.925 208.055 92.215 208.285 ;
        RECT 93.765 208.240 94.055 208.285 ;
        RECT 98.810 208.240 99.130 208.300 ;
        RECT 99.745 208.240 100.035 208.285 ;
        RECT 93.765 208.100 100.035 208.240 ;
        RECT 93.765 208.055 94.055 208.100 ;
        RECT 92.000 207.900 92.140 208.055 ;
        RECT 98.810 208.040 99.130 208.100 ;
        RECT 99.745 208.055 100.035 208.100 ;
        RECT 55.125 207.760 67.300 207.900 ;
        RECT 91.080 207.760 92.140 207.900 ;
        RECT 95.145 207.900 95.435 207.945 ;
        RECT 96.510 207.900 96.830 207.960 ;
        RECT 95.145 207.760 96.830 207.900 ;
        RECT 55.125 207.715 55.415 207.760 ;
        RECT 60.170 207.700 60.490 207.760 ;
        RECT 53.745 207.560 54.035 207.605 ;
        RECT 54.190 207.560 54.510 207.620 ;
        RECT 53.745 207.420 54.510 207.560 ;
        RECT 53.745 207.375 54.035 207.420 ;
        RECT 54.190 207.360 54.510 207.420 ;
        RECT 55.570 207.360 55.890 207.620 ;
        RECT 65.230 207.560 65.550 207.620 ;
        RECT 68.465 207.560 68.755 207.605 ;
        RECT 65.230 207.420 68.755 207.560 ;
        RECT 65.230 207.360 65.550 207.420 ;
        RECT 68.465 207.375 68.755 207.420 ;
        RECT 69.370 207.360 69.690 207.620 ;
        RECT 71.670 207.560 71.990 207.620 ;
        RECT 84.105 207.560 84.395 207.605 ;
        RECT 91.080 207.560 91.220 207.760 ;
        RECT 95.145 207.715 95.435 207.760 ;
        RECT 96.510 207.700 96.830 207.760 ;
        RECT 102.045 207.900 102.335 207.945 ;
        RECT 106.630 207.900 106.950 207.960 ;
        RECT 102.045 207.760 106.950 207.900 ;
        RECT 102.045 207.715 102.335 207.760 ;
        RECT 106.630 207.700 106.950 207.760 ;
        RECT 71.670 207.420 91.220 207.560 ;
        RECT 93.290 207.560 93.610 207.620 ;
        RECT 96.985 207.560 97.275 207.605 ;
        RECT 93.290 207.420 97.275 207.560 ;
        RECT 71.670 207.360 71.990 207.420 ;
        RECT 84.105 207.375 84.395 207.420 ;
        RECT 93.290 207.360 93.610 207.420 ;
        RECT 96.985 207.375 97.275 207.420 ;
        RECT 104.330 207.360 104.650 207.620 ;
        RECT 17.320 206.740 147.040 207.220 ;
        RECT 56.505 206.540 56.795 206.585 ;
        RECT 56.950 206.540 57.270 206.600 ;
        RECT 56.505 206.400 57.270 206.540 ;
        RECT 56.505 206.355 56.795 206.400 ;
        RECT 56.950 206.340 57.270 206.400 ;
        RECT 89.610 206.540 89.930 206.600 ;
        RECT 97.430 206.540 97.750 206.600 ;
        RECT 89.610 206.400 97.750 206.540 ;
        RECT 89.610 206.340 89.930 206.400 ;
        RECT 97.430 206.340 97.750 206.400 ;
        RECT 103.410 206.540 103.730 206.600 ;
        RECT 104.345 206.540 104.635 206.585 ;
        RECT 103.410 206.400 104.635 206.540 ;
        RECT 103.410 206.340 103.730 206.400 ;
        RECT 104.345 206.355 104.635 206.400 ;
        RECT 50.970 206.200 51.290 206.260 ;
        RECT 52.825 206.200 53.115 206.245 ;
        RECT 50.970 206.060 53.115 206.200 ;
        RECT 50.970 206.000 51.290 206.060 ;
        RECT 52.825 206.015 53.115 206.060 ;
        RECT 59.250 206.200 59.540 206.245 ;
        RECT 60.820 206.200 61.110 206.245 ;
        RECT 62.920 206.200 63.210 206.245 ;
        RECT 59.250 206.060 63.210 206.200 ;
        RECT 59.250 206.015 59.540 206.060 ;
        RECT 60.820 206.015 61.110 206.060 ;
        RECT 62.920 206.015 63.210 206.060 ;
        RECT 67.070 206.200 67.360 206.245 ;
        RECT 68.640 206.200 68.930 206.245 ;
        RECT 70.740 206.200 71.030 206.245 ;
        RECT 67.070 206.060 71.030 206.200 ;
        RECT 67.070 206.015 67.360 206.060 ;
        RECT 68.640 206.015 68.930 206.060 ;
        RECT 70.740 206.015 71.030 206.060 ;
        RECT 85.470 206.200 85.760 206.245 ;
        RECT 87.040 206.200 87.330 206.245 ;
        RECT 89.140 206.200 89.430 206.245 ;
        RECT 85.470 206.060 89.430 206.200 ;
        RECT 85.470 206.015 85.760 206.060 ;
        RECT 87.040 206.015 87.330 206.060 ;
        RECT 89.140 206.015 89.430 206.060 ;
        RECT 90.570 206.200 90.860 206.245 ;
        RECT 92.670 206.200 92.960 206.245 ;
        RECT 94.240 206.200 94.530 206.245 ;
        RECT 90.570 206.060 94.530 206.200 ;
        RECT 90.570 206.015 90.860 206.060 ;
        RECT 92.670 206.015 92.960 206.060 ;
        RECT 94.240 206.015 94.530 206.060 ;
        RECT 97.930 206.200 98.220 206.245 ;
        RECT 100.030 206.200 100.320 206.245 ;
        RECT 101.600 206.200 101.890 206.245 ;
        RECT 97.930 206.060 101.890 206.200 ;
        RECT 97.930 206.015 98.220 206.060 ;
        RECT 100.030 206.015 100.320 206.060 ;
        RECT 101.600 206.015 101.890 206.060 ;
        RECT 53.270 205.860 53.590 205.920 ;
        RECT 54.205 205.860 54.495 205.905 ;
        RECT 53.270 205.720 54.495 205.860 ;
        RECT 53.270 205.660 53.590 205.720 ;
        RECT 54.205 205.675 54.495 205.720 ;
        RECT 58.815 205.860 59.105 205.905 ;
        RECT 61.335 205.860 61.625 205.905 ;
        RECT 62.525 205.860 62.815 205.905 ;
        RECT 58.815 205.720 62.815 205.860 ;
        RECT 58.815 205.675 59.105 205.720 ;
        RECT 61.335 205.675 61.625 205.720 ;
        RECT 62.525 205.675 62.815 205.720 ;
        RECT 66.635 205.860 66.925 205.905 ;
        RECT 69.155 205.860 69.445 205.905 ;
        RECT 70.345 205.860 70.635 205.905 ;
        RECT 66.635 205.720 70.635 205.860 ;
        RECT 66.635 205.675 66.925 205.720 ;
        RECT 69.155 205.675 69.445 205.720 ;
        RECT 70.345 205.675 70.635 205.720 ;
        RECT 85.035 205.860 85.325 205.905 ;
        RECT 87.555 205.860 87.845 205.905 ;
        RECT 88.745 205.860 89.035 205.905 ;
        RECT 85.035 205.720 89.035 205.860 ;
        RECT 85.035 205.675 85.325 205.720 ;
        RECT 87.555 205.675 87.845 205.720 ;
        RECT 88.745 205.675 89.035 205.720 ;
        RECT 90.965 205.860 91.255 205.905 ;
        RECT 92.155 205.860 92.445 205.905 ;
        RECT 94.675 205.860 94.965 205.905 ;
        RECT 90.965 205.720 94.965 205.860 ;
        RECT 90.965 205.675 91.255 205.720 ;
        RECT 92.155 205.675 92.445 205.720 ;
        RECT 94.675 205.675 94.965 205.720 ;
        RECT 98.325 205.860 98.615 205.905 ;
        RECT 99.515 205.860 99.805 205.905 ;
        RECT 102.035 205.860 102.325 205.905 ;
        RECT 98.325 205.720 102.325 205.860 ;
        RECT 98.325 205.675 98.615 205.720 ;
        RECT 99.515 205.675 99.805 205.720 ;
        RECT 102.035 205.675 102.325 205.720 ;
        RECT 52.365 205.520 52.655 205.565 ;
        RECT 54.650 205.520 54.970 205.580 ;
        RECT 52.365 205.380 54.970 205.520 ;
        RECT 52.365 205.335 52.655 205.380 ;
        RECT 54.650 205.320 54.970 205.380 ;
        RECT 55.570 205.520 55.890 205.580 ;
        RECT 62.070 205.520 62.360 205.565 ;
        RECT 55.570 205.380 62.360 205.520 ;
        RECT 55.570 205.320 55.890 205.380 ;
        RECT 62.070 205.335 62.360 205.380 ;
        RECT 63.405 205.520 63.695 205.565 ;
        RECT 65.690 205.520 66.010 205.580 ;
        RECT 71.225 205.520 71.515 205.565 ;
        RECT 89.625 205.520 89.915 205.565 ;
        RECT 90.085 205.520 90.375 205.565 ;
        RECT 63.405 205.380 71.515 205.520 ;
        RECT 63.405 205.335 63.695 205.380 ;
        RECT 65.690 205.320 66.010 205.380 ;
        RECT 71.225 205.335 71.515 205.380 ;
        RECT 80.500 205.380 90.375 205.520 ;
        RECT 69.370 205.180 69.690 205.240 ;
        RECT 69.890 205.180 70.180 205.225 ;
        RECT 69.370 205.040 70.180 205.180 ;
        RECT 69.370 204.980 69.690 205.040 ;
        RECT 69.890 204.995 70.180 205.040 ;
        RECT 80.500 204.900 80.640 205.380 ;
        RECT 89.625 205.335 89.915 205.380 ;
        RECT 90.085 205.335 90.375 205.380 ;
        RECT 96.510 205.520 96.830 205.580 ;
        RECT 97.445 205.520 97.735 205.565 ;
        RECT 96.510 205.380 97.735 205.520 ;
        RECT 96.510 205.320 96.830 205.380 ;
        RECT 97.445 205.335 97.735 205.380 ;
        RECT 85.470 205.180 85.790 205.240 ;
        RECT 88.290 205.180 88.580 205.225 ;
        RECT 85.470 205.040 88.580 205.180 ;
        RECT 85.470 204.980 85.790 205.040 ;
        RECT 88.290 204.995 88.580 205.040 ;
        RECT 91.420 205.180 91.710 205.225 ;
        RECT 91.910 205.180 92.230 205.240 ;
        RECT 91.420 205.040 92.230 205.180 ;
        RECT 91.420 204.995 91.710 205.040 ;
        RECT 91.910 204.980 92.230 205.040 ;
        RECT 98.780 205.180 99.070 205.225 ;
        RECT 100.650 205.180 100.970 205.240 ;
        RECT 98.780 205.040 100.970 205.180 ;
        RECT 98.780 204.995 99.070 205.040 ;
        RECT 100.650 204.980 100.970 205.040 ;
        RECT 103.410 205.180 103.730 205.240 ;
        RECT 104.805 205.180 105.095 205.225 ;
        RECT 103.410 205.040 105.095 205.180 ;
        RECT 103.410 204.980 103.730 205.040 ;
        RECT 104.805 204.995 105.095 205.040 ;
        RECT 106.645 205.180 106.935 205.225 ;
        RECT 107.090 205.180 107.410 205.240 ;
        RECT 106.645 205.040 107.410 205.180 ;
        RECT 106.645 204.995 106.935 205.040 ;
        RECT 107.090 204.980 107.410 205.040 ;
        RECT 49.130 204.640 49.450 204.900 ;
        RECT 64.310 204.640 64.630 204.900 ;
        RECT 80.410 204.640 80.730 204.900 ;
        RECT 82.710 204.640 83.030 204.900 ;
        RECT 96.970 204.640 97.290 204.900 ;
        RECT 17.320 204.020 147.040 204.500 ;
        RECT 49.130 203.820 49.450 203.880 ;
        RECT 45.080 203.680 49.450 203.820 ;
        RECT 45.080 203.185 45.220 203.680 ;
        RECT 49.130 203.620 49.450 203.680 ;
        RECT 68.450 203.620 68.770 203.880 ;
        RECT 79.965 203.820 80.255 203.865 ;
        RECT 85.930 203.820 86.250 203.880 ;
        RECT 79.965 203.680 86.250 203.820 ;
        RECT 79.965 203.635 80.255 203.680 ;
        RECT 85.930 203.620 86.250 203.680 ;
        RECT 87.310 203.820 87.630 203.880 ;
        RECT 87.310 203.680 90.760 203.820 ;
        RECT 87.310 203.620 87.630 203.680 ;
        RECT 45.450 203.480 45.770 203.540 ;
        RECT 86.390 203.480 86.710 203.540 ;
        RECT 90.085 203.480 90.375 203.525 ;
        RECT 45.450 203.340 53.960 203.480 ;
        RECT 45.450 203.280 45.770 203.340 ;
        RECT 46.460 203.185 46.600 203.340 ;
        RECT 45.005 202.955 45.295 203.185 ;
        RECT 45.925 202.955 46.215 203.185 ;
        RECT 46.385 202.955 46.675 203.185 ;
        RECT 47.720 203.140 48.010 203.185 ;
        RECT 50.510 203.140 50.830 203.200 ;
        RECT 53.820 203.185 53.960 203.340 ;
        RECT 72.220 203.340 80.640 203.480 ;
        RECT 47.720 203.000 50.830 203.140 ;
        RECT 47.720 202.955 48.010 203.000 ;
        RECT 46.000 202.460 46.140 202.955 ;
        RECT 50.510 202.940 50.830 203.000 ;
        RECT 53.745 202.955 54.035 203.185 ;
        RECT 54.190 203.140 54.510 203.200 ;
        RECT 55.025 203.140 55.315 203.185 ;
        RECT 54.190 203.000 55.315 203.140 ;
        RECT 54.190 202.940 54.510 203.000 ;
        RECT 55.025 202.955 55.315 203.000 ;
        RECT 65.245 203.140 65.535 203.185 ;
        RECT 66.150 203.140 66.470 203.200 ;
        RECT 65.245 203.000 66.470 203.140 ;
        RECT 65.245 202.955 65.535 203.000 ;
        RECT 66.150 202.940 66.470 203.000 ;
        RECT 69.370 202.940 69.690 203.200 ;
        RECT 70.305 203.140 70.595 203.185 ;
        RECT 71.210 203.140 71.530 203.200 ;
        RECT 70.305 203.000 71.530 203.140 ;
        RECT 70.305 202.955 70.595 203.000 ;
        RECT 71.210 202.940 71.530 203.000 ;
        RECT 71.670 202.940 71.990 203.200 ;
        RECT 47.265 202.800 47.555 202.845 ;
        RECT 48.455 202.800 48.745 202.845 ;
        RECT 50.975 202.800 51.265 202.845 ;
        RECT 47.265 202.660 51.265 202.800 ;
        RECT 47.265 202.615 47.555 202.660 ;
        RECT 48.455 202.615 48.745 202.660 ;
        RECT 50.975 202.615 51.265 202.660 ;
        RECT 54.625 202.800 54.915 202.845 ;
        RECT 55.815 202.800 56.105 202.845 ;
        RECT 58.335 202.800 58.625 202.845 ;
        RECT 63.865 202.800 64.155 202.845 ;
        RECT 54.625 202.660 58.625 202.800 ;
        RECT 54.625 202.615 54.915 202.660 ;
        RECT 55.815 202.615 56.105 202.660 ;
        RECT 58.335 202.615 58.625 202.660 ;
        RECT 60.720 202.660 64.155 202.800 ;
        RECT 46.870 202.460 47.160 202.505 ;
        RECT 48.970 202.460 49.260 202.505 ;
        RECT 50.540 202.460 50.830 202.505 ;
        RECT 54.230 202.460 54.520 202.505 ;
        RECT 56.330 202.460 56.620 202.505 ;
        RECT 57.900 202.460 58.190 202.505 ;
        RECT 46.000 202.320 46.600 202.460 ;
        RECT 45.910 201.920 46.230 202.180 ;
        RECT 46.460 202.120 46.600 202.320 ;
        RECT 46.870 202.320 50.830 202.460 ;
        RECT 46.870 202.275 47.160 202.320 ;
        RECT 48.970 202.275 49.260 202.320 ;
        RECT 50.540 202.275 50.830 202.320 ;
        RECT 52.900 202.320 53.960 202.460 ;
        RECT 52.900 202.120 53.040 202.320 ;
        RECT 46.460 201.980 53.040 202.120 ;
        RECT 53.270 201.920 53.590 202.180 ;
        RECT 53.820 202.120 53.960 202.320 ;
        RECT 54.230 202.320 58.190 202.460 ;
        RECT 54.230 202.275 54.520 202.320 ;
        RECT 56.330 202.275 56.620 202.320 ;
        RECT 57.900 202.275 58.190 202.320 ;
        RECT 59.710 202.460 60.030 202.520 ;
        RECT 60.720 202.505 60.860 202.660 ;
        RECT 63.865 202.615 64.155 202.660 ;
        RECT 65.690 202.800 66.010 202.860 ;
        RECT 72.220 202.800 72.360 203.340 ;
        RECT 80.500 203.200 80.640 203.340 ;
        RECT 86.390 203.340 90.375 203.480 ;
        RECT 90.620 203.480 90.760 203.680 ;
        RECT 91.910 203.620 92.230 203.880 ;
        RECT 96.985 203.820 97.275 203.865 ;
        RECT 107.090 203.820 107.410 203.880 ;
        RECT 96.985 203.680 107.410 203.820 ;
        RECT 96.985 203.635 97.275 203.680 ;
        RECT 107.090 203.620 107.410 203.680 ;
        RECT 96.510 203.480 96.830 203.540 ;
        RECT 90.620 203.340 92.600 203.480 ;
        RECT 86.390 203.280 86.710 203.340 ;
        RECT 90.085 203.295 90.375 203.340 ;
        RECT 92.460 203.200 92.600 203.340 ;
        RECT 96.510 203.340 108.240 203.480 ;
        RECT 96.510 203.280 96.830 203.340 ;
        RECT 72.605 203.170 72.895 203.185 ;
        RECT 72.605 203.140 73.740 203.170 ;
        RECT 74.345 203.140 74.635 203.185 ;
        RECT 72.605 203.030 74.635 203.140 ;
        RECT 72.605 202.955 72.895 203.030 ;
        RECT 73.600 203.000 74.635 203.030 ;
        RECT 74.345 202.955 74.635 203.000 ;
        RECT 80.410 202.940 80.730 203.200 ;
        RECT 81.790 203.185 82.110 203.200 ;
        RECT 89.610 203.185 89.930 203.200 ;
        RECT 81.760 202.955 82.110 203.185 ;
        RECT 88.705 202.955 88.995 203.185 ;
        RECT 89.445 202.955 89.930 203.185 ;
        RECT 81.790 202.940 82.110 202.955 ;
        RECT 73.065 202.800 73.355 202.845 ;
        RECT 65.690 202.660 73.355 202.800 ;
        RECT 65.690 202.600 66.010 202.660 ;
        RECT 73.065 202.615 73.355 202.660 ;
        RECT 73.945 202.800 74.235 202.845 ;
        RECT 75.135 202.800 75.425 202.845 ;
        RECT 77.655 202.800 77.945 202.845 ;
        RECT 73.945 202.660 77.945 202.800 ;
        RECT 73.945 202.615 74.235 202.660 ;
        RECT 75.135 202.615 75.425 202.660 ;
        RECT 77.655 202.615 77.945 202.660 ;
        RECT 81.305 202.800 81.595 202.845 ;
        RECT 82.495 202.800 82.785 202.845 ;
        RECT 85.015 202.800 85.305 202.845 ;
        RECT 81.305 202.660 85.305 202.800 ;
        RECT 88.780 202.800 88.920 202.955 ;
        RECT 89.610 202.940 89.930 202.955 ;
        RECT 90.530 202.940 90.850 203.200 ;
        RECT 90.990 203.185 91.310 203.200 ;
        RECT 90.990 203.140 91.320 203.185 ;
        RECT 92.370 203.140 92.690 203.200 ;
        RECT 93.305 203.140 93.595 203.185 ;
        RECT 90.990 203.000 91.505 203.140 ;
        RECT 92.370 203.000 93.595 203.140 ;
        RECT 90.990 202.955 91.320 203.000 ;
        RECT 90.990 202.940 91.310 202.955 ;
        RECT 92.370 202.940 92.690 203.000 ;
        RECT 93.305 202.955 93.595 203.000 ;
        RECT 95.145 203.140 95.435 203.185 ;
        RECT 97.430 203.140 97.750 203.200 ;
        RECT 95.145 203.000 97.750 203.140 ;
        RECT 95.145 202.955 95.435 203.000 ;
        RECT 97.430 202.940 97.750 203.000 ;
        RECT 98.810 202.940 99.130 203.200 ;
        RECT 100.665 203.140 100.955 203.185 ;
        RECT 104.330 203.140 104.650 203.200 ;
        RECT 100.665 203.000 104.650 203.140 ;
        RECT 100.665 202.955 100.955 203.000 ;
        RECT 104.330 202.940 104.650 203.000 ;
        RECT 106.630 203.185 106.950 203.200 ;
        RECT 108.100 203.185 108.240 203.340 ;
        RECT 106.630 203.140 106.980 203.185 ;
        RECT 106.630 203.000 107.145 203.140 ;
        RECT 106.630 202.955 106.980 203.000 ;
        RECT 108.025 202.955 108.315 203.185 ;
        RECT 106.630 202.940 106.950 202.955 ;
        RECT 92.845 202.800 93.135 202.845 ;
        RECT 88.780 202.660 93.135 202.800 ;
        RECT 81.305 202.615 81.595 202.660 ;
        RECT 82.495 202.615 82.785 202.660 ;
        RECT 85.015 202.615 85.305 202.660 ;
        RECT 92.845 202.615 93.135 202.660 ;
        RECT 95.590 202.800 95.910 202.860 ;
        RECT 98.365 202.800 98.655 202.845 ;
        RECT 95.590 202.660 98.655 202.800 ;
        RECT 95.590 202.600 95.910 202.660 ;
        RECT 98.365 202.615 98.655 202.660 ;
        RECT 100.205 202.800 100.495 202.845 ;
        RECT 102.950 202.800 103.270 202.860 ;
        RECT 100.205 202.660 103.270 202.800 ;
        RECT 100.205 202.615 100.495 202.660 ;
        RECT 60.645 202.460 60.935 202.505 ;
        RECT 59.710 202.320 60.935 202.460 ;
        RECT 59.710 202.260 60.030 202.320 ;
        RECT 60.645 202.275 60.935 202.320 ;
        RECT 73.550 202.460 73.840 202.505 ;
        RECT 75.650 202.460 75.940 202.505 ;
        RECT 77.220 202.460 77.510 202.505 ;
        RECT 73.550 202.320 77.510 202.460 ;
        RECT 73.550 202.275 73.840 202.320 ;
        RECT 75.650 202.275 75.940 202.320 ;
        RECT 77.220 202.275 77.510 202.320 ;
        RECT 80.910 202.460 81.200 202.505 ;
        RECT 83.010 202.460 83.300 202.505 ;
        RECT 84.580 202.460 84.870 202.505 ;
        RECT 80.910 202.320 84.870 202.460 ;
        RECT 80.910 202.275 81.200 202.320 ;
        RECT 83.010 202.275 83.300 202.320 ;
        RECT 84.580 202.275 84.870 202.320 ;
        RECT 93.290 202.460 93.610 202.520 ;
        RECT 95.680 202.460 95.820 202.600 ;
        RECT 93.290 202.320 95.820 202.460 ;
        RECT 98.440 202.460 98.580 202.615 ;
        RECT 102.950 202.600 103.270 202.660 ;
        RECT 103.435 202.800 103.725 202.845 ;
        RECT 105.955 202.800 106.245 202.845 ;
        RECT 107.145 202.800 107.435 202.845 ;
        RECT 103.435 202.660 107.435 202.800 ;
        RECT 103.435 202.615 103.725 202.660 ;
        RECT 105.955 202.615 106.245 202.660 ;
        RECT 107.145 202.615 107.435 202.660 ;
        RECT 99.730 202.460 100.050 202.520 ;
        RECT 101.125 202.460 101.415 202.505 ;
        RECT 98.440 202.320 101.415 202.460 ;
        RECT 93.290 202.260 93.610 202.320 ;
        RECT 99.730 202.260 100.050 202.320 ;
        RECT 101.125 202.275 101.415 202.320 ;
        RECT 103.870 202.460 104.160 202.505 ;
        RECT 105.440 202.460 105.730 202.505 ;
        RECT 107.540 202.460 107.830 202.505 ;
        RECT 103.870 202.320 107.830 202.460 ;
        RECT 103.870 202.275 104.160 202.320 ;
        RECT 105.440 202.275 105.730 202.320 ;
        RECT 107.540 202.275 107.830 202.320 ;
        RECT 55.110 202.120 55.430 202.180 ;
        RECT 53.820 201.980 55.430 202.120 ;
        RECT 55.110 201.920 55.430 201.980 ;
        RECT 61.090 201.920 61.410 202.180 ;
        RECT 87.325 202.120 87.615 202.165 ;
        RECT 89.150 202.120 89.470 202.180 ;
        RECT 87.325 201.980 89.470 202.120 ;
        RECT 87.325 201.935 87.615 201.980 ;
        RECT 89.150 201.920 89.470 201.980 ;
        RECT 90.530 202.120 90.850 202.180 ;
        RECT 95.145 202.120 95.435 202.165 ;
        RECT 96.970 202.120 97.290 202.180 ;
        RECT 90.530 201.980 97.290 202.120 ;
        RECT 90.530 201.920 90.850 201.980 ;
        RECT 95.145 201.935 95.435 201.980 ;
        RECT 96.970 201.920 97.290 201.980 ;
        RECT 97.445 202.120 97.735 202.165 ;
        RECT 98.350 202.120 98.670 202.180 ;
        RECT 97.445 201.980 98.670 202.120 ;
        RECT 97.445 201.935 97.735 201.980 ;
        RECT 98.350 201.920 98.670 201.980 ;
        RECT 17.320 201.300 147.040 201.780 ;
        RECT 53.730 201.100 54.050 201.160 ;
        RECT 55.585 201.100 55.875 201.145 ;
        RECT 53.730 200.960 55.875 201.100 ;
        RECT 53.730 200.900 54.050 200.960 ;
        RECT 55.585 200.915 55.875 200.960 ;
        RECT 60.185 201.100 60.475 201.145 ;
        RECT 60.630 201.100 60.950 201.160 ;
        RECT 60.185 200.960 60.950 201.100 ;
        RECT 60.185 200.915 60.475 200.960 ;
        RECT 60.630 200.900 60.950 200.960 ;
        RECT 61.105 200.915 61.395 201.145 ;
        RECT 64.785 201.100 65.075 201.145 ;
        RECT 68.910 201.100 69.230 201.160 ;
        RECT 64.785 200.960 69.230 201.100 ;
        RECT 64.785 200.915 65.075 200.960 ;
        RECT 46.410 200.760 46.700 200.805 ;
        RECT 48.510 200.760 48.800 200.805 ;
        RECT 50.080 200.760 50.370 200.805 ;
        RECT 46.410 200.620 50.370 200.760 ;
        RECT 46.410 200.575 46.700 200.620 ;
        RECT 48.510 200.575 48.800 200.620 ;
        RECT 50.080 200.575 50.370 200.620 ;
        RECT 59.710 200.760 60.030 200.820 ;
        RECT 61.180 200.760 61.320 200.915 ;
        RECT 68.910 200.900 69.230 200.960 ;
        RECT 69.370 201.100 69.690 201.160 ;
        RECT 73.065 201.100 73.355 201.145 ;
        RECT 69.370 200.960 73.355 201.100 ;
        RECT 69.370 200.900 69.690 200.960 ;
        RECT 73.065 200.915 73.355 200.960 ;
        RECT 81.790 201.100 82.110 201.160 ;
        RECT 82.725 201.100 83.015 201.145 ;
        RECT 81.790 200.960 83.015 201.100 ;
        RECT 81.790 200.900 82.110 200.960 ;
        RECT 82.725 200.915 83.015 200.960 ;
        RECT 86.390 200.900 86.710 201.160 ;
        RECT 90.990 200.900 91.310 201.160 ;
        RECT 100.650 200.900 100.970 201.160 ;
        RECT 59.710 200.620 61.320 200.760 ;
        RECT 66.190 200.760 66.480 200.805 ;
        RECT 68.290 200.760 68.580 200.805 ;
        RECT 69.860 200.760 70.150 200.805 ;
        RECT 66.190 200.620 70.150 200.760 ;
        RECT 59.710 200.560 60.030 200.620 ;
        RECT 66.190 200.575 66.480 200.620 ;
        RECT 68.290 200.575 68.580 200.620 ;
        RECT 69.860 200.575 70.150 200.620 ;
        RECT 70.750 200.760 71.070 200.820 ;
        RECT 74.905 200.760 75.195 200.805 ;
        RECT 70.750 200.620 75.195 200.760 ;
        RECT 70.750 200.560 71.070 200.620 ;
        RECT 74.905 200.575 75.195 200.620 ;
        RECT 90.085 200.575 90.375 200.805 ;
        RECT 92.370 200.760 92.690 200.820 ;
        RECT 92.370 200.620 97.660 200.760 ;
        RECT 43.610 200.420 43.930 200.480 ;
        RECT 45.450 200.420 45.770 200.480 ;
        RECT 45.925 200.420 46.215 200.465 ;
        RECT 43.610 200.280 46.215 200.420 ;
        RECT 43.610 200.220 43.930 200.280 ;
        RECT 45.450 200.220 45.770 200.280 ;
        RECT 45.925 200.235 46.215 200.280 ;
        RECT 46.805 200.420 47.095 200.465 ;
        RECT 47.995 200.420 48.285 200.465 ;
        RECT 50.515 200.420 50.805 200.465 ;
        RECT 46.805 200.280 50.805 200.420 ;
        RECT 46.805 200.235 47.095 200.280 ;
        RECT 47.995 200.235 48.285 200.280 ;
        RECT 50.515 200.235 50.805 200.280 ;
        RECT 59.265 200.420 59.555 200.465 ;
        RECT 60.170 200.420 60.490 200.480 ;
        RECT 62.930 200.420 63.250 200.480 ;
        RECT 59.265 200.280 63.250 200.420 ;
        RECT 59.265 200.235 59.555 200.280 ;
        RECT 60.170 200.220 60.490 200.280 ;
        RECT 62.930 200.220 63.250 200.280 ;
        RECT 65.690 200.220 66.010 200.480 ;
        RECT 66.585 200.420 66.875 200.465 ;
        RECT 67.775 200.420 68.065 200.465 ;
        RECT 70.295 200.420 70.585 200.465 ;
        RECT 66.585 200.280 70.585 200.420 ;
        RECT 66.585 200.235 66.875 200.280 ;
        RECT 67.775 200.235 68.065 200.280 ;
        RECT 70.295 200.235 70.585 200.280 ;
        RECT 83.645 200.420 83.935 200.465 ;
        RECT 90.160 200.420 90.300 200.575 ;
        RECT 92.370 200.560 92.690 200.620 ;
        RECT 83.645 200.280 93.520 200.420 ;
        RECT 83.645 200.235 83.935 200.280 ;
        RECT 53.270 200.080 53.590 200.140 ;
        RECT 54.190 200.080 54.510 200.140 ;
        RECT 53.270 199.940 54.510 200.080 ;
        RECT 53.270 199.880 53.590 199.940 ;
        RECT 54.190 199.880 54.510 199.940 ;
        RECT 55.585 200.080 55.875 200.125 ;
        RECT 61.090 200.080 61.410 200.140 ;
        RECT 55.585 199.940 61.410 200.080 ;
        RECT 55.585 199.895 55.875 199.940 ;
        RECT 61.090 199.880 61.410 199.940 ;
        RECT 61.550 200.080 61.870 200.140 ;
        RECT 63.405 200.080 63.695 200.125 ;
        RECT 64.310 200.080 64.630 200.140 ;
        RECT 61.550 199.940 64.630 200.080 ;
        RECT 61.550 199.880 61.870 199.940 ;
        RECT 63.405 199.895 63.695 199.940 ;
        RECT 64.310 199.880 64.630 199.940 ;
        RECT 71.670 200.080 71.990 200.140 ;
        RECT 73.065 200.080 73.355 200.125 ;
        RECT 71.670 199.940 73.355 200.080 ;
        RECT 71.670 199.880 71.990 199.940 ;
        RECT 73.065 199.895 73.355 199.940 ;
        RECT 73.985 200.080 74.275 200.125 ;
        RECT 82.710 200.080 83.030 200.140 ;
        RECT 73.985 199.940 83.030 200.080 ;
        RECT 73.985 199.895 74.275 199.940 ;
        RECT 82.710 199.880 83.030 199.940 ;
        RECT 84.105 200.080 84.395 200.125 ;
        RECT 86.390 200.080 86.710 200.140 ;
        RECT 84.105 199.940 86.710 200.080 ;
        RECT 84.105 199.895 84.395 199.940 ;
        RECT 86.390 199.880 86.710 199.940 ;
        RECT 89.150 199.880 89.470 200.140 ;
        RECT 90.530 200.080 90.850 200.140 ;
        RECT 91.005 200.080 91.295 200.125 ;
        RECT 90.530 199.940 91.295 200.080 ;
        RECT 90.530 199.880 90.850 199.940 ;
        RECT 91.005 199.895 91.295 199.940 ;
        RECT 92.830 199.880 93.150 200.140 ;
        RECT 93.380 200.125 93.520 200.280 ;
        RECT 97.520 200.125 97.660 200.620 ;
        RECT 98.810 200.560 99.130 200.820 ;
        RECT 99.285 200.420 99.575 200.465 ;
        RECT 108.010 200.420 108.330 200.480 ;
        RECT 99.285 200.280 108.330 200.420 ;
        RECT 99.285 200.235 99.575 200.280 ;
        RECT 108.010 200.220 108.330 200.280 ;
        RECT 93.305 199.895 93.595 200.125 ;
        RECT 97.445 199.895 97.735 200.125 ;
        RECT 45.910 199.740 46.230 199.800 ;
        RECT 47.150 199.740 47.440 199.785 ;
        RECT 54.650 199.740 54.970 199.800 ;
        RECT 56.490 199.740 56.810 199.800 ;
        RECT 45.910 199.600 47.440 199.740 ;
        RECT 45.910 199.540 46.230 199.600 ;
        RECT 47.150 199.555 47.440 199.600 ;
        RECT 52.900 199.600 56.810 199.740 ;
        RECT 52.900 199.445 53.040 199.600 ;
        RECT 54.650 199.540 54.970 199.600 ;
        RECT 56.490 199.540 56.810 199.600 ;
        RECT 56.950 199.740 57.270 199.800 ;
        RECT 57.425 199.740 57.715 199.785 ;
        RECT 56.950 199.600 57.715 199.740 ;
        RECT 56.950 199.540 57.270 199.600 ;
        RECT 57.425 199.555 57.715 199.600 ;
        RECT 57.885 199.740 58.175 199.785 ;
        RECT 59.250 199.740 59.570 199.800 ;
        RECT 57.885 199.600 59.570 199.740 ;
        RECT 57.885 199.555 58.175 199.600 ;
        RECT 59.250 199.540 59.570 199.600 ;
        RECT 59.710 199.740 60.030 199.800 ;
        RECT 67.070 199.785 67.390 199.800 ;
        RECT 62.025 199.740 62.315 199.785 ;
        RECT 59.710 199.600 62.315 199.740 ;
        RECT 59.710 199.540 60.030 199.600 ;
        RECT 62.025 199.555 62.315 199.600 ;
        RECT 67.040 199.555 67.390 199.785 ;
        RECT 89.240 199.740 89.380 199.880 ;
        RECT 94.225 199.740 94.515 199.785 ;
        RECT 89.240 199.600 94.515 199.740 ;
        RECT 97.520 199.740 97.660 199.895 ;
        RECT 98.350 199.880 98.670 200.140 ;
        RECT 99.730 199.880 100.050 200.140 ;
        RECT 103.410 199.740 103.730 199.800 ;
        RECT 97.520 199.600 103.730 199.740 ;
        RECT 94.225 199.555 94.515 199.600 ;
        RECT 67.070 199.540 67.390 199.555 ;
        RECT 103.410 199.540 103.730 199.600 ;
        RECT 52.825 199.215 53.115 199.445 ;
        RECT 58.330 199.400 58.650 199.460 ;
        RECT 60.975 199.400 61.265 199.445 ;
        RECT 58.330 199.260 61.265 199.400 ;
        RECT 58.330 199.200 58.650 199.260 ;
        RECT 60.975 199.215 61.265 199.260 ;
        RECT 66.150 199.400 66.470 199.460 ;
        RECT 68.450 199.400 68.770 199.460 ;
        RECT 72.605 199.400 72.895 199.445 ;
        RECT 66.150 199.260 72.895 199.400 ;
        RECT 66.150 199.200 66.470 199.260 ;
        RECT 68.450 199.200 68.770 199.260 ;
        RECT 72.605 199.215 72.895 199.260 ;
        RECT 85.930 199.200 86.250 199.460 ;
        RECT 95.145 199.400 95.435 199.445 ;
        RECT 95.590 199.400 95.910 199.460 ;
        RECT 95.145 199.260 95.910 199.400 ;
        RECT 95.145 199.215 95.435 199.260 ;
        RECT 95.590 199.200 95.910 199.260 ;
        RECT 17.320 198.580 147.040 199.060 ;
        RECT 50.510 198.380 50.830 198.440 ;
        RECT 50.985 198.380 51.275 198.425 ;
        RECT 50.510 198.240 51.275 198.380 ;
        RECT 50.510 198.180 50.830 198.240 ;
        RECT 50.985 198.195 51.275 198.240 ;
        RECT 62.930 198.380 63.250 198.440 ;
        RECT 67.415 198.380 67.705 198.425 ;
        RECT 62.930 198.240 67.705 198.380 ;
        RECT 62.930 198.180 63.250 198.240 ;
        RECT 67.415 198.195 67.705 198.240 ;
        RECT 64.860 197.900 65.920 198.040 ;
        RECT 50.525 197.700 50.815 197.745 ;
        RECT 50.970 197.700 51.290 197.760 ;
        RECT 50.525 197.560 51.290 197.700 ;
        RECT 50.525 197.515 50.815 197.560 ;
        RECT 50.970 197.500 51.290 197.560 ;
        RECT 51.445 197.700 51.735 197.745 ;
        RECT 52.350 197.700 52.670 197.760 ;
        RECT 51.445 197.560 52.670 197.700 ;
        RECT 51.445 197.515 51.735 197.560 ;
        RECT 52.350 197.500 52.670 197.560 ;
        RECT 56.045 197.700 56.335 197.745 ;
        RECT 56.490 197.700 56.810 197.760 ;
        RECT 59.710 197.700 60.030 197.760 ;
        RECT 64.860 197.700 65.000 197.900 ;
        RECT 56.045 197.560 60.030 197.700 ;
        RECT 56.045 197.515 56.335 197.560 ;
        RECT 56.490 197.500 56.810 197.560 ;
        RECT 59.710 197.500 60.030 197.560 ;
        RECT 63.940 197.560 65.000 197.700 ;
        RECT 52.440 197.360 52.580 197.500 ;
        RECT 63.940 197.405 64.080 197.560 ;
        RECT 65.230 197.500 65.550 197.760 ;
        RECT 65.780 197.700 65.920 197.900 ;
        RECT 68.450 197.840 68.770 198.100 ;
        RECT 89.610 198.040 89.930 198.100 ;
        RECT 86.480 197.900 89.930 198.040 ;
        RECT 65.780 197.560 69.600 197.700 ;
        RECT 63.865 197.360 64.155 197.405 ;
        RECT 68.910 197.360 69.230 197.420 ;
        RECT 52.440 197.220 64.155 197.360 ;
        RECT 63.865 197.175 64.155 197.220 ;
        RECT 64.860 197.220 69.230 197.360 ;
        RECT 50.510 197.020 50.830 197.080 ;
        RECT 59.250 197.020 59.570 197.080 ;
        RECT 64.860 197.065 65.000 197.220 ;
        RECT 68.910 197.160 69.230 197.220 ;
        RECT 50.510 196.880 59.570 197.020 ;
        RECT 50.510 196.820 50.830 196.880 ;
        RECT 59.250 196.820 59.570 196.880 ;
        RECT 64.785 196.835 65.075 197.065 ;
        RECT 65.245 197.020 65.535 197.065 ;
        RECT 67.070 197.020 67.390 197.080 ;
        RECT 65.245 196.880 67.390 197.020 ;
        RECT 69.460 197.020 69.600 197.560 ;
        RECT 70.750 197.500 71.070 197.760 ;
        RECT 86.480 197.745 86.620 197.900 ;
        RECT 89.610 197.840 89.930 197.900 ;
        RECT 86.405 197.515 86.695 197.745 ;
        RECT 87.785 197.700 88.075 197.745 ;
        RECT 89.150 197.700 89.470 197.760 ;
        RECT 87.785 197.560 89.470 197.700 ;
        RECT 87.785 197.515 88.075 197.560 ;
        RECT 89.150 197.500 89.470 197.560 ;
        RECT 94.210 197.700 94.530 197.760 ;
        RECT 95.145 197.700 95.435 197.745 ;
        RECT 94.210 197.560 95.435 197.700 ;
        RECT 94.210 197.500 94.530 197.560 ;
        RECT 95.145 197.515 95.435 197.560 ;
        RECT 96.050 197.500 96.370 197.760 ;
        RECT 108.010 197.700 108.330 197.760 ;
        RECT 114.005 197.700 114.295 197.745 ;
        RECT 108.010 197.560 114.295 197.700 ;
        RECT 108.010 197.500 108.330 197.560 ;
        RECT 114.005 197.515 114.295 197.560 ;
        RECT 108.470 197.360 108.790 197.420 ;
        RECT 110.785 197.360 111.075 197.405 ;
        RECT 108.470 197.220 111.075 197.360 ;
        RECT 108.470 197.160 108.790 197.220 ;
        RECT 110.785 197.175 111.075 197.220 ;
        RECT 69.845 197.020 70.135 197.065 ;
        RECT 72.590 197.020 72.910 197.080 ;
        RECT 69.460 196.880 72.910 197.020 ;
        RECT 65.245 196.835 65.535 196.880 ;
        RECT 51.430 196.680 51.750 196.740 ;
        RECT 55.585 196.680 55.875 196.725 ;
        RECT 51.430 196.540 55.875 196.680 ;
        RECT 64.860 196.680 65.000 196.835 ;
        RECT 67.070 196.820 67.390 196.880 ;
        RECT 69.845 196.835 70.135 196.880 ;
        RECT 72.590 196.820 72.910 196.880 ;
        RECT 66.625 196.680 66.915 196.725 ;
        RECT 64.860 196.540 66.915 196.680 ;
        RECT 51.430 196.480 51.750 196.540 ;
        RECT 55.585 196.495 55.875 196.540 ;
        RECT 66.625 196.495 66.915 196.540 ;
        RECT 67.530 196.480 67.850 196.740 ;
        RECT 80.870 196.680 81.190 196.740 ;
        RECT 85.010 196.680 85.330 196.740 ;
        RECT 85.485 196.680 85.775 196.725 ;
        RECT 80.870 196.540 85.775 196.680 ;
        RECT 80.870 196.480 81.190 196.540 ;
        RECT 85.010 196.480 85.330 196.540 ;
        RECT 85.485 196.495 85.775 196.540 ;
        RECT 87.325 196.680 87.615 196.725 ;
        RECT 91.450 196.680 91.770 196.740 ;
        RECT 87.325 196.540 91.770 196.680 ;
        RECT 87.325 196.495 87.615 196.540 ;
        RECT 91.450 196.480 91.770 196.540 ;
        RECT 94.670 196.680 94.990 196.740 ;
        RECT 95.145 196.680 95.435 196.725 ;
        RECT 94.670 196.540 95.435 196.680 ;
        RECT 94.670 196.480 94.990 196.540 ;
        RECT 95.145 196.495 95.435 196.540 ;
        RECT 17.320 195.860 147.040 196.340 ;
        RECT 61.550 195.660 61.870 195.720 ;
        RECT 67.530 195.660 67.850 195.720 ;
        RECT 61.550 195.520 67.850 195.660 ;
        RECT 61.550 195.460 61.870 195.520 ;
        RECT 67.530 195.460 67.850 195.520 ;
        RECT 81.330 195.660 81.650 195.720 ;
        RECT 85.930 195.660 86.250 195.720 ;
        RECT 93.305 195.660 93.595 195.705 ;
        RECT 81.330 195.520 93.595 195.660 ;
        RECT 81.330 195.460 81.650 195.520 ;
        RECT 85.930 195.460 86.250 195.520 ;
        RECT 93.305 195.475 93.595 195.520 ;
        RECT 95.590 195.460 95.910 195.720 ;
        RECT 96.050 195.660 96.370 195.720 ;
        RECT 97.890 195.660 98.210 195.720 ;
        RECT 103.425 195.660 103.715 195.705 ;
        RECT 96.050 195.520 103.715 195.660 ;
        RECT 96.050 195.460 96.370 195.520 ;
        RECT 97.890 195.460 98.210 195.520 ;
        RECT 103.425 195.475 103.715 195.520 ;
        RECT 42.690 195.320 43.010 195.380 ;
        RECT 59.265 195.320 59.555 195.365 ;
        RECT 60.630 195.320 60.950 195.380 ;
        RECT 42.690 195.180 58.560 195.320 ;
        RECT 42.690 195.120 43.010 195.180 ;
        RECT 52.810 194.980 53.130 195.040 ;
        RECT 56.965 194.980 57.255 195.025 ;
        RECT 52.810 194.840 57.255 194.980 ;
        RECT 52.810 194.780 53.130 194.840 ;
        RECT 56.965 194.795 57.255 194.840 ;
        RECT 21.530 194.640 21.850 194.700 ;
        RECT 26.130 194.640 26.450 194.700 ;
        RECT 21.530 194.500 26.450 194.640 ;
        RECT 21.530 194.440 21.850 194.500 ;
        RECT 26.130 194.440 26.450 194.500 ;
        RECT 26.605 194.640 26.895 194.685 ;
        RECT 32.110 194.640 32.430 194.700 ;
        RECT 26.605 194.500 32.430 194.640 ;
        RECT 26.605 194.455 26.895 194.500 ;
        RECT 32.110 194.440 32.430 194.500 ;
        RECT 54.190 194.640 54.510 194.700 ;
        RECT 56.505 194.640 56.795 194.685 ;
        RECT 54.190 194.500 56.795 194.640 ;
        RECT 54.190 194.440 54.510 194.500 ;
        RECT 56.505 194.455 56.795 194.500 ;
        RECT 27.525 194.300 27.815 194.345 ;
        RECT 28.890 194.300 29.210 194.360 ;
        RECT 27.525 194.160 29.210 194.300 ;
        RECT 27.525 194.115 27.815 194.160 ;
        RECT 28.890 194.100 29.210 194.160 ;
        RECT 39.470 194.100 39.790 194.360 ;
        RECT 53.730 194.100 54.050 194.360 ;
        RECT 54.665 194.300 54.955 194.345 ;
        RECT 56.030 194.300 56.350 194.360 ;
        RECT 54.665 194.160 56.350 194.300 ;
        RECT 54.665 194.115 54.955 194.160 ;
        RECT 56.030 194.100 56.350 194.160 ;
        RECT 27.050 193.760 27.370 194.020 ;
        RECT 39.930 193.760 40.250 194.020 ;
        RECT 55.110 193.960 55.430 194.020 ;
        RECT 55.585 193.960 55.875 194.005 ;
        RECT 55.110 193.820 55.875 193.960 ;
        RECT 56.580 193.960 56.720 194.455 ;
        RECT 57.040 194.300 57.180 194.795 ;
        RECT 57.885 194.640 58.175 194.685 ;
        RECT 58.420 194.640 58.560 195.180 ;
        RECT 59.265 195.180 60.950 195.320 ;
        RECT 59.265 195.135 59.555 195.180 ;
        RECT 60.630 195.120 60.950 195.180 ;
        RECT 80.410 195.320 80.730 195.380 ;
        RECT 82.750 195.320 83.040 195.365 ;
        RECT 84.850 195.320 85.140 195.365 ;
        RECT 86.420 195.320 86.710 195.365 ;
        RECT 80.410 195.180 82.480 195.320 ;
        RECT 80.410 195.120 80.730 195.180 ;
        RECT 58.790 194.780 59.110 195.040 ;
        RECT 81.330 194.780 81.650 195.040 ;
        RECT 82.340 195.025 82.480 195.180 ;
        RECT 82.750 195.180 86.710 195.320 ;
        RECT 82.750 195.135 83.040 195.180 ;
        RECT 84.850 195.135 85.140 195.180 ;
        RECT 86.420 195.135 86.710 195.180 ;
        RECT 89.165 195.320 89.455 195.365 ;
        RECT 97.010 195.320 97.300 195.365 ;
        RECT 99.110 195.320 99.400 195.365 ;
        RECT 100.680 195.320 100.970 195.365 ;
        RECT 89.165 195.180 92.600 195.320 ;
        RECT 89.165 195.135 89.455 195.180 ;
        RECT 92.460 195.025 92.600 195.180 ;
        RECT 97.010 195.180 100.970 195.320 ;
        RECT 97.010 195.135 97.300 195.180 ;
        RECT 99.110 195.135 99.400 195.180 ;
        RECT 100.680 195.135 100.970 195.180 ;
        RECT 82.265 194.795 82.555 195.025 ;
        RECT 83.145 194.980 83.435 195.025 ;
        RECT 84.335 194.980 84.625 195.025 ;
        RECT 86.855 194.980 87.145 195.025 ;
        RECT 83.145 194.840 87.145 194.980 ;
        RECT 83.145 194.795 83.435 194.840 ;
        RECT 84.335 194.795 84.625 194.840 ;
        RECT 86.855 194.795 87.145 194.840 ;
        RECT 92.385 194.980 92.675 195.025 ;
        RECT 94.685 194.980 94.975 195.025 ;
        RECT 92.385 194.840 94.975 194.980 ;
        RECT 92.385 194.795 92.675 194.840 ;
        RECT 94.685 194.795 94.975 194.840 ;
        RECT 96.510 194.780 96.830 195.040 ;
        RECT 97.405 194.980 97.695 195.025 ;
        RECT 98.595 194.980 98.885 195.025 ;
        RECT 101.115 194.980 101.405 195.025 ;
        RECT 97.405 194.840 101.405 194.980 ;
        RECT 103.500 194.980 103.640 195.475 ;
        RECT 111.230 195.320 111.520 195.365 ;
        RECT 112.800 195.320 113.090 195.365 ;
        RECT 114.900 195.320 115.190 195.365 ;
        RECT 111.230 195.180 115.190 195.320 ;
        RECT 111.230 195.135 111.520 195.180 ;
        RECT 112.800 195.135 113.090 195.180 ;
        RECT 114.900 195.135 115.190 195.180 ;
        RECT 106.645 194.980 106.935 195.025 ;
        RECT 103.500 194.840 106.935 194.980 ;
        RECT 97.405 194.795 97.695 194.840 ;
        RECT 98.595 194.795 98.885 194.840 ;
        RECT 101.115 194.795 101.405 194.840 ;
        RECT 106.645 194.795 106.935 194.840 ;
        RECT 110.795 194.980 111.085 195.025 ;
        RECT 113.315 194.980 113.605 195.025 ;
        RECT 114.505 194.980 114.795 195.025 ;
        RECT 110.795 194.840 114.795 194.980 ;
        RECT 110.795 194.795 111.085 194.840 ;
        RECT 113.315 194.795 113.605 194.840 ;
        RECT 114.505 194.795 114.795 194.840 ;
        RECT 60.645 194.640 60.935 194.685 ;
        RECT 62.470 194.640 62.790 194.700 ;
        RECT 57.885 194.500 62.790 194.640 ;
        RECT 57.885 194.455 58.175 194.500 ;
        RECT 60.645 194.455 60.935 194.500 ;
        RECT 62.470 194.440 62.790 194.500 ;
        RECT 79.950 194.440 80.270 194.700 ;
        RECT 80.425 194.640 80.715 194.685 ;
        RECT 80.870 194.640 81.190 194.700 ;
        RECT 89.625 194.640 89.915 194.685 ;
        RECT 80.425 194.500 81.190 194.640 ;
        RECT 80.425 194.455 80.715 194.500 ;
        RECT 80.870 194.440 81.190 194.500 ;
        RECT 82.800 194.500 89.915 194.640 ;
        RECT 59.265 194.300 59.555 194.345 ;
        RECT 57.040 194.160 59.555 194.300 ;
        RECT 59.265 194.115 59.555 194.160 ;
        RECT 82.250 194.300 82.570 194.360 ;
        RECT 82.800 194.300 82.940 194.500 ;
        RECT 89.625 194.455 89.915 194.500 ;
        RECT 91.450 194.640 91.770 194.700 ;
        RECT 96.065 194.640 96.355 194.685 ;
        RECT 91.450 194.500 96.355 194.640 ;
        RECT 91.450 194.440 91.770 194.500 ;
        RECT 96.065 194.455 96.355 194.500 ;
        RECT 108.010 194.640 108.330 194.700 ;
        RECT 115.385 194.640 115.675 194.685 ;
        RECT 108.010 194.500 115.675 194.640 ;
        RECT 108.010 194.440 108.330 194.500 ;
        RECT 115.385 194.455 115.675 194.500 ;
        RECT 82.250 194.160 82.940 194.300 ;
        RECT 83.600 194.300 83.890 194.345 ;
        RECT 85.930 194.300 86.250 194.360 ;
        RECT 83.600 194.160 86.250 194.300 ;
        RECT 82.250 194.100 82.570 194.160 ;
        RECT 83.600 194.115 83.890 194.160 ;
        RECT 85.930 194.100 86.250 194.160 ;
        RECT 97.860 194.300 98.150 194.345 ;
        RECT 99.270 194.300 99.590 194.360 ;
        RECT 106.170 194.300 106.490 194.360 ;
        RECT 97.860 194.160 99.590 194.300 ;
        RECT 97.860 194.115 98.150 194.160 ;
        RECT 99.270 194.100 99.590 194.160 ;
        RECT 101.660 194.160 106.490 194.300 ;
        RECT 101.660 194.020 101.800 194.160 ;
        RECT 106.170 194.100 106.490 194.160 ;
        RECT 114.160 194.300 114.450 194.345 ;
        RECT 114.910 194.300 115.230 194.360 ;
        RECT 114.160 194.160 115.230 194.300 ;
        RECT 114.160 194.115 114.450 194.160 ;
        RECT 114.910 194.100 115.230 194.160 ;
        RECT 58.330 193.960 58.650 194.020 ;
        RECT 60.185 193.960 60.475 194.005 ;
        RECT 56.580 193.820 60.475 193.960 ;
        RECT 55.110 193.760 55.430 193.820 ;
        RECT 55.585 193.775 55.875 193.820 ;
        RECT 58.330 193.760 58.650 193.820 ;
        RECT 60.185 193.775 60.475 193.820 ;
        RECT 81.345 193.960 81.635 194.005 ;
        RECT 82.710 193.960 83.030 194.020 ;
        RECT 81.345 193.820 83.030 193.960 ;
        RECT 81.345 193.775 81.635 193.820 ;
        RECT 82.710 193.760 83.030 193.820 ;
        RECT 94.210 193.960 94.530 194.020 ;
        RECT 101.570 193.960 101.890 194.020 ;
        RECT 94.210 193.820 101.890 193.960 ;
        RECT 94.210 193.760 94.530 193.820 ;
        RECT 101.570 193.760 101.890 193.820 ;
        RECT 103.870 193.760 104.190 194.020 ;
        RECT 108.470 193.760 108.790 194.020 ;
        RECT 17.320 193.140 147.040 193.620 ;
        RECT 19.705 192.940 19.995 192.985 ;
        RECT 39.470 192.940 39.790 193.000 ;
        RECT 19.705 192.800 39.790 192.940 ;
        RECT 19.705 192.755 19.995 192.800 ;
        RECT 39.470 192.740 39.790 192.800 ;
        RECT 51.430 192.740 51.750 193.000 ;
        RECT 52.810 192.940 53.130 193.000 ;
        RECT 54.665 192.940 54.955 192.985 ;
        RECT 55.110 192.940 55.430 193.000 ;
        RECT 52.810 192.800 53.500 192.940 ;
        RECT 52.810 192.740 53.130 192.800 ;
        RECT 21.530 192.400 21.850 192.660 ;
        RECT 43.610 192.600 43.930 192.660 ;
        RECT 25.300 192.460 43.930 192.600 ;
        RECT 25.300 192.320 25.440 192.460 ;
        RECT 18.770 192.060 19.090 192.320 ;
        RECT 25.210 192.060 25.530 192.320 ;
        RECT 25.670 192.260 25.990 192.320 ;
        RECT 32.660 192.305 32.800 192.460 ;
        RECT 43.610 192.400 43.930 192.460 ;
        RECT 46.370 192.600 46.690 192.660 ;
        RECT 50.985 192.600 51.275 192.645 ;
        RECT 51.890 192.600 52.210 192.660 ;
        RECT 53.360 192.645 53.500 192.800 ;
        RECT 54.665 192.800 55.430 192.940 ;
        RECT 54.665 192.755 54.955 192.800 ;
        RECT 55.110 192.740 55.430 192.800 ;
        RECT 55.585 192.940 55.875 192.985 ;
        RECT 79.950 192.940 80.270 193.000 ;
        RECT 81.805 192.940 82.095 192.985 ;
        RECT 55.585 192.800 56.260 192.940 ;
        RECT 55.585 192.755 55.875 192.800 ;
        RECT 46.370 192.460 52.210 192.600 ;
        RECT 46.370 192.400 46.690 192.460 ;
        RECT 26.505 192.260 26.795 192.305 ;
        RECT 25.670 192.120 26.795 192.260 ;
        RECT 25.670 192.060 25.990 192.120 ;
        RECT 26.505 192.075 26.795 192.120 ;
        RECT 32.585 192.075 32.875 192.305 ;
        RECT 33.920 192.260 34.210 192.305 ;
        RECT 35.790 192.260 36.110 192.320 ;
        RECT 33.920 192.120 36.110 192.260 ;
        RECT 33.920 192.075 34.210 192.120 ;
        RECT 35.790 192.060 36.110 192.120 ;
        RECT 39.945 192.075 40.235 192.305 ;
        RECT 26.105 191.920 26.395 191.965 ;
        RECT 27.295 191.920 27.585 191.965 ;
        RECT 29.815 191.920 30.105 191.965 ;
        RECT 26.105 191.780 30.105 191.920 ;
        RECT 26.105 191.735 26.395 191.780 ;
        RECT 27.295 191.735 27.585 191.780 ;
        RECT 29.815 191.735 30.105 191.780 ;
        RECT 33.465 191.920 33.755 191.965 ;
        RECT 34.655 191.920 34.945 191.965 ;
        RECT 37.175 191.920 37.465 191.965 ;
        RECT 33.465 191.780 37.465 191.920 ;
        RECT 33.465 191.735 33.755 191.780 ;
        RECT 34.655 191.735 34.945 191.780 ;
        RECT 37.175 191.735 37.465 191.780 ;
        RECT 23.385 191.580 23.675 191.625 ;
        RECT 24.750 191.580 25.070 191.640 ;
        RECT 23.385 191.440 25.070 191.580 ;
        RECT 23.385 191.395 23.675 191.440 ;
        RECT 24.750 191.380 25.070 191.440 ;
        RECT 25.710 191.580 26.000 191.625 ;
        RECT 27.810 191.580 28.100 191.625 ;
        RECT 29.380 191.580 29.670 191.625 ;
        RECT 25.710 191.440 29.670 191.580 ;
        RECT 25.710 191.395 26.000 191.440 ;
        RECT 27.810 191.395 28.100 191.440 ;
        RECT 29.380 191.395 29.670 191.440 ;
        RECT 32.110 191.380 32.430 191.640 ;
        RECT 33.070 191.580 33.360 191.625 ;
        RECT 35.170 191.580 35.460 191.625 ;
        RECT 36.740 191.580 37.030 191.625 ;
        RECT 33.070 191.440 37.030 191.580 ;
        RECT 33.070 191.395 33.360 191.440 ;
        RECT 35.170 191.395 35.460 191.440 ;
        RECT 36.740 191.395 37.030 191.440 ;
        RECT 39.485 191.580 39.775 191.625 ;
        RECT 40.020 191.580 40.160 192.075 ;
        RECT 40.850 192.060 41.170 192.320 ;
        RECT 42.705 192.260 42.995 192.305 ;
        RECT 44.990 192.260 45.310 192.320 ;
        RECT 45.480 192.305 45.740 192.350 ;
        RECT 48.760 192.305 48.900 192.460 ;
        RECT 50.985 192.415 51.275 192.460 ;
        RECT 51.890 192.400 52.210 192.460 ;
        RECT 53.285 192.415 53.575 192.645 ;
        RECT 56.120 192.600 56.260 192.800 ;
        RECT 79.950 192.800 82.095 192.940 ;
        RECT 79.950 192.740 80.270 192.800 ;
        RECT 81.805 192.755 82.095 192.800 ;
        RECT 85.930 192.740 86.250 193.000 ;
        RECT 94.210 192.740 94.530 193.000 ;
        RECT 95.590 192.940 95.910 193.000 ;
        RECT 97.445 192.940 97.735 192.985 ;
        RECT 95.590 192.800 97.735 192.940 ;
        RECT 95.590 192.740 95.910 192.800 ;
        RECT 97.445 192.755 97.735 192.800 ;
        RECT 77.205 192.600 77.495 192.645 ;
        RECT 78.570 192.600 78.890 192.660 ;
        RECT 80.410 192.600 80.730 192.660 ;
        RECT 89.610 192.600 89.930 192.660 ;
        RECT 96.970 192.600 97.290 192.660 ;
        RECT 54.740 192.460 56.260 192.600 ;
        RECT 56.580 192.460 64.540 192.600 ;
        RECT 42.705 192.120 45.310 192.260 ;
        RECT 42.705 192.075 42.995 192.120 ;
        RECT 44.990 192.060 45.310 192.120 ;
        RECT 45.465 192.260 45.755 192.305 ;
        RECT 48.225 192.260 48.515 192.305 ;
        RECT 45.465 192.120 48.515 192.260 ;
        RECT 45.465 192.075 45.755 192.120 ;
        RECT 48.225 192.075 48.515 192.120 ;
        RECT 48.685 192.075 48.975 192.305 ;
        RECT 52.825 192.260 53.115 192.305 ;
        RECT 54.190 192.260 54.510 192.320 ;
        RECT 52.825 192.120 54.510 192.260 ;
        RECT 52.825 192.075 53.115 192.120 ;
        RECT 45.480 192.030 45.740 192.075 ;
        RECT 54.190 192.060 54.510 192.120 ;
        RECT 43.150 191.920 43.470 191.980 ;
        RECT 43.625 191.920 43.915 191.965 ;
        RECT 43.150 191.780 43.915 191.920 ;
        RECT 43.150 191.720 43.470 191.780 ;
        RECT 43.625 191.735 43.915 191.780 ;
        RECT 51.890 191.920 52.210 191.980 ;
        RECT 54.740 191.920 54.880 192.460 ;
        RECT 55.125 192.260 55.415 192.305 ;
        RECT 56.580 192.260 56.720 192.460 ;
        RECT 55.125 192.120 56.720 192.260 ;
        RECT 55.125 192.075 55.415 192.120 ;
        RECT 56.965 192.075 57.255 192.305 ;
        RECT 51.890 191.780 54.880 191.920 ;
        RECT 51.890 191.720 52.210 191.780 ;
        RECT 40.390 191.580 40.710 191.640 ;
        RECT 39.485 191.440 40.710 191.580 ;
        RECT 39.485 191.395 39.775 191.440 ;
        RECT 40.390 191.380 40.710 191.440 ;
        RECT 53.745 191.580 54.035 191.625 ;
        RECT 54.650 191.580 54.970 191.640 ;
        RECT 53.745 191.440 54.970 191.580 ;
        RECT 53.745 191.395 54.035 191.440 ;
        RECT 54.650 191.380 54.970 191.440 ;
        RECT 56.505 191.580 56.795 191.625 ;
        RECT 57.040 191.580 57.180 192.075 ;
        RECT 58.790 192.060 59.110 192.320 ;
        RECT 59.250 192.060 59.570 192.320 ;
        RECT 61.550 192.060 61.870 192.320 ;
        RECT 64.400 192.305 64.540 192.460 ;
        RECT 77.205 192.460 87.540 192.600 ;
        RECT 77.205 192.415 77.495 192.460 ;
        RECT 78.570 192.400 78.890 192.460 ;
        RECT 80.410 192.400 80.730 192.460 ;
        RECT 62.485 192.260 62.775 192.305 ;
        RECT 64.325 192.260 64.615 192.305 ;
        RECT 66.610 192.260 66.930 192.320 ;
        RECT 62.485 192.120 64.080 192.260 ;
        RECT 62.485 192.075 62.775 192.120 ;
        RECT 57.410 191.920 57.730 191.980 ;
        RECT 59.340 191.920 59.480 192.060 ;
        RECT 57.410 191.780 59.480 191.920 ;
        RECT 57.410 191.720 57.730 191.780 ;
        RECT 62.930 191.720 63.250 191.980 ;
        RECT 63.940 191.920 64.080 192.120 ;
        RECT 64.325 192.120 66.930 192.260 ;
        RECT 64.325 192.075 64.615 192.120 ;
        RECT 66.610 192.060 66.930 192.120 ;
        RECT 68.910 192.260 69.230 192.320 ;
        RECT 74.445 192.260 74.735 192.305 ;
        RECT 68.910 192.120 74.735 192.260 ;
        RECT 68.910 192.060 69.230 192.120 ;
        RECT 74.445 192.075 74.735 192.120 ;
        RECT 80.870 192.060 81.190 192.320 ;
        RECT 82.250 192.060 82.570 192.320 ;
        RECT 82.710 192.060 83.030 192.320 ;
        RECT 87.400 192.305 87.540 192.460 ;
        RECT 89.610 192.460 97.290 192.600 ;
        RECT 97.520 192.600 97.660 192.755 ;
        RECT 99.270 192.740 99.590 193.000 ;
        RECT 102.950 192.740 103.270 193.000 ;
        RECT 107.550 192.940 107.870 193.000 ;
        RECT 112.625 192.940 112.915 192.985 ;
        RECT 107.550 192.800 112.915 192.940 ;
        RECT 107.550 192.740 107.870 192.800 ;
        RECT 112.625 192.755 112.915 192.800 ;
        RECT 114.910 192.740 115.230 193.000 ;
        RECT 103.870 192.600 104.190 192.660 ;
        RECT 97.520 192.460 101.340 192.600 ;
        RECT 89.610 192.400 89.930 192.460 ;
        RECT 96.970 192.400 97.290 192.460 ;
        RECT 87.325 192.075 87.615 192.305 ;
        RECT 88.660 192.260 88.950 192.305 ;
        RECT 92.370 192.260 92.690 192.320 ;
        RECT 88.660 192.120 92.690 192.260 ;
        RECT 88.660 192.075 88.950 192.120 ;
        RECT 92.370 192.060 92.690 192.120 ;
        RECT 94.670 192.260 94.990 192.320 ;
        RECT 99.270 192.260 99.590 192.320 ;
        RECT 101.200 192.305 101.340 192.460 ;
        RECT 101.660 192.460 104.190 192.600 ;
        RECT 101.660 192.305 101.800 192.460 ;
        RECT 103.870 192.400 104.190 192.460 ;
        RECT 100.205 192.260 100.495 192.305 ;
        RECT 94.670 192.120 99.040 192.260 ;
        RECT 94.670 192.060 94.990 192.120 ;
        RECT 66.150 191.920 66.470 191.980 ;
        RECT 63.940 191.780 66.470 191.920 ;
        RECT 66.150 191.720 66.470 191.780 ;
        RECT 67.070 191.920 67.390 191.980 ;
        RECT 72.605 191.920 72.895 191.965 ;
        RECT 75.350 191.920 75.670 191.980 ;
        RECT 67.070 191.780 75.670 191.920 ;
        RECT 67.070 191.720 67.390 191.780 ;
        RECT 72.605 191.735 72.895 191.780 ;
        RECT 75.350 191.720 75.670 191.780 ;
        RECT 88.205 191.920 88.495 191.965 ;
        RECT 89.395 191.920 89.685 191.965 ;
        RECT 91.915 191.920 92.205 191.965 ;
        RECT 88.205 191.780 92.205 191.920 ;
        RECT 88.205 191.735 88.495 191.780 ;
        RECT 89.395 191.735 89.685 191.780 ;
        RECT 91.915 191.735 92.205 191.780 ;
        RECT 98.365 191.735 98.655 191.965 ;
        RECT 65.230 191.580 65.550 191.640 ;
        RECT 56.505 191.440 65.550 191.580 ;
        RECT 56.505 191.395 56.795 191.440 ;
        RECT 65.230 191.380 65.550 191.440 ;
        RECT 87.810 191.580 88.100 191.625 ;
        RECT 89.910 191.580 90.200 191.625 ;
        RECT 91.480 191.580 91.770 191.625 ;
        RECT 87.810 191.440 91.770 191.580 ;
        RECT 87.810 191.395 88.100 191.440 ;
        RECT 89.910 191.395 90.200 191.440 ;
        RECT 91.480 191.395 91.770 191.440 ;
        RECT 98.440 191.300 98.580 191.735 ;
        RECT 98.900 191.580 99.040 192.120 ;
        RECT 99.270 192.120 100.495 192.260 ;
        RECT 99.270 192.060 99.590 192.120 ;
        RECT 100.205 192.075 100.495 192.120 ;
        RECT 101.125 192.075 101.415 192.305 ;
        RECT 101.585 192.075 101.875 192.305 ;
        RECT 102.490 192.060 102.810 192.320 ;
        RECT 104.345 192.260 104.635 192.305 ;
        RECT 103.040 192.120 104.635 192.260 ;
        RECT 99.730 191.920 100.050 191.980 ;
        RECT 103.040 191.920 103.180 192.120 ;
        RECT 104.345 192.075 104.635 192.120 ;
        RECT 106.170 192.060 106.490 192.320 ;
        RECT 113.085 192.260 113.375 192.305 ;
        RECT 120.890 192.260 121.210 192.320 ;
        RECT 113.085 192.120 121.210 192.260 ;
        RECT 113.085 192.075 113.375 192.120 ;
        RECT 120.890 192.060 121.210 192.120 ;
        RECT 99.730 191.780 103.180 191.920 ;
        RECT 99.730 191.720 100.050 191.780 ;
        RECT 103.870 191.720 104.190 191.980 ;
        RECT 104.790 191.720 105.110 191.980 ;
        RECT 105.250 191.720 105.570 191.980 ;
        RECT 107.090 191.920 107.410 191.980 ;
        RECT 111.705 191.920 111.995 191.965 ;
        RECT 107.090 191.780 111.995 191.920 ;
        RECT 107.090 191.720 107.410 191.780 ;
        RECT 111.705 191.735 111.995 191.780 ;
        RECT 100.665 191.580 100.955 191.625 ;
        RECT 98.900 191.440 100.955 191.580 ;
        RECT 100.665 191.395 100.955 191.440 ;
        RECT 23.830 191.040 24.150 191.300 ;
        RECT 39.930 191.040 40.250 191.300 ;
        RECT 41.785 191.240 42.075 191.285 ;
        RECT 42.690 191.240 43.010 191.300 ;
        RECT 41.785 191.100 43.010 191.240 ;
        RECT 41.785 191.055 42.075 191.100 ;
        RECT 42.690 191.040 43.010 191.100 ;
        RECT 48.225 191.240 48.515 191.285 ;
        RECT 49.145 191.240 49.435 191.285 ;
        RECT 48.225 191.100 49.435 191.240 ;
        RECT 48.225 191.055 48.515 191.100 ;
        RECT 49.145 191.055 49.435 191.100 ;
        RECT 52.350 191.040 52.670 191.300 ;
        RECT 53.270 191.240 53.590 191.300 ;
        RECT 56.950 191.240 57.270 191.300 ;
        RECT 53.270 191.100 57.270 191.240 ;
        RECT 53.270 191.040 53.590 191.100 ;
        RECT 56.950 191.040 57.270 191.100 ;
        RECT 57.410 191.040 57.730 191.300 ;
        RECT 60.170 191.040 60.490 191.300 ;
        RECT 60.645 191.240 60.935 191.285 ;
        RECT 61.090 191.240 61.410 191.300 ;
        RECT 60.645 191.100 61.410 191.240 ;
        RECT 60.645 191.055 60.935 191.100 ;
        RECT 61.090 191.040 61.410 191.100 ;
        RECT 63.850 191.040 64.170 191.300 ;
        RECT 69.830 191.040 70.150 191.300 ;
        RECT 73.510 191.040 73.830 191.300 ;
        RECT 94.670 191.240 94.990 191.300 ;
        RECT 95.145 191.240 95.435 191.285 ;
        RECT 94.670 191.100 95.435 191.240 ;
        RECT 94.670 191.040 94.990 191.100 ;
        RECT 95.145 191.055 95.435 191.100 ;
        RECT 98.350 191.240 98.670 191.300 ;
        RECT 106.630 191.240 106.950 191.300 ;
        RECT 98.350 191.100 106.950 191.240 ;
        RECT 98.350 191.040 98.670 191.100 ;
        RECT 106.630 191.040 106.950 191.100 ;
        RECT 17.320 190.420 147.040 190.900 ;
        RECT 35.790 190.020 36.110 190.280 ;
        RECT 36.725 190.035 37.015 190.265 ;
        RECT 48.685 190.220 48.975 190.265 ;
        RECT 57.410 190.220 57.730 190.280 ;
        RECT 63.405 190.220 63.695 190.265 ;
        RECT 48.685 190.080 63.695 190.220 ;
        RECT 48.685 190.035 48.975 190.080 ;
        RECT 22.030 189.880 22.320 189.925 ;
        RECT 24.130 189.880 24.420 189.925 ;
        RECT 25.700 189.880 25.990 189.925 ;
        RECT 22.030 189.740 25.990 189.880 ;
        RECT 22.030 189.695 22.320 189.740 ;
        RECT 24.130 189.695 24.420 189.740 ;
        RECT 25.700 189.695 25.990 189.740 ;
        RECT 29.365 189.880 29.655 189.925 ;
        RECT 36.800 189.880 36.940 190.035 ;
        RECT 57.410 190.020 57.730 190.080 ;
        RECT 63.405 190.035 63.695 190.080 ;
        RECT 66.150 190.020 66.470 190.280 ;
        RECT 66.610 190.020 66.930 190.280 ;
        RECT 75.350 190.220 75.670 190.280 ;
        RECT 77.205 190.220 77.495 190.265 ;
        RECT 75.350 190.080 77.495 190.220 ;
        RECT 75.350 190.020 75.670 190.080 ;
        RECT 77.205 190.035 77.495 190.080 ;
        RECT 91.450 190.020 91.770 190.280 ;
        RECT 92.370 190.020 92.690 190.280 ;
        RECT 96.065 190.220 96.355 190.265 ;
        RECT 104.790 190.220 105.110 190.280 ;
        RECT 108.025 190.220 108.315 190.265 ;
        RECT 92.920 190.080 95.820 190.220 ;
        RECT 29.365 189.740 36.940 189.880 ;
        RECT 29.365 189.695 29.655 189.740 ;
        RECT 40.390 189.680 40.710 189.940 ;
        RECT 46.370 189.880 46.690 189.940 ;
        RECT 57.870 189.880 58.190 189.940 ;
        RECT 58.345 189.880 58.635 189.925 ;
        RECT 63.850 189.880 64.170 189.940 ;
        RECT 69.370 189.880 69.690 189.940 ;
        RECT 44.160 189.740 46.690 189.880 ;
        RECT 22.425 189.540 22.715 189.585 ;
        RECT 23.615 189.540 23.905 189.585 ;
        RECT 26.135 189.540 26.425 189.585 ;
        RECT 40.480 189.540 40.620 189.680 ;
        RECT 44.160 189.585 44.300 189.740 ;
        RECT 46.370 189.680 46.690 189.740 ;
        RECT 49.680 189.740 53.040 189.880 ;
        RECT 22.425 189.400 26.425 189.540 ;
        RECT 22.425 189.355 22.715 189.400 ;
        RECT 23.615 189.355 23.905 189.400 ;
        RECT 26.135 189.355 26.425 189.400 ;
        RECT 28.980 189.400 40.620 189.540 ;
        RECT 28.980 189.260 29.120 189.400 ;
        RECT 21.545 189.200 21.835 189.245 ;
        RECT 25.210 189.200 25.530 189.260 ;
        RECT 21.545 189.060 25.530 189.200 ;
        RECT 21.545 189.015 21.835 189.060 ;
        RECT 25.210 189.000 25.530 189.060 ;
        RECT 28.890 189.000 29.210 189.260 ;
        RECT 29.825 189.200 30.115 189.245 ;
        RECT 29.825 189.060 31.420 189.200 ;
        RECT 29.825 189.015 30.115 189.060 ;
        RECT 22.910 188.905 23.230 188.920 ;
        RECT 22.880 188.675 23.230 188.905 ;
        RECT 22.910 188.660 23.230 188.675 ;
        RECT 26.130 188.860 26.450 188.920 ;
        RECT 29.900 188.860 30.040 189.015 ;
        RECT 26.130 188.720 30.040 188.860 ;
        RECT 26.130 188.660 26.450 188.720 ;
        RECT 28.430 188.320 28.750 188.580 ;
        RECT 30.730 188.320 31.050 188.580 ;
        RECT 31.280 188.520 31.420 189.060 ;
        RECT 31.650 189.000 31.970 189.260 ;
        RECT 32.570 189.000 32.890 189.260 ;
        RECT 33.120 189.245 33.260 189.400 ;
        RECT 44.085 189.355 44.375 189.585 ;
        RECT 44.545 189.540 44.835 189.585 ;
        RECT 45.910 189.540 46.230 189.600 ;
        RECT 44.545 189.400 46.230 189.540 ;
        RECT 44.545 189.355 44.835 189.400 ;
        RECT 45.910 189.340 46.230 189.400 ;
        RECT 33.045 189.200 33.335 189.245 ;
        RECT 33.505 189.200 33.795 189.245 ;
        RECT 33.045 189.060 33.795 189.200 ;
        RECT 33.045 189.015 33.335 189.060 ;
        RECT 33.505 189.015 33.795 189.060 ;
        RECT 33.950 189.200 34.270 189.260 ;
        RECT 34.425 189.200 34.715 189.245 ;
        RECT 33.950 189.060 38.320 189.200 ;
        RECT 33.950 189.000 34.270 189.060 ;
        RECT 34.425 189.015 34.715 189.060 ;
        RECT 32.110 188.860 32.430 188.920 ;
        RECT 35.345 188.860 35.635 188.905 ;
        RECT 36.565 188.860 36.855 188.905 ;
        RECT 32.110 188.720 33.260 188.860 ;
        RECT 32.110 188.660 32.430 188.720 ;
        RECT 32.570 188.520 32.890 188.580 ;
        RECT 31.280 188.380 32.890 188.520 ;
        RECT 33.120 188.520 33.260 188.720 ;
        RECT 35.345 188.720 36.855 188.860 ;
        RECT 35.345 188.675 35.635 188.720 ;
        RECT 36.565 188.675 36.855 188.720 ;
        RECT 37.645 188.675 37.935 188.905 ;
        RECT 38.180 188.860 38.320 189.060 ;
        RECT 39.010 189.000 39.330 189.260 ;
        RECT 40.405 189.200 40.695 189.245 ;
        RECT 40.850 189.200 41.170 189.260 ;
        RECT 42.705 189.200 42.995 189.245 ;
        RECT 40.405 189.060 42.995 189.200 ;
        RECT 40.405 189.015 40.695 189.060 ;
        RECT 40.850 189.000 41.170 189.060 ;
        RECT 42.705 189.015 42.995 189.060 ;
        RECT 43.150 189.200 43.470 189.260 ;
        RECT 49.680 189.245 49.820 189.740 ;
        RECT 50.510 189.340 50.830 189.600 ;
        RECT 48.685 189.200 48.975 189.245 ;
        RECT 43.150 189.060 48.975 189.200 ;
        RECT 41.310 188.860 41.630 188.920 ;
        RECT 38.180 188.720 41.630 188.860 ;
        RECT 37.720 188.520 37.860 188.675 ;
        RECT 41.310 188.660 41.630 188.720 ;
        RECT 33.120 188.380 37.860 188.520 ;
        RECT 42.780 188.520 42.920 189.015 ;
        RECT 43.150 189.000 43.470 189.060 ;
        RECT 48.685 189.015 48.975 189.060 ;
        RECT 49.605 189.015 49.895 189.245 ;
        RECT 50.065 189.200 50.355 189.245 ;
        RECT 50.600 189.200 50.740 189.340 ;
        RECT 51.445 189.200 51.735 189.245 ;
        RECT 52.350 189.200 52.670 189.260 ;
        RECT 50.065 189.060 50.740 189.200 ;
        RECT 51.060 189.060 52.670 189.200 ;
        RECT 52.900 189.200 53.040 189.740 ;
        RECT 53.360 189.740 56.260 189.880 ;
        RECT 53.360 189.585 53.500 189.740 ;
        RECT 53.285 189.355 53.575 189.585 ;
        RECT 53.745 189.540 54.035 189.585 ;
        RECT 55.570 189.540 55.890 189.600 ;
        RECT 53.745 189.400 55.890 189.540 ;
        RECT 56.120 189.540 56.260 189.740 ;
        RECT 57.870 189.740 58.635 189.880 ;
        RECT 57.870 189.680 58.190 189.740 ;
        RECT 58.345 189.695 58.635 189.740 ;
        RECT 58.880 189.740 64.170 189.880 ;
        RECT 58.880 189.540 59.020 189.740 ;
        RECT 63.850 189.680 64.170 189.740 ;
        RECT 66.700 189.740 69.690 189.880 ;
        RECT 56.120 189.400 59.020 189.540 ;
        RECT 53.745 189.355 54.035 189.400 ;
        RECT 55.570 189.340 55.890 189.400 ;
        RECT 60.630 189.340 60.950 189.600 ;
        RECT 62.025 189.540 62.315 189.585 ;
        RECT 66.700 189.540 66.840 189.740 ;
        RECT 69.370 189.680 69.690 189.740 ;
        RECT 70.790 189.880 71.080 189.925 ;
        RECT 72.890 189.880 73.180 189.925 ;
        RECT 74.460 189.880 74.750 189.925 ;
        RECT 92.920 189.880 93.060 190.080 ;
        RECT 70.790 189.740 74.750 189.880 ;
        RECT 70.790 189.695 71.080 189.740 ;
        RECT 72.890 189.695 73.180 189.740 ;
        RECT 74.460 189.695 74.750 189.740 ;
        RECT 91.540 189.740 93.060 189.880 ;
        RECT 62.025 189.400 66.840 189.540 ;
        RECT 62.025 189.355 62.315 189.400 ;
        RECT 67.070 189.340 67.390 189.600 ;
        RECT 71.185 189.540 71.475 189.585 ;
        RECT 72.375 189.540 72.665 189.585 ;
        RECT 74.895 189.540 75.185 189.585 ;
        RECT 71.185 189.400 75.185 189.540 ;
        RECT 71.185 189.355 71.475 189.400 ;
        RECT 72.375 189.355 72.665 189.400 ;
        RECT 74.895 189.355 75.185 189.400 ;
        RECT 52.900 189.060 53.500 189.200 ;
        RECT 50.065 189.015 50.355 189.060 ;
        RECT 45.450 188.660 45.770 188.920 ;
        RECT 46.370 188.660 46.690 188.920 ;
        RECT 48.760 188.860 48.900 189.015 ;
        RECT 51.060 188.860 51.200 189.060 ;
        RECT 51.445 189.015 51.735 189.060 ;
        RECT 52.350 189.000 52.670 189.060 ;
        RECT 48.760 188.720 51.200 188.860 ;
        RECT 53.360 188.860 53.500 189.060 ;
        RECT 54.190 189.000 54.510 189.260 ;
        RECT 54.665 189.200 54.955 189.245 ;
        RECT 55.110 189.200 55.430 189.260 ;
        RECT 54.665 189.060 55.430 189.200 ;
        RECT 54.665 189.015 54.955 189.060 ;
        RECT 55.110 189.000 55.430 189.060 ;
        RECT 57.410 189.000 57.730 189.260 ;
        RECT 59.250 189.200 59.570 189.260 ;
        RECT 63.405 189.200 63.695 189.245 ;
        RECT 59.250 189.060 63.695 189.200 ;
        RECT 59.250 189.000 59.570 189.060 ;
        RECT 63.405 189.015 63.695 189.060 ;
        RECT 65.230 189.000 65.550 189.260 ;
        RECT 65.690 189.000 66.010 189.260 ;
        RECT 68.910 189.000 69.230 189.260 ;
        RECT 69.830 189.000 70.150 189.260 ;
        RECT 70.305 189.015 70.595 189.245 ;
        RECT 71.640 189.015 71.930 189.245 ;
        RECT 78.570 189.200 78.890 189.260 ;
        RECT 73.830 189.060 78.890 189.200 ;
        RECT 56.965 188.860 57.255 188.905 ;
        RECT 53.360 188.720 57.255 188.860 ;
        RECT 56.965 188.675 57.255 188.720 ;
        RECT 58.345 188.860 58.635 188.905 ;
        RECT 58.345 188.720 62.700 188.860 ;
        RECT 58.345 188.675 58.635 188.720 ;
        RECT 45.540 188.520 45.680 188.660 ;
        RECT 42.780 188.380 45.680 188.520 ;
        RECT 46.830 188.520 47.150 188.580 ;
        RECT 47.305 188.520 47.595 188.565 ;
        RECT 46.830 188.380 47.595 188.520 ;
        RECT 32.570 188.320 32.890 188.380 ;
        RECT 46.830 188.320 47.150 188.380 ;
        RECT 47.305 188.335 47.595 188.380 ;
        RECT 52.365 188.520 52.655 188.565 ;
        RECT 53.270 188.520 53.590 188.580 ;
        RECT 52.365 188.380 53.590 188.520 ;
        RECT 52.365 188.335 52.655 188.380 ;
        RECT 53.270 188.320 53.590 188.380 ;
        RECT 55.585 188.520 55.875 188.565 ;
        RECT 56.490 188.520 56.810 188.580 ;
        RECT 55.585 188.380 56.810 188.520 ;
        RECT 55.585 188.335 55.875 188.380 ;
        RECT 56.490 188.320 56.810 188.380 ;
        RECT 61.090 188.320 61.410 188.580 ;
        RECT 62.560 188.565 62.700 188.720 ;
        RECT 62.485 188.335 62.775 188.565 ;
        RECT 69.370 188.320 69.690 188.580 ;
        RECT 70.380 188.520 70.520 189.015 ;
        RECT 71.210 188.860 71.530 188.920 ;
        RECT 71.760 188.860 71.900 189.015 ;
        RECT 71.210 188.720 71.900 188.860 ;
        RECT 71.210 188.660 71.530 188.720 ;
        RECT 73.830 188.520 73.970 189.060 ;
        RECT 78.570 189.000 78.890 189.060 ;
        RECT 85.010 189.000 85.330 189.260 ;
        RECT 86.405 189.015 86.695 189.245 ;
        RECT 86.480 188.860 86.620 189.015 ;
        RECT 89.150 189.000 89.470 189.260 ;
        RECT 90.085 189.015 90.375 189.245 ;
        RECT 89.625 188.860 89.915 188.905 ;
        RECT 86.480 188.720 89.915 188.860 ;
        RECT 90.160 188.860 90.300 189.015 ;
        RECT 90.530 189.000 90.850 189.260 ;
        RECT 91.540 189.245 91.680 189.740 ;
        RECT 94.670 189.680 94.990 189.940 ;
        RECT 95.680 189.880 95.820 190.080 ;
        RECT 96.065 190.080 105.110 190.220 ;
        RECT 96.065 190.035 96.355 190.080 ;
        RECT 104.790 190.020 105.110 190.080 ;
        RECT 105.340 190.080 108.315 190.220 ;
        RECT 99.730 189.880 100.050 189.940 ;
        RECT 105.340 189.880 105.480 190.080 ;
        RECT 108.025 190.035 108.315 190.080 ;
        RECT 108.470 189.880 108.790 189.940 ;
        RECT 95.680 189.740 100.050 189.880 ;
        RECT 99.730 189.680 100.050 189.740 ;
        RECT 103.960 189.740 105.480 189.880 ;
        RECT 107.180 189.740 108.790 189.880 ;
        RECT 94.760 189.540 94.900 189.680 ;
        RECT 96.050 189.540 96.370 189.600 ;
        RECT 92.920 189.400 94.900 189.540 ;
        RECT 95.220 189.400 96.370 189.540 ;
        RECT 92.920 189.245 93.060 189.400 ;
        RECT 91.465 189.015 91.755 189.245 ;
        RECT 92.845 189.015 93.135 189.245 ;
        RECT 93.305 189.015 93.595 189.245 ;
        RECT 93.765 189.200 94.055 189.245 ;
        RECT 94.210 189.200 94.530 189.260 ;
        RECT 93.765 189.060 94.530 189.200 ;
        RECT 93.765 189.015 94.055 189.060 ;
        RECT 93.380 188.860 93.520 189.015 ;
        RECT 94.210 189.000 94.530 189.060 ;
        RECT 94.685 189.200 94.975 189.245 ;
        RECT 95.220 189.200 95.360 189.400 ;
        RECT 96.050 189.340 96.370 189.400 ;
        RECT 100.190 189.540 100.510 189.600 ;
        RECT 103.960 189.540 104.100 189.740 ;
        RECT 107.180 189.540 107.320 189.740 ;
        RECT 108.470 189.680 108.790 189.740 ;
        RECT 100.190 189.400 104.100 189.540 ;
        RECT 100.190 189.340 100.510 189.400 ;
        RECT 94.685 189.060 95.360 189.200 ;
        RECT 95.590 189.200 95.910 189.260 ;
        RECT 96.985 189.200 97.275 189.245 ;
        RECT 95.590 189.060 97.275 189.200 ;
        RECT 94.685 189.015 94.975 189.060 ;
        RECT 95.590 189.000 95.910 189.060 ;
        RECT 96.985 189.015 97.275 189.060 ;
        RECT 97.445 189.200 97.735 189.245 ;
        RECT 98.350 189.200 98.670 189.260 ;
        RECT 97.445 189.060 98.670 189.200 ;
        RECT 97.445 189.015 97.735 189.060 ;
        RECT 98.350 189.000 98.670 189.060 ;
        RECT 98.810 189.000 99.130 189.260 ;
        RECT 99.285 189.200 99.575 189.245 ;
        RECT 101.110 189.200 101.430 189.260 ;
        RECT 102.950 189.245 103.270 189.260 ;
        RECT 103.960 189.245 104.100 189.400 ;
        RECT 104.880 189.400 107.320 189.540 ;
        RECT 107.550 189.540 107.870 189.600 ;
        RECT 113.085 189.540 113.375 189.585 ;
        RECT 107.550 189.400 113.375 189.540 ;
        RECT 104.880 189.245 105.020 189.400 ;
        RECT 107.550 189.340 107.870 189.400 ;
        RECT 113.085 189.355 113.375 189.400 ;
        RECT 99.285 189.060 101.430 189.200 ;
        RECT 99.285 189.015 99.575 189.060 ;
        RECT 101.110 189.000 101.430 189.060 ;
        RECT 102.940 189.015 103.270 189.245 ;
        RECT 103.885 189.015 104.175 189.245 ;
        RECT 104.800 189.015 105.090 189.245 ;
        RECT 105.265 189.015 105.555 189.245 ;
        RECT 102.950 189.000 103.270 189.015 ;
        RECT 97.890 188.860 98.210 188.920 ;
        RECT 100.650 188.860 100.970 188.920 ;
        RECT 90.160 188.720 90.760 188.860 ;
        RECT 93.380 188.720 94.900 188.860 ;
        RECT 89.625 188.675 89.915 188.720 ;
        RECT 70.380 188.380 73.970 188.520 ;
        RECT 84.090 188.320 84.410 188.580 ;
        RECT 85.930 188.320 86.250 188.580 ;
        RECT 90.620 188.520 90.760 188.720 ;
        RECT 94.760 188.580 94.900 188.720 ;
        RECT 97.890 188.720 100.970 188.860 ;
        RECT 97.890 188.660 98.210 188.720 ;
        RECT 100.650 188.660 100.970 188.720 ;
        RECT 94.210 188.520 94.530 188.580 ;
        RECT 90.620 188.380 94.530 188.520 ;
        RECT 94.210 188.320 94.530 188.380 ;
        RECT 94.670 188.320 94.990 188.580 ;
        RECT 95.605 188.520 95.895 188.565 ;
        RECT 96.050 188.520 96.370 188.580 ;
        RECT 95.605 188.380 96.370 188.520 ;
        RECT 95.605 188.335 95.895 188.380 ;
        RECT 96.050 188.320 96.370 188.380 ;
        RECT 100.190 188.520 100.510 188.580 ;
        RECT 101.200 188.520 101.340 189.000 ;
        RECT 101.570 188.660 101.890 188.920 ;
        RECT 103.425 188.675 103.715 188.905 ;
        RECT 105.340 188.860 105.480 189.015 ;
        RECT 105.710 189.000 106.030 189.260 ;
        RECT 106.630 189.200 106.950 189.260 ;
        RECT 108.025 189.200 108.315 189.245 ;
        RECT 106.630 189.060 108.315 189.200 ;
        RECT 106.630 189.000 106.950 189.060 ;
        RECT 108.025 189.015 108.315 189.060 ;
        RECT 108.945 189.015 109.235 189.245 ;
        RECT 106.185 188.860 106.475 188.905 ;
        RECT 109.020 188.860 109.160 189.015 ;
        RECT 117.210 189.000 117.530 189.260 ;
        RECT 123.205 189.200 123.495 189.245 ;
        RECT 124.570 189.200 124.890 189.260 ;
        RECT 123.205 189.060 124.890 189.200 ;
        RECT 123.205 189.015 123.495 189.060 ;
        RECT 124.570 189.000 124.890 189.060 ;
        RECT 125.030 189.000 125.350 189.260 ;
        RECT 105.340 188.720 106.475 188.860 ;
        RECT 106.185 188.675 106.475 188.720 ;
        RECT 106.720 188.720 109.160 188.860 ;
        RECT 112.165 188.860 112.455 188.905 ;
        RECT 118.130 188.860 118.450 188.920 ;
        RECT 112.165 188.720 118.450 188.860 ;
        RECT 100.190 188.380 101.340 188.520 ;
        RECT 100.190 188.320 100.510 188.380 ;
        RECT 102.030 188.320 102.350 188.580 ;
        RECT 102.490 188.520 102.810 188.580 ;
        RECT 103.500 188.520 103.640 188.675 ;
        RECT 105.250 188.520 105.570 188.580 ;
        RECT 106.720 188.520 106.860 188.720 ;
        RECT 112.165 188.675 112.455 188.720 ;
        RECT 118.130 188.660 118.450 188.720 ;
        RECT 123.665 188.675 123.955 188.905 ;
        RECT 124.125 188.860 124.415 188.905 ;
        RECT 126.870 188.860 127.190 188.920 ;
        RECT 124.125 188.720 127.190 188.860 ;
        RECT 124.125 188.675 124.415 188.720 ;
        RECT 102.490 188.380 106.860 188.520 ;
        RECT 102.490 188.320 102.810 188.380 ;
        RECT 105.250 188.320 105.570 188.380 ;
        RECT 110.310 188.320 110.630 188.580 ;
        RECT 112.625 188.520 112.915 188.565 ;
        RECT 114.465 188.520 114.755 188.565 ;
        RECT 112.625 188.380 114.755 188.520 ;
        RECT 112.625 188.335 112.915 188.380 ;
        RECT 114.465 188.335 114.755 188.380 ;
        RECT 122.270 188.320 122.590 188.580 ;
        RECT 123.740 188.520 123.880 188.675 ;
        RECT 126.870 188.660 127.190 188.720 ;
        RECT 131.930 188.520 132.250 188.580 ;
        RECT 123.740 188.380 132.250 188.520 ;
        RECT 131.930 188.320 132.250 188.380 ;
        RECT 17.320 187.700 147.040 188.180 ;
        RECT 19.245 187.500 19.535 187.545 ;
        RECT 21.530 187.500 21.850 187.560 ;
        RECT 19.245 187.360 21.850 187.500 ;
        RECT 19.245 187.315 19.535 187.360 ;
        RECT 21.530 187.300 21.850 187.360 ;
        RECT 25.210 187.300 25.530 187.560 ;
        RECT 27.525 187.500 27.815 187.545 ;
        RECT 28.890 187.500 29.210 187.560 ;
        RECT 43.150 187.500 43.470 187.560 ;
        RECT 27.525 187.360 29.210 187.500 ;
        RECT 27.525 187.315 27.815 187.360 ;
        RECT 28.890 187.300 29.210 187.360 ;
        RECT 37.720 187.360 43.470 187.500 ;
        RECT 23.830 187.160 24.150 187.220 ;
        RECT 24.810 187.160 25.100 187.205 ;
        RECT 23.830 187.020 25.100 187.160 ;
        RECT 23.830 186.960 24.150 187.020 ;
        RECT 24.810 186.975 25.100 187.020 ;
        RECT 25.300 186.820 25.440 187.300 ;
        RECT 27.985 187.160 28.275 187.205 ;
        RECT 31.650 187.160 31.970 187.220 ;
        RECT 37.720 187.160 37.860 187.360 ;
        RECT 43.150 187.300 43.470 187.360 ;
        RECT 51.890 187.300 52.210 187.560 ;
        RECT 54.190 187.300 54.510 187.560 ;
        RECT 54.650 187.300 54.970 187.560 ;
        RECT 55.110 187.500 55.430 187.560 ;
        RECT 60.630 187.500 60.950 187.560 ;
        RECT 55.110 187.360 60.950 187.500 ;
        RECT 55.110 187.300 55.430 187.360 ;
        RECT 27.985 187.020 31.970 187.160 ;
        RECT 27.985 186.975 28.275 187.020 ;
        RECT 31.650 186.960 31.970 187.020 ;
        RECT 33.580 187.020 37.860 187.160 ;
        RECT 26.145 186.820 26.435 186.865 ;
        RECT 25.300 186.680 26.435 186.820 ;
        RECT 26.145 186.635 26.435 186.680 ;
        RECT 28.430 186.820 28.750 186.880 ;
        RECT 33.580 186.865 33.720 187.020 ;
        RECT 28.430 186.680 32.340 186.820 ;
        RECT 28.430 186.620 28.750 186.680 ;
        RECT 21.555 186.480 21.845 186.525 ;
        RECT 24.075 186.480 24.365 186.525 ;
        RECT 25.265 186.480 25.555 186.525 ;
        RECT 21.555 186.340 25.555 186.480 ;
        RECT 21.555 186.295 21.845 186.340 ;
        RECT 24.075 186.295 24.365 186.340 ;
        RECT 25.265 186.295 25.555 186.340 ;
        RECT 28.890 186.480 29.210 186.540 ;
        RECT 30.745 186.480 31.035 186.525 ;
        RECT 28.890 186.340 31.035 186.480 ;
        RECT 28.890 186.280 29.210 186.340 ;
        RECT 30.745 186.295 31.035 186.340 ;
        RECT 31.190 186.280 31.510 186.540 ;
        RECT 32.200 186.525 32.340 186.680 ;
        RECT 33.505 186.635 33.795 186.865 ;
        RECT 34.425 186.820 34.715 186.865 ;
        RECT 35.790 186.820 36.110 186.880 ;
        RECT 34.425 186.680 36.110 186.820 ;
        RECT 34.425 186.635 34.715 186.680 ;
        RECT 31.665 186.295 31.955 186.525 ;
        RECT 32.125 186.480 32.415 186.525 ;
        RECT 34.500 186.480 34.640 186.635 ;
        RECT 35.790 186.620 36.110 186.680 ;
        RECT 37.170 186.620 37.490 186.880 ;
        RECT 37.720 186.865 37.860 187.020 ;
        RECT 39.945 187.160 40.235 187.205 ;
        RECT 45.465 187.160 45.755 187.205 ;
        RECT 39.945 187.020 45.755 187.160 ;
        RECT 39.945 186.975 40.235 187.020 ;
        RECT 45.465 186.975 45.755 187.020 ;
        RECT 46.830 186.960 47.150 187.220 ;
        RECT 53.730 187.160 54.050 187.220 ;
        RECT 51.060 187.020 54.050 187.160 ;
        RECT 51.060 186.880 51.200 187.020 ;
        RECT 53.730 186.960 54.050 187.020 ;
        RECT 37.645 186.820 37.935 186.865 ;
        RECT 38.550 186.820 38.870 186.880 ;
        RECT 37.645 186.680 38.870 186.820 ;
        RECT 37.645 186.635 37.935 186.680 ;
        RECT 38.550 186.620 38.870 186.680 ;
        RECT 39.025 186.820 39.315 186.865 ;
        RECT 39.470 186.820 39.790 186.880 ;
        RECT 39.025 186.680 39.790 186.820 ;
        RECT 39.025 186.635 39.315 186.680 ;
        RECT 39.470 186.620 39.790 186.680 ;
        RECT 40.390 186.620 40.710 186.880 ;
        RECT 40.865 186.635 41.155 186.865 ;
        RECT 41.310 186.820 41.630 186.880 ;
        RECT 43.625 186.820 43.915 186.865 ;
        RECT 41.310 186.680 43.915 186.820 ;
        RECT 39.930 186.480 40.250 186.540 ;
        RECT 32.125 186.340 34.640 186.480 ;
        RECT 35.420 186.340 40.250 186.480 ;
        RECT 40.940 186.480 41.080 186.635 ;
        RECT 41.310 186.620 41.630 186.680 ;
        RECT 43.625 186.635 43.915 186.680 ;
        RECT 44.395 186.820 44.685 186.865 ;
        RECT 44.990 186.820 45.310 186.880 ;
        RECT 45.925 186.820 46.215 186.865 ;
        RECT 44.395 186.635 44.760 186.820 ;
        RECT 43.150 186.480 43.470 186.540 ;
        RECT 40.940 186.340 43.470 186.480 ;
        RECT 44.620 186.480 44.760 186.635 ;
        RECT 44.990 186.680 46.215 186.820 ;
        RECT 44.990 186.620 45.310 186.680 ;
        RECT 45.925 186.635 46.215 186.680 ;
        RECT 50.970 186.620 51.290 186.880 ;
        RECT 51.905 186.635 52.195 186.865 ;
        RECT 46.370 186.480 46.690 186.540 ;
        RECT 44.620 186.340 46.690 186.480 ;
        RECT 51.980 186.480 52.120 186.635 ;
        RECT 52.350 186.620 52.670 186.880 ;
        RECT 55.570 186.620 55.890 186.880 ;
        RECT 56.045 186.820 56.335 186.865 ;
        RECT 56.950 186.820 57.270 186.880 ;
        RECT 56.045 186.680 57.270 186.820 ;
        RECT 56.045 186.635 56.335 186.680 ;
        RECT 56.950 186.620 57.270 186.680 ;
        RECT 57.410 186.620 57.730 186.880 ;
        RECT 58.880 186.865 59.020 187.360 ;
        RECT 60.630 187.300 60.950 187.360 ;
        RECT 61.090 187.300 61.410 187.560 ;
        RECT 71.210 187.300 71.530 187.560 ;
        RECT 78.570 187.300 78.890 187.560 ;
        RECT 85.930 187.500 86.250 187.560 ;
        RECT 87.785 187.500 88.075 187.545 ;
        RECT 90.530 187.500 90.850 187.560 ;
        RECT 85.930 187.360 90.850 187.500 ;
        RECT 85.930 187.300 86.250 187.360 ;
        RECT 87.785 187.315 88.075 187.360 ;
        RECT 90.530 187.300 90.850 187.360 ;
        RECT 98.810 187.500 99.130 187.560 ;
        RECT 100.665 187.500 100.955 187.545 ;
        RECT 98.810 187.360 100.955 187.500 ;
        RECT 98.810 187.300 99.130 187.360 ;
        RECT 100.665 187.315 100.955 187.360 ;
        RECT 101.110 187.500 101.430 187.560 ;
        RECT 103.870 187.500 104.190 187.560 ;
        RECT 104.345 187.500 104.635 187.545 ;
        RECT 101.110 187.360 103.640 187.500 ;
        RECT 101.110 187.300 101.430 187.360 ;
        RECT 60.170 187.160 60.490 187.220 ;
        RECT 62.025 187.160 62.315 187.205 ;
        RECT 60.170 187.020 62.315 187.160 ;
        RECT 60.170 186.960 60.490 187.020 ;
        RECT 62.025 186.975 62.315 187.020 ;
        RECT 72.590 186.960 72.910 187.220 ;
        RECT 78.660 187.160 78.800 187.300 ;
        RECT 82.220 187.160 82.510 187.205 ;
        RECT 84.090 187.160 84.410 187.220 ;
        RECT 78.660 187.020 80.180 187.160 ;
        RECT 57.885 186.635 58.175 186.865 ;
        RECT 58.805 186.635 59.095 186.865 ;
        RECT 52.825 186.480 53.115 186.525 ;
        RECT 57.960 186.480 58.100 186.635 ;
        RECT 59.250 186.620 59.570 186.880 ;
        RECT 59.710 186.620 60.030 186.880 ;
        RECT 61.550 186.620 61.870 186.880 ;
        RECT 62.945 186.635 63.235 186.865 ;
        RECT 69.370 186.820 69.690 186.880 ;
        RECT 71.225 186.820 71.515 186.865 ;
        RECT 69.370 186.680 71.515 186.820 ;
        RECT 61.090 186.480 61.410 186.540 ;
        RECT 51.980 186.340 56.260 186.480 ;
        RECT 57.960 186.340 61.410 186.480 ;
        RECT 32.125 186.295 32.415 186.340 ;
        RECT 21.990 186.140 22.280 186.185 ;
        RECT 23.560 186.140 23.850 186.185 ;
        RECT 25.660 186.140 25.950 186.185 ;
        RECT 21.990 186.000 25.950 186.140 ;
        RECT 21.990 185.955 22.280 186.000 ;
        RECT 23.560 185.955 23.850 186.000 ;
        RECT 25.660 185.955 25.950 186.000 ;
        RECT 29.365 186.140 29.655 186.185 ;
        RECT 31.740 186.140 31.880 186.295 ;
        RECT 32.570 186.140 32.890 186.200 ;
        RECT 34.870 186.140 35.190 186.200 ;
        RECT 35.420 186.185 35.560 186.340 ;
        RECT 39.930 186.280 40.250 186.340 ;
        RECT 43.150 186.280 43.470 186.340 ;
        RECT 46.370 186.280 46.690 186.340 ;
        RECT 52.825 186.295 53.115 186.340 ;
        RECT 56.120 186.200 56.260 186.340 ;
        RECT 61.090 186.280 61.410 186.340 ;
        RECT 29.365 186.000 35.190 186.140 ;
        RECT 29.365 185.955 29.655 186.000 ;
        RECT 32.570 185.940 32.890 186.000 ;
        RECT 34.870 185.940 35.190 186.000 ;
        RECT 35.345 185.955 35.635 186.185 ;
        RECT 36.265 186.140 36.555 186.185 ;
        RECT 40.850 186.140 41.170 186.200 ;
        RECT 36.265 186.000 41.170 186.140 ;
        RECT 36.265 185.955 36.555 186.000 ;
        RECT 40.850 185.940 41.170 186.000 ;
        RECT 56.030 185.940 56.350 186.200 ;
        RECT 57.870 186.140 58.190 186.200 ;
        RECT 63.020 186.140 63.160 186.635 ;
        RECT 69.370 186.620 69.690 186.680 ;
        RECT 71.225 186.635 71.515 186.680 ;
        RECT 71.685 186.820 71.975 186.865 ;
        RECT 73.510 186.820 73.830 186.880 ;
        RECT 80.040 186.865 80.180 187.020 ;
        RECT 82.220 187.020 84.410 187.160 ;
        RECT 82.220 186.975 82.510 187.020 ;
        RECT 84.090 186.960 84.410 187.020 ;
        RECT 99.285 187.160 99.575 187.205 ;
        RECT 102.490 187.160 102.810 187.220 ;
        RECT 99.285 187.020 102.810 187.160 ;
        RECT 103.500 187.160 103.640 187.360 ;
        RECT 103.870 187.360 104.635 187.500 ;
        RECT 103.870 187.300 104.190 187.360 ;
        RECT 104.345 187.315 104.635 187.360 ;
        RECT 105.250 187.300 105.570 187.560 ;
        RECT 120.890 187.300 121.210 187.560 ;
        RECT 123.205 187.500 123.495 187.545 ;
        RECT 125.965 187.500 126.255 187.545 ;
        RECT 127.330 187.500 127.650 187.560 ;
        RECT 123.205 187.360 127.650 187.500 ;
        RECT 123.205 187.315 123.495 187.360 ;
        RECT 125.965 187.315 126.255 187.360 ;
        RECT 127.330 187.300 127.650 187.360 ;
        RECT 108.900 187.160 109.190 187.205 ;
        RECT 110.310 187.160 110.630 187.220 ;
        RECT 103.500 187.020 105.020 187.160 ;
        RECT 99.285 186.975 99.575 187.020 ;
        RECT 102.490 186.960 102.810 187.020 ;
        RECT 71.685 186.680 73.830 186.820 ;
        RECT 71.685 186.635 71.975 186.680 ;
        RECT 73.510 186.620 73.830 186.680 ;
        RECT 78.685 186.820 78.975 186.865 ;
        RECT 79.965 186.820 80.255 186.865 ;
        RECT 80.885 186.820 81.175 186.865 ;
        RECT 78.685 186.680 79.720 186.820 ;
        RECT 78.685 186.635 78.975 186.680 ;
        RECT 75.375 186.480 75.665 186.525 ;
        RECT 77.895 186.480 78.185 186.525 ;
        RECT 79.085 186.480 79.375 186.525 ;
        RECT 75.375 186.340 79.375 186.480 ;
        RECT 79.580 186.480 79.720 186.680 ;
        RECT 79.965 186.680 81.175 186.820 ;
        RECT 79.965 186.635 80.255 186.680 ;
        RECT 80.885 186.635 81.175 186.680 ;
        RECT 97.905 186.820 98.195 186.865 ;
        RECT 98.350 186.820 98.670 186.880 ;
        RECT 97.905 186.680 98.670 186.820 ;
        RECT 97.905 186.635 98.195 186.680 ;
        RECT 98.350 186.620 98.670 186.680 ;
        RECT 98.810 186.620 99.130 186.880 ;
        RECT 99.745 186.820 100.035 186.865 ;
        RECT 101.570 186.820 101.890 186.880 ;
        RECT 99.745 186.680 101.890 186.820 ;
        RECT 99.745 186.635 100.035 186.680 ;
        RECT 101.570 186.620 101.890 186.680 ;
        RECT 102.030 186.620 102.350 186.880 ;
        RECT 104.880 186.865 105.020 187.020 ;
        RECT 108.900 187.020 110.630 187.160 ;
        RECT 108.900 186.975 109.190 187.020 ;
        RECT 110.310 186.960 110.630 187.020 ;
        RECT 123.650 187.160 123.970 187.220 ;
        RECT 123.650 187.020 133.080 187.160 ;
        RECT 123.650 186.960 123.970 187.020 ;
        RECT 102.965 186.810 103.255 186.865 ;
        RECT 103.500 186.810 104.560 186.820 ;
        RECT 102.965 186.680 104.560 186.810 ;
        RECT 102.965 186.670 103.640 186.680 ;
        RECT 102.965 186.635 103.255 186.670 ;
        RECT 81.765 186.480 82.055 186.525 ;
        RECT 82.955 186.480 83.245 186.525 ;
        RECT 85.475 186.480 85.765 186.525 ;
        RECT 79.580 186.340 81.100 186.480 ;
        RECT 75.375 186.295 75.665 186.340 ;
        RECT 77.895 186.295 78.185 186.340 ;
        RECT 79.085 186.295 79.375 186.340 ;
        RECT 67.070 186.140 67.390 186.200 ;
        RECT 57.870 186.000 63.160 186.140 ;
        RECT 63.480 186.000 67.390 186.140 ;
        RECT 57.870 185.940 58.190 186.000 ;
        RECT 26.130 185.800 26.450 185.860 ;
        RECT 26.605 185.800 26.895 185.845 ;
        RECT 26.130 185.660 26.895 185.800 ;
        RECT 26.130 185.600 26.450 185.660 ;
        RECT 26.605 185.615 26.895 185.660 ;
        RECT 27.510 185.800 27.830 185.860 ;
        RECT 29.825 185.800 30.115 185.845 ;
        RECT 27.510 185.660 30.115 185.800 ;
        RECT 27.510 185.600 27.830 185.660 ;
        RECT 29.825 185.615 30.115 185.660 ;
        RECT 31.190 185.800 31.510 185.860 ;
        RECT 33.505 185.800 33.795 185.845 ;
        RECT 37.170 185.800 37.490 185.860 ;
        RECT 31.190 185.660 37.490 185.800 ;
        RECT 31.190 185.600 31.510 185.660 ;
        RECT 33.505 185.615 33.795 185.660 ;
        RECT 37.170 185.600 37.490 185.660 ;
        RECT 38.565 185.800 38.855 185.845 ;
        RECT 40.390 185.800 40.710 185.860 ;
        RECT 38.565 185.660 40.710 185.800 ;
        RECT 38.565 185.615 38.855 185.660 ;
        RECT 40.390 185.600 40.710 185.660 ;
        RECT 41.785 185.800 42.075 185.845 ;
        RECT 42.690 185.800 43.010 185.860 ;
        RECT 41.785 185.660 43.010 185.800 ;
        RECT 41.785 185.615 42.075 185.660 ;
        RECT 42.690 185.600 43.010 185.660 ;
        RECT 50.510 185.800 50.830 185.860 ;
        RECT 52.365 185.800 52.655 185.845 ;
        RECT 50.510 185.660 52.655 185.800 ;
        RECT 50.510 185.600 50.830 185.660 ;
        RECT 52.365 185.615 52.655 185.660 ;
        RECT 56.965 185.800 57.255 185.845 ;
        RECT 63.480 185.800 63.620 186.000 ;
        RECT 67.070 185.940 67.390 186.000 ;
        RECT 75.810 186.140 76.100 186.185 ;
        RECT 77.380 186.140 77.670 186.185 ;
        RECT 79.480 186.140 79.770 186.185 ;
        RECT 75.810 186.000 79.770 186.140 ;
        RECT 75.810 185.955 76.100 186.000 ;
        RECT 77.380 185.955 77.670 186.000 ;
        RECT 79.480 185.955 79.770 186.000 ;
        RECT 56.965 185.660 63.620 185.800 ;
        RECT 56.965 185.615 57.255 185.660 ;
        RECT 63.850 185.600 64.170 185.860 ;
        RECT 69.830 185.800 70.150 185.860 ;
        RECT 73.065 185.800 73.355 185.845 ;
        RECT 69.830 185.660 73.355 185.800 ;
        RECT 80.960 185.800 81.100 186.340 ;
        RECT 81.765 186.340 85.765 186.480 ;
        RECT 81.765 186.295 82.055 186.340 ;
        RECT 82.955 186.295 83.245 186.340 ;
        RECT 85.475 186.295 85.765 186.340 ;
        RECT 100.650 186.480 100.970 186.540 ;
        RECT 102.505 186.480 102.795 186.525 ;
        RECT 103.425 186.480 103.715 186.525 ;
        RECT 100.650 186.340 102.795 186.480 ;
        RECT 100.650 186.280 100.970 186.340 ;
        RECT 102.505 186.295 102.795 186.340 ;
        RECT 103.040 186.340 103.715 186.480 ;
        RECT 104.420 186.480 104.560 186.680 ;
        RECT 104.805 186.635 105.095 186.865 ;
        RECT 107.565 186.820 107.855 186.865 ;
        RECT 108.010 186.820 108.330 186.880 ;
        RECT 107.565 186.680 108.330 186.820 ;
        RECT 107.565 186.635 107.855 186.680 ;
        RECT 108.010 186.620 108.330 186.680 ;
        RECT 122.745 186.820 123.035 186.865 ;
        RECT 125.490 186.820 125.810 186.880 ;
        RECT 122.745 186.680 125.810 186.820 ;
        RECT 122.745 186.635 123.035 186.680 ;
        RECT 125.490 186.620 125.810 186.680 ;
        RECT 131.585 186.820 131.875 186.865 ;
        RECT 132.390 186.820 132.710 186.880 ;
        RECT 132.940 186.865 133.080 187.020 ;
        RECT 131.585 186.680 132.710 186.820 ;
        RECT 131.585 186.635 131.875 186.680 ;
        RECT 132.390 186.620 132.710 186.680 ;
        RECT 132.865 186.635 133.155 186.865 ;
        RECT 134.230 186.620 134.550 186.880 ;
        RECT 106.630 186.480 106.950 186.540 ;
        RECT 104.420 186.340 106.950 186.480 ;
        RECT 81.370 186.140 81.660 186.185 ;
        RECT 83.470 186.140 83.760 186.185 ;
        RECT 85.040 186.140 85.330 186.185 ;
        RECT 81.370 186.000 85.330 186.140 ;
        RECT 81.370 185.955 81.660 186.000 ;
        RECT 83.470 185.955 83.760 186.000 ;
        RECT 85.040 185.955 85.330 186.000 ;
        RECT 82.250 185.800 82.570 185.860 ;
        RECT 80.960 185.660 82.570 185.800 ;
        RECT 103.040 185.800 103.180 186.340 ;
        RECT 103.425 186.295 103.715 186.340 ;
        RECT 106.630 186.280 106.950 186.340 ;
        RECT 108.445 186.480 108.735 186.525 ;
        RECT 109.635 186.480 109.925 186.525 ;
        RECT 112.155 186.480 112.445 186.525 ;
        RECT 108.445 186.340 112.445 186.480 ;
        RECT 108.445 186.295 108.735 186.340 ;
        RECT 109.635 186.295 109.925 186.340 ;
        RECT 112.155 186.295 112.445 186.340 ;
        RECT 120.890 186.480 121.210 186.540 ;
        RECT 123.665 186.480 123.955 186.525 ;
        RECT 120.890 186.340 123.955 186.480 ;
        RECT 120.890 186.280 121.210 186.340 ;
        RECT 123.665 186.295 123.955 186.340 ;
        RECT 128.275 186.480 128.565 186.525 ;
        RECT 130.795 186.480 131.085 186.525 ;
        RECT 131.985 186.480 132.275 186.525 ;
        RECT 128.275 186.340 132.275 186.480 ;
        RECT 128.275 186.295 128.565 186.340 ;
        RECT 130.795 186.295 131.085 186.340 ;
        RECT 131.985 186.295 132.275 186.340 ;
        RECT 108.050 186.140 108.340 186.185 ;
        RECT 110.150 186.140 110.440 186.185 ;
        RECT 111.720 186.140 112.010 186.185 ;
        RECT 108.050 186.000 112.010 186.140 ;
        RECT 108.050 185.955 108.340 186.000 ;
        RECT 110.150 185.955 110.440 186.000 ;
        RECT 111.720 185.955 112.010 186.000 ;
        RECT 128.710 186.140 129.000 186.185 ;
        RECT 130.280 186.140 130.570 186.185 ;
        RECT 132.380 186.140 132.670 186.185 ;
        RECT 128.710 186.000 132.670 186.140 ;
        RECT 128.710 185.955 129.000 186.000 ;
        RECT 130.280 185.955 130.570 186.000 ;
        RECT 132.380 185.955 132.670 186.000 ;
        RECT 132.850 186.140 133.170 186.200 ;
        RECT 133.325 186.140 133.615 186.185 ;
        RECT 132.850 186.000 133.615 186.140 ;
        RECT 132.850 185.940 133.170 186.000 ;
        RECT 133.325 185.955 133.615 186.000 ;
        RECT 114.465 185.800 114.755 185.845 ;
        RECT 117.210 185.800 117.530 185.860 ;
        RECT 103.040 185.660 117.530 185.800 ;
        RECT 69.830 185.600 70.150 185.660 ;
        RECT 73.065 185.615 73.355 185.660 ;
        RECT 82.250 185.600 82.570 185.660 ;
        RECT 114.465 185.615 114.755 185.660 ;
        RECT 117.210 185.600 117.530 185.660 ;
        RECT 17.320 184.980 147.040 185.460 ;
        RECT 22.910 184.580 23.230 184.840 ;
        RECT 23.845 184.595 24.135 184.825 ;
        RECT 23.920 184.440 24.060 184.595 ;
        RECT 27.050 184.580 27.370 184.840 ;
        RECT 35.330 184.780 35.650 184.840 ;
        RECT 39.010 184.780 39.330 184.840 ;
        RECT 35.330 184.640 39.330 184.780 ;
        RECT 35.330 184.580 35.650 184.640 ;
        RECT 39.010 184.580 39.330 184.640 ;
        RECT 59.265 184.780 59.555 184.825 ;
        RECT 61.550 184.780 61.870 184.840 ;
        RECT 96.510 184.780 96.830 184.840 ;
        RECT 99.730 184.780 100.050 184.840 ;
        RECT 59.265 184.640 61.870 184.780 ;
        RECT 59.265 184.595 59.555 184.640 ;
        RECT 61.550 184.580 61.870 184.640 ;
        RECT 95.220 184.640 100.050 184.780 ;
        RECT 43.150 184.440 43.470 184.500 ;
        RECT 23.920 184.300 29.120 184.440 ;
        RECT 26.130 184.100 26.450 184.160 ;
        RECT 28.980 184.145 29.120 184.300 ;
        RECT 41.860 184.300 43.470 184.440 ;
        RECT 28.905 184.100 29.195 184.145 ;
        RECT 39.025 184.100 39.315 184.145 ;
        RECT 41.860 184.100 42.000 184.300 ;
        RECT 43.150 184.240 43.470 184.300 ;
        RECT 45.910 184.440 46.230 184.500 ;
        RECT 50.970 184.440 51.290 184.500 ;
        RECT 45.910 184.300 51.290 184.440 ;
        RECT 45.910 184.240 46.230 184.300 ;
        RECT 50.970 184.240 51.290 184.300 ;
        RECT 52.350 184.440 52.670 184.500 ;
        RECT 52.825 184.440 53.115 184.485 ;
        RECT 55.570 184.440 55.890 184.500 ;
        RECT 69.830 184.440 70.150 184.500 ;
        RECT 52.350 184.300 58.560 184.440 ;
        RECT 52.350 184.240 52.670 184.300 ;
        RECT 52.825 184.255 53.115 184.300 ;
        RECT 55.570 184.240 55.890 184.300 ;
        RECT 43.625 184.100 43.915 184.145 ;
        RECT 26.130 183.960 28.660 184.100 ;
        RECT 26.130 183.900 26.450 183.960 ;
        RECT 27.510 183.760 27.830 183.820 ;
        RECT 28.520 183.805 28.660 183.960 ;
        RECT 28.905 183.960 29.305 184.100 ;
        RECT 39.025 183.960 41.540 184.100 ;
        RECT 41.860 183.960 43.915 184.100 ;
        RECT 28.905 183.915 29.195 183.960 ;
        RECT 39.025 183.915 39.315 183.960 ;
        RECT 24.380 183.620 27.830 183.760 ;
        RECT 23.765 183.420 24.055 183.465 ;
        RECT 24.380 183.420 24.520 183.620 ;
        RECT 27.510 183.560 27.830 183.620 ;
        RECT 28.445 183.575 28.735 183.805 ;
        RECT 35.790 183.760 36.110 183.820 ;
        RECT 35.790 183.620 38.320 183.760 ;
        RECT 35.790 183.560 36.110 183.620 ;
        RECT 23.765 183.280 24.520 183.420 ;
        RECT 24.750 183.420 25.070 183.480 ;
        RECT 27.985 183.420 28.275 183.465 ;
        RECT 32.110 183.420 32.430 183.480 ;
        RECT 24.750 183.280 32.430 183.420 ;
        RECT 23.765 183.235 24.055 183.280 ;
        RECT 24.750 183.220 25.070 183.280 ;
        RECT 27.985 183.235 28.275 183.280 ;
        RECT 32.110 183.220 32.430 183.280 ;
        RECT 37.170 183.420 37.490 183.480 ;
        RECT 37.645 183.420 37.935 183.465 ;
        RECT 37.170 183.280 37.935 183.420 ;
        RECT 38.180 183.420 38.320 183.620 ;
        RECT 38.550 183.560 38.870 183.820 ;
        RECT 39.470 183.805 39.790 183.820 ;
        RECT 39.470 183.760 39.800 183.805 ;
        RECT 39.470 183.620 40.160 183.760 ;
        RECT 39.470 183.575 39.800 183.620 ;
        RECT 39.470 183.560 39.790 183.575 ;
        RECT 39.025 183.420 39.315 183.465 ;
        RECT 38.180 183.280 39.315 183.420 ;
        RECT 40.020 183.420 40.160 183.620 ;
        RECT 40.390 183.560 40.710 183.820 ;
        RECT 41.400 183.805 41.540 183.960 ;
        RECT 43.625 183.915 43.915 183.960 ;
        RECT 45.005 184.100 45.295 184.145 ;
        RECT 50.065 184.100 50.355 184.145 ;
        RECT 57.410 184.100 57.730 184.160 ;
        RECT 45.005 183.960 50.355 184.100 ;
        RECT 45.005 183.915 45.295 183.960 ;
        RECT 50.065 183.915 50.355 183.960 ;
        RECT 51.060 183.960 57.730 184.100 ;
        RECT 41.325 183.575 41.615 183.805 ;
        RECT 42.230 183.760 42.550 183.820 ;
        RECT 42.705 183.760 42.995 183.805 ;
        RECT 42.230 183.620 42.995 183.760 ;
        RECT 42.230 183.560 42.550 183.620 ;
        RECT 42.705 183.575 42.995 183.620 ;
        RECT 46.370 183.560 46.690 183.820 ;
        RECT 51.060 183.805 51.200 183.960 ;
        RECT 57.410 183.900 57.730 183.960 ;
        RECT 50.985 183.575 51.275 183.805 ;
        RECT 40.850 183.420 41.170 183.480 ;
        RECT 45.910 183.420 46.230 183.480 ;
        RECT 40.020 183.280 46.230 183.420 ;
        RECT 37.170 183.220 37.490 183.280 ;
        RECT 37.645 183.235 37.935 183.280 ;
        RECT 39.025 183.235 39.315 183.280 ;
        RECT 40.850 183.220 41.170 183.280 ;
        RECT 45.910 183.220 46.230 183.280 ;
        RECT 25.670 183.080 25.990 183.140 ;
        RECT 26.145 183.080 26.435 183.125 ;
        RECT 25.670 182.940 26.435 183.080 ;
        RECT 25.670 182.880 25.990 182.940 ;
        RECT 26.145 182.895 26.435 182.940 ;
        RECT 26.985 183.080 27.275 183.125 ;
        RECT 30.730 183.080 31.050 183.140 ;
        RECT 26.985 182.940 31.050 183.080 ;
        RECT 26.985 182.895 27.275 182.940 ;
        RECT 30.730 182.880 31.050 182.940 ;
        RECT 41.310 182.880 41.630 183.140 ;
        RECT 41.770 182.880 42.090 183.140 ;
        RECT 44.990 183.080 45.310 183.140 ;
        RECT 51.060 183.080 51.200 183.575 ;
        RECT 56.490 183.560 56.810 183.820 ;
        RECT 56.950 183.760 57.270 183.820 ;
        RECT 58.420 183.805 58.560 184.300 ;
        RECT 59.800 184.300 70.150 184.440 ;
        RECT 57.885 183.760 58.175 183.805 ;
        RECT 56.950 183.620 58.175 183.760 ;
        RECT 56.950 183.560 57.270 183.620 ;
        RECT 57.885 183.575 58.175 183.620 ;
        RECT 58.345 183.575 58.635 183.805 ;
        RECT 54.650 183.420 54.970 183.480 ;
        RECT 57.425 183.420 57.715 183.465 ;
        RECT 54.650 183.280 57.715 183.420 ;
        RECT 57.960 183.420 58.100 183.575 ;
        RECT 59.800 183.420 59.940 184.300 ;
        RECT 69.830 184.240 70.150 184.300 ;
        RECT 73.510 184.240 73.830 184.500 ;
        RECT 75.365 184.440 75.655 184.485 ;
        RECT 81.790 184.440 82.110 184.500 ;
        RECT 75.365 184.300 82.110 184.440 ;
        RECT 75.365 184.255 75.655 184.300 ;
        RECT 81.790 184.240 82.110 184.300 ;
        RECT 62.930 184.100 63.250 184.160 ;
        RECT 60.720 183.960 63.250 184.100 ;
        RECT 60.170 183.760 60.490 183.820 ;
        RECT 60.720 183.805 60.860 183.960 ;
        RECT 62.930 183.900 63.250 183.960 ;
        RECT 73.065 184.100 73.355 184.145 ;
        RECT 73.600 184.100 73.740 184.240 ;
        RECT 73.065 183.960 73.740 184.100 ;
        RECT 77.665 184.100 77.955 184.145 ;
        RECT 81.330 184.100 81.650 184.160 ;
        RECT 95.220 184.145 95.360 184.640 ;
        RECT 96.510 184.580 96.830 184.640 ;
        RECT 99.730 184.580 100.050 184.640 ;
        RECT 101.570 184.780 101.890 184.840 ;
        RECT 102.045 184.780 102.335 184.825 ;
        RECT 101.570 184.640 102.335 184.780 ;
        RECT 101.570 184.580 101.890 184.640 ;
        RECT 102.045 184.595 102.335 184.640 ;
        RECT 102.950 184.780 103.270 184.840 ;
        RECT 114.910 184.780 115.230 184.840 ;
        RECT 102.950 184.640 115.230 184.780 ;
        RECT 102.950 184.580 103.270 184.640 ;
        RECT 114.910 184.580 115.230 184.640 ;
        RECT 118.130 184.580 118.450 184.840 ;
        RECT 125.030 184.780 125.350 184.840 ;
        RECT 125.505 184.780 125.795 184.825 ;
        RECT 125.030 184.640 125.795 184.780 ;
        RECT 125.030 184.580 125.350 184.640 ;
        RECT 125.505 184.595 125.795 184.640 ;
        RECT 131.930 184.580 132.250 184.840 ;
        RECT 132.390 184.780 132.710 184.840 ;
        RECT 133.785 184.780 134.075 184.825 ;
        RECT 132.390 184.640 134.075 184.780 ;
        RECT 132.390 184.580 132.710 184.640 ;
        RECT 133.785 184.595 134.075 184.640 ;
        RECT 95.630 184.440 95.920 184.485 ;
        RECT 97.730 184.440 98.020 184.485 ;
        RECT 99.300 184.440 99.590 184.485 ;
        RECT 95.630 184.300 99.590 184.440 ;
        RECT 95.630 184.255 95.920 184.300 ;
        RECT 97.730 184.255 98.020 184.300 ;
        RECT 99.300 184.255 99.590 184.300 ;
        RECT 108.510 184.440 108.800 184.485 ;
        RECT 110.610 184.440 110.900 184.485 ;
        RECT 112.180 184.440 112.470 184.485 ;
        RECT 108.510 184.300 112.470 184.440 ;
        RECT 108.510 184.255 108.800 184.300 ;
        RECT 110.610 184.255 110.900 184.300 ;
        RECT 112.180 184.255 112.470 184.300 ;
        RECT 77.665 183.960 81.650 184.100 ;
        RECT 73.065 183.915 73.355 183.960 ;
        RECT 77.665 183.915 77.955 183.960 ;
        RECT 81.330 183.900 81.650 183.960 ;
        RECT 95.145 183.915 95.435 184.145 ;
        RECT 96.025 184.100 96.315 184.145 ;
        RECT 97.215 184.100 97.505 184.145 ;
        RECT 99.735 184.100 100.025 184.145 ;
        RECT 96.025 183.960 100.025 184.100 ;
        RECT 96.025 183.915 96.315 183.960 ;
        RECT 97.215 183.915 97.505 183.960 ;
        RECT 99.735 183.915 100.025 183.960 ;
        RECT 103.410 184.100 103.730 184.160 ;
        RECT 105.265 184.100 105.555 184.145 ;
        RECT 107.550 184.100 107.870 184.160 ;
        RECT 103.410 183.960 107.870 184.100 ;
        RECT 103.410 183.900 103.730 183.960 ;
        RECT 105.265 183.915 105.555 183.960 ;
        RECT 107.550 183.900 107.870 183.960 ;
        RECT 108.010 183.900 108.330 184.160 ;
        RECT 108.905 184.100 109.195 184.145 ;
        RECT 110.095 184.100 110.385 184.145 ;
        RECT 112.615 184.100 112.905 184.145 ;
        RECT 108.905 183.960 112.905 184.100 ;
        RECT 108.905 183.915 109.195 183.960 ;
        RECT 110.095 183.915 110.385 183.960 ;
        RECT 112.615 183.915 112.905 183.960 ;
        RECT 120.890 183.900 121.210 184.160 ;
        RECT 127.330 183.900 127.650 184.160 ;
        RECT 132.020 184.100 132.160 184.580 ;
        RECT 132.390 184.100 132.710 184.160 ;
        RECT 132.020 183.960 136.760 184.100 ;
        RECT 132.390 183.900 132.710 183.960 ;
        RECT 60.645 183.760 60.935 183.805 ;
        RECT 60.170 183.620 60.935 183.760 ;
        RECT 60.170 183.560 60.490 183.620 ;
        RECT 60.645 183.575 60.935 183.620 ;
        RECT 61.565 183.760 61.855 183.805 ;
        RECT 62.010 183.760 62.330 183.820 ;
        RECT 61.565 183.620 62.330 183.760 ;
        RECT 61.565 183.575 61.855 183.620 ;
        RECT 62.010 183.560 62.330 183.620 ;
        RECT 69.830 183.760 70.150 183.820 ;
        RECT 71.210 183.760 71.530 183.820 ;
        RECT 73.525 183.760 73.815 183.805 ;
        RECT 69.830 183.620 73.815 183.760 ;
        RECT 69.830 183.560 70.150 183.620 ;
        RECT 71.210 183.560 71.530 183.620 ;
        RECT 73.525 183.575 73.815 183.620 ;
        RECT 94.210 183.760 94.530 183.820 ;
        RECT 95.590 183.760 95.910 183.820 ;
        RECT 94.210 183.620 95.910 183.760 ;
        RECT 94.210 183.560 94.530 183.620 ;
        RECT 95.590 183.560 95.910 183.620 ;
        RECT 118.590 183.760 118.910 183.820 ;
        RECT 122.285 183.760 122.575 183.805 ;
        RECT 118.590 183.620 122.575 183.760 ;
        RECT 118.590 183.560 118.910 183.620 ;
        RECT 122.285 183.575 122.575 183.620 ;
        RECT 131.010 183.560 131.330 183.820 ;
        RECT 133.770 183.760 134.090 183.820 ;
        RECT 136.620 183.805 136.760 183.960 ;
        RECT 134.705 183.760 134.995 183.805 ;
        RECT 133.770 183.620 134.995 183.760 ;
        RECT 133.770 183.560 134.090 183.620 ;
        RECT 134.705 183.575 134.995 183.620 ;
        RECT 136.545 183.575 136.835 183.805 ;
        RECT 57.960 183.280 59.940 183.420 ;
        RECT 80.870 183.420 81.190 183.480 ;
        RECT 81.345 183.420 81.635 183.465 ;
        RECT 86.850 183.420 87.170 183.480 ;
        RECT 80.870 183.280 87.170 183.420 ;
        RECT 54.650 183.220 54.970 183.280 ;
        RECT 57.425 183.235 57.715 183.280 ;
        RECT 80.870 183.220 81.190 183.280 ;
        RECT 81.345 183.235 81.635 183.280 ;
        RECT 86.850 183.220 87.170 183.280 ;
        RECT 96.480 183.420 96.770 183.465 ;
        RECT 104.345 183.420 104.635 183.465 ;
        RECT 108.470 183.420 108.790 183.480 ;
        RECT 109.250 183.420 109.540 183.465 ;
        RECT 96.480 183.280 102.720 183.420 ;
        RECT 96.480 183.235 96.770 183.280 ;
        RECT 44.990 182.940 51.200 183.080 ;
        RECT 54.190 183.080 54.510 183.140 ;
        RECT 59.250 183.080 59.570 183.140 ;
        RECT 59.725 183.080 60.015 183.125 ;
        RECT 54.190 182.940 60.015 183.080 ;
        RECT 44.990 182.880 45.310 182.940 ;
        RECT 54.190 182.880 54.510 182.940 ;
        RECT 59.250 182.880 59.570 182.940 ;
        RECT 59.725 182.895 60.015 182.940 ;
        RECT 61.550 183.080 61.870 183.140 ;
        RECT 66.150 183.080 66.470 183.140 ;
        RECT 61.550 182.940 66.470 183.080 ;
        RECT 61.550 182.880 61.870 182.940 ;
        RECT 66.150 182.880 66.470 182.940 ;
        RECT 90.990 183.080 91.310 183.140 ;
        RECT 102.580 183.125 102.720 183.280 ;
        RECT 104.345 183.280 108.240 183.420 ;
        RECT 104.345 183.235 104.635 183.280 ;
        RECT 91.465 183.080 91.755 183.125 ;
        RECT 90.990 182.940 91.755 183.080 ;
        RECT 90.990 182.880 91.310 182.940 ;
        RECT 91.465 182.895 91.755 182.940 ;
        RECT 102.505 182.895 102.795 183.125 ;
        RECT 104.805 183.080 105.095 183.125 ;
        RECT 106.630 183.080 106.950 183.140 ;
        RECT 104.805 182.940 106.950 183.080 ;
        RECT 108.100 183.080 108.240 183.280 ;
        RECT 108.470 183.280 109.540 183.420 ;
        RECT 108.470 183.220 108.790 183.280 ;
        RECT 109.250 183.235 109.540 183.280 ;
        RECT 130.565 183.420 130.855 183.465 ;
        RECT 135.165 183.420 135.455 183.465 ;
        RECT 130.565 183.280 135.455 183.420 ;
        RECT 130.565 183.235 130.855 183.280 ;
        RECT 135.165 183.235 135.455 183.280 ;
        RECT 135.625 183.235 135.915 183.465 ;
        RECT 116.290 183.080 116.610 183.140 ;
        RECT 108.100 182.940 116.610 183.080 ;
        RECT 104.805 182.895 105.095 182.940 ;
        RECT 106.630 182.880 106.950 182.940 ;
        RECT 116.290 182.880 116.610 182.940 ;
        RECT 119.970 182.880 120.290 183.140 ;
        RECT 120.445 183.080 120.735 183.125 ;
        RECT 127.790 183.080 128.110 183.140 ;
        RECT 120.445 182.940 128.110 183.080 ;
        RECT 120.445 182.895 120.735 182.940 ;
        RECT 127.790 182.880 128.110 182.940 ;
        RECT 130.090 183.080 130.410 183.140 ;
        RECT 135.700 183.080 135.840 183.235 ;
        RECT 130.090 182.940 135.840 183.080 ;
        RECT 130.090 182.880 130.410 182.940 ;
        RECT 17.320 182.260 147.040 182.740 ;
        RECT 35.330 182.060 35.650 182.120 ;
        RECT 36.250 182.060 36.570 182.120 ;
        RECT 35.330 181.920 36.570 182.060 ;
        RECT 35.330 181.860 35.650 181.920 ;
        RECT 36.250 181.860 36.570 181.920 ;
        RECT 44.070 182.060 44.390 182.120 ;
        RECT 65.230 182.060 65.550 182.120 ;
        RECT 44.070 181.920 65.550 182.060 ;
        RECT 44.070 181.860 44.390 181.920 ;
        RECT 65.230 181.860 65.550 181.920 ;
        RECT 66.165 182.060 66.455 182.105 ;
        RECT 71.670 182.060 71.990 182.120 ;
        RECT 66.165 181.920 71.990 182.060 ;
        RECT 66.165 181.875 66.455 181.920 ;
        RECT 71.670 181.860 71.990 181.920 ;
        RECT 72.130 182.105 72.450 182.120 ;
        RECT 72.130 182.060 72.565 182.105 ;
        RECT 73.510 182.060 73.830 182.120 ;
        RECT 81.790 182.060 82.110 182.120 ;
        RECT 72.130 181.920 73.830 182.060 ;
        RECT 72.130 181.875 72.565 181.920 ;
        RECT 72.130 181.860 72.450 181.875 ;
        RECT 73.510 181.860 73.830 181.920 ;
        RECT 80.960 181.920 82.110 182.060 ;
        RECT 35.790 181.720 36.110 181.780 ;
        RECT 38.565 181.720 38.855 181.765 ;
        RECT 41.770 181.720 42.090 181.780 ;
        RECT 35.790 181.580 37.400 181.720 ;
        RECT 35.790 181.520 36.110 181.580 ;
        RECT 24.765 181.195 25.055 181.425 ;
        RECT 25.670 181.380 25.990 181.440 ;
        RECT 35.330 181.380 35.650 181.440 ;
        RECT 37.260 181.425 37.400 181.580 ;
        RECT 38.565 181.580 39.240 181.720 ;
        RECT 38.565 181.535 38.855 181.580 ;
        RECT 39.100 181.425 39.240 181.580 ;
        RECT 40.480 181.580 42.090 181.720 ;
        RECT 36.265 181.380 36.555 181.425 ;
        RECT 25.670 181.240 35.650 181.380 ;
        RECT 24.840 181.040 24.980 181.195 ;
        RECT 25.670 181.180 25.990 181.240 ;
        RECT 35.330 181.180 35.650 181.240 ;
        RECT 35.880 181.240 36.555 181.380 ;
        RECT 35.880 181.100 36.020 181.240 ;
        RECT 36.265 181.195 36.555 181.240 ;
        RECT 36.725 181.195 37.015 181.425 ;
        RECT 37.185 181.195 37.475 181.425 ;
        RECT 39.025 181.195 39.315 181.425 ;
        RECT 26.130 181.040 26.450 181.100 ;
        RECT 24.840 180.900 26.450 181.040 ;
        RECT 26.130 180.840 26.450 180.900 ;
        RECT 35.790 180.840 36.110 181.100 ;
        RECT 36.800 181.040 36.940 181.195 ;
        RECT 39.930 181.180 40.250 181.440 ;
        RECT 40.480 181.425 40.620 181.580 ;
        RECT 41.770 181.520 42.090 181.580 ;
        RECT 56.965 181.720 57.255 181.765 ;
        RECT 59.725 181.720 60.015 181.765 ;
        RECT 60.170 181.720 60.490 181.780 ;
        RECT 63.850 181.720 64.170 181.780 ;
        RECT 64.325 181.720 64.615 181.765 ;
        RECT 56.965 181.580 60.490 181.720 ;
        RECT 56.965 181.535 57.255 181.580 ;
        RECT 59.725 181.535 60.015 181.580 ;
        RECT 60.170 181.520 60.490 181.580 ;
        RECT 61.180 181.580 63.160 181.720 ;
        RECT 40.405 181.195 40.695 181.425 ;
        RECT 40.865 181.380 41.155 181.425 ;
        RECT 41.310 181.380 41.630 181.440 ;
        RECT 42.690 181.380 43.010 181.440 ;
        RECT 40.865 181.240 43.010 181.380 ;
        RECT 40.865 181.195 41.155 181.240 ;
        RECT 41.310 181.180 41.630 181.240 ;
        RECT 42.690 181.180 43.010 181.240 ;
        RECT 43.625 181.380 43.915 181.425 ;
        RECT 47.750 181.380 48.070 181.440 ;
        RECT 43.625 181.240 48.070 181.380 ;
        RECT 43.625 181.195 43.915 181.240 ;
        RECT 47.750 181.180 48.070 181.240 ;
        RECT 50.985 181.380 51.275 181.425 ;
        RECT 52.810 181.380 53.130 181.440 ;
        RECT 50.985 181.240 53.130 181.380 ;
        RECT 50.985 181.195 51.275 181.240 ;
        RECT 52.810 181.180 53.130 181.240 ;
        RECT 54.205 181.380 54.495 181.425 ;
        RECT 55.570 181.380 55.890 181.440 ;
        RECT 54.205 181.240 55.890 181.380 ;
        RECT 54.205 181.195 54.495 181.240 ;
        RECT 39.470 181.040 39.790 181.100 ;
        RECT 36.800 180.900 39.790 181.040 ;
        RECT 39.470 180.840 39.790 180.900 ;
        RECT 47.305 181.040 47.595 181.085 ;
        RECT 54.280 181.040 54.420 181.195 ;
        RECT 55.570 181.180 55.890 181.240 ;
        RECT 56.505 181.380 56.795 181.425 ;
        RECT 57.410 181.380 57.730 181.440 ;
        RECT 56.505 181.240 57.730 181.380 ;
        RECT 56.505 181.195 56.795 181.240 ;
        RECT 57.410 181.180 57.730 181.240 ;
        RECT 58.805 181.195 59.095 181.425 ;
        RECT 47.305 180.900 54.420 181.040 ;
        RECT 47.305 180.855 47.595 180.900 ;
        RECT 34.870 180.700 35.190 180.760 ;
        RECT 36.710 180.700 37.030 180.760 ;
        RECT 34.870 180.560 37.030 180.700 ;
        RECT 34.870 180.500 35.190 180.560 ;
        RECT 36.710 180.500 37.030 180.560 ;
        RECT 46.370 180.700 46.690 180.760 ;
        RECT 58.880 180.700 59.020 181.195 ;
        RECT 60.630 181.180 60.950 181.440 ;
        RECT 59.710 181.040 60.030 181.100 ;
        RECT 61.180 181.085 61.320 181.580 ;
        RECT 62.010 181.180 62.330 181.440 ;
        RECT 61.105 181.040 61.395 181.085 ;
        RECT 59.710 180.900 61.395 181.040 ;
        RECT 59.710 180.840 60.030 180.900 ;
        RECT 61.105 180.855 61.395 180.900 ;
        RECT 62.100 180.700 62.240 181.180 ;
        RECT 46.370 180.560 62.240 180.700 ;
        RECT 63.020 180.700 63.160 181.580 ;
        RECT 63.850 181.580 64.615 181.720 ;
        RECT 63.850 181.520 64.170 181.580 ;
        RECT 64.325 181.535 64.615 181.580 ;
        RECT 64.785 181.720 65.075 181.765 ;
        RECT 65.690 181.720 66.010 181.780 ;
        RECT 67.545 181.720 67.835 181.765 ;
        RECT 64.785 181.580 67.835 181.720 ;
        RECT 64.785 181.535 65.075 181.580 ;
        RECT 65.690 181.520 66.010 181.580 ;
        RECT 67.545 181.535 67.835 181.580 ;
        RECT 69.845 181.720 70.135 181.765 ;
        RECT 71.225 181.720 71.515 181.765 ;
        RECT 69.845 181.580 70.520 181.720 ;
        RECT 69.845 181.535 70.135 181.580 ;
        RECT 70.380 181.440 70.520 181.580 ;
        RECT 71.225 181.580 74.200 181.720 ;
        RECT 71.225 181.535 71.515 181.580 ;
        RECT 63.390 181.180 63.710 181.440 ;
        RECT 65.230 181.180 65.550 181.440 ;
        RECT 66.610 181.180 66.930 181.440 ;
        RECT 69.385 181.370 69.675 181.425 ;
        RECT 69.385 181.230 70.060 181.370 ;
        RECT 69.385 181.195 69.675 181.230 ;
        RECT 66.150 181.040 66.470 181.100 ;
        RECT 68.465 181.040 68.755 181.085 ;
        RECT 66.150 180.900 68.755 181.040 ;
        RECT 69.920 181.040 70.060 181.230 ;
        RECT 70.290 181.180 70.610 181.440 ;
        RECT 70.765 181.380 71.055 181.425 ;
        RECT 73.525 181.380 73.815 181.425 ;
        RECT 70.765 181.240 73.815 181.380 ;
        RECT 70.765 181.195 71.055 181.240 ;
        RECT 73.525 181.195 73.815 181.240 ;
        RECT 74.060 181.100 74.200 181.580 ;
        RECT 80.960 181.425 81.100 181.920 ;
        RECT 81.790 181.860 82.110 181.920 ;
        RECT 90.990 181.860 91.310 182.120 ;
        RECT 94.670 182.060 94.990 182.120 ;
        RECT 95.605 182.060 95.895 182.105 ;
        RECT 94.670 181.920 95.895 182.060 ;
        RECT 94.670 181.860 94.990 181.920 ;
        RECT 95.605 181.875 95.895 181.920 ;
        RECT 106.630 181.860 106.950 182.120 ;
        RECT 108.470 181.860 108.790 182.120 ;
        RECT 110.325 182.060 110.615 182.105 ;
        RECT 111.690 182.060 112.010 182.120 ;
        RECT 110.325 181.920 112.010 182.060 ;
        RECT 110.325 181.875 110.615 181.920 ;
        RECT 111.690 181.860 112.010 181.920 ;
        RECT 116.290 181.860 116.610 182.120 ;
        RECT 118.590 181.860 118.910 182.120 ;
        RECT 127.790 181.860 128.110 182.120 ;
        RECT 133.770 181.860 134.090 182.120 ;
        RECT 134.230 181.860 134.550 182.120 ;
        RECT 81.345 181.720 81.635 181.765 ;
        RECT 82.250 181.720 82.570 181.780 ;
        RECT 81.345 181.580 82.570 181.720 ;
        RECT 81.345 181.535 81.635 181.580 ;
        RECT 82.250 181.520 82.570 181.580 ;
        RECT 108.010 181.720 108.330 181.780 ;
        RECT 123.650 181.720 123.970 181.780 ;
        RECT 108.010 181.580 123.970 181.720 ;
        RECT 108.010 181.520 108.330 181.580 ;
        RECT 79.965 181.195 80.255 181.425 ;
        RECT 80.885 181.195 81.175 181.425 ;
        RECT 81.805 181.195 82.095 181.425 ;
        RECT 90.545 181.380 90.835 181.425 ;
        RECT 96.510 181.380 96.830 181.440 ;
        RECT 90.545 181.240 96.830 181.380 ;
        RECT 90.545 181.195 90.835 181.240 ;
        RECT 72.130 181.040 72.450 181.100 ;
        RECT 73.970 181.040 74.290 181.100 ;
        RECT 76.285 181.040 76.575 181.085 ;
        RECT 69.920 180.900 72.450 181.040 ;
        RECT 66.150 180.840 66.470 180.900 ;
        RECT 68.465 180.855 68.755 180.900 ;
        RECT 72.130 180.840 72.450 180.900 ;
        RECT 73.140 180.900 76.575 181.040 ;
        RECT 80.040 181.040 80.180 181.195 ;
        RECT 81.330 181.040 81.650 181.100 ;
        RECT 80.040 180.900 81.650 181.040 ;
        RECT 73.140 180.700 73.280 180.900 ;
        RECT 73.970 180.840 74.290 180.900 ;
        RECT 76.285 180.855 76.575 180.900 ;
        RECT 81.330 180.840 81.650 180.900 ;
        RECT 63.020 180.560 73.280 180.700 ;
        RECT 73.510 180.700 73.830 180.760 ;
        RECT 81.880 180.700 82.020 181.195 ;
        RECT 96.510 181.180 96.830 181.240 ;
        RECT 96.970 181.380 97.290 181.440 ;
        RECT 97.445 181.380 97.735 181.425 ;
        RECT 99.745 181.380 100.035 181.425 ;
        RECT 96.970 181.240 97.735 181.380 ;
        RECT 96.970 181.180 97.290 181.240 ;
        RECT 97.445 181.195 97.735 181.240 ;
        RECT 97.980 181.240 100.035 181.380 ;
        RECT 97.980 181.100 98.120 181.240 ;
        RECT 99.745 181.195 100.035 181.240 ;
        RECT 102.030 181.380 102.350 181.440 ;
        RECT 103.425 181.380 103.715 181.425 ;
        RECT 102.030 181.240 103.715 181.380 ;
        RECT 102.030 181.180 102.350 181.240 ;
        RECT 103.425 181.195 103.715 181.240 ;
        RECT 110.785 181.380 111.075 181.425 ;
        RECT 112.625 181.380 112.915 181.425 ;
        RECT 110.785 181.240 112.915 181.380 ;
        RECT 110.785 181.195 111.075 181.240 ;
        RECT 112.625 181.195 112.915 181.240 ;
        RECT 114.910 181.380 115.230 181.440 ;
        RECT 115.385 181.380 115.675 181.425 ;
        RECT 114.910 181.240 115.675 181.380 ;
        RECT 114.910 181.180 115.230 181.240 ;
        RECT 115.385 181.195 115.675 181.240 ;
        RECT 117.210 181.380 117.530 181.440 ;
        RECT 120.980 181.425 121.120 181.580 ;
        RECT 123.650 181.520 123.970 181.580 ;
        RECT 118.145 181.380 118.435 181.425 ;
        RECT 117.210 181.240 118.435 181.380 ;
        RECT 117.210 181.180 117.530 181.240 ;
        RECT 118.145 181.195 118.435 181.240 ;
        RECT 120.905 181.195 121.195 181.425 ;
        RECT 122.240 181.380 122.530 181.425 ;
        RECT 124.110 181.380 124.430 181.440 ;
        RECT 122.240 181.240 124.430 181.380 ;
        RECT 127.880 181.380 128.020 181.860 ;
        RECT 128.710 181.720 129.030 181.780 ;
        RECT 132.865 181.720 133.155 181.765 ;
        RECT 128.710 181.580 133.155 181.720 ;
        RECT 128.710 181.520 129.030 181.580 ;
        RECT 132.865 181.535 133.155 181.580 ;
        RECT 131.025 181.380 131.315 181.425 ;
        RECT 127.880 181.240 131.315 181.380 ;
        RECT 122.240 181.195 122.530 181.240 ;
        RECT 124.110 181.180 124.430 181.240 ;
        RECT 131.025 181.195 131.315 181.240 ;
        RECT 131.930 181.180 132.250 181.440 ;
        RECT 139.865 181.380 140.155 181.425 ;
        RECT 140.670 181.380 140.990 181.440 ;
        RECT 139.865 181.240 140.990 181.380 ;
        RECT 139.865 181.195 140.155 181.240 ;
        RECT 140.670 181.180 140.990 181.240 ;
        RECT 91.925 180.855 92.215 181.085 ;
        RECT 73.510 180.560 82.020 180.700 ;
        RECT 92.000 180.700 92.140 180.855 ;
        RECT 97.890 180.840 98.210 181.100 ;
        RECT 98.825 181.040 99.115 181.085 ;
        RECT 100.190 181.040 100.510 181.100 ;
        RECT 98.825 180.900 100.510 181.040 ;
        RECT 98.825 180.855 99.115 180.900 ;
        RECT 100.190 180.840 100.510 180.900 ;
        RECT 107.550 181.040 107.870 181.100 ;
        RECT 111.245 181.040 111.535 181.085 ;
        RECT 107.550 180.900 111.535 181.040 ;
        RECT 107.550 180.840 107.870 180.900 ;
        RECT 111.245 180.855 111.535 180.900 ;
        RECT 119.525 180.855 119.815 181.085 ;
        RECT 121.785 181.040 122.075 181.085 ;
        RECT 122.975 181.040 123.265 181.085 ;
        RECT 125.495 181.040 125.785 181.085 ;
        RECT 121.785 180.900 125.785 181.040 ;
        RECT 121.785 180.855 122.075 180.900 ;
        RECT 122.975 180.855 123.265 180.900 ;
        RECT 125.495 180.855 125.785 180.900 ;
        RECT 136.555 181.040 136.845 181.085 ;
        RECT 139.075 181.040 139.365 181.085 ;
        RECT 140.265 181.040 140.555 181.085 ;
        RECT 136.555 180.900 140.555 181.040 ;
        RECT 136.555 180.855 136.845 180.900 ;
        RECT 139.075 180.855 139.365 180.900 ;
        RECT 140.265 180.855 140.555 180.900 ;
        RECT 141.145 180.855 141.435 181.085 ;
        RECT 103.410 180.700 103.730 180.760 ;
        RECT 92.000 180.560 103.730 180.700 ;
        RECT 46.370 180.500 46.690 180.560 ;
        RECT 73.510 180.500 73.830 180.560 ;
        RECT 103.410 180.500 103.730 180.560 ;
        RECT 116.290 180.700 116.610 180.760 ;
        RECT 119.600 180.700 119.740 180.855 ;
        RECT 120.890 180.700 121.210 180.760 ;
        RECT 116.290 180.560 121.210 180.700 ;
        RECT 116.290 180.500 116.610 180.560 ;
        RECT 120.890 180.500 121.210 180.560 ;
        RECT 121.390 180.700 121.680 180.745 ;
        RECT 123.490 180.700 123.780 180.745 ;
        RECT 125.060 180.700 125.350 180.745 ;
        RECT 121.390 180.560 125.350 180.700 ;
        RECT 121.390 180.515 121.680 180.560 ;
        RECT 123.490 180.515 123.780 180.560 ;
        RECT 125.060 180.515 125.350 180.560 ;
        RECT 136.990 180.700 137.280 180.745 ;
        RECT 138.560 180.700 138.850 180.745 ;
        RECT 140.660 180.700 140.950 180.745 ;
        RECT 136.990 180.560 140.950 180.700 ;
        RECT 136.990 180.515 137.280 180.560 ;
        RECT 138.560 180.515 138.850 180.560 ;
        RECT 140.660 180.515 140.950 180.560 ;
        RECT 25.225 180.360 25.515 180.405 ;
        RECT 29.350 180.360 29.670 180.420 ;
        RECT 25.225 180.220 29.670 180.360 ;
        RECT 25.225 180.175 25.515 180.220 ;
        RECT 29.350 180.160 29.670 180.220 ;
        RECT 39.470 180.360 39.790 180.420 ;
        RECT 42.245 180.360 42.535 180.405 ;
        RECT 39.470 180.220 42.535 180.360 ;
        RECT 39.470 180.160 39.790 180.220 ;
        RECT 42.245 180.175 42.535 180.220 ;
        RECT 58.330 180.160 58.650 180.420 ;
        RECT 60.170 180.360 60.490 180.420 ;
        RECT 60.645 180.360 60.935 180.405 ;
        RECT 60.170 180.220 60.935 180.360 ;
        RECT 60.170 180.160 60.490 180.220 ;
        RECT 60.645 180.175 60.935 180.220 ;
        RECT 62.470 180.360 62.790 180.420 ;
        RECT 62.945 180.360 63.235 180.405 ;
        RECT 62.470 180.220 63.235 180.360 ;
        RECT 62.470 180.160 62.790 180.220 ;
        RECT 62.945 180.175 63.235 180.220 ;
        RECT 70.750 180.160 71.070 180.420 ;
        RECT 71.210 180.360 71.530 180.420 ;
        RECT 72.145 180.360 72.435 180.405 ;
        RECT 71.210 180.220 72.435 180.360 ;
        RECT 71.210 180.160 71.530 180.220 ;
        RECT 72.145 180.175 72.435 180.220 ;
        RECT 72.590 180.360 72.910 180.420 ;
        RECT 73.065 180.360 73.355 180.405 ;
        RECT 72.590 180.220 73.355 180.360 ;
        RECT 72.590 180.160 72.910 180.220 ;
        RECT 73.065 180.175 73.355 180.220 ;
        RECT 85.930 180.360 86.250 180.420 ;
        RECT 88.705 180.360 88.995 180.405 ;
        RECT 85.930 180.220 88.995 180.360 ;
        RECT 85.930 180.160 86.250 180.220 ;
        RECT 88.705 180.175 88.995 180.220 ;
        RECT 102.490 180.360 102.810 180.420 ;
        RECT 102.965 180.360 103.255 180.405 ;
        RECT 102.490 180.220 103.255 180.360 ;
        RECT 102.490 180.160 102.810 180.220 ;
        RECT 102.965 180.175 103.255 180.220 ;
        RECT 128.250 180.160 128.570 180.420 ;
        RECT 137.450 180.360 137.770 180.420 ;
        RECT 141.220 180.360 141.360 180.855 ;
        RECT 137.450 180.220 141.360 180.360 ;
        RECT 137.450 180.160 137.770 180.220 ;
        RECT 17.320 179.540 147.040 180.020 ;
        RECT 23.385 179.340 23.675 179.385 ;
        RECT 32.110 179.340 32.430 179.400 ;
        RECT 23.385 179.200 32.430 179.340 ;
        RECT 23.385 179.155 23.675 179.200 ;
        RECT 32.110 179.140 32.430 179.200 ;
        RECT 41.785 179.340 42.075 179.385 ;
        RECT 42.230 179.340 42.550 179.400 ;
        RECT 80.870 179.340 81.190 179.400 ;
        RECT 41.785 179.200 42.550 179.340 ;
        RECT 41.785 179.155 42.075 179.200 ;
        RECT 42.230 179.140 42.550 179.200 ;
        RECT 55.200 179.200 81.190 179.340 ;
        RECT 24.750 179.000 25.070 179.060 ;
        RECT 27.970 179.000 28.290 179.060 ;
        RECT 31.190 179.000 31.510 179.060 ;
        RECT 54.190 179.000 54.510 179.060 ;
        RECT 24.750 178.860 31.510 179.000 ;
        RECT 24.750 178.800 25.070 178.860 ;
        RECT 27.970 178.800 28.290 178.860 ;
        RECT 31.190 178.800 31.510 178.860 ;
        RECT 43.240 178.860 54.510 179.000 ;
        RECT 24.840 178.660 24.980 178.800 ;
        RECT 24.380 178.520 24.980 178.660 ;
        RECT 26.605 178.660 26.895 178.705 ;
        RECT 30.270 178.660 30.590 178.720 ;
        RECT 43.240 178.660 43.380 178.860 ;
        RECT 54.190 178.800 54.510 178.860 ;
        RECT 26.605 178.520 30.590 178.660 ;
        RECT 24.380 178.025 24.520 178.520 ;
        RECT 26.605 178.475 26.895 178.520 ;
        RECT 30.270 178.460 30.590 178.520 ;
        RECT 36.340 178.520 43.380 178.660 ;
        RECT 43.610 178.660 43.930 178.720 ;
        RECT 44.085 178.660 44.375 178.705 ;
        RECT 52.810 178.660 53.130 178.720 ;
        RECT 43.610 178.520 53.130 178.660 ;
        RECT 24.765 178.320 25.055 178.365 ;
        RECT 26.130 178.320 26.450 178.380 ;
        RECT 24.765 178.180 26.450 178.320 ;
        RECT 24.765 178.135 25.055 178.180 ;
        RECT 26.130 178.120 26.450 178.180 ;
        RECT 27.050 178.120 27.370 178.380 ;
        RECT 27.525 178.320 27.815 178.365 ;
        RECT 28.445 178.320 28.735 178.365 ;
        RECT 27.525 178.180 28.735 178.320 ;
        RECT 27.525 178.135 27.815 178.180 ;
        RECT 28.445 178.135 28.735 178.180 ;
        RECT 24.305 177.795 24.595 178.025 ;
        RECT 25.670 177.780 25.990 178.040 ;
        RECT 28.520 177.980 28.660 178.135 ;
        RECT 29.350 178.120 29.670 178.380 ;
        RECT 34.885 178.320 35.175 178.365 ;
        RECT 35.330 178.320 35.650 178.380 ;
        RECT 34.885 178.180 35.650 178.320 ;
        RECT 34.885 178.135 35.175 178.180 ;
        RECT 35.330 178.120 35.650 178.180 ;
        RECT 35.790 178.120 36.110 178.380 ;
        RECT 36.340 178.365 36.480 178.520 ;
        RECT 43.610 178.460 43.930 178.520 ;
        RECT 44.085 178.475 44.375 178.520 ;
        RECT 52.810 178.460 53.130 178.520 ;
        RECT 36.265 178.135 36.555 178.365 ;
        RECT 36.710 178.120 37.030 178.380 ;
        RECT 37.630 178.320 37.950 178.380 ;
        RECT 38.550 178.320 38.870 178.380 ;
        RECT 37.630 178.180 38.870 178.320 ;
        RECT 37.630 178.120 37.950 178.180 ;
        RECT 38.550 178.120 38.870 178.180 ;
        RECT 39.485 178.135 39.775 178.365 ;
        RECT 35.880 177.980 36.020 178.120 ;
        RECT 39.025 177.980 39.315 178.025 ;
        RECT 28.520 177.840 35.560 177.980 ;
        RECT 35.880 177.840 39.315 177.980 ;
        RECT 39.560 177.980 39.700 178.135 ;
        RECT 39.930 178.120 40.250 178.380 ;
        RECT 41.785 178.320 42.075 178.365 ;
        RECT 44.530 178.320 44.850 178.380 ;
        RECT 41.785 178.180 44.850 178.320 ;
        RECT 41.785 178.135 42.075 178.180 ;
        RECT 44.530 178.120 44.850 178.180 ;
        RECT 47.750 178.320 48.070 178.380 ;
        RECT 55.200 178.320 55.340 179.200 ;
        RECT 80.870 179.140 81.190 179.200 ;
        RECT 92.845 179.340 93.135 179.385 ;
        RECT 97.890 179.340 98.210 179.400 ;
        RECT 92.845 179.200 98.210 179.340 ;
        RECT 92.845 179.155 93.135 179.200 ;
        RECT 97.890 179.140 98.210 179.200 ;
        RECT 116.765 179.340 117.055 179.385 ;
        RECT 118.590 179.340 118.910 179.400 ;
        RECT 116.765 179.200 118.910 179.340 ;
        RECT 116.765 179.155 117.055 179.200 ;
        RECT 118.590 179.140 118.910 179.200 ;
        RECT 124.110 179.140 124.430 179.400 ;
        RECT 126.870 179.340 127.190 179.400 ;
        RECT 127.345 179.340 127.635 179.385 ;
        RECT 126.870 179.200 127.635 179.340 ;
        RECT 126.870 179.140 127.190 179.200 ;
        RECT 127.345 179.155 127.635 179.200 ;
        RECT 129.185 179.340 129.475 179.385 ;
        RECT 132.850 179.340 133.170 179.400 ;
        RECT 129.185 179.200 133.170 179.340 ;
        RECT 129.185 179.155 129.475 179.200 ;
        RECT 57.870 178.800 58.190 179.060 ;
        RECT 62.930 178.800 63.250 179.060 ;
        RECT 63.390 179.000 63.710 179.060 ;
        RECT 64.785 179.000 65.075 179.045 ;
        RECT 63.390 178.860 65.075 179.000 ;
        RECT 63.390 178.800 63.710 178.860 ;
        RECT 64.785 178.815 65.075 178.860 ;
        RECT 72.145 179.000 72.435 179.045 ;
        RECT 76.730 179.000 77.020 179.045 ;
        RECT 78.300 179.000 78.590 179.045 ;
        RECT 80.400 179.000 80.690 179.045 ;
        RECT 72.145 178.860 76.040 179.000 ;
        RECT 72.145 178.815 72.435 178.860 ;
        RECT 58.345 178.660 58.635 178.705 ;
        RECT 61.105 178.660 61.395 178.705 ;
        RECT 57.040 178.520 58.100 178.660 ;
        RECT 57.040 178.365 57.180 178.520 ;
        RECT 47.750 178.180 55.340 178.320 ;
        RECT 47.750 178.120 48.070 178.180 ;
        RECT 56.965 178.135 57.255 178.365 ;
        RECT 57.425 178.135 57.715 178.365 ;
        RECT 57.960 178.320 58.100 178.520 ;
        RECT 58.345 178.520 61.395 178.660 ;
        RECT 63.020 178.660 63.160 178.800 ;
        RECT 66.610 178.660 66.930 178.720 ;
        RECT 63.020 178.520 66.930 178.660 ;
        RECT 58.345 178.475 58.635 178.520 ;
        RECT 61.105 178.475 61.395 178.520 ;
        RECT 66.610 178.460 66.930 178.520 ;
        RECT 72.590 178.460 72.910 178.720 ;
        RECT 59.710 178.320 60.030 178.380 ;
        RECT 57.960 178.180 60.030 178.320 ;
        RECT 40.390 177.980 40.710 178.040 ;
        RECT 39.560 177.840 40.710 177.980 ;
        RECT 22.450 177.440 22.770 177.700 ;
        RECT 23.305 177.640 23.595 177.685 ;
        RECT 28.445 177.640 28.735 177.685 ;
        RECT 23.305 177.500 28.735 177.640 ;
        RECT 35.420 177.640 35.560 177.840 ;
        RECT 39.025 177.795 39.315 177.840 ;
        RECT 40.390 177.780 40.710 177.840 ;
        RECT 53.270 177.980 53.590 178.040 ;
        RECT 57.500 177.980 57.640 178.135 ;
        RECT 59.710 178.120 60.030 178.180 ;
        RECT 60.170 178.120 60.490 178.380 ;
        RECT 60.630 178.120 60.950 178.380 ;
        RECT 61.550 178.120 61.870 178.380 ;
        RECT 62.470 178.120 62.790 178.380 ;
        RECT 63.405 178.135 63.695 178.365 ;
        RECT 58.330 177.980 58.650 178.040 ;
        RECT 58.805 177.980 59.095 178.025 ;
        RECT 53.270 177.840 59.095 177.980 ;
        RECT 63.480 177.980 63.620 178.135 ;
        RECT 63.850 178.120 64.170 178.380 ;
        RECT 70.750 178.320 71.070 178.380 ;
        RECT 72.145 178.320 72.435 178.365 ;
        RECT 70.750 178.180 72.435 178.320 ;
        RECT 75.900 178.320 76.040 178.860 ;
        RECT 76.730 178.860 80.690 179.000 ;
        RECT 76.730 178.815 77.020 178.860 ;
        RECT 78.300 178.815 78.590 178.860 ;
        RECT 80.400 178.815 80.690 178.860 ;
        RECT 85.050 179.000 85.340 179.045 ;
        RECT 87.150 179.000 87.440 179.045 ;
        RECT 88.720 179.000 89.010 179.045 ;
        RECT 85.050 178.860 89.010 179.000 ;
        RECT 85.050 178.815 85.340 178.860 ;
        RECT 87.150 178.815 87.440 178.860 ;
        RECT 88.720 178.815 89.010 178.860 ;
        RECT 91.465 179.000 91.755 179.045 ;
        RECT 94.670 179.000 94.990 179.060 ;
        RECT 91.465 178.860 94.990 179.000 ;
        RECT 91.465 178.815 91.755 178.860 ;
        RECT 94.670 178.800 94.990 178.860 ;
        RECT 95.590 179.000 95.880 179.045 ;
        RECT 97.160 179.000 97.450 179.045 ;
        RECT 99.260 179.000 99.550 179.045 ;
        RECT 95.590 178.860 99.550 179.000 ;
        RECT 95.590 178.815 95.880 178.860 ;
        RECT 97.160 178.815 97.450 178.860 ;
        RECT 99.260 178.815 99.550 178.860 ;
        RECT 119.510 179.000 119.800 179.045 ;
        RECT 121.080 179.000 121.370 179.045 ;
        RECT 123.180 179.000 123.470 179.045 ;
        RECT 119.510 178.860 123.470 179.000 ;
        RECT 119.510 178.815 119.800 178.860 ;
        RECT 121.080 178.815 121.370 178.860 ;
        RECT 123.180 178.815 123.470 178.860 ;
        RECT 126.410 179.000 126.730 179.060 ;
        RECT 129.260 179.000 129.400 179.155 ;
        RECT 132.850 179.140 133.170 179.200 ;
        RECT 140.670 179.340 140.990 179.400 ;
        RECT 141.145 179.340 141.435 179.385 ;
        RECT 140.670 179.200 141.435 179.340 ;
        RECT 140.670 179.140 140.990 179.200 ;
        RECT 141.145 179.155 141.435 179.200 ;
        RECT 126.410 178.860 129.400 179.000 ;
        RECT 129.630 179.000 129.950 179.060 ;
        RECT 131.470 179.000 131.790 179.060 ;
        RECT 129.630 178.860 131.790 179.000 ;
        RECT 126.410 178.800 126.730 178.860 ;
        RECT 129.630 178.800 129.950 178.860 ;
        RECT 131.470 178.800 131.790 178.860 ;
        RECT 134.270 179.000 134.560 179.045 ;
        RECT 136.370 179.000 136.660 179.045 ;
        RECT 137.940 179.000 138.230 179.045 ;
        RECT 134.270 178.860 138.230 179.000 ;
        RECT 134.270 178.815 134.560 178.860 ;
        RECT 136.370 178.815 136.660 178.860 ;
        RECT 137.940 178.815 138.230 178.860 ;
        RECT 76.295 178.660 76.585 178.705 ;
        RECT 78.815 178.660 79.105 178.705 ;
        RECT 80.005 178.660 80.295 178.705 ;
        RECT 76.295 178.520 80.295 178.660 ;
        RECT 76.295 178.475 76.585 178.520 ;
        RECT 78.815 178.475 79.105 178.520 ;
        RECT 80.005 178.475 80.295 178.520 ;
        RECT 85.445 178.660 85.735 178.705 ;
        RECT 86.635 178.660 86.925 178.705 ;
        RECT 89.155 178.660 89.445 178.705 ;
        RECT 85.445 178.520 89.445 178.660 ;
        RECT 85.445 178.475 85.735 178.520 ;
        RECT 86.635 178.475 86.925 178.520 ;
        RECT 89.155 178.475 89.445 178.520 ;
        RECT 95.155 178.660 95.445 178.705 ;
        RECT 97.675 178.660 97.965 178.705 ;
        RECT 98.865 178.660 99.155 178.705 ;
        RECT 95.155 178.520 99.155 178.660 ;
        RECT 95.155 178.475 95.445 178.520 ;
        RECT 97.675 178.475 97.965 178.520 ;
        RECT 98.865 178.475 99.155 178.520 ;
        RECT 99.730 178.460 100.050 178.720 ;
        RECT 102.490 178.460 102.810 178.720 ;
        RECT 102.965 178.660 103.255 178.705 ;
        RECT 103.410 178.660 103.730 178.720 ;
        RECT 102.965 178.520 103.730 178.660 ;
        RECT 102.965 178.475 103.255 178.520 ;
        RECT 79.550 178.320 79.840 178.365 ;
        RECT 75.900 178.180 79.840 178.320 ;
        RECT 70.750 178.120 71.070 178.180 ;
        RECT 72.145 178.135 72.435 178.180 ;
        RECT 79.550 178.135 79.840 178.180 ;
        RECT 80.885 178.320 81.175 178.365 ;
        RECT 81.330 178.320 81.650 178.380 ;
        RECT 84.565 178.320 84.855 178.365 ;
        RECT 101.110 178.320 101.430 178.380 ;
        RECT 103.040 178.320 103.180 178.475 ;
        RECT 103.410 178.460 103.730 178.520 ;
        RECT 119.075 178.660 119.365 178.705 ;
        RECT 121.595 178.660 121.885 178.705 ;
        RECT 122.785 178.660 123.075 178.705 ;
        RECT 119.075 178.520 123.075 178.660 ;
        RECT 119.075 178.475 119.365 178.520 ;
        RECT 121.595 178.475 121.885 178.520 ;
        RECT 122.785 178.475 123.075 178.520 ;
        RECT 123.650 178.660 123.970 178.720 ;
        RECT 127.330 178.660 127.650 178.720 ;
        RECT 133.785 178.660 134.075 178.705 ;
        RECT 123.650 178.520 134.075 178.660 ;
        RECT 123.650 178.460 123.970 178.520 ;
        RECT 127.330 178.460 127.650 178.520 ;
        RECT 133.785 178.475 134.075 178.520 ;
        RECT 134.665 178.660 134.955 178.705 ;
        RECT 135.855 178.660 136.145 178.705 ;
        RECT 138.375 178.660 138.665 178.705 ;
        RECT 134.665 178.520 138.665 178.660 ;
        RECT 134.665 178.475 134.955 178.520 ;
        RECT 135.855 178.475 136.145 178.520 ;
        RECT 138.375 178.475 138.665 178.520 ;
        RECT 138.920 178.520 143.200 178.660 ;
        RECT 80.885 178.180 86.620 178.320 ;
        RECT 80.885 178.135 81.175 178.180 ;
        RECT 81.330 178.120 81.650 178.180 ;
        RECT 84.565 178.135 84.855 178.180 ;
        RECT 86.480 178.040 86.620 178.180 ;
        RECT 101.110 178.180 103.180 178.320 ;
        RECT 108.945 178.320 109.235 178.365 ;
        RECT 110.310 178.320 110.630 178.380 ;
        RECT 108.945 178.180 110.630 178.320 ;
        RECT 101.110 178.120 101.430 178.180 ;
        RECT 108.945 178.135 109.235 178.180 ;
        RECT 110.310 178.120 110.630 178.180 ;
        RECT 110.770 178.120 111.090 178.380 ;
        RECT 122.270 178.365 122.590 178.380 ;
        RECT 122.270 178.135 122.620 178.365 ;
        RECT 125.045 178.320 125.335 178.365 ;
        RECT 126.885 178.320 127.175 178.365 ;
        RECT 128.250 178.320 128.570 178.380 ;
        RECT 125.045 178.180 126.640 178.320 ;
        RECT 125.045 178.135 125.335 178.180 ;
        RECT 122.270 178.120 122.590 178.135 ;
        RECT 66.610 177.980 66.930 178.040 ;
        RECT 63.480 177.840 66.930 177.980 ;
        RECT 53.270 177.780 53.590 177.840 ;
        RECT 58.330 177.780 58.650 177.840 ;
        RECT 58.805 177.795 59.095 177.840 ;
        RECT 66.610 177.780 66.930 177.840 ;
        RECT 73.510 177.780 73.830 178.040 ;
        RECT 85.930 178.025 86.250 178.040 ;
        RECT 85.900 177.980 86.250 178.025 ;
        RECT 85.735 177.840 86.250 177.980 ;
        RECT 85.900 177.795 86.250 177.840 ;
        RECT 85.930 177.780 86.250 177.795 ;
        RECT 86.390 177.780 86.710 178.040 ;
        RECT 98.520 177.980 98.810 178.025 ;
        RECT 98.520 177.840 100.420 177.980 ;
        RECT 98.520 177.795 98.810 177.840 ;
        RECT 37.630 177.640 37.950 177.700 ;
        RECT 35.420 177.500 37.950 177.640 ;
        RECT 23.305 177.455 23.595 177.500 ;
        RECT 28.445 177.455 28.735 177.500 ;
        RECT 37.630 177.440 37.950 177.500 ;
        RECT 38.090 177.440 38.410 177.700 ;
        RECT 42.705 177.640 42.995 177.685 ;
        RECT 45.450 177.640 45.770 177.700 ;
        RECT 42.705 177.500 45.770 177.640 ;
        RECT 42.705 177.455 42.995 177.500 ;
        RECT 45.450 177.440 45.770 177.500 ;
        RECT 73.970 177.440 74.290 177.700 ;
        RECT 100.280 177.685 100.420 177.840 ;
        RECT 109.405 177.795 109.695 178.025 ;
        RECT 109.865 177.980 110.155 178.025 ;
        RECT 115.830 177.980 116.150 178.040 ;
        RECT 125.490 177.980 125.810 178.040 ;
        RECT 109.865 177.840 116.150 177.980 ;
        RECT 109.865 177.795 110.155 177.840 ;
        RECT 100.205 177.455 100.495 177.685 ;
        RECT 102.045 177.640 102.335 177.685 ;
        RECT 107.550 177.640 107.870 177.700 ;
        RECT 102.045 177.500 107.870 177.640 ;
        RECT 102.045 177.455 102.335 177.500 ;
        RECT 107.550 177.440 107.870 177.500 ;
        RECT 108.025 177.640 108.315 177.685 ;
        RECT 108.470 177.640 108.790 177.700 ;
        RECT 108.025 177.500 108.790 177.640 ;
        RECT 109.480 177.640 109.620 177.795 ;
        RECT 115.830 177.780 116.150 177.840 ;
        RECT 122.130 177.840 125.810 177.980 ;
        RECT 112.150 177.640 112.470 177.700 ;
        RECT 122.130 177.640 122.270 177.840 ;
        RECT 125.490 177.780 125.810 177.840 ;
        RECT 125.950 177.780 126.270 178.040 ;
        RECT 126.500 177.980 126.640 178.180 ;
        RECT 126.885 178.180 128.570 178.320 ;
        RECT 126.885 178.135 127.175 178.180 ;
        RECT 128.250 178.120 128.570 178.180 ;
        RECT 128.725 178.135 129.015 178.365 ;
        RECT 127.790 177.980 128.110 178.040 ;
        RECT 126.500 177.840 128.110 177.980 ;
        RECT 128.800 177.980 128.940 178.135 ;
        RECT 129.170 178.120 129.490 178.380 ;
        RECT 129.630 178.120 129.950 178.380 ;
        RECT 131.930 178.120 132.250 178.380 ;
        RECT 133.860 178.320 134.000 178.475 ;
        RECT 137.450 178.320 137.770 178.380 ;
        RECT 133.860 178.180 137.770 178.320 ;
        RECT 137.450 178.120 137.770 178.180 ;
        RECT 129.720 177.980 129.860 178.120 ;
        RECT 130.550 178.025 130.870 178.040 ;
        RECT 128.800 177.840 129.860 177.980 ;
        RECT 127.790 177.780 128.110 177.840 ;
        RECT 130.435 177.795 130.870 178.025 ;
        RECT 131.025 177.795 131.315 178.025 ;
        RECT 131.485 177.980 131.775 178.025 ;
        RECT 132.390 177.980 132.710 178.040 ;
        RECT 131.485 177.840 132.710 177.980 ;
        RECT 131.485 177.795 131.775 177.840 ;
        RECT 130.550 177.780 130.870 177.795 ;
        RECT 109.480 177.500 122.270 177.640 ;
        RECT 129.170 177.640 129.490 177.700 ;
        RECT 131.100 177.640 131.240 177.795 ;
        RECT 132.390 177.780 132.710 177.840 ;
        RECT 132.865 177.980 133.155 178.025 ;
        RECT 135.010 177.980 135.300 178.025 ;
        RECT 132.865 177.840 135.300 177.980 ;
        RECT 132.865 177.795 133.155 177.840 ;
        RECT 135.010 177.795 135.300 177.840 ;
        RECT 135.610 177.980 135.930 178.040 ;
        RECT 138.920 177.980 139.060 178.520 ;
        RECT 142.050 178.120 142.370 178.380 ;
        RECT 143.060 178.365 143.200 178.520 ;
        RECT 142.985 178.135 143.275 178.365 ;
        RECT 143.890 178.120 144.210 178.380 ;
        RECT 142.525 177.980 142.815 178.025 ;
        RECT 135.610 177.840 139.060 177.980 ;
        RECT 139.380 177.840 142.815 177.980 ;
        RECT 135.610 177.780 135.930 177.840 ;
        RECT 129.170 177.500 131.240 177.640 ;
        RECT 132.480 177.640 132.620 177.780 ;
        RECT 139.380 177.640 139.520 177.840 ;
        RECT 142.525 177.795 142.815 177.840 ;
        RECT 132.480 177.500 139.520 177.640 ;
        RECT 108.025 177.455 108.315 177.500 ;
        RECT 108.470 177.440 108.790 177.500 ;
        RECT 112.150 177.440 112.470 177.500 ;
        RECT 129.170 177.440 129.490 177.500 ;
        RECT 140.670 177.440 140.990 177.700 ;
        RECT 17.320 176.820 147.040 177.300 ;
        RECT 30.270 176.665 30.590 176.680 ;
        RECT 26.605 176.435 26.895 176.665 ;
        RECT 30.205 176.435 30.590 176.665 ;
        RECT 21.040 176.280 21.330 176.325 ;
        RECT 22.450 176.280 22.770 176.340 ;
        RECT 21.040 176.140 22.770 176.280 ;
        RECT 26.680 176.280 26.820 176.435 ;
        RECT 30.270 176.420 30.590 176.435 ;
        RECT 32.110 176.420 32.430 176.680 ;
        RECT 39.010 176.620 39.330 176.680 ;
        RECT 38.180 176.480 39.330 176.620 ;
        RECT 27.050 176.280 27.370 176.340 ;
        RECT 28.065 176.280 28.355 176.325 ;
        RECT 26.680 176.140 27.370 176.280 ;
        RECT 21.040 176.095 21.330 176.140 ;
        RECT 22.450 176.080 22.770 176.140 ;
        RECT 27.050 176.080 27.370 176.140 ;
        RECT 27.600 176.140 28.355 176.280 ;
        RECT 26.130 175.940 26.450 176.000 ;
        RECT 27.600 175.940 27.740 176.140 ;
        RECT 28.065 176.095 28.355 176.140 ;
        RECT 31.190 176.080 31.510 176.340 ;
        RECT 26.130 175.800 27.740 175.940 ;
        RECT 26.130 175.740 26.450 175.800 ;
        RECT 31.665 175.755 31.955 175.985 ;
        RECT 37.185 175.940 37.475 175.985 ;
        RECT 37.630 175.940 37.950 176.000 ;
        RECT 38.180 175.985 38.320 176.480 ;
        RECT 39.010 176.420 39.330 176.480 ;
        RECT 39.930 176.620 40.250 176.680 ;
        RECT 40.865 176.620 41.155 176.665 ;
        RECT 39.930 176.480 41.155 176.620 ;
        RECT 39.930 176.420 40.250 176.480 ;
        RECT 40.865 176.435 41.155 176.480 ;
        RECT 60.170 176.620 60.490 176.680 ;
        RECT 61.565 176.620 61.855 176.665 ;
        RECT 60.170 176.480 61.855 176.620 ;
        RECT 60.170 176.420 60.490 176.480 ;
        RECT 61.565 176.435 61.855 176.480 ;
        RECT 62.010 176.620 62.330 176.680 ;
        RECT 63.850 176.620 64.170 176.680 ;
        RECT 110.310 176.620 110.630 176.680 ;
        RECT 113.990 176.620 114.310 176.680 ;
        RECT 62.010 176.480 64.540 176.620 ;
        RECT 62.010 176.420 62.330 176.480 ;
        RECT 63.850 176.420 64.170 176.480 ;
        RECT 38.550 176.280 38.870 176.340 ;
        RECT 44.990 176.280 45.310 176.340 ;
        RECT 38.550 176.140 41.540 176.280 ;
        RECT 38.550 176.080 38.870 176.140 ;
        RECT 39.100 175.985 39.240 176.140 ;
        RECT 41.400 175.985 41.540 176.140 ;
        RECT 42.320 176.140 45.310 176.280 ;
        RECT 42.320 175.985 42.460 176.140 ;
        RECT 44.990 176.080 45.310 176.140 ;
        RECT 60.630 176.280 60.950 176.340 ;
        RECT 62.945 176.280 63.235 176.325 ;
        RECT 60.630 176.140 63.235 176.280 ;
        RECT 60.630 176.080 60.950 176.140 ;
        RECT 62.945 176.095 63.235 176.140 ;
        RECT 64.400 176.280 64.540 176.480 ;
        RECT 110.310 176.480 114.310 176.620 ;
        RECT 110.310 176.420 110.630 176.480 ;
        RECT 113.990 176.420 114.310 176.480 ;
        RECT 124.125 176.620 124.415 176.665 ;
        RECT 125.950 176.620 126.270 176.680 ;
        RECT 129.630 176.620 129.950 176.680 ;
        RECT 131.930 176.620 132.250 176.680 ;
        RECT 124.125 176.480 126.270 176.620 ;
        RECT 124.125 176.435 124.415 176.480 ;
        RECT 125.950 176.420 126.270 176.480 ;
        RECT 126.960 176.480 129.950 176.620 ;
        RECT 66.150 176.280 66.470 176.340 ;
        RECT 64.400 176.140 66.470 176.280 ;
        RECT 37.185 175.800 37.950 175.940 ;
        RECT 37.185 175.755 37.475 175.800 ;
        RECT 19.705 175.415 19.995 175.645 ;
        RECT 20.585 175.600 20.875 175.645 ;
        RECT 21.775 175.600 22.065 175.645 ;
        RECT 24.295 175.600 24.585 175.645 ;
        RECT 20.585 175.460 24.585 175.600 ;
        RECT 20.585 175.415 20.875 175.460 ;
        RECT 21.775 175.415 22.065 175.460 ;
        RECT 24.295 175.415 24.585 175.460 ;
        RECT 19.780 174.920 19.920 175.415 ;
        RECT 20.190 175.260 20.480 175.305 ;
        RECT 22.290 175.260 22.580 175.305 ;
        RECT 23.860 175.260 24.150 175.305 ;
        RECT 20.190 175.120 24.150 175.260 ;
        RECT 20.190 175.075 20.480 175.120 ;
        RECT 22.290 175.075 22.580 175.120 ;
        RECT 23.860 175.075 24.150 175.120 ;
        RECT 26.590 175.260 26.910 175.320 ;
        RECT 28.905 175.260 29.195 175.305 ;
        RECT 31.740 175.260 31.880 175.755 ;
        RECT 37.630 175.740 37.950 175.800 ;
        RECT 38.105 175.755 38.395 175.985 ;
        RECT 39.025 175.755 39.315 175.985 ;
        RECT 39.945 175.755 40.235 175.985 ;
        RECT 41.325 175.755 41.615 175.985 ;
        RECT 42.245 175.755 42.535 175.985 ;
        RECT 42.690 175.940 43.010 176.000 ;
        RECT 44.545 175.940 44.835 175.985 ;
        RECT 42.690 175.800 44.835 175.940 ;
        RECT 34.870 175.600 35.190 175.660 ;
        RECT 38.565 175.600 38.855 175.645 ;
        RECT 34.870 175.460 38.855 175.600 ;
        RECT 40.020 175.600 40.160 175.755 ;
        RECT 40.390 175.600 40.710 175.660 ;
        RECT 42.320 175.600 42.460 175.755 ;
        RECT 42.690 175.740 43.010 175.800 ;
        RECT 44.545 175.755 44.835 175.800 ;
        RECT 45.450 175.740 45.770 176.000 ;
        RECT 45.910 175.740 46.230 176.000 ;
        RECT 61.105 175.755 61.395 175.985 ;
        RECT 40.020 175.460 42.460 175.600 ;
        RECT 61.180 175.600 61.320 175.755 ;
        RECT 62.010 175.740 62.330 176.000 ;
        RECT 63.390 175.940 63.710 176.000 ;
        RECT 64.400 175.985 64.540 176.140 ;
        RECT 66.150 176.080 66.470 176.140 ;
        RECT 126.410 176.080 126.730 176.340 ;
        RECT 63.865 175.940 64.155 175.985 ;
        RECT 63.390 175.800 64.155 175.940 ;
        RECT 63.390 175.740 63.710 175.800 ;
        RECT 63.865 175.755 64.155 175.800 ;
        RECT 64.325 175.755 64.615 175.985 ;
        RECT 65.245 175.755 65.535 175.985 ;
        RECT 65.705 175.940 65.995 175.985 ;
        RECT 66.610 175.940 66.930 176.000 ;
        RECT 65.705 175.800 66.930 175.940 ;
        RECT 65.705 175.755 65.995 175.800 ;
        RECT 63.480 175.600 63.620 175.740 ;
        RECT 61.180 175.460 63.620 175.600 ;
        RECT 65.320 175.600 65.460 175.755 ;
        RECT 66.610 175.740 66.930 175.800 ;
        RECT 72.590 175.940 72.910 176.000 ;
        RECT 78.125 175.940 78.415 175.985 ;
        RECT 72.590 175.800 78.415 175.940 ;
        RECT 72.590 175.740 72.910 175.800 ;
        RECT 78.125 175.755 78.415 175.800 ;
        RECT 79.045 175.755 79.335 175.985 ;
        RECT 88.660 175.940 88.950 175.985 ;
        RECT 94.670 175.940 94.990 176.000 ;
        RECT 88.660 175.800 94.990 175.940 ;
        RECT 88.660 175.755 88.950 175.800 ;
        RECT 73.050 175.600 73.370 175.660 ;
        RECT 74.445 175.600 74.735 175.645 ;
        RECT 65.320 175.460 74.735 175.600 ;
        RECT 34.870 175.400 35.190 175.460 ;
        RECT 38.565 175.415 38.855 175.460 ;
        RECT 40.390 175.400 40.710 175.460 ;
        RECT 73.050 175.400 73.370 175.460 ;
        RECT 74.445 175.415 74.735 175.460 ;
        RECT 77.665 175.600 77.955 175.645 ;
        RECT 79.120 175.600 79.260 175.755 ;
        RECT 94.670 175.740 94.990 175.800 ;
        RECT 98.350 175.740 98.670 176.000 ;
        RECT 99.730 175.940 100.050 176.000 ;
        RECT 106.645 175.940 106.935 175.985 ;
        RECT 108.010 175.940 108.330 176.000 ;
        RECT 99.730 175.800 108.330 175.940 ;
        RECT 99.730 175.740 100.050 175.800 ;
        RECT 106.645 175.755 106.935 175.800 ;
        RECT 108.010 175.740 108.330 175.800 ;
        RECT 110.310 175.940 110.630 176.000 ;
        RECT 110.785 175.940 111.075 175.985 ;
        RECT 110.310 175.800 111.075 175.940 ;
        RECT 110.310 175.740 110.630 175.800 ;
        RECT 110.785 175.755 111.075 175.800 ;
        RECT 111.230 175.740 111.550 176.000 ;
        RECT 125.045 175.755 125.335 175.985 ;
        RECT 125.965 175.940 126.255 175.985 ;
        RECT 126.960 175.940 127.100 176.480 ;
        RECT 129.630 176.420 129.950 176.480 ;
        RECT 130.640 176.480 132.250 176.620 ;
        RECT 127.505 176.280 127.795 176.325 ;
        RECT 129.170 176.280 129.490 176.340 ;
        RECT 127.505 176.140 129.490 176.280 ;
        RECT 127.505 176.095 127.795 176.140 ;
        RECT 129.170 176.080 129.490 176.140 ;
        RECT 125.965 175.800 127.100 175.940 ;
        RECT 125.965 175.755 126.255 175.800 ;
        RECT 128.725 175.755 129.015 175.985 ;
        RECT 129.705 175.940 129.995 175.985 ;
        RECT 130.640 175.940 130.780 176.480 ;
        RECT 131.930 176.420 132.250 176.480 ;
        RECT 132.850 176.420 133.170 176.680 ;
        RECT 135.165 176.620 135.455 176.665 ;
        RECT 135.610 176.620 135.930 176.680 ;
        RECT 135.165 176.480 135.930 176.620 ;
        RECT 135.165 176.435 135.455 176.480 ;
        RECT 135.610 176.420 135.930 176.480 ;
        RECT 132.940 176.280 133.080 176.420 ;
        RECT 143.890 176.280 144.210 176.340 ;
        RECT 131.100 176.140 144.210 176.280 ;
        RECT 131.100 175.985 131.240 176.140 ;
        RECT 143.890 176.080 144.210 176.140 ;
        RECT 129.705 175.800 130.780 175.940 ;
        RECT 129.705 175.755 129.995 175.800 ;
        RECT 131.025 175.755 131.315 175.985 ;
        RECT 131.470 175.940 131.790 176.000 ;
        RECT 131.945 175.940 132.235 175.985 ;
        RECT 131.470 175.800 132.235 175.940 ;
        RECT 77.665 175.460 79.260 175.600 ;
        RECT 86.390 175.600 86.710 175.660 ;
        RECT 87.325 175.600 87.615 175.645 ;
        RECT 86.390 175.460 87.615 175.600 ;
        RECT 77.665 175.415 77.955 175.460 ;
        RECT 86.390 175.400 86.710 175.460 ;
        RECT 87.325 175.415 87.615 175.460 ;
        RECT 88.205 175.600 88.495 175.645 ;
        RECT 89.395 175.600 89.685 175.645 ;
        RECT 91.915 175.600 92.205 175.645 ;
        RECT 88.205 175.460 92.205 175.600 ;
        RECT 88.205 175.415 88.495 175.460 ;
        RECT 89.395 175.415 89.685 175.460 ;
        RECT 91.915 175.415 92.205 175.460 ;
        RECT 95.130 175.600 95.450 175.660 ;
        RECT 99.820 175.600 99.960 175.740 ;
        RECT 95.130 175.460 99.960 175.600 ;
        RECT 95.130 175.400 95.450 175.460 ;
        RECT 101.585 175.415 101.875 175.645 ;
        RECT 26.590 175.120 31.880 175.260 ;
        RECT 39.930 175.260 40.250 175.320 ;
        RECT 45.005 175.260 45.295 175.305 ;
        RECT 39.930 175.120 45.295 175.260 ;
        RECT 26.590 175.060 26.910 175.120 ;
        RECT 28.905 175.075 29.195 175.120 ;
        RECT 39.930 175.060 40.250 175.120 ;
        RECT 45.005 175.075 45.295 175.120 ;
        RECT 87.810 175.260 88.100 175.305 ;
        RECT 89.910 175.260 90.200 175.305 ;
        RECT 91.480 175.260 91.770 175.305 ;
        RECT 87.810 175.120 91.770 175.260 ;
        RECT 87.810 175.075 88.100 175.120 ;
        RECT 89.910 175.075 90.200 175.120 ;
        RECT 91.480 175.075 91.770 175.120 ;
        RECT 94.225 175.260 94.515 175.305 ;
        RECT 96.970 175.260 97.290 175.320 ;
        RECT 101.660 175.260 101.800 175.415 ;
        RECT 105.250 175.400 105.570 175.660 ;
        RECT 123.650 175.600 123.970 175.660 ;
        RECT 125.120 175.600 125.260 175.755 ;
        RECT 128.250 175.600 128.570 175.660 ;
        RECT 123.650 175.460 128.570 175.600 ;
        RECT 123.650 175.400 123.970 175.460 ;
        RECT 128.250 175.400 128.570 175.460 ;
        RECT 94.225 175.120 101.800 175.260 ;
        RECT 112.165 175.260 112.455 175.305 ;
        RECT 115.370 175.260 115.690 175.320 ;
        RECT 128.800 175.260 128.940 175.755 ;
        RECT 131.470 175.740 131.790 175.800 ;
        RECT 131.945 175.755 132.235 175.800 ;
        RECT 133.770 175.740 134.090 176.000 ;
        RECT 134.245 175.940 134.535 175.985 ;
        RECT 134.690 175.940 135.010 176.000 ;
        RECT 134.245 175.800 135.010 175.940 ;
        RECT 134.245 175.755 134.535 175.800 ;
        RECT 134.690 175.740 135.010 175.800 ;
        RECT 136.530 175.740 136.850 176.000 ;
        RECT 137.450 175.740 137.770 176.000 ;
        RECT 137.910 175.740 138.230 176.000 ;
        RECT 138.830 175.985 139.150 176.000 ;
        RECT 138.800 175.755 139.150 175.985 ;
        RECT 138.830 175.740 139.150 175.755 ;
        RECT 130.550 175.600 130.870 175.660 ;
        RECT 132.865 175.600 133.155 175.645 ;
        RECT 130.550 175.460 133.155 175.600 ;
        RECT 130.550 175.400 130.870 175.460 ;
        RECT 132.865 175.415 133.155 175.460 ;
        RECT 133.310 175.600 133.630 175.660 ;
        RECT 138.000 175.600 138.140 175.740 ;
        RECT 133.310 175.460 138.140 175.600 ;
        RECT 138.345 175.600 138.635 175.645 ;
        RECT 139.535 175.600 139.825 175.645 ;
        RECT 142.055 175.600 142.345 175.645 ;
        RECT 138.345 175.460 142.345 175.600 ;
        RECT 133.310 175.400 133.630 175.460 ;
        RECT 138.345 175.415 138.635 175.460 ;
        RECT 139.535 175.415 139.825 175.460 ;
        RECT 142.055 175.415 142.345 175.460 ;
        RECT 112.165 175.120 115.690 175.260 ;
        RECT 94.225 175.075 94.515 175.120 ;
        RECT 96.970 175.060 97.290 175.120 ;
        RECT 112.165 175.075 112.455 175.120 ;
        RECT 115.370 175.060 115.690 175.120 ;
        RECT 127.420 175.120 128.940 175.260 ;
        RECT 25.210 174.920 25.530 174.980 ;
        RECT 19.780 174.780 25.530 174.920 ;
        RECT 25.210 174.720 25.530 174.780 ;
        RECT 25.670 174.920 25.990 174.980 ;
        RECT 27.985 174.920 28.275 174.965 ;
        RECT 25.670 174.780 28.275 174.920 ;
        RECT 25.670 174.720 25.990 174.780 ;
        RECT 27.985 174.735 28.275 174.780 ;
        RECT 29.350 174.720 29.670 174.980 ;
        RECT 29.810 174.920 30.130 174.980 ;
        RECT 30.285 174.920 30.575 174.965 ;
        RECT 29.810 174.780 30.575 174.920 ;
        RECT 29.810 174.720 30.130 174.780 ;
        RECT 30.285 174.735 30.575 174.780 ;
        RECT 38.550 174.920 38.870 174.980 ;
        RECT 41.325 174.920 41.615 174.965 ;
        RECT 38.550 174.780 41.615 174.920 ;
        RECT 38.550 174.720 38.870 174.780 ;
        RECT 41.325 174.735 41.615 174.780 ;
        RECT 43.610 174.720 43.930 174.980 ;
        RECT 78.110 174.720 78.430 174.980 ;
        RECT 95.145 174.920 95.435 174.965 ;
        RECT 96.050 174.920 96.370 174.980 ;
        RECT 95.145 174.780 96.370 174.920 ;
        RECT 95.145 174.735 95.435 174.780 ;
        RECT 96.050 174.720 96.370 174.780 ;
        RECT 97.430 174.920 97.750 174.980 ;
        RECT 98.825 174.920 99.115 174.965 ;
        RECT 97.430 174.780 99.115 174.920 ;
        RECT 97.430 174.720 97.750 174.780 ;
        RECT 98.825 174.735 99.115 174.780 ;
        RECT 102.505 174.920 102.795 174.965 ;
        RECT 102.950 174.920 103.270 174.980 ;
        RECT 102.505 174.780 103.270 174.920 ;
        RECT 102.505 174.735 102.795 174.780 ;
        RECT 102.950 174.720 103.270 174.780 ;
        RECT 105.710 174.920 106.030 174.980 ;
        RECT 109.405 174.920 109.695 174.965 ;
        RECT 105.710 174.780 109.695 174.920 ;
        RECT 105.710 174.720 106.030 174.780 ;
        RECT 109.405 174.735 109.695 174.780 ;
        RECT 126.870 174.920 127.190 174.980 ;
        RECT 127.420 174.965 127.560 175.120 ;
        RECT 127.345 174.920 127.635 174.965 ;
        RECT 126.870 174.780 127.635 174.920 ;
        RECT 126.870 174.720 127.190 174.780 ;
        RECT 127.345 174.735 127.635 174.780 ;
        RECT 127.790 174.920 128.110 174.980 ;
        RECT 128.265 174.920 128.555 174.965 ;
        RECT 127.790 174.780 128.555 174.920 ;
        RECT 128.800 174.920 128.940 175.120 ;
        RECT 129.645 175.260 129.935 175.305 ;
        RECT 130.090 175.260 130.410 175.320 ;
        RECT 129.645 175.120 130.410 175.260 ;
        RECT 129.645 175.075 129.935 175.120 ;
        RECT 130.090 175.060 130.410 175.120 ;
        RECT 132.390 175.260 132.710 175.320 ;
        RECT 135.610 175.260 135.930 175.320 ;
        RECT 132.390 175.120 135.930 175.260 ;
        RECT 132.390 175.060 132.710 175.120 ;
        RECT 135.610 175.060 135.930 175.120 ;
        RECT 137.950 175.260 138.240 175.305 ;
        RECT 140.050 175.260 140.340 175.305 ;
        RECT 141.620 175.260 141.910 175.305 ;
        RECT 137.950 175.120 141.910 175.260 ;
        RECT 137.950 175.075 138.240 175.120 ;
        RECT 140.050 175.075 140.340 175.120 ;
        RECT 141.620 175.075 141.910 175.120 ;
        RECT 131.930 174.920 132.250 174.980 ;
        RECT 136.070 174.920 136.390 174.980 ;
        RECT 128.800 174.780 136.390 174.920 ;
        RECT 127.790 174.720 128.110 174.780 ;
        RECT 128.265 174.735 128.555 174.780 ;
        RECT 131.930 174.720 132.250 174.780 ;
        RECT 136.070 174.720 136.390 174.780 ;
        RECT 136.530 174.920 136.850 174.980 ;
        RECT 144.365 174.920 144.655 174.965 ;
        RECT 136.530 174.780 144.655 174.920 ;
        RECT 136.530 174.720 136.850 174.780 ;
        RECT 144.365 174.735 144.655 174.780 ;
        RECT 17.320 174.100 147.040 174.580 ;
        RECT 22.005 173.900 22.295 173.945 ;
        RECT 25.670 173.900 25.990 173.960 ;
        RECT 22.005 173.760 25.990 173.900 ;
        RECT 22.005 173.715 22.295 173.760 ;
        RECT 25.670 173.700 25.990 173.760 ;
        RECT 45.005 173.900 45.295 173.945 ;
        RECT 45.910 173.900 46.230 173.960 ;
        RECT 45.005 173.760 46.230 173.900 ;
        RECT 45.005 173.715 45.295 173.760 ;
        RECT 45.910 173.700 46.230 173.760 ;
        RECT 65.230 173.900 65.550 173.960 ;
        RECT 66.610 173.900 66.930 173.960 ;
        RECT 65.230 173.760 66.930 173.900 ;
        RECT 65.230 173.700 65.550 173.760 ;
        RECT 66.610 173.700 66.930 173.760 ;
        RECT 73.050 173.700 73.370 173.960 ;
        RECT 93.305 173.900 93.595 173.945 ;
        RECT 98.350 173.900 98.670 173.960 ;
        RECT 93.305 173.760 98.670 173.900 ;
        RECT 93.305 173.715 93.595 173.760 ;
        RECT 98.350 173.700 98.670 173.760 ;
        RECT 114.925 173.900 115.215 173.945 ;
        RECT 115.370 173.900 115.690 173.960 ;
        RECT 114.925 173.760 115.690 173.900 ;
        RECT 114.925 173.715 115.215 173.760 ;
        RECT 115.370 173.700 115.690 173.760 ;
        RECT 123.650 173.700 123.970 173.960 ;
        RECT 129.170 173.900 129.490 173.960 ;
        RECT 133.785 173.900 134.075 173.945 ;
        RECT 129.170 173.760 134.075 173.900 ;
        RECT 129.170 173.700 129.490 173.760 ;
        RECT 133.785 173.715 134.075 173.760 ;
        RECT 135.085 173.760 137.220 173.900 ;
        RECT 24.750 173.560 25.040 173.605 ;
        RECT 26.320 173.560 26.610 173.605 ;
        RECT 28.420 173.560 28.710 173.605 ;
        RECT 24.750 173.420 28.710 173.560 ;
        RECT 24.750 173.375 25.040 173.420 ;
        RECT 26.320 173.375 26.610 173.420 ;
        RECT 28.420 173.375 28.710 173.420 ;
        RECT 38.550 173.360 38.870 173.620 ;
        RECT 39.025 173.560 39.315 173.605 ;
        RECT 39.930 173.560 40.250 173.620 ;
        RECT 46.385 173.560 46.675 173.605 ;
        RECT 39.025 173.420 40.250 173.560 ;
        RECT 39.025 173.375 39.315 173.420 ;
        RECT 39.930 173.360 40.250 173.420 ;
        RECT 41.860 173.420 46.675 173.560 ;
        RECT 41.860 173.265 42.000 173.420 ;
        RECT 24.315 173.220 24.605 173.265 ;
        RECT 26.835 173.220 27.125 173.265 ;
        RECT 28.025 173.220 28.315 173.265 ;
        RECT 24.315 173.080 28.315 173.220 ;
        RECT 24.315 173.035 24.605 173.080 ;
        RECT 26.835 173.035 27.125 173.080 ;
        RECT 28.025 173.035 28.315 173.080 ;
        RECT 41.785 173.035 42.075 173.265 ;
        RECT 43.610 173.020 43.930 173.280 ;
        RECT 25.210 172.880 25.530 172.940 ;
        RECT 28.905 172.880 29.195 172.925 ;
        RECT 25.210 172.740 29.195 172.880 ;
        RECT 25.210 172.680 25.530 172.740 ;
        RECT 28.905 172.695 29.195 172.740 ;
        RECT 38.090 172.680 38.410 172.940 ;
        RECT 39.470 172.680 39.790 172.940 ;
        RECT 42.245 172.880 42.535 172.925 ;
        RECT 43.150 172.880 43.470 172.940 ;
        RECT 45.540 172.925 45.680 173.420 ;
        RECT 46.385 173.375 46.675 173.420 ;
        RECT 49.130 173.560 49.420 173.605 ;
        RECT 50.700 173.560 50.990 173.605 ;
        RECT 52.800 173.560 53.090 173.605 ;
        RECT 49.130 173.420 53.090 173.560 ;
        RECT 49.130 173.375 49.420 173.420 ;
        RECT 50.700 173.375 50.990 173.420 ;
        RECT 52.800 173.375 53.090 173.420 ;
        RECT 58.330 173.560 58.650 173.620 ;
        RECT 68.005 173.560 68.295 173.605 ;
        RECT 72.605 173.560 72.895 173.605 ;
        RECT 58.330 173.420 68.295 173.560 ;
        RECT 58.330 173.360 58.650 173.420 ;
        RECT 68.005 173.375 68.295 173.420 ;
        RECT 68.540 173.420 72.895 173.560 ;
        RECT 48.695 173.220 48.985 173.265 ;
        RECT 51.215 173.220 51.505 173.265 ;
        RECT 52.405 173.220 52.695 173.265 ;
        RECT 68.540 173.220 68.680 173.420 ;
        RECT 72.605 173.375 72.895 173.420 ;
        RECT 48.695 173.080 52.695 173.220 ;
        RECT 48.695 173.035 48.985 173.080 ;
        RECT 51.215 173.035 51.505 173.080 ;
        RECT 52.405 173.035 52.695 173.080 ;
        RECT 66.700 173.080 68.680 173.220 ;
        RECT 70.765 173.220 71.055 173.265 ;
        RECT 73.140 173.220 73.280 173.700 ;
        RECT 75.810 173.560 76.100 173.605 ;
        RECT 77.380 173.560 77.670 173.605 ;
        RECT 79.480 173.560 79.770 173.605 ;
        RECT 75.810 173.420 79.770 173.560 ;
        RECT 75.810 173.375 76.100 173.420 ;
        RECT 77.380 173.375 77.670 173.420 ;
        RECT 79.480 173.375 79.770 173.420 ;
        RECT 86.890 173.560 87.180 173.605 ;
        RECT 88.990 173.560 89.280 173.605 ;
        RECT 90.560 173.560 90.850 173.605 ;
        RECT 86.890 173.420 90.850 173.560 ;
        RECT 86.890 173.375 87.180 173.420 ;
        RECT 88.990 173.375 89.280 173.420 ;
        RECT 90.560 173.375 90.850 173.420 ;
        RECT 108.510 173.560 108.800 173.605 ;
        RECT 110.610 173.560 110.900 173.605 ;
        RECT 112.180 173.560 112.470 173.605 ;
        RECT 133.310 173.560 133.630 173.620 ;
        RECT 108.510 173.420 112.470 173.560 ;
        RECT 108.510 173.375 108.800 173.420 ;
        RECT 110.610 173.375 110.900 173.420 ;
        RECT 112.180 173.375 112.470 173.420 ;
        RECT 131.560 173.420 133.630 173.560 ;
        RECT 70.765 173.080 73.280 173.220 ;
        RECT 75.375 173.220 75.665 173.265 ;
        RECT 77.895 173.220 78.185 173.265 ;
        RECT 79.085 173.220 79.375 173.265 ;
        RECT 75.375 173.080 79.375 173.220 ;
        RECT 66.700 172.940 66.840 173.080 ;
        RECT 70.765 173.035 71.055 173.080 ;
        RECT 75.375 173.035 75.665 173.080 ;
        RECT 77.895 173.035 78.185 173.080 ;
        RECT 79.085 173.035 79.375 173.080 ;
        RECT 87.285 173.220 87.575 173.265 ;
        RECT 88.475 173.220 88.765 173.265 ;
        RECT 90.995 173.220 91.285 173.265 ;
        RECT 87.285 173.080 91.285 173.220 ;
        RECT 87.285 173.035 87.575 173.080 ;
        RECT 88.475 173.035 88.765 173.080 ;
        RECT 90.995 173.035 91.285 173.080 ;
        RECT 96.050 173.020 96.370 173.280 ;
        RECT 96.985 173.220 97.275 173.265 ;
        RECT 98.350 173.220 98.670 173.280 ;
        RECT 101.110 173.220 101.430 173.280 ;
        RECT 96.985 173.080 101.430 173.220 ;
        RECT 96.985 173.035 97.275 173.080 ;
        RECT 98.350 173.020 98.670 173.080 ;
        RECT 101.110 173.020 101.430 173.080 ;
        RECT 102.950 173.020 103.270 173.280 ;
        RECT 103.885 173.220 104.175 173.265 ;
        RECT 103.885 173.080 107.780 173.220 ;
        RECT 103.885 173.035 104.175 173.080 ;
        RECT 44.545 172.880 44.835 172.925 ;
        RECT 42.245 172.740 44.835 172.880 ;
        RECT 42.245 172.695 42.535 172.740 ;
        RECT 43.150 172.680 43.470 172.740 ;
        RECT 44.545 172.695 44.835 172.740 ;
        RECT 45.465 172.880 45.755 172.925 ;
        RECT 48.210 172.880 48.530 172.940 ;
        RECT 45.465 172.740 48.530 172.880 ;
        RECT 45.465 172.695 45.755 172.740 ;
        RECT 48.210 172.680 48.530 172.740 ;
        RECT 52.810 172.880 53.130 172.940 ;
        RECT 53.285 172.880 53.575 172.925 ;
        RECT 66.610 172.880 66.930 172.940 ;
        RECT 52.810 172.740 53.575 172.880 ;
        RECT 52.810 172.680 53.130 172.740 ;
        RECT 53.285 172.695 53.575 172.740 ;
        RECT 65.780 172.740 66.930 172.880 ;
        RECT 27.680 172.540 27.970 172.585 ;
        RECT 29.350 172.540 29.670 172.600 ;
        RECT 27.680 172.400 29.670 172.540 ;
        RECT 27.680 172.355 27.970 172.400 ;
        RECT 29.350 172.340 29.670 172.400 ;
        RECT 43.610 172.540 43.930 172.600 ;
        RECT 51.890 172.585 52.210 172.600 ;
        RECT 44.085 172.540 44.375 172.585 ;
        RECT 43.610 172.400 44.375 172.540 ;
        RECT 43.610 172.340 43.930 172.400 ;
        RECT 44.085 172.355 44.375 172.400 ;
        RECT 51.890 172.355 52.240 172.585 ;
        RECT 61.090 172.540 61.410 172.600 ;
        RECT 65.085 172.540 65.375 172.585 ;
        RECT 65.780 172.540 65.920 172.740 ;
        RECT 66.610 172.680 66.930 172.740 ;
        RECT 68.450 172.680 68.770 172.940 ;
        RECT 69.385 172.695 69.675 172.925 ;
        RECT 71.685 172.880 71.975 172.925 ;
        RECT 72.590 172.880 72.910 172.940 ;
        RECT 71.685 172.740 72.910 172.880 ;
        RECT 71.685 172.695 71.975 172.740 ;
        RECT 61.090 172.400 65.920 172.540 ;
        RECT 66.150 172.540 66.470 172.600 ;
        RECT 67.085 172.540 67.375 172.585 ;
        RECT 66.150 172.400 67.375 172.540 ;
        RECT 51.890 172.340 52.210 172.355 ;
        RECT 61.090 172.340 61.410 172.400 ;
        RECT 65.085 172.355 65.375 172.400 ;
        RECT 66.150 172.340 66.470 172.400 ;
        RECT 67.085 172.355 67.375 172.400 ;
        RECT 67.990 172.340 68.310 172.600 ;
        RECT 69.460 172.540 69.600 172.695 ;
        RECT 72.590 172.680 72.910 172.740 ;
        RECT 79.965 172.880 80.255 172.925 ;
        RECT 83.630 172.880 83.950 172.940 ;
        RECT 86.390 172.880 86.710 172.940 ;
        RECT 79.965 172.740 86.710 172.880 ;
        RECT 79.965 172.695 80.255 172.740 ;
        RECT 83.630 172.680 83.950 172.740 ;
        RECT 86.390 172.680 86.710 172.740 ;
        RECT 105.710 172.680 106.030 172.940 ;
        RECT 106.630 172.680 106.950 172.940 ;
        RECT 107.640 172.880 107.780 173.080 ;
        RECT 108.010 173.020 108.330 173.280 ;
        RECT 108.905 173.220 109.195 173.265 ;
        RECT 110.095 173.220 110.385 173.265 ;
        RECT 112.615 173.220 112.905 173.265 ;
        RECT 108.905 173.080 112.905 173.220 ;
        RECT 108.905 173.035 109.195 173.080 ;
        RECT 110.095 173.035 110.385 173.080 ;
        RECT 112.615 173.035 112.905 173.080 ;
        RECT 114.450 172.880 114.770 172.940 ;
        RECT 107.640 172.740 114.770 172.880 ;
        RECT 114.450 172.680 114.770 172.740 ;
        RECT 123.205 172.695 123.495 172.925 ;
        RECT 123.650 172.880 123.970 172.940 ;
        RECT 124.125 172.880 124.415 172.925 ;
        RECT 123.650 172.740 124.415 172.880 ;
        RECT 68.540 172.400 69.600 172.540 ;
        RECT 74.430 172.540 74.750 172.600 ;
        RECT 78.630 172.540 78.920 172.585 ;
        RECT 74.430 172.400 78.920 172.540 ;
        RECT 40.390 172.000 40.710 172.260 ;
        RECT 40.865 172.200 41.155 172.245 ;
        RECT 41.310 172.200 41.630 172.260 ;
        RECT 40.865 172.060 41.630 172.200 ;
        RECT 40.865 172.015 41.155 172.060 ;
        RECT 41.310 172.000 41.630 172.060 ;
        RECT 63.390 172.200 63.710 172.260 ;
        RECT 64.325 172.200 64.615 172.245 ;
        RECT 63.390 172.060 64.615 172.200 ;
        RECT 63.390 172.000 63.710 172.060 ;
        RECT 64.325 172.015 64.615 172.060 ;
        RECT 67.530 172.200 67.850 172.260 ;
        RECT 68.540 172.200 68.680 172.400 ;
        RECT 74.430 172.340 74.750 172.400 ;
        RECT 78.630 172.355 78.920 172.400 ;
        RECT 87.740 172.540 88.030 172.585 ;
        RECT 106.185 172.540 106.475 172.585 ;
        RECT 109.250 172.540 109.540 172.585 ;
        RECT 87.740 172.400 93.980 172.540 ;
        RECT 87.740 172.355 88.030 172.400 ;
        RECT 67.530 172.060 68.680 172.200 ;
        RECT 67.530 172.000 67.850 172.060 ;
        RECT 68.910 172.000 69.230 172.260 ;
        RECT 93.840 172.245 93.980 172.400 ;
        RECT 106.185 172.400 109.540 172.540 ;
        RECT 123.280 172.540 123.420 172.695 ;
        RECT 123.650 172.680 123.970 172.740 ;
        RECT 124.125 172.695 124.415 172.740 ;
        RECT 128.250 172.880 128.570 172.940 ;
        RECT 131.560 172.925 131.700 173.420 ;
        RECT 133.310 173.360 133.630 173.420 ;
        RECT 135.085 173.220 135.225 173.760 ;
        RECT 136.070 173.560 136.390 173.620 ;
        RECT 136.070 173.420 136.760 173.560 ;
        RECT 136.070 173.360 136.390 173.420 ;
        RECT 134.780 173.080 135.225 173.220 ;
        RECT 130.565 172.880 130.855 172.925 ;
        RECT 128.250 172.740 130.855 172.880 ;
        RECT 128.250 172.680 128.570 172.740 ;
        RECT 130.565 172.695 130.855 172.740 ;
        RECT 131.485 172.695 131.775 172.925 ;
        RECT 131.930 172.680 132.250 172.940 ;
        RECT 132.865 172.880 133.155 172.925 ;
        RECT 133.310 172.880 133.630 172.940 ;
        RECT 132.865 172.740 133.630 172.880 ;
        RECT 132.865 172.695 133.155 172.740 ;
        RECT 133.310 172.680 133.630 172.740 ;
        RECT 133.770 172.680 134.090 172.940 ;
        RECT 134.230 172.880 134.550 172.940 ;
        RECT 134.780 172.925 134.920 173.080 ;
        RECT 134.705 172.880 134.995 172.925 ;
        RECT 134.230 172.740 134.995 172.880 ;
        RECT 134.230 172.680 134.550 172.740 ;
        RECT 134.705 172.695 134.995 172.740 ;
        RECT 135.610 172.880 135.930 172.940 ;
        RECT 136.085 172.880 136.375 172.925 ;
        RECT 135.610 172.740 136.375 172.880 ;
        RECT 136.620 172.880 136.760 173.420 ;
        RECT 137.080 173.220 137.220 173.760 ;
        RECT 138.830 173.700 139.150 173.960 ;
        RECT 137.910 173.560 138.230 173.620 ;
        RECT 137.910 173.420 140.440 173.560 ;
        RECT 137.910 173.360 138.230 173.420 ;
        RECT 139.765 173.220 140.055 173.265 ;
        RECT 137.080 173.080 140.055 173.220 ;
        RECT 139.765 173.035 140.055 173.080 ;
        RECT 140.300 173.220 140.440 173.420 ;
        RECT 141.145 173.220 141.435 173.265 ;
        RECT 140.300 173.080 141.435 173.220 ;
        RECT 137.465 172.880 137.755 172.925 ;
        RECT 136.620 172.740 137.755 172.880 ;
        RECT 135.610 172.680 135.930 172.740 ;
        RECT 136.085 172.695 136.375 172.740 ;
        RECT 137.465 172.695 137.755 172.740 ;
        RECT 125.490 172.540 125.810 172.600 ;
        RECT 132.405 172.540 132.695 172.585 ;
        RECT 137.005 172.540 137.295 172.585 ;
        RECT 123.280 172.400 131.700 172.540 ;
        RECT 106.185 172.355 106.475 172.400 ;
        RECT 109.250 172.355 109.540 172.400 ;
        RECT 125.490 172.340 125.810 172.400 ;
        RECT 93.765 172.015 94.055 172.245 ;
        RECT 95.590 172.000 95.910 172.260 ;
        RECT 96.050 172.200 96.370 172.260 ;
        RECT 100.665 172.200 100.955 172.245 ;
        RECT 96.050 172.060 100.955 172.200 ;
        RECT 96.050 172.000 96.370 172.060 ;
        RECT 100.665 172.015 100.955 172.060 ;
        RECT 102.505 172.200 102.795 172.245 ;
        RECT 113.990 172.200 114.310 172.260 ;
        RECT 102.505 172.060 114.310 172.200 ;
        RECT 102.505 172.015 102.795 172.060 ;
        RECT 113.990 172.000 114.310 172.060 ;
        RECT 124.110 172.200 124.430 172.260 ;
        RECT 126.410 172.200 126.730 172.260 ;
        RECT 128.250 172.200 128.570 172.260 ;
        RECT 124.110 172.060 128.570 172.200 ;
        RECT 124.110 172.000 124.430 172.060 ;
        RECT 126.410 172.000 126.730 172.060 ;
        RECT 128.250 172.000 128.570 172.060 ;
        RECT 128.710 172.200 129.030 172.260 ;
        RECT 131.025 172.200 131.315 172.245 ;
        RECT 128.710 172.060 131.315 172.200 ;
        RECT 131.560 172.200 131.700 172.400 ;
        RECT 132.405 172.400 137.295 172.540 ;
        RECT 137.540 172.540 137.680 172.695 ;
        RECT 137.910 172.680 138.230 172.940 ;
        RECT 140.300 172.925 140.440 173.080 ;
        RECT 141.145 173.035 141.435 173.080 ;
        RECT 140.225 172.695 140.515 172.925 ;
        RECT 140.670 172.680 140.990 172.940 ;
        RECT 141.605 172.695 141.895 172.925 ;
        RECT 138.370 172.540 138.690 172.600 ;
        RECT 141.680 172.540 141.820 172.695 ;
        RECT 137.540 172.400 141.820 172.540 ;
        RECT 132.405 172.355 132.695 172.400 ;
        RECT 137.005 172.355 137.295 172.400 ;
        RECT 138.370 172.340 138.690 172.400 ;
        RECT 132.850 172.200 133.170 172.260 ;
        RECT 131.560 172.060 133.170 172.200 ;
        RECT 128.710 172.000 129.030 172.060 ;
        RECT 131.025 172.015 131.315 172.060 ;
        RECT 132.850 172.000 133.170 172.060 ;
        RECT 17.320 171.380 147.040 171.860 ;
        RECT 37.170 170.980 37.490 171.240 ;
        RECT 38.090 170.980 38.410 171.240 ;
        RECT 39.930 171.180 40.250 171.240 ;
        RECT 40.405 171.180 40.695 171.225 ;
        RECT 39.930 171.040 40.695 171.180 ;
        RECT 39.930 170.980 40.250 171.040 ;
        RECT 40.405 170.995 40.695 171.040 ;
        RECT 43.610 170.980 43.930 171.240 ;
        RECT 51.890 171.180 52.210 171.240 ;
        RECT 52.365 171.180 52.655 171.225 ;
        RECT 51.890 171.040 52.655 171.180 ;
        RECT 51.890 170.980 52.210 171.040 ;
        RECT 52.365 170.995 52.655 171.040 ;
        RECT 56.950 171.180 57.270 171.240 ;
        RECT 67.530 171.180 67.850 171.240 ;
        RECT 56.950 171.040 67.850 171.180 ;
        RECT 56.950 170.980 57.270 171.040 ;
        RECT 67.530 170.980 67.850 171.040 ;
        RECT 67.990 171.180 68.310 171.240 ;
        RECT 69.385 171.180 69.675 171.225 ;
        RECT 78.110 171.180 78.430 171.240 ;
        RECT 67.990 171.040 69.675 171.180 ;
        RECT 67.990 170.980 68.310 171.040 ;
        RECT 69.385 170.995 69.675 171.040 ;
        RECT 74.520 171.040 78.430 171.180 ;
        RECT 39.485 170.840 39.775 170.885 ;
        RECT 66.150 170.840 66.470 170.900 ;
        RECT 37.720 170.700 39.775 170.840 ;
        RECT 34.870 170.300 35.190 170.560 ;
        RECT 36.250 170.500 36.570 170.560 ;
        RECT 37.200 170.500 37.490 170.545 ;
        RECT 37.720 170.500 37.860 170.700 ;
        RECT 39.485 170.655 39.775 170.700 ;
        RECT 60.720 170.700 66.470 170.840 ;
        RECT 67.620 170.840 67.760 170.980 ;
        RECT 73.065 170.840 73.355 170.885 ;
        RECT 73.510 170.840 73.830 170.900 ;
        RECT 67.620 170.700 73.830 170.840 ;
        RECT 36.250 170.360 37.860 170.500 ;
        RECT 36.250 170.300 36.570 170.360 ;
        RECT 37.200 170.315 37.490 170.360 ;
        RECT 38.550 170.300 38.870 170.560 ;
        RECT 40.390 170.500 40.710 170.560 ;
        RECT 45.005 170.500 45.295 170.545 ;
        RECT 40.390 170.360 45.295 170.500 ;
        RECT 40.390 170.300 40.710 170.360 ;
        RECT 45.005 170.315 45.295 170.360 ;
        RECT 48.210 170.300 48.530 170.560 ;
        RECT 51.445 170.500 51.735 170.545 ;
        RECT 50.140 170.360 51.735 170.500 ;
        RECT 44.530 169.960 44.850 170.220 ;
        RECT 45.450 170.160 45.770 170.220 ;
        RECT 46.385 170.160 46.675 170.205 ;
        RECT 45.450 170.020 46.675 170.160 ;
        RECT 45.450 169.960 45.770 170.020 ;
        RECT 46.385 169.975 46.675 170.020 ;
        RECT 46.830 169.960 47.150 170.220 ;
        RECT 48.670 169.960 48.990 170.220 ;
        RECT 50.140 170.205 50.280 170.360 ;
        RECT 51.445 170.315 51.735 170.360 ;
        RECT 58.330 170.300 58.650 170.560 ;
        RECT 60.720 170.545 60.860 170.700 ;
        RECT 66.150 170.640 66.470 170.700 ;
        RECT 73.065 170.655 73.355 170.700 ;
        RECT 73.510 170.640 73.830 170.700 ;
        RECT 60.645 170.315 60.935 170.545 ;
        RECT 62.945 170.500 63.235 170.545 ;
        RECT 65.245 170.500 65.535 170.545 ;
        RECT 62.945 170.360 65.535 170.500 ;
        RECT 62.945 170.315 63.235 170.360 ;
        RECT 65.245 170.315 65.535 170.360 ;
        RECT 66.610 170.500 66.930 170.560 ;
        RECT 74.520 170.545 74.660 171.040 ;
        RECT 78.110 170.980 78.430 171.040 ;
        RECT 94.670 171.180 94.990 171.240 ;
        RECT 95.145 171.180 95.435 171.225 ;
        RECT 94.670 171.040 95.435 171.180 ;
        RECT 94.670 170.980 94.990 171.040 ;
        RECT 95.145 170.995 95.435 171.040 ;
        RECT 97.430 170.980 97.750 171.240 ;
        RECT 108.470 171.180 108.790 171.240 ;
        RECT 110.770 171.180 111.090 171.240 ;
        RECT 114.910 171.180 115.230 171.240 ;
        RECT 108.470 171.040 109.465 171.180 ;
        RECT 108.470 170.980 108.790 171.040 ;
        RECT 83.630 170.840 83.950 170.900 ;
        RECT 109.325 170.885 109.465 171.040 ;
        RECT 110.770 171.040 115.230 171.180 ;
        RECT 110.770 170.980 111.090 171.040 ;
        RECT 114.910 170.980 115.230 171.040 ;
        RECT 126.410 171.180 126.730 171.240 ;
        RECT 129.170 171.180 129.490 171.240 ;
        RECT 126.410 171.040 127.100 171.180 ;
        RECT 126.410 170.980 126.730 171.040 ;
        RECT 77.740 170.700 83.950 170.840 ;
        RECT 77.740 170.545 77.880 170.700 ;
        RECT 83.630 170.640 83.950 170.700 ;
        RECT 109.250 170.655 109.540 170.885 ;
        RECT 126.960 170.840 127.100 171.040 ;
        RECT 127.880 171.040 129.490 171.180 ;
        RECT 127.345 170.840 127.635 170.885 ;
        RECT 126.960 170.700 127.635 170.840 ;
        RECT 127.345 170.655 127.635 170.700 ;
        RECT 66.610 170.370 73.970 170.500 ;
        RECT 66.610 170.360 74.200 170.370 ;
        RECT 66.610 170.300 66.930 170.360 ;
        RECT 73.830 170.230 74.200 170.360 ;
        RECT 74.445 170.315 74.735 170.545 ;
        RECT 77.665 170.315 77.955 170.545 ;
        RECT 78.110 170.500 78.430 170.560 ;
        RECT 78.945 170.500 79.235 170.545 ;
        RECT 78.110 170.360 79.235 170.500 ;
        RECT 78.110 170.300 78.430 170.360 ;
        RECT 78.945 170.315 79.235 170.360 ;
        RECT 96.970 170.300 97.290 170.560 ;
        RECT 100.650 170.500 100.970 170.560 ;
        RECT 101.125 170.500 101.415 170.545 ;
        RECT 100.650 170.360 101.415 170.500 ;
        RECT 100.650 170.300 100.970 170.360 ;
        RECT 101.125 170.315 101.415 170.360 ;
        RECT 105.265 170.500 105.555 170.545 ;
        RECT 108.010 170.500 108.330 170.560 ;
        RECT 105.265 170.360 108.330 170.500 ;
        RECT 105.265 170.315 105.555 170.360 ;
        RECT 108.010 170.300 108.330 170.360 ;
        RECT 115.370 170.500 115.690 170.560 ;
        RECT 117.670 170.500 117.990 170.560 ;
        RECT 118.145 170.500 118.435 170.545 ;
        RECT 115.370 170.360 118.435 170.500 ;
        RECT 115.370 170.300 115.690 170.360 ;
        RECT 117.670 170.300 117.990 170.360 ;
        RECT 118.145 170.315 118.435 170.360 ;
        RECT 118.590 170.300 118.910 170.560 ;
        RECT 126.410 170.300 126.730 170.560 ;
        RECT 127.880 170.545 128.020 171.040 ;
        RECT 129.170 170.980 129.490 171.040 ;
        RECT 129.630 171.180 129.950 171.240 ;
        RECT 133.310 171.180 133.630 171.240 ;
        RECT 136.085 171.180 136.375 171.225 ;
        RECT 129.630 171.040 132.160 171.180 ;
        RECT 129.630 170.980 129.950 171.040 ;
        RECT 130.550 170.840 130.870 170.900 ;
        RECT 128.800 170.700 130.870 170.840 ;
        RECT 127.805 170.315 128.095 170.545 ;
        RECT 128.250 170.300 128.570 170.560 ;
        RECT 50.065 169.975 50.355 170.205 ;
        RECT 50.510 169.960 50.830 170.220 ;
        RECT 56.950 169.960 57.270 170.220 ;
        RECT 61.090 169.960 61.410 170.220 ;
        RECT 63.390 169.960 63.710 170.220 ;
        RECT 65.690 170.160 66.010 170.220 ;
        RECT 68.005 170.160 68.295 170.205 ;
        RECT 72.145 170.160 72.435 170.205 ;
        RECT 65.690 170.020 68.295 170.160 ;
        RECT 65.690 169.960 66.010 170.020 ;
        RECT 68.005 169.975 68.295 170.020 ;
        RECT 69.000 170.020 72.435 170.160 ;
        RECT 57.885 169.820 58.175 169.865 ;
        RECT 63.480 169.820 63.620 169.960 ;
        RECT 57.885 169.680 63.620 169.820 ;
        RECT 64.785 169.820 65.075 169.865 ;
        RECT 68.450 169.820 68.770 169.880 ;
        RECT 64.785 169.680 68.770 169.820 ;
        RECT 57.885 169.635 58.175 169.680 ;
        RECT 64.785 169.635 65.075 169.680 ;
        RECT 68.450 169.620 68.770 169.680 ;
        RECT 35.345 169.480 35.635 169.525 ;
        RECT 39.010 169.480 39.330 169.540 ;
        RECT 45.910 169.480 46.230 169.540 ;
        RECT 53.270 169.480 53.590 169.540 ;
        RECT 35.345 169.340 53.590 169.480 ;
        RECT 35.345 169.295 35.635 169.340 ;
        RECT 39.010 169.280 39.330 169.340 ;
        RECT 45.910 169.280 46.230 169.340 ;
        RECT 53.270 169.280 53.590 169.340 ;
        RECT 58.330 169.280 58.650 169.540 ;
        RECT 58.790 169.480 59.110 169.540 ;
        RECT 59.265 169.480 59.555 169.525 ;
        RECT 58.790 169.340 59.555 169.480 ;
        RECT 58.790 169.280 59.110 169.340 ;
        RECT 59.265 169.295 59.555 169.340 ;
        RECT 65.230 169.480 65.550 169.540 ;
        RECT 69.000 169.480 69.140 170.020 ;
        RECT 72.145 169.975 72.435 170.020 ;
        RECT 74.060 169.865 74.200 170.230 ;
        RECT 78.545 170.160 78.835 170.205 ;
        RECT 79.735 170.160 80.025 170.205 ;
        RECT 82.255 170.160 82.545 170.205 ;
        RECT 78.545 170.020 82.545 170.160 ;
        RECT 78.545 169.975 78.835 170.020 ;
        RECT 79.735 169.975 80.025 170.020 ;
        RECT 82.255 169.975 82.545 170.020 ;
        RECT 98.350 169.960 98.670 170.220 ;
        RECT 108.905 170.160 109.195 170.205 ;
        RECT 110.095 170.160 110.385 170.205 ;
        RECT 112.615 170.160 112.905 170.205 ;
        RECT 108.905 170.020 112.905 170.160 ;
        RECT 108.905 169.975 109.195 170.020 ;
        RECT 110.095 169.975 110.385 170.020 ;
        RECT 112.615 169.975 112.905 170.020 ;
        RECT 73.985 169.635 74.275 169.865 ;
        RECT 74.430 169.620 74.750 169.880 ;
        RECT 78.150 169.820 78.440 169.865 ;
        RECT 80.250 169.820 80.540 169.865 ;
        RECT 81.820 169.820 82.110 169.865 ;
        RECT 78.150 169.680 82.110 169.820 ;
        RECT 78.150 169.635 78.440 169.680 ;
        RECT 80.250 169.635 80.540 169.680 ;
        RECT 81.820 169.635 82.110 169.680 ;
        RECT 108.510 169.820 108.800 169.865 ;
        RECT 110.610 169.820 110.900 169.865 ;
        RECT 112.180 169.820 112.470 169.865 ;
        RECT 115.460 169.820 115.600 170.300 ;
        RECT 116.305 169.975 116.595 170.205 ;
        RECT 119.525 170.160 119.815 170.205 ;
        RECT 128.800 170.160 128.940 170.700 ;
        RECT 130.550 170.640 130.870 170.700 ;
        RECT 129.245 170.315 129.535 170.545 ;
        RECT 119.525 170.020 128.940 170.160 ;
        RECT 129.260 170.160 129.400 170.315 ;
        RECT 131.470 170.160 131.790 170.220 ;
        RECT 129.260 170.020 131.790 170.160 ;
        RECT 119.525 169.975 119.815 170.020 ;
        RECT 108.510 169.680 112.470 169.820 ;
        RECT 108.510 169.635 108.800 169.680 ;
        RECT 110.610 169.635 110.900 169.680 ;
        RECT 112.180 169.635 112.470 169.680 ;
        RECT 112.700 169.680 115.600 169.820 ;
        RECT 116.380 169.820 116.520 169.975 ;
        RECT 130.180 169.880 130.320 170.020 ;
        RECT 131.470 169.960 131.790 170.020 ;
        RECT 118.130 169.820 118.450 169.880 ;
        RECT 116.380 169.680 118.450 169.820 ;
        RECT 65.230 169.340 69.140 169.480 ;
        RECT 65.230 169.280 65.550 169.340 ;
        RECT 84.550 169.280 84.870 169.540 ;
        RECT 107.090 169.480 107.410 169.540 ;
        RECT 112.700 169.480 112.840 169.680 ;
        RECT 118.130 169.620 118.450 169.680 ;
        RECT 126.425 169.820 126.715 169.865 ;
        RECT 129.630 169.820 129.950 169.880 ;
        RECT 126.425 169.680 129.950 169.820 ;
        RECT 126.425 169.635 126.715 169.680 ;
        RECT 129.630 169.620 129.950 169.680 ;
        RECT 130.090 169.620 130.410 169.880 ;
        RECT 107.090 169.340 112.840 169.480 ;
        RECT 128.265 169.480 128.555 169.525 ;
        RECT 131.010 169.480 131.330 169.540 ;
        RECT 128.265 169.340 131.330 169.480 ;
        RECT 131.560 169.480 131.700 169.960 ;
        RECT 132.020 169.820 132.160 171.040 ;
        RECT 133.310 171.040 136.375 171.180 ;
        RECT 133.310 170.980 133.630 171.040 ;
        RECT 136.085 170.995 136.375 171.040 ;
        RECT 143.890 170.840 144.210 170.900 ;
        RECT 137.080 170.700 144.210 170.840 ;
        RECT 132.405 170.315 132.695 170.545 ;
        RECT 132.850 170.500 133.170 170.560 ;
        RECT 133.325 170.500 133.615 170.545 ;
        RECT 132.850 170.360 133.615 170.500 ;
        RECT 132.480 170.160 132.620 170.315 ;
        RECT 132.850 170.300 133.170 170.360 ;
        RECT 133.325 170.315 133.615 170.360 ;
        RECT 133.770 170.300 134.090 170.560 ;
        RECT 134.230 170.300 134.550 170.560 ;
        RECT 134.690 170.300 135.010 170.560 ;
        RECT 137.080 170.545 137.220 170.700 ;
        RECT 143.890 170.640 144.210 170.700 ;
        RECT 137.005 170.315 137.295 170.545 ;
        RECT 138.370 170.300 138.690 170.560 ;
        RECT 139.305 170.500 139.595 170.545 ;
        RECT 140.670 170.500 140.990 170.560 ;
        RECT 139.195 170.360 140.990 170.500 ;
        RECT 139.305 170.315 139.595 170.360 ;
        RECT 133.860 170.160 134.000 170.300 ;
        RECT 135.150 170.160 135.470 170.220 ;
        RECT 137.925 170.160 138.215 170.205 ;
        RECT 139.380 170.160 139.520 170.315 ;
        RECT 140.670 170.300 140.990 170.360 ;
        RECT 132.480 170.020 133.080 170.160 ;
        RECT 133.860 170.020 134.875 170.160 ;
        RECT 132.940 169.880 133.080 170.020 ;
        RECT 132.390 169.820 132.710 169.880 ;
        RECT 132.020 169.680 132.710 169.820 ;
        RECT 132.390 169.620 132.710 169.680 ;
        RECT 132.850 169.620 133.170 169.880 ;
        RECT 134.735 169.820 134.875 170.020 ;
        RECT 135.150 170.020 139.520 170.160 ;
        RECT 135.150 169.960 135.470 170.020 ;
        RECT 137.925 169.975 138.215 170.020 ;
        RECT 136.990 169.820 137.310 169.880 ;
        RECT 138.385 169.820 138.675 169.865 ;
        RECT 134.735 169.680 138.675 169.820 ;
        RECT 136.990 169.620 137.310 169.680 ;
        RECT 138.385 169.635 138.675 169.680 ;
        RECT 135.150 169.480 135.470 169.540 ;
        RECT 131.560 169.340 135.470 169.480 ;
        RECT 107.090 169.280 107.410 169.340 ;
        RECT 128.265 169.295 128.555 169.340 ;
        RECT 131.010 169.280 131.330 169.340 ;
        RECT 135.150 169.280 135.470 169.340 ;
        RECT 135.610 169.280 135.930 169.540 ;
        RECT 17.320 168.660 147.040 169.140 ;
        RECT 34.885 168.460 35.175 168.505 ;
        RECT 36.250 168.460 36.570 168.520 ;
        RECT 34.885 168.320 36.570 168.460 ;
        RECT 34.885 168.275 35.175 168.320 ;
        RECT 36.250 168.260 36.570 168.320 ;
        RECT 36.725 168.460 37.015 168.505 ;
        RECT 37.170 168.460 37.490 168.520 ;
        RECT 36.725 168.320 37.490 168.460 ;
        RECT 36.725 168.275 37.015 168.320 ;
        RECT 37.170 168.260 37.490 168.320 ;
        RECT 39.470 168.460 39.790 168.520 ;
        RECT 43.625 168.460 43.915 168.505 ;
        RECT 39.470 168.320 43.915 168.460 ;
        RECT 39.470 168.260 39.790 168.320 ;
        RECT 43.625 168.275 43.915 168.320 ;
        RECT 44.530 168.460 44.850 168.520 ;
        RECT 45.925 168.460 46.215 168.505 ;
        RECT 44.530 168.320 46.215 168.460 ;
        RECT 44.530 168.260 44.850 168.320 ;
        RECT 45.925 168.275 46.215 168.320 ;
        RECT 47.305 168.460 47.595 168.505 ;
        RECT 47.750 168.460 48.070 168.520 ;
        RECT 47.305 168.320 48.070 168.460 ;
        RECT 47.305 168.275 47.595 168.320 ;
        RECT 47.750 168.260 48.070 168.320 ;
        RECT 48.225 168.460 48.515 168.505 ;
        RECT 48.670 168.460 48.990 168.520 ;
        RECT 48.225 168.320 48.990 168.460 ;
        RECT 48.225 168.275 48.515 168.320 ;
        RECT 48.670 168.260 48.990 168.320 ;
        RECT 65.690 168.260 66.010 168.520 ;
        RECT 95.130 168.460 95.450 168.520 ;
        RECT 93.380 168.320 95.450 168.460 ;
        RECT 29.350 168.120 29.670 168.180 ;
        RECT 33.505 168.120 33.795 168.165 ;
        RECT 38.550 168.120 38.870 168.180 ;
        RECT 46.830 168.120 47.150 168.180 ;
        RECT 49.145 168.120 49.435 168.165 ;
        RECT 27.600 167.980 33.260 168.120 ;
        RECT 27.600 167.825 27.740 167.980 ;
        RECT 29.350 167.920 29.670 167.980 ;
        RECT 27.525 167.595 27.815 167.825 ;
        RECT 33.120 167.780 33.260 167.980 ;
        RECT 33.505 167.980 38.870 168.120 ;
        RECT 33.505 167.935 33.795 167.980 ;
        RECT 38.550 167.920 38.870 167.980 ;
        RECT 41.860 167.980 46.140 168.120 ;
        RECT 34.425 167.780 34.715 167.825 ;
        RECT 33.120 167.640 34.715 167.780 ;
        RECT 24.765 167.440 25.055 167.485 ;
        RECT 24.765 167.300 25.900 167.440 ;
        RECT 24.765 167.255 25.055 167.300 ;
        RECT 25.760 167.145 25.900 167.300 ;
        RECT 26.590 167.240 26.910 167.500 ;
        RECT 30.745 167.255 31.035 167.485 ;
        RECT 32.585 167.410 32.875 167.485 ;
        RECT 33.120 167.410 33.260 167.640 ;
        RECT 34.425 167.595 34.715 167.640 ;
        RECT 34.885 167.595 35.175 167.825 ;
        RECT 33.950 167.440 34.270 167.500 ;
        RECT 34.960 167.440 35.100 167.595 ;
        RECT 36.265 167.440 36.555 167.485 ;
        RECT 32.585 167.270 33.260 167.410 ;
        RECT 33.580 167.300 34.270 167.440 ;
        RECT 32.585 167.255 32.875 167.270 ;
        RECT 25.685 167.100 25.975 167.145 ;
        RECT 27.510 167.100 27.830 167.160 ;
        RECT 25.685 166.960 27.830 167.100 ;
        RECT 25.685 166.915 25.975 166.960 ;
        RECT 27.510 166.900 27.830 166.960 ;
        RECT 21.070 166.760 21.390 166.820 ;
        RECT 24.305 166.760 24.595 166.805 ;
        RECT 21.070 166.620 24.595 166.760 ;
        RECT 21.070 166.560 21.390 166.620 ;
        RECT 24.305 166.575 24.595 166.620 ;
        RECT 28.890 166.760 29.210 166.820 ;
        RECT 30.820 166.760 30.960 167.255 ;
        RECT 31.650 166.900 31.970 167.160 ;
        RECT 32.125 167.100 32.415 167.145 ;
        RECT 33.580 167.100 33.720 167.300 ;
        RECT 33.950 167.240 34.270 167.300 ;
        RECT 34.500 167.300 36.555 167.440 ;
        RECT 32.125 166.960 33.720 167.100 ;
        RECT 32.125 166.915 32.415 166.960 ;
        RECT 34.500 166.760 34.640 167.300 ;
        RECT 36.265 167.255 36.555 167.300 ;
        RECT 37.185 167.440 37.475 167.485 ;
        RECT 41.860 167.440 42.000 167.980 ;
        RECT 44.545 167.780 44.835 167.825 ;
        RECT 45.450 167.780 45.770 167.840 ;
        RECT 44.545 167.640 45.770 167.780 ;
        RECT 46.000 167.780 46.140 167.980 ;
        RECT 46.830 167.980 49.435 168.120 ;
        RECT 46.830 167.920 47.150 167.980 ;
        RECT 49.145 167.935 49.435 167.980 ;
        RECT 58.830 168.120 59.120 168.165 ;
        RECT 60.930 168.120 61.220 168.165 ;
        RECT 62.500 168.120 62.790 168.165 ;
        RECT 58.830 167.980 62.790 168.120 ;
        RECT 58.830 167.935 59.120 167.980 ;
        RECT 60.930 167.935 61.220 167.980 ;
        RECT 62.500 167.935 62.790 167.980 ;
        RECT 65.245 168.120 65.535 168.165 ;
        RECT 66.150 168.120 66.470 168.180 ;
        RECT 65.245 167.980 66.470 168.120 ;
        RECT 65.245 167.935 65.535 167.980 ;
        RECT 66.150 167.920 66.470 167.980 ;
        RECT 68.450 168.120 68.740 168.165 ;
        RECT 70.020 168.120 70.310 168.165 ;
        RECT 72.120 168.120 72.410 168.165 ;
        RECT 68.450 167.980 72.410 168.120 ;
        RECT 68.450 167.935 68.740 167.980 ;
        RECT 70.020 167.935 70.310 167.980 ;
        RECT 72.120 167.935 72.410 167.980 ;
        RECT 52.350 167.780 52.670 167.840 ;
        RECT 46.000 167.640 52.670 167.780 ;
        RECT 44.545 167.595 44.835 167.640 ;
        RECT 45.450 167.580 45.770 167.640 ;
        RECT 52.350 167.580 52.670 167.640 ;
        RECT 55.570 167.780 55.890 167.840 ;
        RECT 58.345 167.780 58.635 167.825 ;
        RECT 55.570 167.640 58.635 167.780 ;
        RECT 55.570 167.580 55.890 167.640 ;
        RECT 58.345 167.595 58.635 167.640 ;
        RECT 59.225 167.780 59.515 167.825 ;
        RECT 60.415 167.780 60.705 167.825 ;
        RECT 62.935 167.780 63.225 167.825 ;
        RECT 59.225 167.640 63.225 167.780 ;
        RECT 59.225 167.595 59.515 167.640 ;
        RECT 60.415 167.595 60.705 167.640 ;
        RECT 62.935 167.595 63.225 167.640 ;
        RECT 68.015 167.780 68.305 167.825 ;
        RECT 70.535 167.780 70.825 167.825 ;
        RECT 71.725 167.780 72.015 167.825 ;
        RECT 68.015 167.640 72.015 167.780 ;
        RECT 68.015 167.595 68.305 167.640 ;
        RECT 70.535 167.595 70.825 167.640 ;
        RECT 71.725 167.595 72.015 167.640 ;
        RECT 72.605 167.780 72.895 167.825 ;
        RECT 83.630 167.780 83.950 167.840 ;
        RECT 72.605 167.640 83.950 167.780 ;
        RECT 72.605 167.595 72.895 167.640 ;
        RECT 83.630 167.580 83.950 167.640 ;
        RECT 85.010 167.580 85.330 167.840 ;
        RECT 93.380 167.825 93.520 168.320 ;
        RECT 95.130 168.260 95.450 168.320 ;
        RECT 96.970 168.460 97.290 168.520 ;
        RECT 100.665 168.460 100.955 168.505 ;
        RECT 96.970 168.320 100.955 168.460 ;
        RECT 96.970 168.260 97.290 168.320 ;
        RECT 100.665 168.275 100.955 168.320 ;
        RECT 106.630 168.460 106.950 168.520 ;
        RECT 107.105 168.460 107.395 168.505 ;
        RECT 106.630 168.320 107.395 168.460 ;
        RECT 106.630 168.260 106.950 168.320 ;
        RECT 107.105 168.275 107.395 168.320 ;
        RECT 107.550 168.260 107.870 168.520 ;
        RECT 108.485 168.460 108.775 168.505 ;
        RECT 111.230 168.460 111.550 168.520 ;
        RECT 114.925 168.460 115.215 168.505 ;
        RECT 119.510 168.460 119.830 168.520 ;
        RECT 108.485 168.320 111.550 168.460 ;
        RECT 108.485 168.275 108.775 168.320 ;
        RECT 93.790 168.120 94.080 168.165 ;
        RECT 95.890 168.120 96.180 168.165 ;
        RECT 97.460 168.120 97.750 168.165 ;
        RECT 93.790 167.980 97.750 168.120 ;
        RECT 93.790 167.935 94.080 167.980 ;
        RECT 95.890 167.935 96.180 167.980 ;
        RECT 97.460 167.935 97.750 167.980 ;
        RECT 93.305 167.595 93.595 167.825 ;
        RECT 94.185 167.780 94.475 167.825 ;
        RECT 95.375 167.780 95.665 167.825 ;
        RECT 97.895 167.780 98.185 167.825 ;
        RECT 94.185 167.640 98.185 167.780 ;
        RECT 94.185 167.595 94.475 167.640 ;
        RECT 95.375 167.595 95.665 167.640 ;
        RECT 97.895 167.595 98.185 167.640 ;
        RECT 103.870 167.780 104.190 167.840 ;
        RECT 103.870 167.640 106.860 167.780 ;
        RECT 103.870 167.580 104.190 167.640 ;
        RECT 37.185 167.300 42.000 167.440 ;
        RECT 45.005 167.440 45.295 167.485 ;
        RECT 47.750 167.440 48.070 167.500 ;
        RECT 48.685 167.440 48.975 167.485 ;
        RECT 45.005 167.300 48.975 167.440 ;
        RECT 37.185 167.255 37.475 167.300 ;
        RECT 45.005 167.255 45.295 167.300 ;
        RECT 35.330 167.100 35.650 167.160 ;
        RECT 35.805 167.100 36.095 167.145 ;
        RECT 37.260 167.100 37.400 167.255 ;
        RECT 47.750 167.240 48.070 167.300 ;
        RECT 48.685 167.255 48.975 167.300 ;
        RECT 50.510 167.440 50.830 167.500 ;
        RECT 53.285 167.440 53.575 167.485 ;
        RECT 50.510 167.300 53.575 167.440 ;
        RECT 50.510 167.240 50.830 167.300 ;
        RECT 53.285 167.255 53.575 167.300 ;
        RECT 56.950 167.240 57.270 167.500 ;
        RECT 57.885 167.440 58.175 167.485 ;
        RECT 58.790 167.440 59.110 167.500 ;
        RECT 57.885 167.300 59.110 167.440 ;
        RECT 57.885 167.255 58.175 167.300 ;
        RECT 58.790 167.240 59.110 167.300 ;
        RECT 68.910 167.440 69.230 167.500 ;
        RECT 71.270 167.440 71.560 167.485 ;
        RECT 68.910 167.300 71.560 167.440 ;
        RECT 68.910 167.240 69.230 167.300 ;
        RECT 71.270 167.255 71.560 167.300 ;
        RECT 94.640 167.440 94.930 167.485 ;
        RECT 96.050 167.440 96.370 167.500 ;
        RECT 94.640 167.300 96.370 167.440 ;
        RECT 94.640 167.255 94.930 167.300 ;
        RECT 96.050 167.240 96.370 167.300 ;
        RECT 99.730 167.440 100.050 167.500 ;
        RECT 105.250 167.440 105.570 167.500 ;
        RECT 105.725 167.440 106.015 167.485 ;
        RECT 99.730 167.300 106.015 167.440 ;
        RECT 99.730 167.240 100.050 167.300 ;
        RECT 105.250 167.240 105.570 167.300 ;
        RECT 105.725 167.255 106.015 167.300 ;
        RECT 35.330 166.960 37.400 167.100 ;
        RECT 35.330 166.900 35.650 166.960 ;
        RECT 35.805 166.915 36.095 166.960 ;
        RECT 43.610 166.900 43.930 167.160 ;
        RECT 46.385 167.100 46.675 167.145 ;
        RECT 45.080 166.960 46.675 167.100 ;
        RECT 45.080 166.820 45.220 166.960 ;
        RECT 46.385 166.915 46.675 166.960 ;
        RECT 57.425 167.100 57.715 167.145 ;
        RECT 59.570 167.100 59.860 167.145 ;
        RECT 102.505 167.100 102.795 167.145 ;
        RECT 103.410 167.100 103.730 167.160 ;
        RECT 57.425 166.960 59.860 167.100 ;
        RECT 57.425 166.915 57.715 166.960 ;
        RECT 59.570 166.915 59.860 166.960 ;
        RECT 64.860 166.960 73.970 167.100 ;
        RECT 28.890 166.620 34.640 166.760 ;
        RECT 28.890 166.560 29.210 166.620 ;
        RECT 44.990 166.560 45.310 166.820 ;
        RECT 47.290 166.805 47.610 166.820 ;
        RECT 47.290 166.575 47.675 166.805 ;
        RECT 53.745 166.760 54.035 166.805 ;
        RECT 64.860 166.760 65.000 166.960 ;
        RECT 53.745 166.620 65.000 166.760 ;
        RECT 73.830 166.760 73.970 166.960 ;
        RECT 102.505 166.960 103.730 167.100 ;
        RECT 106.720 167.100 106.860 167.640 ;
        RECT 107.155 167.440 107.445 167.485 ;
        RECT 107.640 167.440 107.780 168.260 ;
        RECT 108.010 168.120 108.330 168.180 ;
        RECT 108.560 168.120 108.700 168.275 ;
        RECT 111.230 168.260 111.550 168.320 ;
        RECT 111.780 168.320 115.215 168.460 ;
        RECT 108.010 167.980 108.700 168.120 ;
        RECT 108.010 167.920 108.330 167.980 ;
        RECT 108.470 167.780 108.790 167.840 ;
        RECT 111.780 167.780 111.920 168.320 ;
        RECT 114.925 168.275 115.215 168.320 ;
        RECT 115.460 168.320 119.830 168.460 ;
        RECT 113.990 167.920 114.310 168.180 ;
        RECT 108.100 167.640 111.920 167.780 ;
        RECT 108.100 167.485 108.240 167.640 ;
        RECT 108.470 167.580 108.790 167.640 ;
        RECT 112.150 167.580 112.470 167.840 ;
        RECT 113.545 167.780 113.835 167.825 ;
        RECT 115.460 167.780 115.600 168.320 ;
        RECT 119.510 168.260 119.830 168.320 ;
        RECT 125.045 168.460 125.335 168.505 ;
        RECT 125.950 168.460 126.270 168.520 ;
        RECT 130.090 168.460 130.410 168.520 ;
        RECT 125.045 168.320 126.270 168.460 ;
        RECT 125.045 168.275 125.335 168.320 ;
        RECT 125.950 168.260 126.270 168.320 ;
        RECT 127.420 168.320 130.410 168.460 ;
        RECT 118.590 168.120 118.910 168.180 ;
        RECT 115.920 167.980 118.910 168.120 ;
        RECT 115.920 167.825 116.060 167.980 ;
        RECT 118.590 167.920 118.910 167.980 ;
        RECT 125.490 168.120 125.810 168.180 ;
        RECT 127.420 168.120 127.560 168.320 ;
        RECT 130.090 168.260 130.410 168.320 ;
        RECT 134.230 168.260 134.550 168.520 ;
        RECT 135.625 168.460 135.915 168.505 ;
        RECT 136.070 168.460 136.390 168.520 ;
        RECT 135.625 168.320 136.390 168.460 ;
        RECT 135.625 168.275 135.915 168.320 ;
        RECT 136.070 168.260 136.390 168.320 ;
        RECT 125.490 167.980 127.560 168.120 ;
        RECT 127.790 168.120 128.110 168.180 ;
        RECT 131.010 168.120 131.330 168.180 ;
        RECT 127.790 167.980 131.330 168.120 ;
        RECT 125.490 167.920 125.810 167.980 ;
        RECT 127.790 167.920 128.110 167.980 ;
        RECT 131.010 167.920 131.330 167.980 ;
        RECT 134.690 168.120 135.010 168.180 ;
        RECT 134.690 167.980 136.300 168.120 ;
        RECT 134.690 167.920 135.010 167.980 ;
        RECT 113.545 167.640 115.600 167.780 ;
        RECT 113.545 167.595 113.835 167.640 ;
        RECT 115.845 167.595 116.135 167.825 ;
        RECT 117.670 167.780 117.990 167.840 ;
        RECT 117.300 167.640 117.990 167.780 ;
        RECT 107.155 167.300 107.780 167.440 ;
        RECT 107.155 167.255 107.445 167.300 ;
        RECT 108.025 167.255 108.315 167.485 ;
        RECT 114.910 167.240 115.230 167.500 ;
        RECT 117.300 167.485 117.440 167.640 ;
        RECT 117.670 167.580 117.990 167.640 ;
        RECT 124.110 167.580 124.430 167.840 ;
        RECT 129.740 167.780 130.030 167.825 ;
        RECT 134.245 167.780 134.535 167.825 ;
        RECT 135.610 167.780 135.930 167.840 ;
        RECT 129.740 167.640 134.000 167.780 ;
        RECT 129.740 167.595 130.030 167.640 ;
        RECT 117.225 167.255 117.515 167.485 ;
        RECT 118.590 167.240 118.910 167.500 ;
        RECT 119.050 167.440 119.370 167.500 ;
        RECT 119.985 167.440 120.275 167.485 ;
        RECT 119.050 167.300 120.275 167.440 ;
        RECT 119.050 167.240 119.370 167.300 ;
        RECT 119.985 167.255 120.275 167.300 ;
        RECT 120.905 167.255 121.195 167.485 ;
        RECT 110.770 167.100 111.090 167.160 ;
        RECT 116.290 167.100 116.610 167.160 ;
        RECT 106.720 166.960 116.610 167.100 ;
        RECT 118.680 167.100 118.820 167.240 ;
        RECT 120.980 167.100 121.120 167.255 ;
        RECT 125.490 167.240 125.810 167.500 ;
        RECT 127.790 167.440 128.110 167.500 ;
        RECT 128.725 167.440 129.015 167.485 ;
        RECT 130.565 167.440 130.855 167.485 ;
        RECT 131.470 167.440 131.790 167.500 ;
        RECT 133.860 167.485 134.000 167.640 ;
        RECT 134.245 167.640 135.930 167.780 ;
        RECT 134.245 167.595 134.535 167.640 ;
        RECT 135.610 167.580 135.930 167.640 ;
        RECT 136.160 167.485 136.300 167.980 ;
        RECT 127.790 167.300 129.015 167.440 ;
        RECT 127.790 167.240 128.110 167.300 ;
        RECT 128.725 167.255 129.015 167.300 ;
        RECT 130.180 167.300 130.855 167.440 ;
        RECT 130.180 167.160 130.320 167.300 ;
        RECT 130.565 167.255 130.855 167.300 ;
        RECT 131.100 167.300 131.790 167.440 ;
        RECT 118.680 166.960 121.120 167.100 ;
        RECT 121.810 167.100 122.130 167.160 ;
        RECT 125.965 167.100 126.255 167.145 ;
        RECT 126.870 167.100 127.190 167.160 ;
        RECT 129.185 167.100 129.475 167.145 ;
        RECT 121.810 166.960 129.475 167.100 ;
        RECT 102.505 166.915 102.795 166.960 ;
        RECT 103.410 166.900 103.730 166.960 ;
        RECT 110.770 166.900 111.090 166.960 ;
        RECT 116.290 166.900 116.610 166.960 ;
        RECT 121.810 166.900 122.130 166.960 ;
        RECT 125.965 166.915 126.255 166.960 ;
        RECT 126.870 166.900 127.190 166.960 ;
        RECT 129.185 166.915 129.475 166.960 ;
        RECT 130.090 166.900 130.410 167.160 ;
        RECT 131.100 167.100 131.240 167.300 ;
        RECT 131.470 167.240 131.790 167.300 ;
        RECT 133.785 167.255 134.075 167.485 ;
        RECT 136.085 167.255 136.375 167.485 ;
        RECT 136.990 167.240 137.310 167.500 ;
        RECT 145.270 167.240 145.590 167.500 ;
        RECT 130.640 166.960 131.240 167.100 ;
        RECT 132.850 167.100 133.170 167.160 ;
        RECT 132.850 166.960 144.580 167.100 ;
        RECT 78.110 166.760 78.430 166.820 ;
        RECT 73.830 166.620 78.430 166.760 ;
        RECT 53.745 166.575 54.035 166.620 ;
        RECT 47.290 166.560 47.610 166.575 ;
        RECT 78.110 166.560 78.430 166.620 ;
        RECT 87.310 166.760 87.630 166.820 ;
        RECT 87.785 166.760 88.075 166.805 ;
        RECT 87.310 166.620 88.075 166.760 ;
        RECT 87.310 166.560 87.630 166.620 ;
        RECT 87.785 166.575 88.075 166.620 ;
        RECT 100.205 166.760 100.495 166.805 ;
        RECT 102.965 166.760 103.255 166.805 ;
        RECT 104.330 166.760 104.650 166.820 ;
        RECT 100.205 166.620 104.650 166.760 ;
        RECT 100.205 166.575 100.495 166.620 ;
        RECT 102.965 166.575 103.255 166.620 ;
        RECT 104.330 166.560 104.650 166.620 ;
        RECT 106.185 166.760 106.475 166.805 ;
        RECT 107.550 166.760 107.870 166.820 ;
        RECT 106.185 166.620 107.870 166.760 ;
        RECT 106.185 166.575 106.475 166.620 ;
        RECT 107.550 166.560 107.870 166.620 ;
        RECT 114.450 166.760 114.770 166.820 ;
        RECT 120.445 166.760 120.735 166.805 ;
        RECT 114.450 166.620 120.735 166.760 ;
        RECT 114.450 166.560 114.770 166.620 ;
        RECT 120.445 166.575 120.735 166.620 ;
        RECT 122.730 166.560 123.050 166.820 ;
        RECT 124.570 166.760 124.890 166.820 ;
        RECT 128.250 166.760 128.570 166.820 ;
        RECT 124.570 166.620 128.570 166.760 ;
        RECT 124.570 166.560 124.890 166.620 ;
        RECT 128.250 166.560 128.570 166.620 ;
        RECT 128.710 166.760 129.030 166.820 ;
        RECT 130.640 166.760 130.780 166.960 ;
        RECT 132.850 166.900 133.170 166.960 ;
        RECT 128.710 166.620 130.780 166.760 ;
        RECT 131.025 166.760 131.315 166.805 ;
        RECT 133.770 166.760 134.090 166.820 ;
        RECT 131.025 166.620 134.090 166.760 ;
        RECT 128.710 166.560 129.030 166.620 ;
        RECT 131.025 166.575 131.315 166.620 ;
        RECT 133.770 166.560 134.090 166.620 ;
        RECT 134.230 166.760 134.550 166.820 ;
        RECT 144.440 166.805 144.580 166.960 ;
        RECT 136.085 166.760 136.375 166.805 ;
        RECT 134.230 166.620 136.375 166.760 ;
        RECT 134.230 166.560 134.550 166.620 ;
        RECT 136.085 166.575 136.375 166.620 ;
        RECT 144.365 166.575 144.655 166.805 ;
        RECT 17.320 165.940 147.040 166.420 ;
        RECT 23.765 165.740 24.055 165.785 ;
        RECT 25.225 165.740 25.515 165.785 ;
        RECT 23.765 165.600 25.515 165.740 ;
        RECT 23.765 165.555 24.055 165.600 ;
        RECT 25.225 165.555 25.515 165.600 ;
        RECT 33.950 165.740 34.270 165.800 ;
        RECT 35.790 165.740 36.110 165.800 ;
        RECT 41.770 165.740 42.090 165.800 ;
        RECT 33.950 165.600 42.090 165.740 ;
        RECT 33.950 165.540 34.270 165.600 ;
        RECT 35.790 165.540 36.110 165.600 ;
        RECT 41.770 165.540 42.090 165.600 ;
        RECT 43.610 165.540 43.930 165.800 ;
        RECT 45.450 165.540 45.770 165.800 ;
        RECT 65.230 165.740 65.550 165.800 ;
        RECT 68.465 165.740 68.755 165.785 ;
        RECT 65.230 165.600 68.755 165.740 ;
        RECT 65.230 165.540 65.550 165.600 ;
        RECT 68.465 165.555 68.755 165.600 ;
        RECT 84.105 165.555 84.395 165.785 ;
        RECT 100.190 165.740 100.510 165.800 ;
        RECT 105.250 165.740 105.570 165.800 ;
        RECT 114.465 165.740 114.755 165.785 ;
        RECT 123.650 165.740 123.970 165.800 ;
        RECT 126.410 165.740 126.730 165.800 ;
        RECT 100.190 165.600 105.020 165.740 ;
        RECT 21.990 165.400 22.310 165.460 ;
        RECT 24.765 165.400 25.055 165.445 ;
        RECT 26.590 165.400 26.910 165.460 ;
        RECT 38.565 165.400 38.855 165.445 ;
        RECT 21.990 165.260 25.055 165.400 ;
        RECT 21.990 165.200 22.310 165.260 ;
        RECT 24.765 165.215 25.055 165.260 ;
        RECT 25.530 165.260 30.040 165.400 ;
        RECT 21.545 165.060 21.835 165.105 ;
        RECT 22.465 165.060 22.755 165.105 ;
        RECT 25.530 165.060 25.670 165.260 ;
        RECT 26.590 165.200 26.910 165.260 ;
        RECT 21.545 164.920 22.220 165.060 ;
        RECT 21.545 164.875 21.835 164.920 ;
        RECT 22.080 164.380 22.220 164.920 ;
        RECT 22.465 164.920 25.670 165.060 ;
        RECT 22.465 164.875 22.755 164.920 ;
        RECT 26.145 164.875 26.435 165.105 ;
        RECT 27.065 165.060 27.355 165.105 ;
        RECT 27.510 165.060 27.830 165.120 ;
        RECT 28.890 165.060 29.210 165.120 ;
        RECT 27.065 164.920 27.830 165.060 ;
        RECT 27.065 164.875 27.355 164.920 ;
        RECT 26.220 164.720 26.360 164.875 ;
        RECT 27.510 164.860 27.830 164.920 ;
        RECT 28.060 164.920 29.210 165.060 ;
        RECT 28.060 164.720 28.200 164.920 ;
        RECT 28.890 164.860 29.210 164.920 ;
        RECT 29.350 164.860 29.670 165.120 ;
        RECT 29.900 165.105 30.040 165.260 ;
        RECT 32.200 165.260 38.855 165.400 ;
        RECT 32.200 165.120 32.340 165.260 ;
        RECT 38.565 165.215 38.855 165.260 ;
        RECT 42.245 165.400 42.535 165.445 ;
        RECT 45.540 165.400 45.680 165.540 ;
        RECT 42.245 165.260 45.680 165.400 ;
        RECT 58.330 165.400 58.650 165.460 ;
        RECT 62.790 165.400 63.080 165.445 ;
        RECT 58.330 165.260 63.080 165.400 ;
        RECT 42.245 165.215 42.535 165.260 ;
        RECT 58.330 165.200 58.650 165.260 ;
        RECT 62.790 165.215 63.080 165.260 ;
        RECT 82.420 165.400 82.710 165.445 ;
        RECT 84.180 165.400 84.320 165.555 ;
        RECT 100.190 165.540 100.510 165.600 ;
        RECT 82.420 165.260 84.320 165.400 ;
        RECT 86.865 165.400 87.155 165.445 ;
        RECT 87.310 165.400 87.630 165.460 ;
        RECT 86.865 165.260 87.630 165.400 ;
        RECT 82.420 165.215 82.710 165.260 ;
        RECT 86.865 165.215 87.155 165.260 ;
        RECT 87.310 165.200 87.630 165.260 ;
        RECT 87.770 165.200 88.090 165.460 ;
        RECT 90.545 165.400 90.835 165.445 ;
        RECT 90.990 165.400 91.310 165.460 ;
        RECT 103.870 165.400 104.190 165.460 ;
        RECT 90.545 165.260 104.190 165.400 ;
        RECT 90.545 165.215 90.835 165.260 ;
        RECT 90.990 165.200 91.310 165.260 ;
        RECT 103.870 165.200 104.190 165.260 ;
        RECT 29.825 164.875 30.115 165.105 ;
        RECT 32.110 164.860 32.430 165.120 ;
        RECT 37.645 165.060 37.935 165.105 ;
        RECT 39.470 165.060 39.790 165.120 ;
        RECT 37.645 164.920 39.790 165.060 ;
        RECT 37.645 164.875 37.935 164.920 ;
        RECT 39.470 164.860 39.790 164.920 ;
        RECT 39.945 165.060 40.235 165.105 ;
        RECT 40.390 165.060 40.710 165.120 ;
        RECT 39.945 164.920 41.540 165.060 ;
        RECT 39.945 164.875 40.235 164.920 ;
        RECT 40.390 164.860 40.710 164.920 ;
        RECT 26.220 164.580 28.200 164.720 ;
        RECT 28.430 164.520 28.750 164.780 ;
        RECT 26.130 164.380 26.450 164.440 ;
        RECT 29.440 164.380 29.580 164.860 ;
        RECT 31.650 164.720 31.970 164.780 ;
        RECT 35.330 164.720 35.650 164.780 ;
        RECT 31.650 164.580 35.650 164.720 ;
        RECT 31.650 164.520 31.970 164.580 ;
        RECT 35.330 164.520 35.650 164.580 ;
        RECT 22.080 164.240 29.580 164.380 ;
        RECT 34.870 164.380 35.190 164.440 ;
        RECT 41.400 164.380 41.540 164.920 ;
        RECT 41.785 164.875 42.075 165.105 ;
        RECT 42.705 165.060 42.995 165.105 ;
        RECT 44.070 165.060 44.390 165.120 ;
        RECT 44.545 165.060 44.835 165.105 ;
        RECT 42.705 164.920 44.835 165.060 ;
        RECT 42.705 164.875 42.995 164.920 ;
        RECT 41.860 164.720 42.000 164.875 ;
        RECT 44.070 164.860 44.390 164.920 ;
        RECT 44.545 164.875 44.835 164.920 ;
        RECT 44.990 164.860 45.310 165.120 ;
        RECT 45.465 165.060 45.755 165.105 ;
        RECT 45.910 165.060 46.230 165.120 ;
        RECT 45.465 164.920 46.230 165.060 ;
        RECT 45.465 164.875 45.755 164.920 ;
        RECT 45.910 164.860 46.230 164.920 ;
        RECT 46.370 164.860 46.690 165.120 ;
        RECT 46.845 164.875 47.135 165.105 ;
        RECT 47.290 165.060 47.610 165.120 ;
        RECT 54.190 165.105 54.510 165.120 ;
        RECT 47.765 165.060 48.055 165.105 ;
        RECT 47.290 164.920 48.055 165.060 ;
        RECT 43.150 164.720 43.470 164.780 ;
        RECT 45.080 164.720 45.220 164.860 ;
        RECT 46.920 164.720 47.060 164.875 ;
        RECT 47.290 164.860 47.610 164.920 ;
        RECT 47.765 164.875 48.055 164.920 ;
        RECT 54.190 164.875 54.540 165.105 ;
        RECT 83.170 165.060 83.490 165.120 ;
        RECT 85.025 165.060 85.315 165.105 ;
        RECT 83.170 164.920 85.315 165.060 ;
        RECT 54.190 164.860 54.510 164.875 ;
        RECT 83.170 164.860 83.490 164.920 ;
        RECT 85.025 164.875 85.315 164.920 ;
        RECT 85.485 164.875 85.775 165.105 ;
        RECT 88.230 165.060 88.550 165.120 ;
        RECT 88.705 165.060 88.995 165.105 ;
        RECT 88.230 164.920 88.995 165.060 ;
        RECT 41.860 164.580 47.060 164.720 ;
        RECT 43.150 164.520 43.470 164.580 ;
        RECT 47.380 164.380 47.520 164.860 ;
        RECT 50.995 164.720 51.285 164.765 ;
        RECT 53.515 164.720 53.805 164.765 ;
        RECT 54.705 164.720 54.995 164.765 ;
        RECT 50.995 164.580 54.995 164.720 ;
        RECT 50.995 164.535 51.285 164.580 ;
        RECT 53.515 164.535 53.805 164.580 ;
        RECT 54.705 164.535 54.995 164.580 ;
        RECT 55.570 164.720 55.890 164.780 ;
        RECT 61.565 164.720 61.855 164.765 ;
        RECT 55.570 164.580 61.855 164.720 ;
        RECT 55.570 164.520 55.890 164.580 ;
        RECT 61.565 164.535 61.855 164.580 ;
        RECT 62.445 164.720 62.735 164.765 ;
        RECT 63.635 164.720 63.925 164.765 ;
        RECT 66.155 164.720 66.445 164.765 ;
        RECT 62.445 164.580 66.445 164.720 ;
        RECT 62.445 164.535 62.735 164.580 ;
        RECT 63.635 164.535 63.925 164.580 ;
        RECT 66.155 164.535 66.445 164.580 ;
        RECT 79.055 164.720 79.345 164.765 ;
        RECT 81.575 164.720 81.865 164.765 ;
        RECT 82.765 164.720 83.055 164.765 ;
        RECT 79.055 164.580 83.055 164.720 ;
        RECT 79.055 164.535 79.345 164.580 ;
        RECT 81.575 164.535 81.865 164.580 ;
        RECT 82.765 164.535 83.055 164.580 ;
        RECT 83.630 164.520 83.950 164.780 ;
        RECT 34.870 164.240 41.080 164.380 ;
        RECT 41.400 164.240 47.520 164.380 ;
        RECT 51.430 164.380 51.720 164.425 ;
        RECT 53.000 164.380 53.290 164.425 ;
        RECT 55.100 164.380 55.390 164.425 ;
        RECT 51.430 164.240 55.390 164.380 ;
        RECT 26.130 164.180 26.450 164.240 ;
        RECT 34.870 164.180 35.190 164.240 ;
        RECT 20.625 164.040 20.915 164.085 ;
        RECT 21.530 164.040 21.850 164.100 ;
        RECT 20.625 163.900 21.850 164.040 ;
        RECT 20.625 163.855 20.915 163.900 ;
        RECT 21.530 163.840 21.850 163.900 ;
        RECT 22.925 164.040 23.215 164.085 ;
        RECT 23.370 164.040 23.690 164.100 ;
        RECT 22.925 163.900 23.690 164.040 ;
        RECT 22.925 163.855 23.215 163.900 ;
        RECT 23.370 163.840 23.690 163.900 ;
        RECT 23.845 164.040 24.135 164.085 ;
        RECT 27.050 164.040 27.370 164.100 ;
        RECT 23.845 163.900 27.370 164.040 ;
        RECT 23.845 163.855 24.135 163.900 ;
        RECT 27.050 163.840 27.370 163.900 ;
        RECT 30.730 163.840 31.050 164.100 ;
        RECT 31.650 163.840 31.970 164.100 ;
        RECT 36.725 164.040 37.015 164.085 ;
        RECT 38.090 164.040 38.410 164.100 ;
        RECT 36.725 163.900 38.410 164.040 ;
        RECT 36.725 163.855 37.015 163.900 ;
        RECT 38.090 163.840 38.410 163.900 ;
        RECT 39.470 163.840 39.790 164.100 ;
        RECT 40.940 164.040 41.080 164.240 ;
        RECT 51.430 164.195 51.720 164.240 ;
        RECT 53.000 164.195 53.290 164.240 ;
        RECT 55.100 164.195 55.390 164.240 ;
        RECT 62.050 164.380 62.340 164.425 ;
        RECT 64.150 164.380 64.440 164.425 ;
        RECT 65.720 164.380 66.010 164.425 ;
        RECT 62.050 164.240 66.010 164.380 ;
        RECT 62.050 164.195 62.340 164.240 ;
        RECT 64.150 164.195 64.440 164.240 ;
        RECT 65.720 164.195 66.010 164.240 ;
        RECT 79.490 164.380 79.780 164.425 ;
        RECT 81.060 164.380 81.350 164.425 ;
        RECT 83.160 164.380 83.450 164.425 ;
        RECT 79.490 164.240 83.450 164.380 ;
        RECT 85.560 164.380 85.700 164.875 ;
        RECT 88.230 164.860 88.550 164.920 ;
        RECT 88.705 164.875 88.995 164.920 ;
        RECT 98.810 164.860 99.130 165.120 ;
        RECT 99.730 164.860 100.050 165.120 ;
        RECT 104.880 165.060 105.020 165.600 ;
        RECT 105.250 165.600 105.940 165.740 ;
        RECT 105.250 165.540 105.570 165.600 ;
        RECT 105.800 165.445 105.940 165.600 ;
        RECT 114.465 165.600 126.730 165.740 ;
        RECT 114.465 165.555 114.755 165.600 ;
        RECT 123.650 165.540 123.970 165.600 ;
        RECT 126.410 165.540 126.730 165.600 ;
        RECT 130.640 165.600 135.840 165.740 ;
        RECT 130.640 165.460 130.780 165.600 ;
        RECT 105.770 165.215 106.060 165.445 ;
        RECT 108.470 165.400 108.790 165.460 ;
        RECT 106.765 165.260 111.000 165.400 ;
        RECT 106.765 165.060 106.905 165.260 ;
        RECT 108.470 165.200 108.790 165.260 ;
        RECT 104.880 164.920 106.905 165.060 ;
        RECT 107.105 165.060 107.395 165.105 ;
        RECT 108.010 165.060 108.330 165.120 ;
        RECT 110.860 165.105 111.000 165.260 ;
        RECT 111.230 165.200 111.550 165.460 ;
        RECT 114.925 165.400 115.215 165.445 ;
        RECT 115.370 165.400 115.690 165.460 ;
        RECT 117.670 165.400 117.990 165.460 ;
        RECT 121.810 165.445 122.130 165.460 ;
        RECT 114.925 165.260 117.990 165.400 ;
        RECT 114.925 165.215 115.215 165.260 ;
        RECT 115.370 165.200 115.690 165.260 ;
        RECT 117.670 165.200 117.990 165.260 ;
        RECT 121.745 165.215 122.130 165.445 ;
        RECT 122.745 165.400 123.035 165.445 ;
        RECT 125.490 165.400 125.810 165.460 ;
        RECT 122.745 165.260 125.810 165.400 ;
        RECT 122.745 165.215 123.035 165.260 ;
        RECT 121.810 165.200 122.130 165.215 ;
        RECT 125.490 165.200 125.810 165.260 ;
        RECT 127.330 165.200 127.650 165.460 ;
        RECT 130.550 165.400 130.870 165.460 ;
        RECT 135.700 165.445 135.840 165.600 ;
        RECT 130.180 165.260 130.870 165.400 ;
        RECT 110.785 165.060 111.075 165.105 ;
        RECT 107.105 164.920 108.330 165.060 ;
        RECT 107.105 164.875 107.395 164.920 ;
        RECT 108.010 164.860 108.330 164.920 ;
        RECT 109.940 164.920 111.075 165.060 ;
        RECT 111.320 165.060 111.460 165.200 ;
        RECT 113.070 165.060 113.390 165.120 ;
        RECT 117.225 165.060 117.515 165.105 ;
        RECT 111.320 164.920 113.390 165.060 ;
        RECT 85.930 164.720 86.250 164.780 ;
        RECT 87.325 164.720 87.615 164.765 ;
        RECT 85.930 164.580 87.615 164.720 ;
        RECT 85.930 164.520 86.250 164.580 ;
        RECT 87.325 164.535 87.615 164.580 ;
        RECT 102.515 164.720 102.805 164.765 ;
        RECT 105.035 164.720 105.325 164.765 ;
        RECT 106.225 164.720 106.515 164.765 ;
        RECT 102.515 164.580 106.515 164.720 ;
        RECT 102.515 164.535 102.805 164.580 ;
        RECT 105.035 164.535 105.325 164.580 ;
        RECT 106.225 164.535 106.515 164.580 ;
        RECT 88.690 164.380 89.010 164.440 ;
        RECT 85.560 164.240 89.010 164.380 ;
        RECT 79.490 164.195 79.780 164.240 ;
        RECT 81.060 164.195 81.350 164.240 ;
        RECT 83.160 164.195 83.450 164.240 ;
        RECT 88.690 164.180 89.010 164.240 ;
        RECT 99.285 164.380 99.575 164.425 ;
        RECT 102.950 164.380 103.240 164.425 ;
        RECT 104.520 164.380 104.810 164.425 ;
        RECT 106.620 164.380 106.910 164.425 ;
        RECT 99.285 164.240 102.720 164.380 ;
        RECT 99.285 164.195 99.575 164.240 ;
        RECT 46.370 164.040 46.690 164.100 ;
        RECT 40.940 163.900 46.690 164.040 ;
        RECT 46.370 163.840 46.690 163.900 ;
        RECT 47.290 163.840 47.610 164.100 ;
        RECT 47.750 164.040 48.070 164.100 ;
        RECT 48.685 164.040 48.975 164.085 ;
        RECT 47.750 163.900 48.975 164.040 ;
        RECT 47.750 163.840 48.070 163.900 ;
        RECT 48.685 163.855 48.975 163.900 ;
        RECT 76.745 164.040 77.035 164.085 ;
        RECT 85.010 164.040 85.330 164.100 ;
        RECT 76.745 163.900 85.330 164.040 ;
        RECT 102.580 164.040 102.720 164.240 ;
        RECT 102.950 164.240 106.910 164.380 ;
        RECT 102.950 164.195 103.240 164.240 ;
        RECT 104.520 164.195 104.810 164.240 ;
        RECT 106.620 164.195 106.910 164.240 ;
        RECT 106.170 164.040 106.490 164.100 ;
        RECT 102.580 163.900 106.490 164.040 ;
        RECT 76.745 163.855 77.035 163.900 ;
        RECT 85.010 163.840 85.330 163.900 ;
        RECT 106.170 163.840 106.490 163.900 ;
        RECT 107.565 164.040 107.855 164.085 ;
        RECT 108.470 164.040 108.790 164.100 ;
        RECT 107.565 163.900 108.790 164.040 ;
        RECT 109.940 164.040 110.080 164.920 ;
        RECT 110.785 164.875 111.075 164.920 ;
        RECT 113.070 164.860 113.390 164.920 ;
        RECT 115.000 164.920 117.515 165.060 ;
        RECT 115.000 164.780 115.140 164.920 ;
        RECT 117.225 164.875 117.515 164.920 ;
        RECT 123.190 164.860 123.510 165.120 ;
        RECT 129.170 164.860 129.490 165.120 ;
        RECT 130.180 165.105 130.320 165.260 ;
        RECT 130.550 165.200 130.870 165.260 ;
        RECT 135.625 165.215 135.915 165.445 ;
        RECT 137.450 165.400 137.770 165.460 ;
        RECT 136.620 165.260 137.770 165.400 ;
        RECT 130.105 164.875 130.395 165.105 ;
        RECT 131.010 164.860 131.330 165.120 ;
        RECT 132.000 164.875 132.290 165.105 ;
        RECT 134.705 165.060 134.995 165.105 ;
        RECT 135.150 165.060 135.470 165.120 ;
        RECT 136.620 165.105 136.760 165.260 ;
        RECT 137.450 165.200 137.770 165.260 ;
        RECT 137.910 165.105 138.230 165.120 ;
        RECT 134.705 164.920 135.470 165.060 ;
        RECT 134.705 164.875 134.995 164.920 ;
        RECT 110.310 164.720 110.630 164.780 ;
        RECT 111.245 164.720 111.535 164.765 ;
        RECT 110.310 164.580 111.535 164.720 ;
        RECT 110.310 164.520 110.630 164.580 ;
        RECT 111.245 164.535 111.535 164.580 ;
        RECT 112.610 164.720 112.930 164.780 ;
        RECT 113.545 164.720 113.835 164.765 ;
        RECT 112.610 164.580 113.835 164.720 ;
        RECT 112.610 164.520 112.930 164.580 ;
        RECT 113.545 164.535 113.835 164.580 ;
        RECT 114.910 164.520 115.230 164.780 ;
        RECT 116.765 164.720 117.055 164.765 ;
        RECT 117.670 164.720 117.990 164.780 ;
        RECT 125.950 164.720 126.270 164.780 ;
        RECT 130.565 164.720 130.855 164.765 ;
        RECT 116.765 164.580 126.270 164.720 ;
        RECT 116.765 164.535 117.055 164.580 ;
        RECT 117.670 164.520 117.990 164.580 ;
        RECT 120.980 164.425 121.120 164.580 ;
        RECT 125.950 164.520 126.270 164.580 ;
        RECT 130.180 164.580 130.855 164.720 ;
        RECT 130.180 164.440 130.320 164.580 ;
        RECT 130.565 164.535 130.855 164.580 ;
        RECT 120.905 164.195 121.195 164.425 ;
        RECT 130.090 164.180 130.410 164.440 ;
        RECT 132.020 164.380 132.160 164.875 ;
        RECT 135.150 164.860 135.470 164.920 ;
        RECT 136.545 164.875 136.835 165.105 ;
        RECT 137.880 164.875 138.230 165.105 ;
        RECT 137.910 164.860 138.230 164.875 ;
        RECT 143.890 164.860 144.210 165.120 ;
        RECT 137.425 164.720 137.715 164.765 ;
        RECT 138.615 164.720 138.905 164.765 ;
        RECT 141.135 164.720 141.425 164.765 ;
        RECT 137.425 164.580 141.425 164.720 ;
        RECT 137.425 164.535 137.715 164.580 ;
        RECT 138.615 164.535 138.905 164.580 ;
        RECT 141.135 164.535 141.425 164.580 ;
        RECT 131.560 164.240 132.160 164.380 ;
        RECT 132.865 164.380 133.155 164.425 ;
        RECT 136.530 164.380 136.850 164.440 ;
        RECT 132.865 164.240 136.850 164.380 ;
        RECT 115.385 164.040 115.675 164.085 ;
        RECT 109.940 163.900 115.675 164.040 ;
        RECT 107.565 163.855 107.855 163.900 ;
        RECT 108.470 163.840 108.790 163.900 ;
        RECT 115.385 163.855 115.675 163.900 ;
        RECT 118.130 163.840 118.450 164.100 ;
        RECT 121.825 164.040 122.115 164.085 ;
        RECT 124.110 164.040 124.430 164.100 ;
        RECT 121.825 163.900 124.430 164.040 ;
        RECT 121.825 163.855 122.115 163.900 ;
        RECT 124.110 163.840 124.430 163.900 ;
        RECT 128.710 164.040 129.030 164.100 ;
        RECT 131.560 164.040 131.700 164.240 ;
        RECT 132.865 164.195 133.155 164.240 ;
        RECT 136.530 164.180 136.850 164.240 ;
        RECT 137.030 164.380 137.320 164.425 ;
        RECT 139.130 164.380 139.420 164.425 ;
        RECT 140.700 164.380 140.990 164.425 ;
        RECT 137.030 164.240 140.990 164.380 ;
        RECT 137.030 164.195 137.320 164.240 ;
        RECT 139.130 164.195 139.420 164.240 ;
        RECT 140.700 164.195 140.990 164.240 ;
        RECT 128.710 163.900 131.700 164.040 ;
        RECT 131.930 164.040 132.250 164.100 ;
        RECT 133.785 164.040 134.075 164.085 ;
        RECT 131.930 163.900 134.075 164.040 ;
        RECT 128.710 163.840 129.030 163.900 ;
        RECT 131.930 163.840 132.250 163.900 ;
        RECT 133.785 163.855 134.075 163.900 ;
        RECT 143.430 163.840 143.750 164.100 ;
        RECT 144.810 163.840 145.130 164.100 ;
        RECT 17.320 163.220 147.040 163.700 ;
        RECT 26.130 162.820 26.450 163.080 ;
        RECT 27.050 162.820 27.370 163.080 ;
        RECT 28.890 162.820 29.210 163.080 ;
        RECT 29.825 163.020 30.115 163.065 ;
        RECT 32.110 163.020 32.430 163.080 ;
        RECT 39.945 163.020 40.235 163.065 ;
        RECT 40.390 163.020 40.710 163.080 ;
        RECT 29.825 162.880 39.240 163.020 ;
        RECT 29.825 162.835 30.115 162.880 ;
        RECT 32.110 162.820 32.430 162.880 ;
        RECT 19.730 162.680 20.020 162.725 ;
        RECT 21.830 162.680 22.120 162.725 ;
        RECT 23.400 162.680 23.690 162.725 ;
        RECT 19.730 162.540 23.690 162.680 ;
        RECT 19.730 162.495 20.020 162.540 ;
        RECT 21.830 162.495 22.120 162.540 ;
        RECT 23.400 162.495 23.690 162.540 ;
        RECT 20.125 162.340 20.415 162.385 ;
        RECT 21.315 162.340 21.605 162.385 ;
        RECT 23.835 162.340 24.125 162.385 ;
        RECT 28.980 162.340 29.120 162.820 ;
        RECT 31.230 162.680 31.520 162.725 ;
        RECT 33.330 162.680 33.620 162.725 ;
        RECT 34.900 162.680 35.190 162.725 ;
        RECT 31.230 162.540 35.190 162.680 ;
        RECT 31.230 162.495 31.520 162.540 ;
        RECT 33.330 162.495 33.620 162.540 ;
        RECT 34.900 162.495 35.190 162.540 ;
        RECT 20.125 162.200 24.125 162.340 ;
        RECT 20.125 162.155 20.415 162.200 ;
        RECT 21.315 162.155 21.605 162.200 ;
        RECT 23.835 162.155 24.125 162.200 ;
        RECT 26.680 162.200 29.120 162.340 ;
        RECT 31.625 162.340 31.915 162.385 ;
        RECT 32.815 162.340 33.105 162.385 ;
        RECT 35.335 162.340 35.625 162.385 ;
        RECT 31.625 162.200 35.625 162.340 ;
        RECT 19.230 161.800 19.550 162.060 ;
        RECT 26.680 162.045 26.820 162.200 ;
        RECT 31.625 162.155 31.915 162.200 ;
        RECT 32.815 162.155 33.105 162.200 ;
        RECT 35.335 162.155 35.625 162.200 ;
        RECT 26.605 161.815 26.895 162.045 ;
        RECT 27.510 162.000 27.830 162.060 ;
        RECT 30.270 162.000 30.590 162.060 ;
        RECT 39.100 162.045 39.240 162.880 ;
        RECT 39.945 162.880 40.710 163.020 ;
        RECT 39.945 162.835 40.235 162.880 ;
        RECT 40.390 162.820 40.710 162.880 ;
        RECT 45.465 163.020 45.755 163.065 ;
        RECT 47.290 163.020 47.610 163.080 ;
        RECT 45.465 162.880 47.610 163.020 ;
        RECT 45.465 162.835 45.755 162.880 ;
        RECT 47.290 162.820 47.610 162.880 ;
        RECT 51.905 163.020 52.195 163.065 ;
        RECT 54.190 163.020 54.510 163.080 ;
        RECT 51.905 162.880 54.510 163.020 ;
        RECT 51.905 162.835 52.195 162.880 ;
        RECT 54.190 162.820 54.510 162.880 ;
        RECT 84.550 163.020 84.870 163.080 ;
        RECT 87.325 163.020 87.615 163.065 ;
        RECT 84.550 162.880 87.615 163.020 ;
        RECT 84.550 162.820 84.870 162.880 ;
        RECT 87.325 162.835 87.615 162.880 ;
        RECT 88.690 163.020 89.010 163.080 ;
        RECT 89.165 163.020 89.455 163.065 ;
        RECT 92.370 163.020 92.690 163.080 ;
        RECT 88.690 162.880 92.690 163.020 ;
        RECT 88.690 162.820 89.010 162.880 ;
        RECT 89.165 162.835 89.455 162.880 ;
        RECT 92.370 162.820 92.690 162.880 ;
        RECT 98.810 163.020 99.130 163.080 ;
        RECT 110.310 163.020 110.630 163.080 ;
        RECT 112.610 163.020 112.930 163.080 ;
        RECT 98.810 162.880 112.930 163.020 ;
        RECT 98.810 162.820 99.130 162.880 ;
        RECT 110.310 162.820 110.630 162.880 ;
        RECT 112.610 162.820 112.930 162.880 ;
        RECT 113.070 162.820 113.390 163.080 ;
        RECT 117.685 163.020 117.975 163.065 ;
        RECT 119.050 163.020 119.370 163.080 ;
        RECT 117.685 162.880 119.370 163.020 ;
        RECT 117.685 162.835 117.975 162.880 ;
        RECT 119.050 162.820 119.370 162.880 ;
        RECT 119.510 163.020 119.830 163.080 ;
        RECT 132.390 163.020 132.710 163.080 ;
        RECT 133.785 163.020 134.075 163.065 ;
        RECT 119.510 162.880 131.700 163.020 ;
        RECT 119.510 162.820 119.830 162.880 ;
        RECT 49.605 162.495 49.895 162.725 ;
        RECT 84.105 162.680 84.395 162.725 ;
        RECT 85.930 162.680 86.250 162.740 ;
        RECT 84.105 162.540 86.250 162.680 ;
        RECT 84.105 162.495 84.395 162.540 ;
        RECT 47.290 162.140 47.610 162.400 ;
        RECT 49.680 162.340 49.820 162.495 ;
        RECT 85.930 162.480 86.250 162.540 ;
        RECT 87.770 162.680 88.090 162.740 ;
        RECT 89.610 162.680 89.930 162.740 ;
        RECT 87.770 162.540 89.930 162.680 ;
        RECT 87.770 162.480 88.090 162.540 ;
        RECT 89.610 162.480 89.930 162.540 ;
        RECT 91.030 162.680 91.320 162.725 ;
        RECT 93.130 162.680 93.420 162.725 ;
        RECT 94.700 162.680 94.990 162.725 ;
        RECT 91.030 162.540 94.990 162.680 ;
        RECT 91.030 162.495 91.320 162.540 ;
        RECT 93.130 162.495 93.420 162.540 ;
        RECT 94.700 162.495 94.990 162.540 ;
        RECT 107.090 162.680 107.410 162.740 ;
        RECT 111.245 162.680 111.535 162.725 ;
        RECT 114.910 162.680 115.230 162.740 ;
        RECT 120.430 162.680 120.750 162.740 ;
        RECT 107.090 162.540 115.230 162.680 ;
        RECT 107.090 162.480 107.410 162.540 ;
        RECT 111.245 162.495 111.535 162.540 ;
        RECT 114.910 162.480 115.230 162.540 ;
        RECT 119.600 162.540 120.750 162.680 ;
        RECT 83.630 162.340 83.950 162.400 ;
        RECT 90.545 162.340 90.835 162.385 ;
        RECT 49.680 162.200 51.200 162.340 ;
        RECT 30.745 162.000 31.035 162.045 ;
        RECT 27.315 161.875 29.200 162.000 ;
        RECT 27.315 161.860 29.425 161.875 ;
        RECT 27.510 161.800 27.830 161.860 ;
        RECT 20.580 161.475 20.870 161.705 ;
        RECT 27.985 161.475 28.275 161.705 ;
        RECT 29.060 161.690 29.425 161.860 ;
        RECT 30.270 161.860 31.035 162.000 ;
        RECT 30.270 161.800 30.590 161.860 ;
        RECT 30.745 161.815 31.035 161.860 ;
        RECT 31.740 161.860 32.800 162.000 ;
        RECT 29.135 161.645 29.425 161.690 ;
        RECT 29.810 161.660 30.130 161.720 ;
        RECT 31.740 161.660 31.880 161.860 ;
        RECT 32.110 161.705 32.430 161.720 ;
        RECT 29.810 161.520 31.880 161.660 ;
        RECT 20.150 161.320 20.470 161.380 ;
        RECT 20.700 161.320 20.840 161.475 ;
        RECT 20.150 161.180 20.840 161.320 ;
        RECT 21.990 161.320 22.310 161.380 ;
        RECT 27.510 161.320 27.830 161.380 ;
        RECT 21.990 161.180 27.830 161.320 ;
        RECT 28.060 161.320 28.200 161.475 ;
        RECT 29.810 161.460 30.130 161.520 ;
        RECT 32.080 161.475 32.430 161.705 ;
        RECT 32.660 161.660 32.800 161.860 ;
        RECT 38.565 161.815 38.855 162.045 ;
        RECT 39.025 161.815 39.315 162.045 ;
        RECT 38.640 161.660 38.780 161.815 ;
        RECT 39.930 161.800 40.250 162.060 ;
        RECT 40.390 162.000 40.710 162.060 ;
        RECT 42.245 162.000 42.535 162.045 ;
        RECT 40.390 161.860 42.535 162.000 ;
        RECT 40.390 161.800 40.710 161.860 ;
        RECT 42.245 161.815 42.535 161.860 ;
        RECT 42.780 161.860 44.760 162.000 ;
        RECT 40.020 161.660 40.160 161.800 ;
        RECT 32.660 161.520 38.320 161.660 ;
        RECT 38.640 161.520 40.160 161.660 ;
        RECT 41.310 161.660 41.630 161.720 ;
        RECT 42.780 161.660 42.920 161.860 ;
        RECT 41.310 161.520 42.920 161.660 ;
        RECT 32.110 161.460 32.430 161.475 ;
        RECT 28.430 161.320 28.750 161.380 ;
        RECT 34.870 161.320 35.190 161.380 ;
        RECT 37.645 161.320 37.935 161.365 ;
        RECT 28.060 161.180 37.935 161.320 ;
        RECT 38.180 161.320 38.320 161.520 ;
        RECT 41.310 161.460 41.630 161.520 ;
        RECT 43.150 161.460 43.470 161.720 ;
        RECT 44.620 161.705 44.760 161.860 ;
        RECT 47.750 161.800 48.070 162.060 ;
        RECT 50.065 162.000 50.355 162.045 ;
        RECT 50.510 162.000 50.830 162.060 ;
        RECT 51.060 162.045 51.200 162.200 ;
        RECT 83.630 162.200 90.835 162.340 ;
        RECT 83.630 162.140 83.950 162.200 ;
        RECT 90.545 162.155 90.835 162.200 ;
        RECT 91.425 162.340 91.715 162.385 ;
        RECT 92.615 162.340 92.905 162.385 ;
        RECT 95.135 162.340 95.425 162.385 ;
        RECT 91.425 162.200 95.425 162.340 ;
        RECT 91.425 162.155 91.715 162.200 ;
        RECT 92.615 162.155 92.905 162.200 ;
        RECT 95.135 162.155 95.425 162.200 ;
        RECT 98.825 162.340 99.115 162.385 ;
        RECT 101.110 162.340 101.430 162.400 ;
        RECT 112.610 162.340 112.930 162.400 ;
        RECT 114.465 162.340 114.755 162.385 ;
        RECT 98.825 162.200 108.240 162.340 ;
        RECT 98.825 162.155 99.115 162.200 ;
        RECT 101.110 162.140 101.430 162.200 ;
        RECT 50.065 161.860 50.830 162.000 ;
        RECT 50.065 161.815 50.355 161.860 ;
        RECT 44.545 161.660 44.835 161.705 ;
        RECT 50.140 161.660 50.280 161.815 ;
        RECT 50.510 161.800 50.830 161.860 ;
        RECT 50.985 161.815 51.275 162.045 ;
        RECT 82.710 161.800 83.030 162.060 ;
        RECT 84.090 161.800 84.410 162.060 ;
        RECT 85.025 161.815 85.315 162.045 ;
        RECT 85.485 162.000 85.775 162.045 ;
        RECT 87.310 162.000 87.630 162.060 ;
        RECT 85.485 161.860 87.630 162.000 ;
        RECT 85.485 161.815 85.775 161.860 ;
        RECT 44.545 161.520 50.280 161.660 ;
        RECT 85.100 161.660 85.240 161.815 ;
        RECT 87.310 161.800 87.630 161.860 ;
        RECT 88.230 162.000 88.550 162.060 ;
        RECT 88.705 162.000 88.995 162.045 ;
        RECT 88.230 161.860 88.995 162.000 ;
        RECT 88.230 161.800 88.550 161.860 ;
        RECT 88.705 161.815 88.995 161.860 ;
        RECT 89.610 161.800 89.930 162.060 ;
        RECT 100.650 162.000 100.970 162.060 ;
        RECT 102.505 162.000 102.795 162.045 ;
        RECT 91.540 161.860 102.795 162.000 ;
        RECT 86.850 161.660 87.170 161.720 ;
        RECT 91.540 161.660 91.680 161.860 ;
        RECT 100.650 161.800 100.970 161.860 ;
        RECT 102.505 161.815 102.795 161.860 ;
        RECT 102.950 162.000 103.270 162.060 ;
        RECT 108.100 162.045 108.240 162.200 ;
        RECT 112.610 162.200 114.755 162.340 ;
        RECT 115.000 162.340 115.140 162.480 ;
        RECT 115.000 162.200 116.060 162.340 ;
        RECT 112.610 162.140 112.930 162.200 ;
        RECT 114.465 162.155 114.755 162.200 ;
        RECT 105.725 162.000 106.015 162.045 ;
        RECT 102.950 161.860 106.015 162.000 ;
        RECT 85.100 161.520 85.700 161.660 ;
        RECT 44.545 161.475 44.835 161.520 ;
        RECT 38.550 161.320 38.870 161.380 ;
        RECT 40.865 161.320 41.155 161.365 ;
        RECT 38.180 161.180 41.155 161.320 ;
        RECT 20.150 161.120 20.470 161.180 ;
        RECT 21.990 161.120 22.310 161.180 ;
        RECT 27.510 161.120 27.830 161.180 ;
        RECT 28.430 161.120 28.750 161.180 ;
        RECT 34.870 161.120 35.190 161.180 ;
        RECT 37.645 161.135 37.935 161.180 ;
        RECT 38.550 161.120 38.870 161.180 ;
        RECT 40.865 161.135 41.155 161.180 ;
        RECT 44.085 161.320 44.375 161.365 ;
        RECT 45.545 161.320 45.835 161.365 ;
        RECT 44.085 161.180 45.835 161.320 ;
        RECT 44.085 161.135 44.375 161.180 ;
        RECT 45.545 161.135 45.835 161.180 ;
        RECT 46.370 161.120 46.690 161.380 ;
        RECT 85.560 161.320 85.700 161.520 ;
        RECT 86.850 161.520 91.680 161.660 ;
        RECT 91.880 161.660 92.170 161.705 ;
        RECT 102.580 161.660 102.720 161.815 ;
        RECT 102.950 161.800 103.270 161.860 ;
        RECT 105.725 161.815 106.015 161.860 ;
        RECT 108.025 161.815 108.315 162.045 ;
        RECT 115.370 161.800 115.690 162.060 ;
        RECT 115.920 162.045 116.060 162.200 ;
        RECT 115.845 161.815 116.135 162.045 ;
        RECT 118.130 162.000 118.450 162.060 ;
        RECT 119.600 162.045 119.740 162.540 ;
        RECT 120.430 162.480 120.750 162.540 ;
        RECT 123.650 162.680 123.970 162.740 ;
        RECT 128.710 162.680 129.030 162.740 ;
        RECT 123.650 162.540 129.030 162.680 ;
        RECT 123.650 162.480 123.970 162.540 ;
        RECT 124.570 162.340 124.890 162.400 ;
        RECT 120.060 162.200 124.890 162.340 ;
        RECT 120.060 162.045 120.200 162.200 ;
        RECT 124.570 162.140 124.890 162.200 ;
        RECT 118.605 162.000 118.895 162.045 ;
        RECT 118.130 161.860 118.895 162.000 ;
        RECT 118.130 161.800 118.450 161.860 ;
        RECT 118.605 161.815 118.895 161.860 ;
        RECT 119.525 161.815 119.815 162.045 ;
        RECT 119.985 161.815 120.275 162.045 ;
        RECT 120.430 162.000 120.750 162.060 ;
        RECT 121.825 162.000 122.115 162.045 ;
        RECT 120.430 161.860 122.115 162.000 ;
        RECT 120.430 161.800 120.750 161.860 ;
        RECT 121.825 161.815 122.115 161.860 ;
        RECT 122.270 162.000 122.590 162.060 ;
        RECT 122.745 162.000 123.035 162.045 ;
        RECT 122.270 161.860 123.035 162.000 ;
        RECT 122.270 161.800 122.590 161.860 ;
        RECT 122.745 161.815 123.035 161.860 ;
        RECT 123.205 162.000 123.495 162.045 ;
        RECT 124.110 162.000 124.430 162.060 ;
        RECT 127.420 162.045 127.560 162.540 ;
        RECT 128.710 162.480 129.030 162.540 ;
        RECT 130.105 162.680 130.395 162.725 ;
        RECT 131.010 162.680 131.330 162.740 ;
        RECT 130.105 162.540 131.330 162.680 ;
        RECT 130.105 162.495 130.395 162.540 ;
        RECT 131.010 162.480 131.330 162.540 ;
        RECT 127.790 162.140 128.110 162.400 ;
        RECT 128.250 162.140 128.570 162.400 ;
        RECT 126.425 162.000 126.715 162.045 ;
        RECT 123.205 161.860 124.430 162.000 ;
        RECT 123.205 161.815 123.495 161.860 ;
        RECT 124.110 161.800 124.430 161.860 ;
        RECT 125.580 161.860 126.715 162.000 ;
        RECT 91.880 161.520 98.120 161.660 ;
        RECT 102.580 161.520 123.420 161.660 ;
        RECT 86.850 161.460 87.170 161.520 ;
        RECT 91.880 161.475 92.170 161.520 ;
        RECT 87.325 161.320 87.615 161.365 ;
        RECT 87.770 161.320 88.090 161.380 ;
        RECT 85.560 161.180 88.090 161.320 ;
        RECT 87.325 161.135 87.615 161.180 ;
        RECT 87.770 161.120 88.090 161.180 ;
        RECT 88.230 161.120 88.550 161.380 ;
        RECT 96.970 161.320 97.290 161.380 ;
        RECT 97.445 161.320 97.735 161.365 ;
        RECT 96.970 161.180 97.735 161.320 ;
        RECT 97.980 161.320 98.120 161.520 ;
        RECT 123.280 161.380 123.420 161.520 ;
        RECT 102.965 161.320 103.255 161.365 ;
        RECT 97.980 161.180 103.255 161.320 ;
        RECT 96.970 161.120 97.290 161.180 ;
        RECT 97.445 161.135 97.735 161.180 ;
        RECT 102.965 161.135 103.255 161.180 ;
        RECT 109.850 161.320 110.170 161.380 ;
        RECT 113.085 161.320 113.375 161.365 ;
        RECT 109.850 161.180 113.375 161.320 ;
        RECT 109.850 161.120 110.170 161.180 ;
        RECT 113.085 161.135 113.375 161.180 ;
        RECT 114.005 161.320 114.295 161.365 ;
        RECT 118.590 161.320 118.910 161.380 ;
        RECT 114.005 161.180 118.910 161.320 ;
        RECT 114.005 161.135 114.295 161.180 ;
        RECT 118.590 161.120 118.910 161.180 ;
        RECT 120.905 161.320 121.195 161.365 ;
        RECT 121.350 161.320 121.670 161.380 ;
        RECT 120.905 161.180 121.670 161.320 ;
        RECT 120.905 161.135 121.195 161.180 ;
        RECT 121.350 161.120 121.670 161.180 ;
        RECT 123.190 161.120 123.510 161.380 ;
        RECT 125.580 161.320 125.720 161.860 ;
        RECT 126.425 161.815 126.715 161.860 ;
        RECT 127.345 161.815 127.635 162.045 ;
        RECT 129.185 162.000 129.475 162.045 ;
        RECT 130.090 162.000 130.410 162.060 ;
        RECT 131.560 162.045 131.700 162.880 ;
        RECT 132.390 162.880 134.075 163.020 ;
        RECT 132.390 162.820 132.710 162.880 ;
        RECT 133.785 162.835 134.075 162.880 ;
        RECT 137.465 163.020 137.755 163.065 ;
        RECT 137.910 163.020 138.230 163.080 ;
        RECT 137.465 162.880 138.230 163.020 ;
        RECT 137.465 162.835 137.755 162.880 ;
        RECT 137.910 162.820 138.230 162.880 ;
        RECT 136.530 162.340 136.850 162.400 ;
        RECT 140.225 162.340 140.515 162.385 ;
        RECT 132.020 162.200 134.920 162.340 ;
        RECT 129.185 161.860 130.410 162.000 ;
        RECT 129.185 161.815 129.475 161.860 ;
        RECT 130.090 161.800 130.410 161.860 ;
        RECT 131.485 161.815 131.775 162.045 ;
        RECT 125.965 161.660 126.255 161.705 ;
        RECT 126.870 161.660 127.190 161.720 ;
        RECT 125.965 161.520 127.190 161.660 ;
        RECT 125.965 161.475 126.255 161.520 ;
        RECT 126.870 161.460 127.190 161.520 ;
        RECT 127.790 161.660 128.110 161.720 ;
        RECT 132.020 161.660 132.160 162.200 ;
        RECT 134.780 162.060 134.920 162.200 ;
        RECT 136.530 162.200 140.515 162.340 ;
        RECT 136.530 162.140 136.850 162.200 ;
        RECT 140.225 162.155 140.515 162.200 ;
        RECT 133.770 161.800 134.090 162.060 ;
        RECT 134.690 161.800 135.010 162.060 ;
        RECT 143.430 162.000 143.750 162.060 ;
        RECT 144.365 162.000 144.655 162.045 ;
        RECT 143.430 161.860 144.655 162.000 ;
        RECT 143.430 161.800 143.750 161.860 ;
        RECT 144.365 161.815 144.655 161.860 ;
        RECT 127.790 161.520 132.160 161.660 ;
        RECT 127.790 161.460 128.110 161.520 ;
        RECT 132.390 161.460 132.710 161.720 ;
        RECT 133.310 161.660 133.630 161.720 ;
        RECT 138.830 161.660 139.150 161.720 ;
        RECT 133.310 161.520 139.150 161.660 ;
        RECT 133.310 161.460 133.630 161.520 ;
        RECT 138.830 161.460 139.150 161.520 ;
        RECT 139.305 161.660 139.595 161.705 ;
        RECT 141.605 161.660 141.895 161.705 ;
        RECT 139.305 161.520 141.895 161.660 ;
        RECT 139.305 161.475 139.595 161.520 ;
        RECT 141.605 161.475 141.895 161.520 ;
        RECT 129.170 161.320 129.490 161.380 ;
        RECT 130.550 161.320 130.870 161.380 ;
        RECT 125.580 161.180 130.870 161.320 ;
        RECT 129.170 161.120 129.490 161.180 ;
        RECT 130.550 161.120 130.870 161.180 ;
        RECT 131.010 161.320 131.330 161.380 ;
        RECT 134.690 161.320 135.010 161.380 ;
        RECT 131.010 161.180 135.010 161.320 ;
        RECT 131.010 161.120 131.330 161.180 ;
        RECT 134.690 161.120 135.010 161.180 ;
        RECT 135.625 161.320 135.915 161.365 ;
        RECT 136.070 161.320 136.390 161.380 ;
        RECT 135.625 161.180 136.390 161.320 ;
        RECT 135.625 161.135 135.915 161.180 ;
        RECT 136.070 161.120 136.390 161.180 ;
        RECT 139.750 161.120 140.070 161.380 ;
        RECT 17.320 160.500 147.040 160.980 ;
        RECT 20.150 160.100 20.470 160.360 ;
        RECT 21.005 160.300 21.295 160.345 ;
        RECT 21.530 160.300 21.850 160.360 ;
        RECT 25.210 160.300 25.530 160.360 ;
        RECT 30.270 160.300 30.590 160.360 ;
        RECT 21.005 160.160 21.850 160.300 ;
        RECT 21.005 160.115 21.295 160.160 ;
        RECT 21.530 160.100 21.850 160.160 ;
        RECT 23.460 160.160 30.590 160.300 ;
        RECT 21.990 159.760 22.310 160.020 ;
        RECT 19.230 159.620 19.550 159.680 ;
        RECT 22.465 159.620 22.755 159.665 ;
        RECT 23.460 159.620 23.600 160.160 ;
        RECT 25.210 160.100 25.530 160.160 ;
        RECT 30.270 160.100 30.590 160.160 ;
        RECT 30.730 160.345 31.050 160.360 ;
        RECT 30.730 160.115 31.115 160.345 ;
        RECT 31.665 160.300 31.955 160.345 ;
        RECT 32.110 160.300 32.430 160.360 ;
        RECT 31.665 160.160 32.430 160.300 ;
        RECT 31.665 160.115 31.955 160.160 ;
        RECT 30.730 160.100 31.050 160.115 ;
        RECT 32.110 160.100 32.430 160.160 ;
        RECT 39.930 160.300 40.250 160.360 ;
        RECT 42.245 160.300 42.535 160.345 ;
        RECT 39.930 160.160 42.535 160.300 ;
        RECT 39.930 160.100 40.250 160.160 ;
        RECT 42.245 160.115 42.535 160.160 ;
        RECT 43.150 160.300 43.470 160.360 ;
        RECT 45.005 160.300 45.295 160.345 ;
        RECT 43.150 160.160 45.295 160.300 ;
        RECT 43.150 160.100 43.470 160.160 ;
        RECT 45.005 160.115 45.295 160.160 ;
        RECT 88.690 160.100 89.010 160.360 ;
        RECT 91.925 160.300 92.215 160.345 ;
        RECT 100.650 160.300 100.970 160.360 ;
        RECT 91.925 160.160 100.970 160.300 ;
        RECT 91.925 160.115 92.215 160.160 ;
        RECT 100.650 160.100 100.970 160.160 ;
        RECT 101.585 160.300 101.875 160.345 ;
        RECT 102.950 160.300 103.270 160.360 ;
        RECT 101.585 160.160 103.270 160.300 ;
        RECT 101.585 160.115 101.875 160.160 ;
        RECT 102.950 160.100 103.270 160.160 ;
        RECT 105.250 160.300 105.570 160.360 ;
        RECT 105.725 160.300 106.015 160.345 ;
        RECT 105.250 160.160 106.015 160.300 ;
        RECT 105.250 160.100 105.570 160.160 ;
        RECT 105.725 160.115 106.015 160.160 ;
        RECT 106.630 160.300 106.950 160.360 ;
        RECT 115.830 160.300 116.150 160.360 ;
        RECT 116.305 160.300 116.595 160.345 ;
        RECT 106.630 160.160 108.470 160.300 ;
        RECT 106.630 160.100 106.950 160.160 ;
        RECT 23.830 160.005 24.150 160.020 ;
        RECT 23.800 159.960 24.150 160.005 ;
        RECT 27.970 159.960 28.290 160.020 ;
        RECT 29.810 159.960 30.130 160.020 ;
        RECT 23.800 159.820 24.300 159.960 ;
        RECT 27.970 159.820 30.130 159.960 ;
        RECT 23.800 159.775 24.150 159.820 ;
        RECT 23.830 159.760 24.150 159.775 ;
        RECT 27.970 159.760 28.290 159.820 ;
        RECT 29.810 159.760 30.130 159.820 ;
        RECT 19.230 159.480 23.600 159.620 ;
        RECT 30.360 159.620 30.500 160.100 ;
        RECT 55.570 159.960 55.890 160.020 ;
        RECT 35.420 159.820 55.890 159.960 ;
        RECT 35.420 159.665 35.560 159.820 ;
        RECT 36.710 159.665 37.030 159.680 ;
        RECT 35.345 159.620 35.635 159.665 ;
        RECT 30.360 159.480 35.635 159.620 ;
        RECT 19.230 159.420 19.550 159.480 ;
        RECT 22.465 159.435 22.755 159.480 ;
        RECT 35.345 159.435 35.635 159.480 ;
        RECT 36.680 159.435 37.030 159.665 ;
        RECT 36.710 159.420 37.030 159.435 ;
        RECT 46.370 159.620 46.690 159.680 ;
        RECT 51.980 159.665 52.120 159.820 ;
        RECT 55.570 159.760 55.890 159.820 ;
        RECT 82.710 159.960 83.030 160.020 ;
        RECT 89.150 159.960 89.470 160.020 ;
        RECT 96.065 159.960 96.355 160.005 ;
        RECT 82.710 159.820 89.470 159.960 ;
        RECT 82.710 159.760 83.030 159.820 ;
        RECT 89.150 159.760 89.470 159.820 ;
        RECT 90.620 159.820 96.355 159.960 ;
        RECT 50.570 159.620 50.860 159.665 ;
        RECT 46.370 159.480 50.860 159.620 ;
        RECT 46.370 159.420 46.690 159.480 ;
        RECT 50.570 159.435 50.860 159.480 ;
        RECT 51.905 159.435 52.195 159.665 ;
        RECT 62.945 159.620 63.235 159.665 ;
        RECT 64.325 159.620 64.615 159.665 ;
        RECT 62.945 159.480 64.615 159.620 ;
        RECT 62.945 159.435 63.235 159.480 ;
        RECT 64.325 159.435 64.615 159.480 ;
        RECT 84.090 159.620 84.410 159.680 ;
        RECT 87.785 159.620 88.075 159.665 ;
        RECT 84.090 159.480 88.075 159.620 ;
        RECT 84.090 159.420 84.410 159.480 ;
        RECT 87.785 159.435 88.075 159.480 ;
        RECT 23.345 159.280 23.635 159.325 ;
        RECT 24.535 159.280 24.825 159.325 ;
        RECT 27.055 159.280 27.345 159.325 ;
        RECT 23.345 159.140 27.345 159.280 ;
        RECT 23.345 159.095 23.635 159.140 ;
        RECT 24.535 159.095 24.825 159.140 ;
        RECT 27.055 159.095 27.345 159.140 ;
        RECT 36.225 159.280 36.515 159.325 ;
        RECT 37.415 159.280 37.705 159.325 ;
        RECT 39.935 159.280 40.225 159.325 ;
        RECT 36.225 159.140 40.225 159.280 ;
        RECT 36.225 159.095 36.515 159.140 ;
        RECT 37.415 159.095 37.705 159.140 ;
        RECT 39.935 159.095 40.225 159.140 ;
        RECT 47.315 159.280 47.605 159.325 ;
        RECT 49.835 159.280 50.125 159.325 ;
        RECT 51.025 159.280 51.315 159.325 ;
        RECT 47.315 159.140 51.315 159.280 ;
        RECT 47.315 159.095 47.605 159.140 ;
        RECT 49.835 159.095 50.125 159.140 ;
        RECT 51.025 159.095 51.315 159.140 ;
        RECT 67.070 159.080 67.390 159.340 ;
        RECT 79.490 159.080 79.810 159.340 ;
        RECT 87.860 159.280 88.000 159.435 ;
        RECT 89.610 159.420 89.930 159.680 ;
        RECT 90.620 159.665 90.760 159.820 ;
        RECT 96.065 159.775 96.355 159.820 ;
        RECT 96.970 159.960 97.290 160.020 ;
        RECT 106.170 159.960 106.490 160.020 ;
        RECT 107.565 159.960 107.855 160.005 ;
        RECT 96.970 159.820 105.020 159.960 ;
        RECT 96.970 159.760 97.290 159.820 ;
        RECT 90.545 159.435 90.835 159.665 ;
        RECT 92.370 159.620 92.690 159.680 ;
        RECT 92.845 159.620 93.135 159.665 ;
        RECT 95.145 159.620 95.435 159.665 ;
        RECT 92.370 159.480 95.435 159.620 ;
        RECT 88.230 159.280 88.550 159.340 ;
        RECT 90.620 159.280 90.760 159.435 ;
        RECT 92.370 159.420 92.690 159.480 ;
        RECT 92.845 159.435 93.135 159.480 ;
        RECT 95.145 159.435 95.435 159.480 ;
        RECT 98.365 159.620 98.655 159.665 ;
        RECT 98.810 159.620 99.130 159.680 ;
        RECT 98.365 159.480 99.130 159.620 ;
        RECT 98.365 159.435 98.655 159.480 ;
        RECT 98.810 159.420 99.130 159.480 ;
        RECT 99.270 159.420 99.590 159.680 ;
        RECT 99.730 159.420 100.050 159.680 ;
        RECT 100.190 159.420 100.510 159.680 ;
        RECT 104.880 159.665 105.020 159.820 ;
        RECT 106.170 159.820 107.855 159.960 ;
        RECT 108.330 159.960 108.470 160.160 ;
        RECT 115.830 160.160 116.595 160.300 ;
        RECT 115.830 160.100 116.150 160.160 ;
        RECT 116.305 160.115 116.595 160.160 ;
        RECT 118.130 160.100 118.450 160.360 ;
        RECT 122.745 160.300 123.035 160.345 ;
        RECT 125.950 160.300 126.270 160.360 ;
        RECT 132.390 160.300 132.710 160.360 ;
        RECT 133.770 160.300 134.090 160.360 ;
        RECT 122.745 160.160 125.720 160.300 ;
        RECT 122.745 160.115 123.035 160.160 ;
        RECT 118.220 159.960 118.360 160.100 ;
        RECT 108.330 159.820 116.060 159.960 ;
        RECT 118.220 159.820 121.120 159.960 ;
        RECT 106.170 159.760 106.490 159.820 ;
        RECT 107.565 159.775 107.855 159.820 ;
        RECT 104.805 159.435 105.095 159.665 ;
        RECT 106.630 159.420 106.950 159.680 ;
        RECT 107.090 159.420 107.410 159.680 ;
        RECT 108.470 159.420 108.790 159.680 ;
        RECT 110.310 159.420 110.630 159.680 ;
        RECT 112.625 159.620 112.915 159.665 ;
        RECT 113.070 159.620 113.390 159.680 ;
        RECT 115.920 159.665 116.060 159.820 ;
        RECT 114.465 159.620 114.755 159.665 ;
        RECT 112.625 159.480 113.390 159.620 ;
        RECT 112.625 159.435 112.915 159.480 ;
        RECT 113.070 159.420 113.390 159.480 ;
        RECT 113.620 159.480 114.755 159.620 ;
        RECT 87.860 159.140 90.760 159.280 ;
        RECT 88.230 159.080 88.550 159.140 ;
        RECT 97.905 159.095 98.195 159.325 ;
        RECT 102.045 159.280 102.335 159.325 ;
        RECT 99.820 159.140 102.335 159.280 ;
        RECT 22.950 158.940 23.240 158.985 ;
        RECT 25.050 158.940 25.340 158.985 ;
        RECT 26.620 158.940 26.910 158.985 ;
        RECT 22.950 158.800 26.910 158.940 ;
        RECT 22.950 158.755 23.240 158.800 ;
        RECT 25.050 158.755 25.340 158.800 ;
        RECT 26.620 158.755 26.910 158.800 ;
        RECT 28.890 158.940 29.210 159.000 ;
        RECT 29.365 158.940 29.655 158.985 ;
        RECT 28.890 158.800 29.655 158.940 ;
        RECT 28.890 158.740 29.210 158.800 ;
        RECT 29.365 158.755 29.655 158.800 ;
        RECT 35.830 158.940 36.120 158.985 ;
        RECT 37.930 158.940 38.220 158.985 ;
        RECT 39.500 158.940 39.790 158.985 ;
        RECT 35.830 158.800 39.790 158.940 ;
        RECT 35.830 158.755 36.120 158.800 ;
        RECT 37.930 158.755 38.220 158.800 ;
        RECT 39.500 158.755 39.790 158.800 ;
        RECT 47.750 158.940 48.040 158.985 ;
        RECT 49.320 158.940 49.610 158.985 ;
        RECT 51.420 158.940 51.710 158.985 ;
        RECT 47.750 158.800 51.710 158.940 ;
        RECT 97.980 158.940 98.120 159.095 ;
        RECT 99.820 158.940 99.960 159.140 ;
        RECT 102.045 159.095 102.335 159.140 ;
        RECT 113.620 159.000 113.760 159.480 ;
        RECT 114.465 159.435 114.755 159.480 ;
        RECT 115.845 159.435 116.135 159.665 ;
        RECT 117.225 159.620 117.515 159.665 ;
        RECT 116.380 159.480 117.515 159.620 ;
        RECT 115.370 159.280 115.690 159.340 ;
        RECT 116.380 159.280 116.520 159.480 ;
        RECT 117.225 159.435 117.515 159.480 ;
        RECT 118.145 159.620 118.435 159.665 ;
        RECT 118.590 159.620 118.910 159.680 ;
        RECT 118.145 159.480 118.910 159.620 ;
        RECT 118.145 159.435 118.435 159.480 ;
        RECT 118.590 159.420 118.910 159.480 ;
        RECT 119.050 159.420 119.370 159.680 ;
        RECT 119.985 159.620 120.275 159.665 ;
        RECT 120.430 159.620 120.750 159.680 ;
        RECT 120.980 159.665 121.120 159.820 ;
        RECT 123.190 159.760 123.510 160.020 ;
        RECT 125.580 159.960 125.720 160.160 ;
        RECT 125.950 160.160 129.860 160.300 ;
        RECT 125.950 160.100 126.270 160.160 ;
        RECT 125.580 159.820 129.400 159.960 ;
        RECT 119.985 159.480 120.750 159.620 ;
        RECT 119.985 159.435 120.275 159.480 ;
        RECT 120.430 159.420 120.750 159.480 ;
        RECT 120.905 159.435 121.195 159.665 ;
        RECT 128.265 159.620 128.555 159.665 ;
        RECT 128.710 159.620 129.030 159.680 ;
        RECT 129.260 159.665 129.400 159.820 ;
        RECT 129.720 159.665 129.860 160.160 ;
        RECT 132.390 160.160 134.090 160.300 ;
        RECT 132.390 160.100 132.710 160.160 ;
        RECT 133.770 160.100 134.090 160.160 ;
        RECT 134.705 160.300 134.995 160.345 ;
        RECT 139.750 160.300 140.070 160.360 ;
        RECT 134.705 160.160 140.070 160.300 ;
        RECT 134.705 160.115 134.995 160.160 ;
        RECT 139.750 160.100 140.070 160.160 ;
        RECT 131.485 159.960 131.775 160.005 ;
        RECT 144.350 159.960 144.670 160.020 ;
        RECT 131.485 159.820 144.670 159.960 ;
        RECT 131.485 159.775 131.775 159.820 ;
        RECT 144.350 159.760 144.670 159.820 ;
        RECT 128.265 159.480 129.030 159.620 ;
        RECT 128.265 159.435 128.555 159.480 ;
        RECT 128.710 159.420 129.030 159.480 ;
        RECT 129.185 159.435 129.475 159.665 ;
        RECT 129.645 159.435 129.935 159.665 ;
        RECT 130.090 159.420 130.410 159.680 ;
        RECT 131.930 159.420 132.250 159.680 ;
        RECT 132.390 159.620 132.710 159.680 ;
        RECT 132.865 159.620 133.155 159.665 ;
        RECT 132.390 159.480 133.155 159.620 ;
        RECT 132.390 159.420 132.710 159.480 ;
        RECT 132.865 159.435 133.155 159.480 ;
        RECT 133.310 159.420 133.630 159.680 ;
        RECT 133.770 159.420 134.090 159.680 ;
        RECT 136.990 159.665 137.310 159.680 ;
        RECT 136.960 159.435 137.310 159.665 ;
        RECT 143.905 159.435 144.195 159.665 ;
        RECT 136.990 159.420 137.310 159.435 ;
        RECT 115.370 159.140 116.520 159.280 ;
        RECT 121.365 159.280 121.655 159.325 ;
        RECT 124.570 159.280 124.890 159.340 ;
        RECT 121.365 159.140 124.890 159.280 ;
        RECT 115.370 159.080 115.690 159.140 ;
        RECT 121.365 159.095 121.655 159.140 ;
        RECT 124.570 159.080 124.890 159.140 ;
        RECT 127.345 159.280 127.635 159.325 ;
        RECT 135.625 159.280 135.915 159.325 ;
        RECT 127.345 159.140 135.915 159.280 ;
        RECT 127.345 159.095 127.635 159.140 ;
        RECT 129.260 159.000 129.400 159.140 ;
        RECT 133.860 159.000 134.000 159.140 ;
        RECT 135.625 159.095 135.915 159.140 ;
        RECT 136.505 159.280 136.795 159.325 ;
        RECT 137.695 159.280 137.985 159.325 ;
        RECT 140.215 159.280 140.505 159.325 ;
        RECT 136.505 159.140 140.505 159.280 ;
        RECT 136.505 159.095 136.795 159.140 ;
        RECT 137.695 159.095 137.985 159.140 ;
        RECT 140.215 159.095 140.505 159.140 ;
        RECT 97.980 158.800 99.960 158.940 ;
        RECT 100.650 158.940 100.970 159.000 ;
        RECT 113.530 158.940 113.850 159.000 ;
        RECT 100.650 158.800 113.850 158.940 ;
        RECT 47.750 158.755 48.040 158.800 ;
        RECT 49.320 158.755 49.610 158.800 ;
        RECT 51.420 158.755 51.710 158.800 ;
        RECT 100.650 158.740 100.970 158.800 ;
        RECT 113.530 158.740 113.850 158.800 ;
        RECT 114.925 158.940 115.215 158.985 ;
        RECT 119.525 158.940 119.815 158.985 ;
        RECT 114.925 158.800 119.280 158.940 ;
        RECT 114.925 158.755 115.215 158.800 ;
        RECT 21.070 158.400 21.390 158.660 ;
        RECT 30.745 158.600 31.035 158.645 ;
        RECT 31.650 158.600 31.970 158.660 ;
        RECT 30.745 158.460 31.970 158.600 ;
        RECT 30.745 158.415 31.035 158.460 ;
        RECT 31.650 158.400 31.970 158.460 ;
        RECT 62.470 158.400 62.790 158.660 ;
        RECT 82.710 158.400 83.030 158.660 ;
        RECT 87.770 158.400 88.090 158.660 ;
        RECT 96.985 158.600 97.275 158.645 ;
        RECT 99.270 158.600 99.590 158.660 ;
        RECT 115.830 158.600 116.150 158.660 ;
        RECT 96.985 158.460 116.150 158.600 ;
        RECT 96.985 158.415 97.275 158.460 ;
        RECT 99.270 158.400 99.590 158.460 ;
        RECT 115.830 158.400 116.150 158.460 ;
        RECT 117.685 158.600 117.975 158.645 ;
        RECT 118.130 158.600 118.450 158.660 ;
        RECT 117.685 158.460 118.450 158.600 ;
        RECT 119.140 158.600 119.280 158.800 ;
        RECT 119.525 158.800 128.940 158.940 ;
        RECT 119.525 158.755 119.815 158.800 ;
        RECT 121.350 158.600 121.670 158.660 ;
        RECT 119.140 158.460 121.670 158.600 ;
        RECT 117.685 158.415 117.975 158.460 ;
        RECT 118.130 158.400 118.450 158.460 ;
        RECT 121.350 158.400 121.670 158.460 ;
        RECT 121.825 158.600 122.115 158.645 ;
        RECT 123.650 158.600 123.970 158.660 ;
        RECT 121.825 158.460 123.970 158.600 ;
        RECT 128.800 158.600 128.940 158.800 ;
        RECT 129.170 158.740 129.490 159.000 ;
        RECT 133.770 158.740 134.090 159.000 ;
        RECT 136.110 158.940 136.400 158.985 ;
        RECT 138.210 158.940 138.500 158.985 ;
        RECT 139.780 158.940 140.070 158.985 ;
        RECT 143.980 158.940 144.120 159.435 ;
        RECT 136.110 158.800 140.070 158.940 ;
        RECT 136.110 158.755 136.400 158.800 ;
        RECT 138.210 158.755 138.500 158.800 ;
        RECT 139.780 158.755 140.070 158.800 ;
        RECT 140.300 158.800 144.120 158.940 ;
        RECT 130.090 158.600 130.410 158.660 ;
        RECT 128.800 158.460 130.410 158.600 ;
        RECT 121.825 158.415 122.115 158.460 ;
        RECT 123.650 158.400 123.970 158.460 ;
        RECT 130.090 158.400 130.410 158.460 ;
        RECT 132.850 158.600 133.170 158.660 ;
        RECT 140.300 158.600 140.440 158.800 ;
        RECT 144.810 158.740 145.130 159.000 ;
        RECT 132.850 158.460 140.440 158.600 ;
        RECT 132.850 158.400 133.170 158.460 ;
        RECT 142.510 158.400 142.830 158.660 ;
        RECT 17.320 157.780 147.040 158.260 ;
        RECT 36.710 157.380 37.030 157.640 ;
        RECT 37.645 157.580 37.935 157.625 ;
        RECT 39.470 157.580 39.790 157.640 ;
        RECT 37.645 157.440 39.790 157.580 ;
        RECT 37.645 157.395 37.935 157.440 ;
        RECT 39.470 157.380 39.790 157.440 ;
        RECT 78.585 157.580 78.875 157.625 ;
        RECT 79.490 157.580 79.810 157.640 ;
        RECT 78.585 157.440 79.810 157.580 ;
        RECT 78.585 157.395 78.875 157.440 ;
        RECT 79.490 157.380 79.810 157.440 ;
        RECT 79.965 157.580 80.255 157.625 ;
        RECT 82.710 157.580 83.030 157.640 ;
        RECT 79.965 157.440 83.030 157.580 ;
        RECT 79.965 157.395 80.255 157.440 ;
        RECT 82.710 157.380 83.030 157.440 ;
        RECT 97.445 157.580 97.735 157.625 ;
        RECT 97.890 157.580 98.210 157.640 ;
        RECT 97.445 157.440 98.210 157.580 ;
        RECT 97.445 157.395 97.735 157.440 ;
        RECT 97.890 157.380 98.210 157.440 ;
        RECT 113.530 157.580 113.850 157.640 ;
        RECT 122.745 157.580 123.035 157.625 ;
        RECT 124.110 157.580 124.430 157.640 ;
        RECT 127.790 157.580 128.110 157.640 ;
        RECT 113.530 157.440 122.500 157.580 ;
        RECT 113.530 157.380 113.850 157.440 ;
        RECT 56.030 157.240 56.350 157.300 ;
        RECT 68.465 157.240 68.755 157.285 ;
        RECT 56.030 157.100 68.755 157.240 ;
        RECT 56.030 157.040 56.350 157.100 ;
        RECT 68.465 157.055 68.755 157.100 ;
        RECT 72.170 157.240 72.460 157.285 ;
        RECT 74.270 157.240 74.560 157.285 ;
        RECT 75.840 157.240 76.130 157.285 ;
        RECT 117.670 157.240 117.990 157.300 ;
        RECT 72.170 157.100 76.130 157.240 ;
        RECT 72.170 157.055 72.460 157.100 ;
        RECT 74.270 157.055 74.560 157.100 ;
        RECT 75.840 157.055 76.130 157.100 ;
        RECT 117.300 157.100 117.990 157.240 ;
        RECT 62.930 156.900 63.250 156.960 ;
        RECT 66.165 156.900 66.455 156.945 ;
        RECT 62.930 156.760 66.455 156.900 ;
        RECT 62.930 156.700 63.250 156.760 ;
        RECT 66.165 156.715 66.455 156.760 ;
        RECT 71.670 156.700 71.990 156.960 ;
        RECT 72.565 156.900 72.855 156.945 ;
        RECT 73.755 156.900 74.045 156.945 ;
        RECT 76.275 156.900 76.565 156.945 ;
        RECT 72.565 156.760 76.565 156.900 ;
        RECT 72.565 156.715 72.855 156.760 ;
        RECT 73.755 156.715 74.045 156.760 ;
        RECT 76.275 156.715 76.565 156.760 ;
        RECT 96.970 156.900 97.290 156.960 ;
        RECT 117.300 156.945 117.440 157.100 ;
        RECT 117.670 157.040 117.990 157.100 ;
        RECT 118.590 157.240 118.910 157.300 ;
        RECT 118.590 157.100 122.040 157.240 ;
        RECT 118.590 157.040 118.910 157.100 ;
        RECT 96.970 156.760 98.580 156.900 ;
        RECT 96.970 156.700 97.290 156.760 ;
        RECT 57.410 156.560 57.730 156.620 ;
        RECT 58.805 156.560 59.095 156.605 ;
        RECT 57.410 156.420 59.095 156.560 ;
        RECT 57.410 156.360 57.730 156.420 ;
        RECT 58.805 156.375 59.095 156.420 ;
        RECT 63.390 156.360 63.710 156.620 ;
        RECT 64.770 156.360 65.090 156.620 ;
        RECT 67.530 156.560 67.850 156.620 ;
        RECT 70.305 156.560 70.595 156.605 ;
        RECT 67.530 156.420 70.595 156.560 ;
        RECT 67.530 156.360 67.850 156.420 ;
        RECT 70.305 156.375 70.595 156.420 ;
        RECT 71.225 156.560 71.515 156.605 ;
        RECT 71.225 156.420 74.200 156.560 ;
        RECT 71.225 156.375 71.515 156.420 ;
        RECT 74.060 156.280 74.200 156.420 ;
        RECT 97.430 156.360 97.750 156.620 ;
        RECT 98.440 156.605 98.580 156.760 ;
        RECT 117.225 156.715 117.515 156.945 ;
        RECT 98.365 156.375 98.655 156.605 ;
        RECT 109.850 156.560 110.170 156.620 ;
        RECT 112.165 156.560 112.455 156.605 ;
        RECT 109.850 156.420 112.455 156.560 ;
        RECT 109.850 156.360 110.170 156.420 ;
        RECT 112.165 156.375 112.455 156.420 ;
        RECT 115.830 156.360 116.150 156.620 ;
        RECT 116.765 156.560 117.055 156.605 ;
        RECT 116.380 156.420 117.055 156.560 ;
        RECT 116.380 156.280 116.520 156.420 ;
        RECT 116.765 156.375 117.055 156.420 ;
        RECT 117.670 156.360 117.990 156.620 ;
        RECT 118.145 156.560 118.435 156.605 ;
        RECT 118.590 156.560 118.910 156.620 ;
        RECT 120.430 156.560 120.750 156.620 ;
        RECT 121.900 156.605 122.040 157.100 ;
        RECT 122.360 156.900 122.500 157.440 ;
        RECT 122.745 157.440 128.110 157.580 ;
        RECT 122.745 157.395 123.035 157.440 ;
        RECT 124.110 157.380 124.430 157.440 ;
        RECT 127.790 157.380 128.110 157.440 ;
        RECT 129.645 157.580 129.935 157.625 ;
        RECT 131.485 157.580 131.775 157.625 ;
        RECT 129.645 157.440 131.240 157.580 ;
        RECT 129.645 157.395 129.935 157.440 ;
        RECT 131.100 157.240 131.240 157.440 ;
        RECT 131.485 157.440 135.840 157.580 ;
        RECT 131.485 157.395 131.775 157.440 ;
        RECT 134.245 157.240 134.535 157.285 ;
        RECT 131.100 157.100 134.535 157.240 ;
        RECT 134.245 157.055 134.535 157.100 ;
        RECT 127.790 156.900 128.110 156.960 ;
        RECT 129.185 156.900 129.475 156.945 ;
        RECT 129.630 156.900 129.950 156.960 ;
        RECT 122.360 156.760 122.960 156.900 ;
        RECT 122.820 156.605 122.960 156.760 ;
        RECT 127.790 156.760 129.950 156.900 ;
        RECT 127.790 156.700 128.110 156.760 ;
        RECT 129.185 156.715 129.475 156.760 ;
        RECT 129.630 156.700 129.950 156.760 ;
        RECT 132.390 156.900 132.710 156.960 ;
        RECT 133.785 156.900 134.075 156.945 ;
        RECT 132.390 156.760 134.075 156.900 ;
        RECT 135.700 156.900 135.840 157.440 ;
        RECT 136.990 157.380 137.310 157.640 ;
        RECT 139.765 156.900 140.055 156.945 ;
        RECT 142.510 156.900 142.830 156.960 ;
        RECT 143.905 156.900 144.195 156.945 ;
        RECT 135.700 156.760 140.055 156.900 ;
        RECT 132.390 156.700 132.710 156.760 ;
        RECT 133.785 156.715 134.075 156.760 ;
        RECT 139.765 156.715 140.055 156.760 ;
        RECT 140.760 156.760 144.195 156.900 ;
        RECT 118.145 156.420 120.750 156.560 ;
        RECT 118.145 156.375 118.435 156.420 ;
        RECT 118.590 156.360 118.910 156.420 ;
        RECT 120.430 156.360 120.750 156.420 ;
        RECT 121.825 156.375 122.115 156.605 ;
        RECT 122.745 156.560 123.035 156.605 ;
        RECT 123.650 156.560 123.970 156.620 ;
        RECT 122.745 156.420 123.970 156.560 ;
        RECT 122.745 156.375 123.035 156.420 ;
        RECT 123.650 156.360 123.970 156.420 ;
        RECT 125.505 156.560 125.795 156.605 ;
        RECT 128.710 156.560 129.030 156.620 ;
        RECT 125.505 156.420 129.030 156.560 ;
        RECT 125.505 156.375 125.795 156.420 ;
        RECT 128.710 156.360 129.030 156.420 ;
        RECT 130.550 156.360 130.870 156.620 ;
        RECT 131.010 156.560 131.330 156.620 ;
        RECT 134.230 156.560 134.550 156.620 ;
        RECT 134.705 156.560 134.995 156.605 ;
        RECT 131.010 156.420 134.995 156.560 ;
        RECT 131.010 156.360 131.330 156.420 ;
        RECT 134.230 156.360 134.550 156.420 ;
        RECT 134.705 156.375 134.995 156.420 ;
        RECT 135.150 156.360 135.470 156.620 ;
        RECT 135.625 156.560 135.915 156.605 ;
        RECT 140.760 156.560 140.900 156.760 ;
        RECT 142.510 156.700 142.830 156.760 ;
        RECT 143.905 156.715 144.195 156.760 ;
        RECT 135.625 156.420 140.900 156.560 ;
        RECT 135.625 156.375 135.915 156.420 ;
        RECT 37.565 156.220 37.855 156.265 ;
        RECT 38.090 156.220 38.410 156.280 ;
        RECT 37.565 156.080 38.410 156.220 ;
        RECT 37.565 156.035 37.855 156.080 ;
        RECT 38.090 156.020 38.410 156.080 ;
        RECT 38.550 156.020 38.870 156.280 ;
        RECT 61.550 156.220 61.870 156.280 ;
        RECT 62.485 156.220 62.775 156.265 ;
        RECT 61.550 156.080 62.775 156.220 ;
        RECT 61.550 156.020 61.870 156.080 ;
        RECT 62.485 156.035 62.775 156.080 ;
        RECT 64.325 156.220 64.615 156.265 ;
        RECT 67.070 156.220 67.390 156.280 ;
        RECT 64.325 156.080 67.390 156.220 ;
        RECT 64.325 156.035 64.615 156.080 ;
        RECT 67.070 156.020 67.390 156.080 ;
        RECT 68.005 156.035 68.295 156.265 ;
        RECT 69.370 156.220 69.690 156.280 ;
        RECT 73.050 156.265 73.370 156.280 ;
        RECT 70.765 156.220 71.055 156.265 ;
        RECT 69.370 156.080 71.055 156.220 ;
        RECT 62.010 155.680 62.330 155.940 ;
        RECT 64.770 155.880 65.090 155.940 ;
        RECT 68.080 155.880 68.220 156.035 ;
        RECT 69.370 156.020 69.690 156.080 ;
        RECT 70.765 156.035 71.055 156.080 ;
        RECT 73.020 156.035 73.370 156.265 ;
        RECT 73.050 156.020 73.370 156.035 ;
        RECT 73.970 156.020 74.290 156.280 ;
        RECT 74.890 156.220 75.210 156.280 ;
        RECT 79.805 156.220 80.095 156.265 ;
        RECT 80.410 156.220 80.730 156.280 ;
        RECT 74.890 156.080 80.730 156.220 ;
        RECT 74.890 156.020 75.210 156.080 ;
        RECT 79.805 156.035 80.095 156.080 ;
        RECT 80.410 156.020 80.730 156.080 ;
        RECT 80.885 156.220 81.175 156.265 ;
        RECT 82.710 156.220 83.030 156.280 ;
        RECT 80.885 156.080 83.030 156.220 ;
        RECT 80.885 156.035 81.175 156.080 ;
        RECT 82.710 156.020 83.030 156.080 ;
        RECT 116.290 156.020 116.610 156.280 ;
        RECT 124.570 156.220 124.890 156.280 ;
        RECT 126.885 156.220 127.175 156.265 ;
        RECT 124.570 156.080 127.175 156.220 ;
        RECT 124.570 156.020 124.890 156.080 ;
        RECT 126.885 156.035 127.175 156.080 ;
        RECT 127.805 156.220 128.095 156.265 ;
        RECT 128.250 156.220 128.570 156.280 ;
        RECT 129.630 156.220 129.950 156.280 ;
        RECT 138.845 156.220 139.135 156.265 ;
        RECT 141.145 156.220 141.435 156.265 ;
        RECT 127.805 156.080 129.400 156.220 ;
        RECT 127.805 156.035 128.095 156.080 ;
        RECT 128.250 156.020 128.570 156.080 ;
        RECT 64.770 155.740 68.220 155.880 ;
        RECT 64.770 155.680 65.090 155.740 ;
        RECT 79.030 155.680 79.350 155.940 ;
        RECT 113.990 155.880 114.310 155.940 ;
        RECT 115.385 155.880 115.675 155.925 ;
        RECT 113.990 155.740 115.675 155.880 ;
        RECT 113.990 155.680 114.310 155.740 ;
        RECT 115.385 155.695 115.675 155.740 ;
        RECT 119.050 155.680 119.370 155.940 ;
        RECT 128.710 155.680 129.030 155.940 ;
        RECT 129.260 155.880 129.400 156.080 ;
        RECT 129.630 156.080 138.600 156.220 ;
        RECT 129.630 156.020 129.950 156.080 ;
        RECT 135.150 155.880 135.470 155.940 ;
        RECT 129.260 155.740 135.470 155.880 ;
        RECT 135.150 155.680 135.470 155.740 ;
        RECT 136.545 155.880 136.835 155.925 ;
        RECT 137.910 155.880 138.230 155.940 ;
        RECT 136.545 155.740 138.230 155.880 ;
        RECT 138.460 155.880 138.600 156.080 ;
        RECT 138.845 156.080 141.435 156.220 ;
        RECT 138.845 156.035 139.135 156.080 ;
        RECT 141.145 156.035 141.435 156.080 ;
        RECT 139.305 155.880 139.595 155.925 ;
        RECT 138.460 155.740 139.595 155.880 ;
        RECT 136.545 155.695 136.835 155.740 ;
        RECT 137.910 155.680 138.230 155.740 ;
        RECT 139.305 155.695 139.595 155.740 ;
        RECT 17.320 155.060 147.040 155.540 ;
        RECT 57.410 154.660 57.730 154.920 ;
        RECT 57.885 154.675 58.175 154.905 ;
        RECT 62.470 154.860 62.790 154.920 ;
        RECT 59.800 154.720 62.790 154.860 ;
        RECT 57.960 154.520 58.100 154.675 ;
        RECT 59.800 154.520 59.940 154.720 ;
        RECT 62.470 154.660 62.790 154.720 ;
        RECT 68.465 154.860 68.755 154.905 ;
        RECT 73.050 154.860 73.370 154.920 ;
        RECT 68.465 154.720 73.370 154.860 ;
        RECT 68.465 154.675 68.755 154.720 ;
        RECT 73.050 154.660 73.370 154.720 ;
        RECT 82.710 154.660 83.030 154.920 ;
        RECT 109.850 154.660 110.170 154.920 ;
        RECT 111.245 154.675 111.535 154.905 ;
        RECT 114.465 154.860 114.755 154.905 ;
        RECT 113.160 154.720 114.755 154.860 ;
        RECT 57.960 154.380 59.940 154.520 ;
        RECT 60.140 154.520 60.430 154.565 ;
        RECT 62.010 154.520 62.330 154.580 ;
        RECT 79.030 154.520 79.350 154.580 ;
        RECT 60.140 154.380 62.330 154.520 ;
        RECT 60.140 154.335 60.430 154.380 ;
        RECT 62.010 154.320 62.330 154.380 ;
        RECT 72.680 154.380 79.350 154.520 ;
        RECT 82.800 154.520 82.940 154.660 ;
        RECT 87.785 154.520 88.075 154.565 ;
        RECT 82.800 154.380 88.075 154.520 ;
        RECT 16.010 154.180 16.330 154.240 ;
        RECT 18.785 154.180 19.075 154.225 ;
        RECT 16.010 154.040 19.075 154.180 ;
        RECT 16.010 153.980 16.330 154.040 ;
        RECT 18.785 153.995 19.075 154.040 ;
        RECT 56.030 153.980 56.350 154.240 ;
        RECT 58.345 153.995 58.635 154.225 ;
        RECT 59.250 154.180 59.570 154.240 ;
        RECT 66.165 154.180 66.455 154.225 ;
        RECT 70.750 154.180 71.070 154.240 ;
        RECT 72.680 154.225 72.820 154.380 ;
        RECT 79.030 154.320 79.350 154.380 ;
        RECT 59.250 154.040 64.080 154.180 ;
        RECT 19.705 153.500 19.995 153.545 ;
        RECT 57.870 153.500 58.190 153.560 ;
        RECT 19.705 153.360 58.190 153.500 ;
        RECT 19.705 153.315 19.995 153.360 ;
        RECT 57.870 153.300 58.190 153.360 ;
        RECT 58.420 153.160 58.560 153.995 ;
        RECT 59.250 153.980 59.570 154.040 ;
        RECT 58.790 153.640 59.110 153.900 ;
        RECT 59.685 153.840 59.975 153.885 ;
        RECT 60.875 153.840 61.165 153.885 ;
        RECT 63.395 153.840 63.685 153.885 ;
        RECT 59.685 153.700 63.685 153.840 ;
        RECT 63.940 153.840 64.080 154.040 ;
        RECT 66.165 154.040 71.070 154.180 ;
        RECT 66.165 153.995 66.455 154.040 ;
        RECT 70.750 153.980 71.070 154.040 ;
        RECT 72.605 153.995 72.895 154.225 ;
        RECT 77.160 154.180 77.450 154.225 ;
        RECT 85.470 154.180 85.790 154.240 ;
        RECT 86.020 154.225 86.160 154.380 ;
        RECT 87.785 154.335 88.075 154.380 ;
        RECT 104.300 154.520 104.590 154.565 ;
        RECT 111.320 154.520 111.460 154.675 ;
        RECT 104.300 154.380 111.460 154.520 ;
        RECT 104.300 154.335 104.590 154.380 ;
        RECT 112.610 154.320 112.930 154.580 ;
        RECT 113.160 154.565 113.300 154.720 ;
        RECT 114.465 154.675 114.755 154.720 ;
        RECT 117.225 154.860 117.515 154.905 ;
        RECT 117.670 154.860 117.990 154.920 ;
        RECT 117.225 154.720 117.990 154.860 ;
        RECT 117.225 154.675 117.515 154.720 ;
        RECT 117.670 154.660 117.990 154.720 ;
        RECT 123.665 154.860 123.955 154.905 ;
        RECT 129.630 154.860 129.950 154.920 ;
        RECT 123.665 154.720 129.950 154.860 ;
        RECT 123.665 154.675 123.955 154.720 ;
        RECT 129.630 154.660 129.950 154.720 ;
        RECT 130.565 154.860 130.855 154.905 ;
        RECT 132.850 154.860 133.170 154.920 ;
        RECT 130.565 154.720 133.170 154.860 ;
        RECT 130.565 154.675 130.855 154.720 ;
        RECT 132.850 154.660 133.170 154.720 ;
        RECT 133.325 154.860 133.615 154.905 ;
        RECT 143.445 154.860 143.735 154.905 ;
        RECT 143.890 154.860 144.210 154.920 ;
        RECT 133.325 154.720 142.280 154.860 ;
        RECT 133.325 154.675 133.615 154.720 ;
        RECT 113.085 154.335 113.375 154.565 ;
        RECT 118.145 154.520 118.435 154.565 ;
        RECT 119.510 154.520 119.830 154.580 ;
        RECT 127.790 154.520 128.110 154.580 ;
        RECT 140.670 154.520 140.990 154.580 ;
        RECT 142.140 154.520 142.280 154.720 ;
        RECT 143.445 154.720 144.210 154.860 ;
        RECT 143.445 154.675 143.735 154.720 ;
        RECT 143.890 154.660 144.210 154.720 ;
        RECT 144.810 154.660 145.130 154.920 ;
        RECT 145.270 154.520 145.590 154.580 ;
        RECT 115.460 154.380 128.110 154.520 ;
        RECT 77.160 154.040 85.790 154.180 ;
        RECT 77.160 153.995 77.450 154.040 ;
        RECT 85.470 153.980 85.790 154.040 ;
        RECT 85.945 153.995 86.235 154.225 ;
        RECT 86.865 153.995 87.155 154.225 ;
        RECT 88.690 154.180 89.010 154.240 ;
        RECT 90.545 154.180 90.835 154.225 ;
        RECT 88.690 154.040 90.835 154.180 ;
        RECT 68.910 153.840 69.230 153.900 ;
        RECT 69.385 153.840 69.675 153.885 ;
        RECT 63.940 153.700 69.675 153.840 ;
        RECT 59.685 153.655 59.975 153.700 ;
        RECT 60.875 153.655 61.165 153.700 ;
        RECT 63.395 153.655 63.685 153.700 ;
        RECT 68.910 153.640 69.230 153.700 ;
        RECT 69.385 153.655 69.675 153.700 ;
        RECT 71.670 153.840 71.990 153.900 ;
        RECT 73.510 153.840 73.830 153.900 ;
        RECT 75.825 153.840 76.115 153.885 ;
        RECT 71.670 153.700 76.115 153.840 ;
        RECT 71.670 153.640 71.990 153.700 ;
        RECT 73.510 153.640 73.830 153.700 ;
        RECT 75.825 153.655 76.115 153.700 ;
        RECT 76.705 153.840 76.995 153.885 ;
        RECT 77.895 153.840 78.185 153.885 ;
        RECT 80.415 153.840 80.705 153.885 ;
        RECT 76.705 153.700 80.705 153.840 ;
        RECT 76.705 153.655 76.995 153.700 ;
        RECT 77.895 153.655 78.185 153.700 ;
        RECT 80.415 153.655 80.705 153.700 ;
        RECT 80.870 153.840 81.190 153.900 ;
        RECT 86.390 153.840 86.710 153.900 ;
        RECT 86.940 153.840 87.080 153.995 ;
        RECT 88.690 153.980 89.010 154.040 ;
        RECT 90.545 153.995 90.835 154.040 ;
        RECT 101.110 154.180 101.430 154.240 ;
        RECT 102.965 154.180 103.255 154.225 ;
        RECT 101.110 154.040 103.255 154.180 ;
        RECT 101.110 153.980 101.430 154.040 ;
        RECT 102.965 153.995 103.255 154.040 ;
        RECT 112.165 153.995 112.455 154.225 ;
        RECT 80.870 153.700 87.080 153.840 ;
        RECT 92.845 153.840 93.135 153.885 ;
        RECT 93.290 153.840 93.610 153.900 ;
        RECT 92.845 153.700 93.610 153.840 ;
        RECT 80.870 153.640 81.190 153.700 ;
        RECT 86.390 153.640 86.710 153.700 ;
        RECT 92.845 153.655 93.135 153.700 ;
        RECT 93.290 153.640 93.610 153.700 ;
        RECT 103.845 153.840 104.135 153.885 ;
        RECT 105.035 153.840 105.325 153.885 ;
        RECT 107.555 153.840 107.845 153.885 ;
        RECT 103.845 153.700 107.845 153.840 ;
        RECT 112.240 153.840 112.380 153.995 ;
        RECT 113.990 153.980 114.310 154.240 ;
        RECT 115.460 153.840 115.600 154.380 ;
        RECT 118.145 154.335 118.435 154.380 ;
        RECT 119.510 154.320 119.830 154.380 ;
        RECT 127.790 154.320 128.110 154.380 ;
        RECT 132.020 154.380 141.820 154.520 ;
        RECT 142.140 154.380 145.590 154.520 ;
        RECT 116.290 153.980 116.610 154.240 ;
        RECT 116.765 153.995 117.055 154.225 ;
        RECT 118.590 154.180 118.910 154.240 ;
        RECT 119.065 154.180 119.355 154.225 ;
        RECT 118.590 154.040 119.355 154.180 ;
        RECT 112.240 153.700 115.600 153.840 ;
        RECT 103.845 153.655 104.135 153.700 ;
        RECT 105.035 153.655 105.325 153.700 ;
        RECT 107.555 153.655 107.845 153.700 ;
        RECT 115.830 153.640 116.150 153.900 ;
        RECT 116.840 153.840 116.980 153.995 ;
        RECT 118.590 153.980 118.910 154.040 ;
        RECT 119.065 153.995 119.355 154.040 ;
        RECT 119.985 154.180 120.275 154.225 ;
        RECT 120.905 154.180 121.195 154.225 ;
        RECT 119.985 154.040 121.195 154.180 ;
        RECT 119.985 153.995 120.275 154.040 ;
        RECT 120.905 153.995 121.195 154.040 ;
        RECT 121.350 154.180 121.670 154.240 ;
        RECT 121.825 154.180 122.115 154.225 ;
        RECT 121.350 154.040 122.115 154.180 ;
        RECT 121.350 153.980 121.670 154.040 ;
        RECT 121.825 153.995 122.115 154.040 ;
        RECT 122.270 153.980 122.590 154.240 ;
        RECT 122.745 154.180 123.035 154.225 ;
        RECT 123.650 154.180 123.970 154.240 ;
        RECT 122.745 154.040 123.970 154.180 ;
        RECT 122.745 153.995 123.035 154.040 ;
        RECT 123.650 153.980 123.970 154.040 ;
        RECT 129.645 154.180 129.935 154.225 ;
        RECT 132.020 154.180 132.160 154.380 ;
        RECT 140.670 154.320 140.990 154.380 ;
        RECT 129.645 154.040 132.160 154.180 ;
        RECT 129.645 153.995 129.935 154.040 ;
        RECT 132.390 153.980 132.710 154.240 ;
        RECT 134.230 153.980 134.550 154.240 ;
        RECT 136.530 153.980 136.850 154.240 ;
        RECT 141.680 154.225 141.820 154.380 ;
        RECT 145.270 154.320 145.590 154.380 ;
        RECT 137.005 154.180 137.295 154.225 ;
        RECT 138.845 154.180 139.135 154.225 ;
        RECT 137.005 154.040 139.135 154.180 ;
        RECT 137.005 153.995 137.295 154.040 ;
        RECT 138.845 153.995 139.135 154.040 ;
        RECT 141.605 153.995 141.895 154.225 ;
        RECT 142.525 154.180 142.815 154.225 ;
        RECT 143.430 154.180 143.750 154.240 ;
        RECT 142.525 154.040 143.750 154.180 ;
        RECT 142.525 153.995 142.815 154.040 ;
        RECT 143.430 153.980 143.750 154.040 ;
        RECT 143.905 154.180 144.195 154.225 ;
        RECT 143.905 154.040 145.040 154.180 ;
        RECT 143.905 153.995 144.195 154.040 ;
        RECT 127.790 153.840 128.110 153.900 ;
        RECT 137.465 153.840 137.755 153.885 ;
        RECT 116.840 153.700 117.440 153.840 ;
        RECT 59.290 153.500 59.580 153.545 ;
        RECT 61.390 153.500 61.680 153.545 ;
        RECT 62.960 153.500 63.250 153.545 ;
        RECT 59.290 153.360 63.250 153.500 ;
        RECT 59.290 153.315 59.580 153.360 ;
        RECT 61.390 153.315 61.680 153.360 ;
        RECT 62.960 153.315 63.250 153.360 ;
        RECT 67.530 153.300 67.850 153.560 ;
        RECT 69.845 153.500 70.135 153.545 ;
        RECT 74.890 153.500 75.210 153.560 ;
        RECT 69.845 153.360 75.210 153.500 ;
        RECT 69.845 153.315 70.135 153.360 ;
        RECT 74.890 153.300 75.210 153.360 ;
        RECT 76.310 153.500 76.600 153.545 ;
        RECT 78.410 153.500 78.700 153.545 ;
        RECT 79.980 153.500 80.270 153.545 ;
        RECT 76.310 153.360 80.270 153.500 ;
        RECT 76.310 153.315 76.600 153.360 ;
        RECT 78.410 153.315 78.700 153.360 ;
        RECT 79.980 153.315 80.270 153.360 ;
        RECT 103.450 153.500 103.740 153.545 ;
        RECT 105.550 153.500 105.840 153.545 ;
        RECT 107.120 153.500 107.410 153.545 ;
        RECT 103.450 153.360 107.410 153.500 ;
        RECT 103.450 153.315 103.740 153.360 ;
        RECT 105.550 153.315 105.840 153.360 ;
        RECT 107.120 153.315 107.410 153.360 ;
        RECT 112.150 153.500 112.470 153.560 ;
        RECT 117.300 153.500 117.440 153.700 ;
        RECT 127.790 153.700 137.755 153.840 ;
        RECT 127.790 153.640 128.110 153.700 ;
        RECT 137.465 153.655 137.755 153.700 ;
        RECT 121.350 153.500 121.670 153.560 ;
        RECT 130.550 153.500 130.870 153.560 ;
        RECT 112.150 153.360 116.980 153.500 ;
        RECT 117.300 153.360 121.670 153.500 ;
        RECT 112.150 153.300 112.470 153.360 ;
        RECT 60.630 153.160 60.950 153.220 ;
        RECT 58.420 153.020 60.950 153.160 ;
        RECT 60.630 152.960 60.950 153.020 ;
        RECT 65.705 153.160 65.995 153.205 ;
        RECT 67.070 153.160 67.390 153.220 ;
        RECT 67.990 153.160 68.310 153.220 ;
        RECT 65.705 153.020 68.310 153.160 ;
        RECT 65.705 152.975 65.995 153.020 ;
        RECT 67.070 152.960 67.390 153.020 ;
        RECT 67.990 152.960 68.310 153.020 ;
        RECT 71.670 152.960 71.990 153.220 ;
        RECT 75.365 153.160 75.655 153.205 ;
        RECT 75.810 153.160 76.130 153.220 ;
        RECT 75.365 153.020 76.130 153.160 ;
        RECT 75.365 152.975 75.655 153.020 ;
        RECT 75.810 152.960 76.130 153.020 ;
        RECT 83.170 152.960 83.490 153.220 ;
        RECT 88.230 152.960 88.550 153.220 ;
        RECT 115.370 152.960 115.690 153.220 ;
        RECT 116.840 153.160 116.980 153.360 ;
        RECT 121.350 153.300 121.670 153.360 ;
        RECT 123.280 153.360 130.870 153.500 ;
        RECT 123.280 153.160 123.420 153.360 ;
        RECT 130.550 153.300 130.870 153.360 ;
        RECT 131.485 153.500 131.775 153.545 ;
        RECT 142.970 153.500 143.290 153.560 ;
        RECT 131.485 153.360 143.290 153.500 ;
        RECT 131.485 153.315 131.775 153.360 ;
        RECT 142.970 153.300 143.290 153.360 ;
        RECT 116.840 153.020 123.420 153.160 ;
        RECT 123.650 153.160 123.970 153.220 ;
        RECT 124.570 153.160 124.890 153.220 ;
        RECT 133.310 153.160 133.630 153.220 ;
        RECT 123.650 153.020 133.630 153.160 ;
        RECT 123.650 152.960 123.970 153.020 ;
        RECT 124.570 152.960 124.890 153.020 ;
        RECT 133.310 152.960 133.630 153.020 ;
        RECT 134.705 153.160 134.995 153.205 ;
        RECT 135.150 153.160 135.470 153.220 ;
        RECT 134.705 153.020 135.470 153.160 ;
        RECT 134.705 152.975 134.995 153.020 ;
        RECT 135.150 152.960 135.470 153.020 ;
        RECT 137.910 153.160 138.230 153.220 ;
        RECT 144.900 153.160 145.040 154.040 ;
        RECT 137.910 153.020 145.040 153.160 ;
        RECT 137.910 152.960 138.230 153.020 ;
        RECT 17.320 152.340 147.040 152.820 ;
        RECT 35.330 152.140 35.650 152.200 ;
        RECT 37.185 152.140 37.475 152.185 ;
        RECT 35.330 152.000 37.475 152.140 ;
        RECT 35.330 151.940 35.650 152.000 ;
        RECT 37.185 151.955 37.475 152.000 ;
        RECT 35.790 151.800 36.110 151.860 ;
        RECT 36.265 151.800 36.555 151.845 ;
        RECT 35.790 151.660 36.555 151.800 ;
        RECT 37.260 151.800 37.400 151.955 ;
        RECT 47.750 151.940 48.070 152.200 ;
        RECT 57.425 152.140 57.715 152.185 ;
        RECT 60.630 152.140 60.950 152.200 ;
        RECT 57.425 152.000 60.950 152.140 ;
        RECT 57.425 151.955 57.715 152.000 ;
        RECT 60.630 151.940 60.950 152.000 ;
        RECT 63.390 152.140 63.710 152.200 ;
        RECT 65.230 152.140 65.550 152.200 ;
        RECT 65.705 152.140 65.995 152.185 ;
        RECT 63.390 152.000 65.995 152.140 ;
        RECT 63.390 151.940 63.710 152.000 ;
        RECT 65.230 151.940 65.550 152.000 ;
        RECT 65.705 151.955 65.995 152.000 ;
        RECT 56.490 151.800 56.810 151.860 ;
        RECT 37.260 151.660 56.810 151.800 ;
        RECT 35.790 151.600 36.110 151.660 ;
        RECT 36.265 151.615 36.555 151.660 ;
        RECT 56.490 151.600 56.810 151.660 ;
        RECT 59.290 151.800 59.580 151.845 ;
        RECT 61.390 151.800 61.680 151.845 ;
        RECT 62.960 151.800 63.250 151.845 ;
        RECT 59.290 151.660 63.250 151.800 ;
        RECT 59.290 151.615 59.580 151.660 ;
        RECT 61.390 151.615 61.680 151.660 ;
        RECT 62.960 151.615 63.250 151.660 ;
        RECT 39.010 151.460 39.330 151.520 ;
        RECT 35.880 151.320 41.080 151.460 ;
        RECT 32.570 151.120 32.890 151.180 ;
        RECT 35.880 151.165 36.020 151.320 ;
        RECT 39.010 151.260 39.330 151.320 ;
        RECT 35.805 151.120 36.095 151.165 ;
        RECT 38.550 151.120 38.870 151.180 ;
        RECT 40.940 151.165 41.080 151.320 ;
        RECT 58.790 151.260 59.110 151.520 ;
        RECT 59.685 151.460 59.975 151.505 ;
        RECT 60.875 151.460 61.165 151.505 ;
        RECT 63.395 151.460 63.685 151.505 ;
        RECT 59.685 151.320 63.685 151.460 ;
        RECT 65.780 151.460 65.920 151.955 ;
        RECT 70.750 151.940 71.070 152.200 ;
        RECT 85.470 151.940 85.790 152.200 ;
        RECT 88.230 152.140 88.550 152.200 ;
        RECT 89.165 152.140 89.455 152.185 ;
        RECT 94.210 152.140 94.530 152.200 ;
        RECT 101.110 152.140 101.430 152.200 ;
        RECT 88.230 152.000 89.455 152.140 ;
        RECT 88.230 151.940 88.550 152.000 ;
        RECT 89.165 151.955 89.455 152.000 ;
        RECT 90.620 152.000 105.940 152.140 ;
        RECT 74.930 151.800 75.220 151.845 ;
        RECT 77.030 151.800 77.320 151.845 ;
        RECT 78.600 151.800 78.890 151.845 ;
        RECT 74.930 151.660 78.890 151.800 ;
        RECT 74.930 151.615 75.220 151.660 ;
        RECT 77.030 151.615 77.320 151.660 ;
        RECT 78.600 151.615 78.890 151.660 ;
        RECT 70.290 151.460 70.610 151.520 ;
        RECT 73.510 151.460 73.830 151.520 ;
        RECT 90.620 151.505 90.760 152.000 ;
        RECT 94.210 151.940 94.530 152.000 ;
        RECT 101.110 151.940 101.430 152.000 ;
        RECT 91.030 151.800 91.320 151.845 ;
        RECT 93.130 151.800 93.420 151.845 ;
        RECT 94.700 151.800 94.990 151.845 ;
        RECT 91.030 151.660 94.990 151.800 ;
        RECT 91.030 151.615 91.320 151.660 ;
        RECT 93.130 151.615 93.420 151.660 ;
        RECT 94.700 151.615 94.990 151.660 ;
        RECT 97.430 151.600 97.750 151.860 ;
        RECT 101.570 151.800 101.860 151.845 ;
        RECT 103.140 151.800 103.430 151.845 ;
        RECT 105.240 151.800 105.530 151.845 ;
        RECT 101.570 151.660 105.530 151.800 ;
        RECT 101.570 151.615 101.860 151.660 ;
        RECT 103.140 151.615 103.430 151.660 ;
        RECT 105.240 151.615 105.530 151.660 ;
        RECT 105.800 151.505 105.940 152.000 ;
        RECT 108.010 151.940 108.330 152.200 ;
        RECT 115.830 152.140 116.150 152.200 ;
        RECT 118.590 152.140 118.910 152.200 ;
        RECT 115.830 152.000 118.910 152.140 ;
        RECT 115.830 151.940 116.150 152.000 ;
        RECT 118.590 151.940 118.910 152.000 ;
        RECT 127.790 151.940 128.110 152.200 ;
        RECT 132.390 152.140 132.710 152.200 ;
        RECT 138.830 152.140 139.150 152.200 ;
        RECT 132.390 152.000 139.150 152.140 ;
        RECT 132.390 151.940 132.710 152.000 ;
        RECT 138.830 151.940 139.150 152.000 ;
        RECT 140.670 151.940 140.990 152.200 ;
        RECT 109.850 151.800 110.170 151.860 ;
        RECT 116.750 151.800 117.070 151.860 ;
        RECT 109.850 151.660 110.540 151.800 ;
        RECT 109.850 151.600 110.170 151.660 ;
        RECT 110.400 151.505 110.540 151.660 ;
        RECT 110.860 151.660 117.070 151.800 ;
        RECT 118.680 151.800 118.820 151.940 ;
        RECT 123.205 151.800 123.495 151.845 ;
        RECT 126.410 151.800 126.730 151.860 ;
        RECT 118.680 151.660 126.730 151.800 ;
        RECT 110.860 151.520 111.000 151.660 ;
        RECT 116.750 151.600 117.070 151.660 ;
        RECT 123.205 151.615 123.495 151.660 ;
        RECT 126.410 151.600 126.730 151.660 ;
        RECT 134.270 151.800 134.560 151.845 ;
        RECT 136.370 151.800 136.660 151.845 ;
        RECT 137.940 151.800 138.230 151.845 ;
        RECT 134.270 151.660 138.230 151.800 ;
        RECT 134.270 151.615 134.560 151.660 ;
        RECT 136.370 151.615 136.660 151.660 ;
        RECT 137.940 151.615 138.230 151.660 ;
        RECT 74.445 151.460 74.735 151.505 ;
        RECT 65.780 151.320 69.140 151.460 ;
        RECT 59.685 151.275 59.975 151.320 ;
        RECT 60.875 151.275 61.165 151.320 ;
        RECT 63.395 151.275 63.685 151.320 ;
        RECT 40.405 151.120 40.695 151.165 ;
        RECT 32.570 150.980 36.095 151.120 ;
        RECT 32.570 150.920 32.890 150.980 ;
        RECT 35.805 150.935 36.095 150.980 ;
        RECT 36.340 150.980 38.870 151.120 ;
        RECT 33.490 150.780 33.810 150.840 ;
        RECT 34.885 150.780 35.175 150.825 ;
        RECT 36.340 150.780 36.480 150.980 ;
        RECT 38.550 150.920 38.870 150.980 ;
        RECT 39.560 150.980 40.695 151.120 ;
        RECT 39.560 150.840 39.700 150.980 ;
        RECT 40.405 150.935 40.695 150.980 ;
        RECT 40.865 150.935 41.155 151.165 ;
        RECT 33.490 150.640 36.480 150.780 ;
        RECT 33.490 150.580 33.810 150.640 ;
        RECT 34.885 150.595 35.175 150.640 ;
        RECT 38.090 150.580 38.410 150.840 ;
        RECT 39.025 150.780 39.315 150.825 ;
        RECT 39.470 150.780 39.790 150.840 ;
        RECT 39.025 150.640 39.790 150.780 ;
        RECT 39.025 150.595 39.315 150.640 ;
        RECT 39.470 150.580 39.790 150.640 ;
        RECT 39.945 150.780 40.235 150.825 ;
        RECT 40.940 150.780 41.080 150.935 ;
        RECT 41.770 150.920 42.090 151.180 ;
        RECT 54.665 151.120 54.955 151.165 ;
        RECT 55.110 151.120 55.430 151.180 ;
        RECT 54.665 150.980 55.430 151.120 ;
        RECT 54.665 150.935 54.955 150.980 ;
        RECT 55.110 150.920 55.430 150.980 ;
        RECT 55.585 151.120 55.875 151.165 ;
        RECT 56.030 151.120 56.350 151.180 ;
        RECT 64.310 151.120 64.630 151.180 ;
        RECT 55.585 150.980 56.350 151.120 ;
        RECT 57.805 150.995 64.630 151.120 ;
        RECT 55.585 150.935 55.875 150.980 ;
        RECT 56.030 150.920 56.350 150.980 ;
        RECT 57.655 150.980 64.630 150.995 ;
        RECT 39.945 150.640 41.080 150.780 ;
        RECT 46.830 150.780 47.150 150.840 ;
        RECT 46.830 150.640 54.880 150.780 ;
        RECT 39.945 150.595 40.235 150.640 ;
        RECT 46.830 150.580 47.150 150.640 ;
        RECT 54.740 150.500 54.880 150.640 ;
        RECT 56.490 150.580 56.810 150.840 ;
        RECT 57.655 150.765 57.945 150.980 ;
        RECT 64.310 150.920 64.630 150.980 ;
        RECT 64.770 151.120 65.090 151.180 ;
        RECT 67.085 151.120 67.375 151.165 ;
        RECT 64.770 150.980 67.375 151.120 ;
        RECT 64.770 150.920 65.090 150.980 ;
        RECT 67.085 150.935 67.375 150.980 ;
        RECT 67.990 150.920 68.310 151.180 ;
        RECT 68.450 150.920 68.770 151.180 ;
        RECT 69.000 151.165 69.140 151.320 ;
        RECT 70.290 151.320 74.735 151.460 ;
        RECT 70.290 151.260 70.610 151.320 ;
        RECT 73.510 151.260 73.830 151.320 ;
        RECT 74.445 151.275 74.735 151.320 ;
        RECT 75.325 151.460 75.615 151.505 ;
        RECT 76.515 151.460 76.805 151.505 ;
        RECT 79.035 151.460 79.325 151.505 ;
        RECT 75.325 151.320 79.325 151.460 ;
        RECT 75.325 151.275 75.615 151.320 ;
        RECT 76.515 151.275 76.805 151.320 ;
        RECT 79.035 151.275 79.325 151.320 ;
        RECT 82.725 151.460 83.015 151.505 ;
        RECT 82.725 151.320 87.080 151.460 ;
        RECT 82.725 151.275 83.015 151.320 ;
        RECT 68.925 150.935 69.215 151.165 ;
        RECT 69.845 150.935 70.135 151.165 ;
        RECT 60.030 150.780 60.320 150.825 ;
        RECT 58.420 150.640 60.320 150.780 ;
        RECT 33.950 150.240 34.270 150.500 ;
        RECT 37.105 150.440 37.395 150.485 ;
        RECT 38.565 150.440 38.855 150.485 ;
        RECT 37.105 150.300 38.855 150.440 ;
        RECT 37.105 150.255 37.395 150.300 ;
        RECT 38.565 150.255 38.855 150.300 ;
        RECT 42.705 150.440 42.995 150.485 ;
        RECT 46.370 150.440 46.690 150.500 ;
        RECT 42.705 150.300 46.690 150.440 ;
        RECT 42.705 150.255 42.995 150.300 ;
        RECT 46.370 150.240 46.690 150.300 ;
        RECT 47.290 150.440 47.610 150.500 ;
        RECT 47.845 150.440 48.135 150.485 ;
        RECT 47.290 150.300 48.135 150.440 ;
        RECT 47.290 150.240 47.610 150.300 ;
        RECT 47.845 150.255 48.135 150.300 ;
        RECT 48.685 150.440 48.975 150.485 ;
        RECT 50.510 150.440 50.830 150.500 ;
        RECT 48.685 150.300 50.830 150.440 ;
        RECT 48.685 150.255 48.975 150.300 ;
        RECT 50.510 150.240 50.830 150.300 ;
        RECT 54.650 150.240 54.970 150.500 ;
        RECT 55.125 150.440 55.415 150.485 ;
        RECT 56.950 150.440 57.270 150.500 ;
        RECT 58.420 150.485 58.560 150.640 ;
        RECT 60.030 150.595 60.320 150.640 ;
        RECT 61.090 150.780 61.410 150.840 ;
        RECT 66.165 150.780 66.455 150.825 ;
        RECT 61.090 150.640 66.455 150.780 ;
        RECT 61.090 150.580 61.410 150.640 ;
        RECT 66.165 150.595 66.455 150.640 ;
        RECT 66.610 150.780 66.930 150.840 ;
        RECT 69.920 150.780 70.060 150.935 ;
        RECT 73.970 150.920 74.290 151.180 ;
        RECT 75.810 151.165 76.130 151.180 ;
        RECT 75.780 151.120 76.130 151.165 ;
        RECT 75.615 150.980 76.130 151.120 ;
        RECT 75.780 150.935 76.130 150.980 ;
        RECT 75.810 150.920 76.130 150.935 ;
        RECT 82.250 150.920 82.570 151.180 ;
        RECT 83.170 150.920 83.490 151.180 ;
        RECT 86.390 150.920 86.710 151.180 ;
        RECT 86.940 151.165 87.080 151.320 ;
        RECT 90.490 151.275 90.780 151.505 ;
        RECT 91.425 151.460 91.715 151.505 ;
        RECT 92.615 151.460 92.905 151.505 ;
        RECT 95.135 151.460 95.425 151.505 ;
        RECT 91.425 151.320 95.425 151.460 ;
        RECT 91.425 151.275 91.715 151.320 ;
        RECT 92.615 151.275 92.905 151.320 ;
        RECT 95.135 151.275 95.425 151.320 ;
        RECT 101.135 151.460 101.425 151.505 ;
        RECT 103.655 151.460 103.945 151.505 ;
        RECT 104.845 151.460 105.135 151.505 ;
        RECT 101.135 151.320 105.135 151.460 ;
        RECT 101.135 151.275 101.425 151.320 ;
        RECT 103.655 151.275 103.945 151.320 ;
        RECT 104.845 151.275 105.135 151.320 ;
        RECT 105.725 151.275 106.015 151.505 ;
        RECT 110.325 151.275 110.615 151.505 ;
        RECT 110.770 151.260 111.090 151.520 ;
        RECT 112.610 151.460 112.930 151.520 ;
        RECT 111.780 151.320 112.930 151.460 ;
        RECT 86.865 150.935 87.155 151.165 ;
        RECT 89.150 151.120 89.470 151.180 ;
        RECT 89.625 151.120 89.915 151.165 ;
        RECT 89.150 150.980 89.915 151.120 ;
        RECT 89.150 150.920 89.470 150.980 ;
        RECT 89.625 150.935 89.915 150.980 ;
        RECT 90.085 151.120 90.375 151.165 ;
        RECT 90.990 151.120 91.310 151.180 ;
        RECT 97.890 151.120 98.210 151.180 ;
        RECT 90.085 150.980 98.210 151.120 ;
        RECT 90.085 150.935 90.375 150.980 ;
        RECT 66.610 150.640 70.060 150.780 ;
        RECT 79.030 150.780 79.350 150.840 ;
        RECT 85.485 150.780 85.775 150.825 ;
        RECT 79.030 150.640 85.775 150.780 ;
        RECT 66.610 150.580 66.930 150.640 ;
        RECT 79.030 150.580 79.350 150.640 ;
        RECT 85.485 150.595 85.775 150.640 ;
        RECT 55.125 150.300 57.270 150.440 ;
        RECT 55.125 150.255 55.415 150.300 ;
        RECT 56.950 150.240 57.270 150.300 ;
        RECT 58.345 150.255 58.635 150.485 ;
        RECT 60.630 150.440 60.950 150.500 ;
        RECT 68.925 150.440 69.215 150.485 ;
        RECT 60.630 150.300 69.215 150.440 ;
        RECT 60.630 150.240 60.950 150.300 ;
        RECT 68.925 150.255 69.215 150.300 ;
        RECT 78.570 150.440 78.890 150.500 ;
        RECT 81.345 150.440 81.635 150.485 ;
        RECT 78.570 150.300 81.635 150.440 ;
        RECT 78.570 150.240 78.890 150.300 ;
        RECT 81.345 150.255 81.635 150.300 ;
        RECT 88.230 150.240 88.550 150.500 ;
        RECT 89.700 150.440 89.840 150.935 ;
        RECT 90.990 150.920 91.310 150.980 ;
        RECT 97.890 150.920 98.210 150.980 ;
        RECT 109.865 151.120 110.155 151.165 ;
        RECT 111.780 151.120 111.920 151.320 ;
        RECT 112.610 151.260 112.930 151.320 ;
        RECT 124.110 151.460 124.430 151.520 ;
        RECT 125.505 151.460 125.795 151.505 ;
        RECT 124.110 151.320 125.795 151.460 ;
        RECT 124.110 151.260 124.430 151.320 ;
        RECT 125.505 151.275 125.795 151.320 ;
        RECT 125.950 151.260 126.270 151.520 ;
        RECT 126.885 151.460 127.175 151.505 ;
        RECT 131.010 151.460 131.330 151.520 ;
        RECT 126.885 151.320 131.330 151.460 ;
        RECT 126.885 151.275 127.175 151.320 ;
        RECT 131.010 151.260 131.330 151.320 ;
        RECT 133.770 151.260 134.090 151.520 ;
        RECT 134.665 151.460 134.955 151.505 ;
        RECT 135.855 151.460 136.145 151.505 ;
        RECT 138.375 151.460 138.665 151.505 ;
        RECT 134.665 151.320 138.665 151.460 ;
        RECT 134.665 151.275 134.955 151.320 ;
        RECT 135.855 151.275 136.145 151.320 ;
        RECT 138.375 151.275 138.665 151.320 ;
        RECT 143.430 151.260 143.750 151.520 ;
        RECT 143.890 151.260 144.210 151.520 ;
        RECT 109.865 150.980 111.920 151.120 ;
        RECT 109.865 150.935 110.155 150.980 ;
        RECT 112.150 150.920 112.470 151.180 ;
        RECT 113.085 151.120 113.375 151.165 ;
        RECT 115.370 151.120 115.690 151.180 ;
        RECT 113.085 150.980 115.690 151.120 ;
        RECT 113.085 150.935 113.375 150.980 ;
        RECT 115.370 150.920 115.690 150.980 ;
        RECT 119.065 151.120 119.355 151.165 ;
        RECT 119.510 151.120 119.830 151.180 ;
        RECT 119.065 150.980 119.830 151.120 ;
        RECT 119.065 150.935 119.355 150.980 ;
        RECT 119.510 150.920 119.830 150.980 ;
        RECT 119.985 151.120 120.275 151.165 ;
        RECT 121.810 151.120 122.130 151.180 ;
        RECT 122.745 151.120 123.035 151.165 ;
        RECT 119.985 150.980 123.035 151.120 ;
        RECT 119.985 150.935 120.275 150.980 ;
        RECT 121.810 150.920 122.130 150.980 ;
        RECT 122.745 150.935 123.035 150.980 ;
        RECT 91.880 150.780 92.170 150.825 ;
        RECT 92.830 150.780 93.150 150.840 ;
        RECT 91.880 150.640 93.150 150.780 ;
        RECT 91.880 150.595 92.170 150.640 ;
        RECT 92.830 150.580 93.150 150.640 ;
        RECT 104.330 150.825 104.650 150.840 ;
        RECT 104.330 150.595 104.680 150.825 ;
        RECT 108.470 150.780 108.790 150.840 ;
        RECT 112.625 150.780 112.915 150.825 ;
        RECT 108.470 150.640 112.915 150.780 ;
        RECT 122.820 150.780 122.960 150.935 ;
        RECT 126.410 150.920 126.730 151.180 ;
        RECT 127.790 151.120 128.110 151.180 ;
        RECT 128.265 151.120 128.555 151.165 ;
        RECT 127.790 150.980 128.555 151.120 ;
        RECT 127.790 150.920 128.110 150.980 ;
        RECT 128.265 150.935 128.555 150.980 ;
        RECT 129.185 151.120 129.475 151.165 ;
        RECT 129.630 151.120 129.950 151.180 ;
        RECT 131.470 151.120 131.790 151.180 ;
        RECT 135.150 151.165 135.470 151.180 ;
        RECT 135.120 151.120 135.470 151.165 ;
        RECT 129.185 150.980 131.790 151.120 ;
        RECT 134.955 150.980 135.470 151.120 ;
        RECT 129.185 150.935 129.475 150.980 ;
        RECT 129.630 150.920 129.950 150.980 ;
        RECT 131.470 150.920 131.790 150.980 ;
        RECT 135.120 150.935 135.470 150.980 ;
        RECT 135.150 150.920 135.470 150.935 ;
        RECT 125.490 150.780 125.810 150.840 ;
        RECT 126.500 150.780 126.640 150.920 ;
        RECT 128.725 150.780 129.015 150.825 ;
        RECT 122.820 150.640 126.180 150.780 ;
        RECT 126.500 150.640 129.015 150.780 ;
        RECT 104.330 150.580 104.650 150.595 ;
        RECT 108.470 150.580 108.790 150.640 ;
        RECT 112.625 150.595 112.915 150.640 ;
        RECT 125.490 150.580 125.810 150.640 ;
        RECT 96.050 150.440 96.370 150.500 ;
        RECT 89.700 150.300 96.370 150.440 ;
        RECT 96.050 150.240 96.370 150.300 ;
        RECT 97.430 150.440 97.750 150.500 ;
        RECT 98.825 150.440 99.115 150.485 ;
        RECT 97.430 150.300 99.115 150.440 ;
        RECT 97.430 150.240 97.750 150.300 ;
        RECT 98.825 150.255 99.115 150.300 ;
        RECT 117.210 150.440 117.530 150.500 ;
        RECT 119.525 150.440 119.815 150.485 ;
        RECT 117.210 150.300 119.815 150.440 ;
        RECT 117.210 150.240 117.530 150.300 ;
        RECT 119.525 150.255 119.815 150.300 ;
        RECT 122.730 150.440 123.050 150.500 ;
        RECT 124.110 150.440 124.430 150.500 ;
        RECT 122.730 150.300 124.430 150.440 ;
        RECT 126.040 150.440 126.180 150.640 ;
        RECT 128.725 150.595 129.015 150.640 ;
        RECT 127.790 150.440 128.110 150.500 ;
        RECT 126.040 150.300 128.110 150.440 ;
        RECT 122.730 150.240 123.050 150.300 ;
        RECT 124.110 150.240 124.430 150.300 ;
        RECT 127.790 150.240 128.110 150.300 ;
        RECT 141.130 150.240 141.450 150.500 ;
        RECT 142.970 150.240 143.290 150.500 ;
        RECT 17.320 149.620 147.040 150.100 ;
        RECT 15.890 149.420 16.310 149.560 ;
        RECT 74.430 149.420 74.750 149.480 ;
        RECT 76.745 149.420 77.035 149.465 ;
        RECT 15.890 149.280 73.970 149.420 ;
        RECT 15.890 149.110 16.310 149.280 ;
        RECT 31.205 149.080 31.495 149.125 ;
        RECT 32.125 149.080 32.415 149.125 ;
        RECT 31.205 148.940 32.415 149.080 ;
        RECT 31.205 148.895 31.495 148.940 ;
        RECT 32.125 148.895 32.415 148.940 ;
        RECT 33.205 149.080 33.495 149.125 ;
        RECT 33.950 149.080 34.270 149.140 ;
        RECT 33.205 148.940 34.270 149.080 ;
        RECT 33.205 148.895 33.495 148.940 ;
        RECT 33.950 148.880 34.270 148.940 ;
        RECT 45.465 149.080 45.755 149.125 ;
        RECT 47.290 149.080 47.610 149.140 ;
        RECT 45.465 148.940 47.610 149.080 ;
        RECT 45.465 148.895 45.755 148.940 ;
        RECT 47.290 148.880 47.610 148.940 ;
        RECT 47.750 149.080 48.070 149.140 ;
        RECT 54.650 149.080 54.970 149.140 ;
        RECT 55.125 149.080 55.415 149.125 ;
        RECT 47.750 148.940 53.960 149.080 ;
        RECT 47.750 148.880 48.070 148.940 ;
        RECT 29.350 148.740 29.670 148.800 ;
        RECT 30.745 148.740 31.035 148.785 ;
        RECT 29.350 148.600 31.035 148.740 ;
        RECT 29.350 148.540 29.670 148.600 ;
        RECT 30.745 148.555 31.035 148.600 ;
        RECT 31.665 148.740 31.955 148.785 ;
        RECT 32.570 148.740 32.890 148.800 ;
        RECT 31.665 148.600 32.890 148.740 ;
        RECT 31.665 148.555 31.955 148.600 ;
        RECT 30.820 148.400 30.960 148.555 ;
        RECT 32.570 148.540 32.890 148.600 ;
        RECT 34.425 148.740 34.715 148.785 ;
        RECT 34.870 148.740 35.190 148.800 ;
        RECT 35.790 148.785 36.110 148.800 ;
        RECT 35.760 148.740 36.110 148.785 ;
        RECT 34.425 148.600 35.190 148.740 ;
        RECT 35.595 148.600 36.110 148.740 ;
        RECT 34.425 148.555 34.715 148.600 ;
        RECT 34.870 148.540 35.190 148.600 ;
        RECT 35.760 148.555 36.110 148.600 ;
        RECT 35.790 148.540 36.110 148.555 ;
        RECT 46.370 148.540 46.690 148.800 ;
        RECT 46.830 148.540 47.150 148.800 ;
        RECT 48.225 148.740 48.515 148.785 ;
        RECT 47.380 148.600 48.515 148.740 ;
        RECT 33.490 148.400 33.810 148.460 ;
        RECT 30.820 148.260 33.810 148.400 ;
        RECT 33.490 148.200 33.810 148.260 ;
        RECT 35.305 148.400 35.595 148.445 ;
        RECT 36.495 148.400 36.785 148.445 ;
        RECT 39.015 148.400 39.305 148.445 ;
        RECT 35.305 148.260 39.305 148.400 ;
        RECT 35.305 148.215 35.595 148.260 ;
        RECT 36.495 148.215 36.785 148.260 ;
        RECT 39.015 148.215 39.305 148.260 ;
        RECT 34.410 148.060 34.730 148.120 ;
        RECT 33.120 147.920 34.730 148.060 ;
        RECT 33.120 147.765 33.260 147.920 ;
        RECT 34.410 147.860 34.730 147.920 ;
        RECT 34.910 148.060 35.200 148.105 ;
        RECT 37.010 148.060 37.300 148.105 ;
        RECT 38.580 148.060 38.870 148.105 ;
        RECT 34.910 147.920 38.870 148.060 ;
        RECT 47.380 148.060 47.520 148.600 ;
        RECT 48.225 148.555 48.515 148.600 ;
        RECT 50.050 148.540 50.370 148.800 ;
        RECT 50.510 148.740 50.830 148.800 ;
        RECT 50.510 148.600 51.025 148.740 ;
        RECT 50.510 148.540 50.830 148.600 ;
        RECT 51.430 148.540 51.750 148.800 ;
        RECT 52.350 148.785 52.670 148.800 ;
        RECT 53.820 148.785 53.960 148.940 ;
        RECT 54.650 148.940 55.415 149.080 ;
        RECT 54.650 148.880 54.970 148.940 ;
        RECT 55.125 148.895 55.415 148.940 ;
        RECT 56.030 149.080 56.350 149.140 ;
        RECT 61.550 149.080 61.870 149.140 ;
        RECT 62.485 149.080 62.775 149.125 ;
        RECT 56.030 148.940 62.775 149.080 ;
        RECT 56.030 148.880 56.350 148.940 ;
        RECT 61.550 148.880 61.870 148.940 ;
        RECT 62.485 148.895 62.775 148.940 ;
        RECT 64.310 148.880 64.630 149.140 ;
        RECT 65.230 148.880 65.550 149.140 ;
        RECT 66.165 149.080 66.455 149.125 ;
        RECT 66.610 149.080 66.930 149.140 ;
        RECT 66.165 148.940 66.930 149.080 ;
        RECT 66.165 148.895 66.455 148.940 ;
        RECT 66.610 148.880 66.930 148.940 ;
        RECT 71.180 149.080 71.470 149.125 ;
        RECT 71.670 149.080 71.990 149.140 ;
        RECT 71.180 148.940 71.990 149.080 ;
        RECT 73.830 149.080 73.970 149.280 ;
        RECT 74.430 149.280 77.035 149.420 ;
        RECT 74.430 149.220 74.750 149.280 ;
        RECT 76.745 149.235 77.035 149.280 ;
        RECT 92.830 149.220 93.150 149.480 ;
        RECT 95.590 149.420 95.910 149.480 ;
        RECT 99.285 149.420 99.575 149.465 ;
        RECT 95.590 149.280 99.575 149.420 ;
        RECT 95.590 149.220 95.910 149.280 ;
        RECT 99.285 149.235 99.575 149.280 ;
        RECT 104.330 149.420 104.650 149.480 ;
        RECT 104.805 149.420 105.095 149.465 ;
        RECT 104.330 149.280 105.095 149.420 ;
        RECT 104.330 149.220 104.650 149.280 ;
        RECT 104.805 149.235 105.095 149.280 ;
        RECT 114.910 149.420 115.230 149.480 ;
        RECT 123.190 149.420 123.510 149.480 ;
        RECT 129.630 149.420 129.950 149.480 ;
        RECT 114.910 149.280 123.510 149.420 ;
        RECT 114.910 149.220 115.230 149.280 ;
        RECT 123.190 149.220 123.510 149.280 ;
        RECT 126.960 149.280 129.950 149.420 ;
        RECT 80.425 149.080 80.715 149.125 ;
        RECT 73.830 148.940 80.715 149.080 ;
        RECT 71.180 148.895 71.470 148.940 ;
        RECT 71.670 148.880 71.990 148.940 ;
        RECT 80.425 148.895 80.715 148.940 ;
        RECT 101.585 149.080 101.875 149.125 ;
        RECT 108.010 149.080 108.330 149.140 ;
        RECT 126.960 149.125 127.100 149.280 ;
        RECT 129.630 149.220 129.950 149.280 ;
        RECT 131.945 149.420 132.235 149.465 ;
        RECT 136.530 149.420 136.850 149.480 ;
        RECT 131.945 149.280 136.850 149.420 ;
        RECT 131.945 149.235 132.235 149.280 ;
        RECT 136.530 149.220 136.850 149.280 ;
        RECT 114.005 149.080 114.295 149.125 ;
        RECT 101.585 148.940 111.000 149.080 ;
        RECT 101.585 148.895 101.875 148.940 ;
        RECT 108.010 148.880 108.330 148.940 ;
        RECT 51.905 148.555 52.195 148.785 ;
        RECT 52.350 148.740 52.680 148.785 ;
        RECT 52.350 148.600 52.865 148.740 ;
        RECT 52.350 148.555 52.680 148.600 ;
        RECT 53.745 148.555 54.035 148.785 ;
        RECT 47.765 148.400 48.055 148.445 ;
        RECT 50.970 148.400 51.290 148.460 ;
        RECT 47.765 148.260 51.290 148.400 ;
        RECT 47.765 148.215 48.055 148.260 ;
        RECT 50.970 148.200 51.290 148.260 ;
        RECT 51.980 148.400 52.120 148.555 ;
        RECT 52.350 148.540 52.670 148.555 ;
        RECT 54.190 148.540 54.510 148.800 ;
        RECT 56.490 148.540 56.810 148.800 ;
        RECT 56.950 148.740 57.270 148.800 ;
        RECT 56.950 148.600 57.465 148.740 ;
        RECT 56.950 148.540 57.270 148.600 ;
        RECT 57.885 148.555 58.175 148.785 ;
        RECT 52.810 148.400 53.130 148.460 ;
        RECT 57.960 148.400 58.100 148.555 ;
        RECT 58.330 148.540 58.650 148.800 ;
        RECT 59.035 148.740 59.325 148.785 ;
        RECT 60.630 148.740 60.950 148.800 ;
        RECT 59.035 148.600 60.950 148.740 ;
        RECT 59.035 148.555 59.325 148.600 ;
        RECT 60.630 148.540 60.950 148.600 ;
        RECT 61.090 148.540 61.410 148.800 ;
        RECT 62.025 148.555 62.315 148.785 ;
        RECT 62.100 148.400 62.240 148.555 ;
        RECT 62.930 148.540 63.250 148.800 ;
        RECT 69.845 148.740 70.135 148.785 ;
        RECT 70.290 148.740 70.610 148.800 ;
        RECT 69.845 148.600 70.610 148.740 ;
        RECT 69.845 148.555 70.135 148.600 ;
        RECT 70.290 148.540 70.610 148.600 ;
        RECT 96.985 148.740 97.275 148.785 ;
        RECT 98.350 148.740 98.670 148.800 ;
        RECT 96.985 148.600 98.670 148.740 ;
        RECT 96.985 148.555 97.275 148.600 ;
        RECT 98.350 148.540 98.670 148.600 ;
        RECT 101.110 148.540 101.430 148.800 ;
        RECT 102.950 148.740 103.270 148.800 ;
        RECT 104.345 148.740 104.635 148.785 ;
        RECT 102.950 148.600 104.635 148.740 ;
        RECT 102.950 148.540 103.270 148.600 ;
        RECT 104.345 148.555 104.635 148.600 ;
        RECT 106.170 148.740 106.490 148.800 ;
        RECT 110.860 148.785 111.000 148.940 ;
        RECT 114.005 148.940 116.980 149.080 ;
        RECT 114.005 148.895 114.295 148.940 ;
        RECT 106.645 148.740 106.935 148.785 ;
        RECT 106.170 148.600 106.935 148.740 ;
        RECT 106.170 148.540 106.490 148.600 ;
        RECT 106.645 148.555 106.935 148.600 ;
        RECT 110.785 148.555 111.075 148.785 ;
        RECT 114.465 148.740 114.755 148.785 ;
        RECT 115.370 148.740 115.690 148.800 ;
        RECT 114.465 148.600 115.690 148.740 ;
        RECT 114.465 148.555 114.755 148.600 ;
        RECT 115.370 148.540 115.690 148.600 ;
        RECT 64.770 148.400 65.090 148.460 ;
        RECT 51.980 148.260 53.130 148.400 ;
        RECT 51.980 148.060 52.120 148.260 ;
        RECT 52.810 148.200 53.130 148.260 ;
        RECT 54.740 148.260 58.100 148.400 ;
        RECT 59.800 148.260 62.240 148.400 ;
        RECT 62.560 148.260 65.090 148.400 ;
        RECT 47.380 147.920 52.120 148.060 ;
        RECT 53.285 148.060 53.575 148.105 ;
        RECT 54.740 148.060 54.880 148.260 ;
        RECT 53.285 147.920 54.880 148.060 ;
        RECT 34.910 147.875 35.200 147.920 ;
        RECT 37.010 147.875 37.300 147.920 ;
        RECT 38.580 147.875 38.870 147.920 ;
        RECT 53.285 147.875 53.575 147.920 ;
        RECT 55.110 147.860 55.430 148.120 ;
        RECT 59.800 148.105 59.940 148.260 ;
        RECT 59.725 147.875 60.015 148.105 ;
        RECT 60.630 148.060 60.950 148.120 ;
        RECT 62.560 148.060 62.700 148.260 ;
        RECT 64.770 148.200 65.090 148.260 ;
        RECT 70.725 148.400 71.015 148.445 ;
        RECT 71.915 148.400 72.205 148.445 ;
        RECT 74.435 148.400 74.725 148.445 ;
        RECT 70.725 148.260 74.725 148.400 ;
        RECT 70.725 148.215 71.015 148.260 ;
        RECT 71.915 148.215 72.205 148.260 ;
        RECT 74.435 148.215 74.725 148.260 ;
        RECT 87.310 148.400 87.630 148.460 ;
        RECT 89.625 148.400 89.915 148.445 ;
        RECT 87.310 148.260 89.915 148.400 ;
        RECT 87.310 148.200 87.630 148.260 ;
        RECT 89.625 148.215 89.915 148.260 ;
        RECT 97.430 148.200 97.750 148.460 ;
        RECT 97.890 148.400 98.210 148.460 ;
        RECT 102.045 148.400 102.335 148.445 ;
        RECT 97.890 148.260 102.335 148.400 ;
        RECT 97.890 148.200 98.210 148.260 ;
        RECT 102.045 148.215 102.335 148.260 ;
        RECT 107.105 148.215 107.395 148.445 ;
        RECT 108.025 148.400 108.315 148.445 ;
        RECT 108.470 148.400 108.790 148.460 ;
        RECT 108.025 148.260 108.790 148.400 ;
        RECT 108.025 148.215 108.315 148.260 ;
        RECT 60.630 147.920 62.700 148.060 ;
        RECT 63.865 148.060 64.155 148.105 ;
        RECT 67.530 148.060 67.850 148.120 ;
        RECT 63.865 147.920 67.850 148.060 ;
        RECT 60.630 147.860 60.950 147.920 ;
        RECT 63.865 147.875 64.155 147.920 ;
        RECT 67.530 147.860 67.850 147.920 ;
        RECT 70.330 148.060 70.620 148.105 ;
        RECT 72.430 148.060 72.720 148.105 ;
        RECT 74.000 148.060 74.290 148.105 ;
        RECT 70.330 147.920 74.290 148.060 ;
        RECT 70.330 147.875 70.620 147.920 ;
        RECT 72.430 147.875 72.720 147.920 ;
        RECT 74.000 147.875 74.290 147.920 ;
        RECT 95.145 148.060 95.435 148.105 ;
        RECT 96.510 148.060 96.830 148.120 ;
        RECT 95.145 147.920 96.830 148.060 ;
        RECT 107.180 148.060 107.320 148.215 ;
        RECT 108.470 148.200 108.790 148.260 ;
        RECT 114.910 148.200 115.230 148.460 ;
        RECT 115.845 148.215 116.135 148.445 ;
        RECT 116.305 148.400 116.595 148.445 ;
        RECT 116.840 148.400 116.980 148.940 ;
        RECT 117.300 148.940 121.120 149.080 ;
        RECT 117.300 148.800 117.440 148.940 ;
        RECT 117.210 148.540 117.530 148.800 ;
        RECT 117.685 148.740 117.975 148.785 ;
        RECT 118.130 148.740 118.450 148.800 ;
        RECT 117.685 148.600 118.450 148.740 ;
        RECT 117.685 148.555 117.975 148.600 ;
        RECT 118.130 148.540 118.450 148.600 ;
        RECT 118.590 148.740 118.910 148.800 ;
        RECT 120.430 148.740 120.750 148.800 ;
        RECT 118.590 148.600 120.750 148.740 ;
        RECT 120.980 148.740 121.120 148.940 ;
        RECT 126.885 148.895 127.175 149.125 ;
        RECT 130.565 149.080 130.855 149.125 ;
        RECT 131.470 149.080 131.790 149.140 ;
        RECT 130.565 148.940 131.790 149.080 ;
        RECT 130.565 148.895 130.855 148.940 ;
        RECT 131.470 148.880 131.790 148.940 ;
        RECT 135.580 149.080 135.870 149.125 ;
        RECT 141.130 149.080 141.450 149.140 ;
        RECT 135.580 148.940 141.450 149.080 ;
        RECT 135.580 148.895 135.870 148.940 ;
        RECT 141.130 148.880 141.450 148.940 ;
        RECT 120.980 148.730 122.040 148.740 ;
        RECT 122.745 148.730 123.035 148.785 ;
        RECT 120.980 148.600 123.035 148.730 ;
        RECT 118.590 148.540 118.910 148.600 ;
        RECT 120.430 148.540 120.750 148.600 ;
        RECT 121.900 148.590 123.035 148.600 ;
        RECT 122.745 148.555 123.035 148.590 ;
        RECT 123.205 148.730 123.495 148.785 ;
        RECT 124.110 148.740 124.430 148.800 ;
        RECT 124.585 148.740 124.875 148.785 ;
        RECT 123.740 148.730 124.875 148.740 ;
        RECT 123.205 148.600 124.875 148.730 ;
        RECT 123.205 148.590 123.880 148.600 ;
        RECT 123.205 148.555 123.495 148.590 ;
        RECT 124.110 148.540 124.430 148.600 ;
        RECT 124.585 148.555 124.875 148.600 ;
        RECT 125.490 148.540 125.810 148.800 ;
        RECT 127.805 148.740 128.095 148.785 ;
        RECT 128.250 148.740 128.570 148.800 ;
        RECT 127.805 148.600 128.570 148.740 ;
        RECT 127.805 148.555 128.095 148.600 ;
        RECT 128.250 148.540 128.570 148.600 ;
        RECT 129.185 148.740 129.475 148.785 ;
        RECT 129.630 148.740 129.950 148.800 ;
        RECT 129.185 148.600 129.950 148.740 ;
        RECT 129.185 148.555 129.475 148.600 ;
        RECT 129.630 148.540 129.950 148.600 ;
        RECT 130.090 148.540 130.410 148.800 ;
        RECT 131.025 148.740 131.315 148.785 ;
        RECT 133.310 148.740 133.630 148.800 ;
        RECT 131.025 148.600 133.630 148.740 ;
        RECT 131.025 148.555 131.315 148.600 ;
        RECT 133.310 148.540 133.630 148.600 ;
        RECT 133.770 148.740 134.090 148.800 ;
        RECT 134.245 148.740 134.535 148.785 ;
        RECT 143.445 148.740 143.735 148.785 ;
        RECT 133.770 148.600 134.535 148.740 ;
        RECT 133.770 148.540 134.090 148.600 ;
        RECT 134.245 148.555 134.535 148.600 ;
        RECT 134.735 148.600 143.735 148.740 ;
        RECT 116.305 148.260 116.980 148.400 ;
        RECT 116.305 148.215 116.595 148.260 ;
        RECT 115.920 148.060 116.060 148.215 ;
        RECT 119.510 148.200 119.830 148.460 ;
        RECT 121.825 148.215 122.115 148.445 ;
        RECT 122.285 148.400 122.575 148.445 ;
        RECT 125.950 148.400 126.270 148.460 ;
        RECT 122.285 148.260 126.270 148.400 ;
        RECT 122.285 148.215 122.575 148.260 ;
        RECT 116.765 148.060 117.055 148.105 ;
        RECT 107.180 147.920 115.140 148.060 ;
        RECT 115.920 147.920 117.055 148.060 ;
        RECT 95.145 147.875 95.435 147.920 ;
        RECT 96.510 147.860 96.830 147.920 ;
        RECT 115.000 147.780 115.140 147.920 ;
        RECT 116.765 147.875 117.055 147.920 ;
        RECT 117.210 148.060 117.530 148.120 ;
        RECT 119.065 148.060 119.355 148.105 ;
        RECT 117.210 147.920 119.355 148.060 ;
        RECT 121.900 148.060 122.040 148.215 ;
        RECT 125.950 148.200 126.270 148.260 ;
        RECT 127.330 148.400 127.650 148.460 ;
        RECT 134.735 148.400 134.875 148.600 ;
        RECT 143.445 148.555 143.735 148.600 ;
        RECT 127.330 148.260 134.875 148.400 ;
        RECT 135.125 148.400 135.415 148.445 ;
        RECT 136.315 148.400 136.605 148.445 ;
        RECT 138.835 148.400 139.125 148.445 ;
        RECT 135.125 148.260 139.125 148.400 ;
        RECT 127.330 148.200 127.650 148.260 ;
        RECT 135.125 148.215 135.415 148.260 ;
        RECT 136.315 148.215 136.605 148.260 ;
        RECT 138.835 148.215 139.125 148.260 ;
        RECT 143.890 148.200 144.210 148.460 ;
        RECT 144.810 148.200 145.130 148.460 ;
        RECT 122.730 148.060 123.050 148.120 ;
        RECT 125.045 148.060 125.335 148.105 ;
        RECT 121.900 147.920 122.500 148.060 ;
        RECT 117.210 147.860 117.530 147.920 ;
        RECT 119.065 147.875 119.355 147.920 ;
        RECT 122.360 147.780 122.500 147.920 ;
        RECT 122.730 147.920 125.335 148.060 ;
        RECT 122.730 147.860 123.050 147.920 ;
        RECT 125.045 147.875 125.335 147.920 ;
        RECT 134.730 148.060 135.020 148.105 ;
        RECT 136.830 148.060 137.120 148.105 ;
        RECT 138.400 148.060 138.690 148.105 ;
        RECT 134.730 147.920 138.690 148.060 ;
        RECT 134.730 147.875 135.020 147.920 ;
        RECT 136.830 147.875 137.120 147.920 ;
        RECT 138.400 147.875 138.690 147.920 ;
        RECT 33.045 147.535 33.335 147.765 ;
        RECT 33.965 147.720 34.255 147.765 ;
        RECT 36.250 147.720 36.570 147.780 ;
        RECT 33.965 147.580 36.570 147.720 ;
        RECT 33.965 147.535 34.255 147.580 ;
        RECT 36.250 147.520 36.570 147.580 ;
        RECT 39.930 147.720 40.250 147.780 ;
        RECT 41.325 147.720 41.615 147.765 ;
        RECT 39.930 147.580 41.615 147.720 ;
        RECT 39.930 147.520 40.250 147.580 ;
        RECT 41.325 147.535 41.615 147.580 ;
        RECT 50.050 147.720 50.370 147.780 ;
        RECT 54.650 147.720 54.970 147.780 ;
        RECT 50.050 147.580 54.970 147.720 ;
        RECT 50.050 147.520 50.370 147.580 ;
        RECT 54.650 147.520 54.970 147.580 ;
        RECT 58.790 147.720 59.110 147.780 ;
        RECT 69.370 147.720 69.690 147.780 ;
        RECT 58.790 147.580 69.690 147.720 ;
        RECT 58.790 147.520 59.110 147.580 ;
        RECT 69.370 147.520 69.690 147.580 ;
        RECT 86.850 147.520 87.170 147.780 ;
        RECT 103.870 147.520 104.190 147.780 ;
        RECT 114.910 147.520 115.230 147.780 ;
        RECT 115.370 147.520 115.690 147.780 ;
        RECT 115.830 147.720 116.150 147.780 ;
        RECT 118.130 147.720 118.450 147.780 ;
        RECT 115.830 147.580 118.450 147.720 ;
        RECT 115.830 147.520 116.150 147.580 ;
        RECT 118.130 147.520 118.450 147.580 ;
        RECT 122.270 147.520 122.590 147.780 ;
        RECT 124.110 147.520 124.430 147.780 ;
        RECT 128.725 147.720 129.015 147.765 ;
        RECT 130.090 147.720 130.410 147.780 ;
        RECT 128.725 147.580 130.410 147.720 ;
        RECT 128.725 147.535 129.015 147.580 ;
        RECT 130.090 147.520 130.410 147.580 ;
        RECT 137.450 147.720 137.770 147.780 ;
        RECT 141.145 147.720 141.435 147.765 ;
        RECT 137.450 147.580 141.435 147.720 ;
        RECT 137.450 147.520 137.770 147.580 ;
        RECT 141.145 147.535 141.435 147.580 ;
        RECT 141.590 147.520 141.910 147.780 ;
        RECT 17.320 146.900 147.040 147.380 ;
        RECT 31.205 146.700 31.495 146.745 ;
        RECT 32.110 146.700 32.430 146.760 ;
        RECT 31.205 146.560 32.430 146.700 ;
        RECT 31.205 146.515 31.495 146.560 ;
        RECT 32.110 146.500 32.430 146.560 ;
        RECT 45.005 146.700 45.295 146.745 ;
        RECT 51.430 146.700 51.750 146.760 ;
        RECT 45.005 146.560 51.750 146.700 ;
        RECT 45.005 146.515 45.295 146.560 ;
        RECT 51.430 146.500 51.750 146.560 ;
        RECT 61.565 146.700 61.855 146.745 ;
        RECT 62.945 146.700 63.235 146.745 ;
        RECT 61.565 146.560 63.235 146.700 ;
        RECT 61.565 146.515 61.855 146.560 ;
        RECT 62.945 146.515 63.235 146.560 ;
        RECT 87.310 146.500 87.630 146.760 ;
        RECT 106.170 146.500 106.490 146.760 ;
        RECT 108.010 146.500 108.330 146.760 ;
        RECT 111.690 146.700 112.010 146.760 ;
        RECT 115.385 146.700 115.675 146.745 ;
        RECT 111.690 146.560 115.675 146.700 ;
        RECT 111.690 146.500 112.010 146.560 ;
        RECT 115.385 146.515 115.675 146.560 ;
        RECT 119.510 146.700 119.830 146.760 ;
        RECT 123.665 146.700 123.955 146.745 ;
        RECT 142.970 146.700 143.290 146.760 ;
        RECT 145.285 146.700 145.575 146.745 ;
        RECT 119.510 146.560 123.955 146.700 ;
        RECT 119.510 146.500 119.830 146.560 ;
        RECT 123.665 146.515 123.955 146.560 ;
        RECT 132.480 146.560 139.060 146.700 ;
        RECT 33.950 146.360 34.240 146.405 ;
        RECT 35.520 146.360 35.810 146.405 ;
        RECT 37.620 146.360 37.910 146.405 ;
        RECT 33.950 146.220 37.910 146.360 ;
        RECT 33.950 146.175 34.240 146.220 ;
        RECT 35.520 146.175 35.810 146.220 ;
        RECT 37.620 146.175 37.910 146.220 ;
        RECT 38.090 146.160 38.410 146.420 ;
        RECT 47.750 146.160 48.070 146.420 ;
        RECT 58.330 146.360 58.650 146.420 ;
        RECT 57.960 146.220 58.650 146.360 ;
        RECT 33.515 146.020 33.805 146.065 ;
        RECT 36.035 146.020 36.325 146.065 ;
        RECT 37.225 146.020 37.515 146.065 ;
        RECT 33.515 145.880 37.515 146.020 ;
        RECT 38.180 146.020 38.320 146.160 ;
        RECT 38.180 145.880 44.300 146.020 ;
        RECT 33.515 145.835 33.805 145.880 ;
        RECT 36.035 145.835 36.325 145.880 ;
        RECT 37.225 145.835 37.515 145.880 ;
        RECT 34.870 145.680 35.190 145.740 ;
        RECT 38.105 145.680 38.395 145.725 ;
        RECT 34.870 145.540 38.395 145.680 ;
        RECT 34.870 145.480 35.190 145.540 ;
        RECT 38.105 145.495 38.395 145.540 ;
        RECT 38.550 145.480 38.870 145.740 ;
        RECT 39.010 145.680 39.330 145.740 ;
        RECT 39.485 145.680 39.775 145.725 ;
        RECT 39.010 145.540 39.775 145.680 ;
        RECT 39.010 145.480 39.330 145.540 ;
        RECT 39.485 145.495 39.775 145.540 ;
        RECT 39.930 145.480 40.250 145.740 ;
        RECT 40.405 145.495 40.695 145.725 ;
        RECT 40.850 145.680 41.170 145.740 ;
        RECT 40.850 145.540 42.000 145.680 ;
        RECT 36.250 145.340 36.570 145.400 ;
        RECT 36.770 145.340 37.060 145.385 ;
        RECT 36.250 145.200 37.060 145.340 ;
        RECT 38.640 145.340 38.780 145.480 ;
        RECT 40.480 145.340 40.620 145.495 ;
        RECT 40.850 145.480 41.170 145.540 ;
        RECT 38.640 145.200 40.620 145.340 ;
        RECT 41.860 145.340 42.000 145.540 ;
        RECT 42.230 145.480 42.550 145.740 ;
        RECT 42.690 145.480 43.010 145.740 ;
        RECT 44.160 145.725 44.300 145.880 ;
        RECT 43.625 145.495 43.915 145.725 ;
        RECT 44.085 145.495 44.375 145.725 ;
        RECT 45.465 145.495 45.755 145.725 ;
        RECT 43.700 145.340 43.840 145.495 ;
        RECT 45.540 145.340 45.680 145.495 ;
        RECT 46.830 145.480 47.150 145.740 ;
        RECT 57.960 145.725 58.100 146.220 ;
        RECT 58.330 146.160 58.650 146.220 ;
        RECT 59.265 146.360 59.555 146.405 ;
        RECT 59.725 146.360 60.015 146.405 ;
        RECT 66.610 146.360 66.930 146.420 ;
        RECT 59.265 146.220 66.930 146.360 ;
        RECT 59.265 146.175 59.555 146.220 ;
        RECT 59.725 146.175 60.015 146.220 ;
        RECT 66.610 146.160 66.930 146.220 ;
        RECT 90.070 146.360 90.360 146.405 ;
        RECT 91.640 146.360 91.930 146.405 ;
        RECT 93.740 146.360 94.030 146.405 ;
        RECT 90.070 146.220 94.030 146.360 ;
        RECT 90.070 146.175 90.360 146.220 ;
        RECT 91.640 146.175 91.930 146.220 ;
        RECT 93.740 146.175 94.030 146.220 ;
        RECT 95.170 146.360 95.460 146.405 ;
        RECT 97.270 146.360 97.560 146.405 ;
        RECT 98.840 146.360 99.130 146.405 ;
        RECT 95.170 146.220 99.130 146.360 ;
        RECT 95.170 146.175 95.460 146.220 ;
        RECT 97.270 146.175 97.560 146.220 ;
        RECT 98.840 146.175 99.130 146.220 ;
        RECT 110.770 146.360 111.060 146.405 ;
        RECT 112.340 146.360 112.630 146.405 ;
        RECT 114.440 146.360 114.730 146.405 ;
        RECT 110.770 146.220 114.730 146.360 ;
        RECT 110.770 146.175 111.060 146.220 ;
        RECT 112.340 146.175 112.630 146.220 ;
        RECT 114.440 146.175 114.730 146.220 ;
        RECT 114.910 146.360 115.230 146.420 ;
        RECT 120.890 146.360 121.210 146.420 ;
        RECT 114.910 146.220 121.210 146.360 ;
        RECT 114.910 146.160 115.230 146.220 ;
        RECT 120.890 146.160 121.210 146.220 ;
        RECT 124.110 146.360 124.430 146.420 ;
        RECT 124.110 146.220 128.020 146.360 ;
        RECT 124.110 146.160 124.430 146.220 ;
        RECT 60.630 146.020 60.950 146.080 ;
        RECT 89.635 146.020 89.925 146.065 ;
        RECT 92.155 146.020 92.445 146.065 ;
        RECT 93.345 146.020 93.635 146.065 ;
        RECT 58.420 145.880 65.000 146.020 ;
        RECT 58.420 145.725 58.560 145.880 ;
        RECT 60.630 145.820 60.950 145.880 ;
        RECT 57.885 145.495 58.175 145.725 ;
        RECT 58.345 145.495 58.635 145.725 ;
        RECT 41.860 145.200 45.680 145.340 ;
        RECT 57.960 145.340 58.100 145.495 ;
        RECT 64.860 145.400 65.000 145.880 ;
        RECT 89.635 145.880 93.635 146.020 ;
        RECT 89.635 145.835 89.925 145.880 ;
        RECT 92.155 145.835 92.445 145.880 ;
        RECT 93.345 145.835 93.635 145.880 ;
        RECT 94.210 146.020 94.530 146.080 ;
        RECT 94.685 146.020 94.975 146.065 ;
        RECT 94.210 145.880 94.975 146.020 ;
        RECT 94.210 145.820 94.530 145.880 ;
        RECT 94.685 145.835 94.975 145.880 ;
        RECT 95.565 146.020 95.855 146.065 ;
        RECT 96.755 146.020 97.045 146.065 ;
        RECT 99.275 146.020 99.565 146.065 ;
        RECT 95.565 145.880 99.565 146.020 ;
        RECT 95.565 145.835 95.855 145.880 ;
        RECT 96.755 145.835 97.045 145.880 ;
        RECT 99.275 145.835 99.565 145.880 ;
        RECT 110.335 146.020 110.625 146.065 ;
        RECT 112.855 146.020 113.145 146.065 ;
        RECT 114.045 146.020 114.335 146.065 ;
        RECT 110.335 145.880 114.335 146.020 ;
        RECT 110.335 145.835 110.625 145.880 ;
        RECT 112.855 145.835 113.145 145.880 ;
        RECT 114.045 145.835 114.335 145.880 ;
        RECT 116.750 146.020 117.070 146.080 ;
        RECT 118.145 146.020 118.435 146.065 ;
        RECT 116.750 145.880 118.435 146.020 ;
        RECT 116.750 145.820 117.070 145.880 ;
        RECT 118.145 145.835 118.435 145.880 ;
        RECT 122.745 146.020 123.035 146.065 ;
        RECT 123.205 146.020 123.495 146.065 ;
        RECT 126.410 146.020 126.730 146.080 ;
        RECT 127.880 146.065 128.020 146.220 ;
        RECT 122.745 145.880 123.495 146.020 ;
        RECT 122.745 145.835 123.035 145.880 ;
        RECT 123.205 145.835 123.495 145.880 ;
        RECT 124.200 145.880 126.730 146.020 ;
        RECT 73.970 145.680 74.290 145.740 ;
        RECT 78.585 145.680 78.875 145.725 ;
        RECT 79.030 145.680 79.350 145.740 ;
        RECT 73.970 145.540 79.350 145.680 ;
        RECT 73.970 145.480 74.290 145.540 ;
        RECT 78.585 145.495 78.875 145.540 ;
        RECT 79.030 145.480 79.350 145.540 ;
        RECT 79.950 145.480 80.270 145.740 ;
        RECT 97.430 145.680 97.750 145.740 ;
        RECT 102.965 145.680 103.255 145.725 ;
        RECT 97.430 145.540 103.255 145.680 ;
        RECT 97.430 145.480 97.750 145.540 ;
        RECT 102.965 145.495 103.255 145.540 ;
        RECT 112.150 145.680 112.470 145.740 ;
        RECT 114.925 145.680 115.215 145.725 ;
        RECT 112.150 145.540 115.215 145.680 ;
        RECT 112.150 145.480 112.470 145.540 ;
        RECT 114.925 145.495 115.215 145.540 ;
        RECT 115.370 145.480 115.690 145.740 ;
        RECT 117.685 145.680 117.975 145.725 ;
        RECT 119.050 145.680 119.370 145.740 ;
        RECT 124.200 145.725 124.340 145.880 ;
        RECT 126.410 145.820 126.730 145.880 ;
        RECT 127.805 145.835 128.095 146.065 ;
        RECT 131.010 146.020 131.330 146.080 ;
        RECT 132.480 146.065 132.620 146.560 ;
        RECT 134.730 146.360 135.020 146.405 ;
        RECT 136.830 146.360 137.120 146.405 ;
        RECT 138.400 146.360 138.690 146.405 ;
        RECT 134.730 146.220 138.690 146.360 ;
        RECT 138.920 146.360 139.060 146.560 ;
        RECT 142.970 146.560 145.575 146.700 ;
        RECT 142.970 146.500 143.290 146.560 ;
        RECT 145.285 146.515 145.575 146.560 ;
        RECT 143.430 146.360 143.750 146.420 ;
        RECT 138.920 146.220 143.750 146.360 ;
        RECT 134.730 146.175 135.020 146.220 ;
        RECT 136.830 146.175 137.120 146.220 ;
        RECT 138.400 146.175 138.690 146.220 ;
        RECT 143.430 146.160 143.750 146.220 ;
        RECT 132.405 146.020 132.695 146.065 ;
        RECT 131.010 145.880 132.695 146.020 ;
        RECT 131.010 145.820 131.330 145.880 ;
        RECT 132.405 145.835 132.695 145.880 ;
        RECT 133.770 146.020 134.090 146.080 ;
        RECT 134.245 146.020 134.535 146.065 ;
        RECT 133.770 145.880 134.535 146.020 ;
        RECT 133.770 145.820 134.090 145.880 ;
        RECT 134.245 145.835 134.535 145.880 ;
        RECT 135.125 146.020 135.415 146.065 ;
        RECT 136.315 146.020 136.605 146.065 ;
        RECT 138.835 146.020 139.125 146.065 ;
        RECT 135.125 145.880 139.125 146.020 ;
        RECT 135.125 145.835 135.415 145.880 ;
        RECT 136.315 145.835 136.605 145.880 ;
        RECT 138.835 145.835 139.125 145.880 ;
        RECT 119.525 145.680 119.815 145.725 ;
        RECT 117.685 145.540 119.815 145.680 ;
        RECT 117.685 145.495 117.975 145.540 ;
        RECT 119.050 145.480 119.370 145.540 ;
        RECT 119.525 145.495 119.815 145.540 ;
        RECT 124.125 145.495 124.415 145.725 ;
        RECT 124.585 145.495 124.875 145.725 ;
        RECT 135.580 145.680 135.870 145.725 ;
        RECT 141.590 145.680 141.910 145.740 ;
        RECT 135.580 145.540 141.910 145.680 ;
        RECT 135.580 145.495 135.870 145.540 ;
        RECT 63.865 145.340 64.155 145.385 ;
        RECT 57.960 145.200 64.155 145.340 ;
        RECT 36.250 145.140 36.570 145.200 ;
        RECT 36.770 145.155 37.060 145.200 ;
        RECT 63.865 145.155 64.155 145.200 ;
        RECT 35.790 145.000 36.110 145.060 ;
        RECT 38.565 145.000 38.855 145.045 ;
        RECT 35.790 144.860 38.855 145.000 ;
        RECT 35.790 144.800 36.110 144.860 ;
        RECT 38.565 144.815 38.855 144.860 ;
        RECT 42.230 145.000 42.550 145.060 ;
        RECT 45.910 145.000 46.230 145.060 ;
        RECT 42.230 144.860 46.230 145.000 ;
        RECT 42.230 144.800 42.550 144.860 ;
        RECT 45.910 144.800 46.230 144.860 ;
        RECT 57.410 145.000 57.730 145.060 ;
        RECT 61.565 145.000 61.855 145.045 ;
        RECT 57.410 144.860 61.855 145.000 ;
        RECT 57.410 144.800 57.730 144.860 ;
        RECT 61.565 144.815 61.855 144.860 ;
        RECT 62.470 144.800 62.790 145.060 ;
        RECT 63.940 145.000 64.080 145.155 ;
        RECT 64.770 145.140 65.090 145.400 ;
        RECT 77.665 145.340 77.955 145.385 ;
        RECT 80.040 145.340 80.180 145.480 ;
        RECT 77.665 145.200 80.180 145.340 ;
        RECT 93.000 145.340 93.290 145.385 ;
        RECT 93.750 145.340 94.070 145.400 ;
        RECT 93.000 145.200 94.070 145.340 ;
        RECT 77.665 145.155 77.955 145.200 ;
        RECT 93.000 145.155 93.290 145.200 ;
        RECT 93.750 145.140 94.070 145.200 ;
        RECT 94.670 145.340 94.990 145.400 ;
        RECT 95.910 145.340 96.200 145.385 ;
        RECT 113.700 145.340 113.990 145.385 ;
        RECT 115.460 145.340 115.600 145.480 ;
        RECT 94.670 145.200 96.200 145.340 ;
        RECT 94.670 145.140 94.990 145.200 ;
        RECT 95.910 145.155 96.200 145.200 ;
        RECT 96.600 145.200 102.260 145.340 ;
        RECT 68.450 145.000 68.770 145.060 ;
        RECT 63.940 144.860 68.770 145.000 ;
        RECT 68.450 144.800 68.770 144.860 ;
        RECT 74.890 145.000 75.210 145.060 ;
        RECT 76.270 145.000 76.590 145.060 ;
        RECT 76.745 145.000 77.035 145.045 ;
        RECT 74.890 144.860 77.035 145.000 ;
        RECT 74.890 144.800 75.210 144.860 ;
        RECT 76.270 144.800 76.590 144.860 ;
        RECT 76.745 144.815 77.035 144.860 ;
        RECT 79.490 144.800 79.810 145.060 ;
        RECT 83.630 145.000 83.950 145.060 ;
        RECT 96.600 145.000 96.740 145.200 ;
        RECT 83.630 144.860 96.740 145.000 ;
        RECT 98.350 145.000 98.670 145.060 ;
        RECT 101.585 145.000 101.875 145.045 ;
        RECT 98.350 144.860 101.875 145.000 ;
        RECT 102.120 145.000 102.260 145.200 ;
        RECT 113.700 145.200 115.600 145.340 ;
        RECT 118.130 145.340 118.450 145.400 ;
        RECT 124.660 145.340 124.800 145.495 ;
        RECT 141.590 145.480 141.910 145.540 ;
        RECT 142.065 145.495 142.355 145.725 ;
        RECT 118.130 145.200 124.800 145.340 ;
        RECT 137.450 145.340 137.770 145.400 ;
        RECT 142.140 145.340 142.280 145.495 ;
        RECT 137.450 145.200 142.280 145.340 ;
        RECT 113.700 145.155 113.990 145.200 ;
        RECT 118.130 145.140 118.450 145.200 ;
        RECT 137.450 145.140 137.770 145.200 ;
        RECT 115.830 145.000 116.150 145.060 ;
        RECT 102.120 144.860 116.150 145.000 ;
        RECT 83.630 144.800 83.950 144.860 ;
        RECT 98.350 144.800 98.670 144.860 ;
        RECT 101.585 144.815 101.875 144.860 ;
        RECT 115.830 144.800 116.150 144.860 ;
        RECT 117.225 145.000 117.515 145.045 ;
        RECT 120.890 145.000 121.210 145.060 ;
        RECT 117.225 144.860 121.210 145.000 ;
        RECT 117.225 144.815 117.515 144.860 ;
        RECT 120.890 144.800 121.210 144.860 ;
        RECT 125.045 145.000 125.335 145.045 ;
        RECT 125.490 145.000 125.810 145.060 ;
        RECT 125.045 144.860 125.810 145.000 ;
        RECT 125.045 144.815 125.335 144.860 ;
        RECT 125.490 144.800 125.810 144.860 ;
        RECT 126.870 144.800 127.190 145.060 ;
        RECT 127.345 145.000 127.635 145.045 ;
        RECT 129.185 145.000 129.475 145.045 ;
        RECT 127.345 144.860 129.475 145.000 ;
        RECT 127.345 144.815 127.635 144.860 ;
        RECT 129.185 144.815 129.475 144.860 ;
        RECT 141.145 145.000 141.435 145.045 ;
        RECT 142.050 145.000 142.370 145.060 ;
        RECT 141.145 144.860 142.370 145.000 ;
        RECT 141.145 144.815 141.435 144.860 ;
        RECT 142.050 144.800 142.370 144.860 ;
        RECT 17.320 144.180 147.040 144.660 ;
        RECT 38.090 143.780 38.410 144.040 ;
        RECT 39.010 143.980 39.330 144.040 ;
        RECT 39.485 143.980 39.775 144.025 ;
        RECT 39.010 143.840 39.775 143.980 ;
        RECT 39.010 143.780 39.330 143.840 ;
        RECT 39.485 143.795 39.775 143.840 ;
        RECT 40.405 143.980 40.695 144.025 ;
        RECT 40.850 143.980 41.170 144.040 ;
        RECT 40.405 143.840 41.170 143.980 ;
        RECT 40.405 143.795 40.695 143.840 ;
        RECT 40.850 143.780 41.170 143.840 ;
        RECT 59.265 143.980 59.555 144.025 ;
        RECT 61.090 143.980 61.410 144.040 ;
        RECT 59.265 143.840 61.410 143.980 ;
        RECT 59.265 143.795 59.555 143.840 ;
        RECT 61.090 143.780 61.410 143.840 ;
        RECT 67.085 143.980 67.375 144.025 ;
        RECT 68.450 143.980 68.770 144.040 ;
        RECT 78.570 143.980 78.890 144.040 ;
        RECT 80.410 143.980 80.730 144.040 ;
        RECT 67.085 143.840 68.770 143.980 ;
        RECT 67.085 143.795 67.375 143.840 ;
        RECT 68.450 143.780 68.770 143.840 ;
        RECT 72.220 143.840 80.730 143.980 ;
        RECT 36.265 143.640 36.555 143.685 ;
        RECT 39.930 143.640 40.250 143.700 ;
        RECT 32.200 143.500 36.555 143.640 ;
        RECT 29.350 142.960 29.670 143.020 ;
        RECT 32.200 143.005 32.340 143.500 ;
        RECT 36.265 143.455 36.555 143.500 ;
        RECT 37.260 143.500 40.250 143.640 ;
        RECT 37.260 143.345 37.400 143.500 ;
        RECT 39.930 143.440 40.250 143.500 ;
        RECT 54.190 143.640 54.510 143.700 ;
        RECT 58.345 143.640 58.635 143.685 ;
        RECT 58.790 143.640 59.110 143.700 ;
        RECT 60.630 143.640 60.950 143.700 ;
        RECT 54.190 143.500 59.110 143.640 ;
        RECT 54.190 143.440 54.510 143.500 ;
        RECT 58.345 143.455 58.635 143.500 ;
        RECT 58.790 143.440 59.110 143.500 ;
        RECT 59.800 143.500 60.950 143.640 ;
        RECT 35.805 143.115 36.095 143.345 ;
        RECT 37.185 143.115 37.475 143.345 ;
        RECT 38.550 143.300 38.870 143.360 ;
        RECT 41.325 143.300 41.615 143.345 ;
        RECT 38.550 143.160 41.615 143.300 ;
        RECT 32.125 142.960 32.415 143.005 ;
        RECT 35.330 142.960 35.650 143.020 ;
        RECT 29.350 142.820 32.415 142.960 ;
        RECT 29.350 142.760 29.670 142.820 ;
        RECT 32.125 142.775 32.415 142.820 ;
        RECT 34.040 142.820 35.650 142.960 ;
        RECT 35.880 142.960 36.020 143.115 ;
        RECT 38.550 143.100 38.870 143.160 ;
        RECT 41.325 143.115 41.615 143.160 ;
        RECT 53.730 143.300 54.050 143.360 ;
        RECT 54.650 143.300 54.970 143.360 ;
        RECT 53.730 143.160 54.970 143.300 ;
        RECT 53.730 143.100 54.050 143.160 ;
        RECT 54.650 143.100 54.970 143.160 ;
        RECT 55.570 143.100 55.890 143.360 ;
        RECT 56.505 143.300 56.795 143.345 ;
        RECT 59.800 143.300 59.940 143.500 ;
        RECT 60.630 143.440 60.950 143.500 ;
        RECT 61.520 143.640 61.810 143.685 ;
        RECT 62.470 143.640 62.790 143.700 ;
        RECT 61.520 143.500 62.790 143.640 ;
        RECT 61.520 143.455 61.810 143.500 ;
        RECT 62.470 143.440 62.790 143.500 ;
        RECT 56.505 143.160 59.940 143.300 ;
        RECT 56.505 143.115 56.795 143.160 ;
        RECT 60.170 143.100 60.490 143.360 ;
        RECT 72.220 143.345 72.360 143.840 ;
        RECT 78.570 143.780 78.890 143.840 ;
        RECT 80.410 143.780 80.730 143.840 ;
        RECT 93.750 143.980 94.070 144.040 ;
        RECT 93.750 143.840 104.100 143.980 ;
        RECT 93.750 143.780 94.070 143.840 ;
        RECT 103.960 143.700 104.100 143.840 ;
        RECT 119.050 143.780 119.370 144.040 ;
        RECT 123.665 143.980 123.955 144.025 ;
        RECT 127.330 143.980 127.650 144.040 ;
        RECT 123.665 143.840 127.650 143.980 ;
        RECT 123.665 143.795 123.955 143.840 ;
        RECT 127.330 143.780 127.650 143.840 ;
        RECT 131.010 143.780 131.330 144.040 ;
        RECT 138.830 143.780 139.150 144.040 ;
        RECT 141.145 143.980 141.435 144.025 ;
        RECT 142.970 143.980 143.290 144.040 ;
        RECT 141.145 143.840 143.290 143.980 ;
        RECT 141.145 143.795 141.435 143.840 ;
        RECT 142.970 143.780 143.290 143.840 ;
        RECT 143.890 143.980 144.210 144.040 ;
        RECT 145.285 143.980 145.575 144.025 ;
        RECT 143.890 143.840 145.575 143.980 ;
        RECT 143.890 143.780 144.210 143.840 ;
        RECT 145.285 143.795 145.575 143.840 ;
        RECT 86.390 143.640 86.710 143.700 ;
        RECT 90.530 143.640 90.850 143.700 ;
        RECT 94.210 143.640 94.530 143.700 ;
        RECT 74.520 143.500 86.710 143.640 ;
        RECT 72.145 143.115 72.435 143.345 ;
        RECT 73.065 143.300 73.355 143.345 ;
        RECT 73.970 143.300 74.290 143.360 ;
        RECT 74.520 143.345 74.660 143.500 ;
        RECT 86.390 143.440 86.710 143.500 ;
        RECT 88.780 143.500 94.530 143.640 ;
        RECT 73.065 143.160 74.290 143.300 ;
        RECT 73.065 143.115 73.355 143.160 ;
        RECT 73.970 143.100 74.290 143.160 ;
        RECT 74.445 143.115 74.735 143.345 ;
        RECT 85.930 143.300 86.250 143.360 ;
        RECT 88.780 143.345 88.920 143.500 ;
        RECT 90.530 143.440 90.850 143.500 ;
        RECT 94.210 143.440 94.530 143.500 ;
        RECT 103.870 143.640 104.190 143.700 ;
        RECT 112.150 143.640 112.470 143.700 ;
        RECT 133.770 143.640 134.090 143.700 ;
        RECT 103.870 143.500 105.940 143.640 ;
        RECT 103.870 143.440 104.190 143.500 ;
        RECT 87.370 143.300 87.660 143.345 ;
        RECT 85.930 143.160 87.660 143.300 ;
        RECT 85.930 143.100 86.250 143.160 ;
        RECT 87.370 143.115 87.660 143.160 ;
        RECT 88.705 143.115 88.995 143.345 ;
        RECT 92.845 143.300 93.135 143.345 ;
        RECT 96.970 143.300 97.290 143.360 ;
        RECT 92.845 143.160 97.290 143.300 ;
        RECT 92.845 143.115 93.135 143.160 ;
        RECT 96.970 143.100 97.290 143.160 ;
        RECT 98.350 143.100 98.670 143.360 ;
        RECT 100.665 143.300 100.955 143.345 ;
        RECT 101.110 143.300 101.430 143.360 ;
        RECT 100.665 143.160 101.430 143.300 ;
        RECT 100.665 143.115 100.955 143.160 ;
        RECT 101.110 143.100 101.430 143.160 ;
        RECT 104.790 143.100 105.110 143.360 ;
        RECT 105.800 143.345 105.940 143.500 ;
        RECT 112.150 143.500 134.090 143.640 ;
        RECT 112.150 143.440 112.470 143.500 ;
        RECT 105.725 143.115 106.015 143.345 ;
        RECT 113.500 143.300 113.790 143.345 ;
        RECT 117.210 143.300 117.530 143.360 ;
        RECT 113.500 143.160 117.530 143.300 ;
        RECT 113.500 143.115 113.790 143.160 ;
        RECT 117.210 143.100 117.530 143.160 ;
        RECT 120.905 143.300 121.195 143.345 ;
        RECT 121.350 143.300 121.670 143.360 ;
        RECT 120.905 143.160 121.670 143.300 ;
        RECT 120.905 143.115 121.195 143.160 ;
        RECT 121.350 143.100 121.670 143.160 ;
        RECT 121.825 143.115 122.115 143.345 ;
        RECT 39.010 142.960 39.330 143.020 ;
        RECT 35.880 142.820 39.330 142.960 ;
        RECT 34.040 142.665 34.180 142.820 ;
        RECT 35.330 142.760 35.650 142.820 ;
        RECT 39.010 142.760 39.330 142.820 ;
        RECT 61.065 142.960 61.355 143.005 ;
        RECT 62.255 142.960 62.545 143.005 ;
        RECT 64.775 142.960 65.065 143.005 ;
        RECT 61.065 142.820 65.065 142.960 ;
        RECT 61.065 142.775 61.355 142.820 ;
        RECT 62.255 142.775 62.545 142.820 ;
        RECT 64.775 142.775 65.065 142.820 ;
        RECT 72.605 142.960 72.895 143.005 ;
        RECT 75.350 142.960 75.670 143.020 ;
        RECT 72.605 142.820 75.670 142.960 ;
        RECT 72.605 142.775 72.895 142.820 ;
        RECT 75.350 142.760 75.670 142.820 ;
        RECT 75.825 142.775 76.115 143.005 ;
        RECT 78.110 142.960 78.430 143.020 ;
        RECT 79.045 142.960 79.335 143.005 ;
        RECT 78.110 142.820 79.335 142.960 ;
        RECT 33.965 142.435 34.255 142.665 ;
        RECT 60.670 142.620 60.960 142.665 ;
        RECT 62.770 142.620 63.060 142.665 ;
        RECT 64.340 142.620 64.630 142.665 ;
        RECT 60.670 142.480 64.630 142.620 ;
        RECT 75.900 142.620 76.040 142.775 ;
        RECT 78.110 142.760 78.430 142.820 ;
        RECT 79.045 142.775 79.335 142.820 ;
        RECT 79.490 142.760 79.810 143.020 ;
        RECT 84.115 142.960 84.405 143.005 ;
        RECT 86.635 142.960 86.925 143.005 ;
        RECT 87.825 142.960 88.115 143.005 ;
        RECT 84.115 142.820 88.115 142.960 ;
        RECT 84.115 142.775 84.405 142.820 ;
        RECT 86.635 142.775 86.925 142.820 ;
        RECT 87.825 142.775 88.115 142.820 ;
        RECT 93.750 142.760 94.070 143.020 ;
        RECT 94.225 142.960 94.515 143.005 ;
        RECT 95.145 142.960 95.435 143.005 ;
        RECT 94.225 142.820 95.435 142.960 ;
        RECT 94.225 142.775 94.515 142.820 ;
        RECT 95.145 142.775 95.435 142.820 ;
        RECT 103.425 142.960 103.715 143.005 ;
        RECT 106.185 142.960 106.475 143.005 ;
        RECT 103.425 142.820 106.475 142.960 ;
        RECT 103.425 142.775 103.715 142.820 ;
        RECT 106.185 142.775 106.475 142.820 ;
        RECT 109.390 142.960 109.710 143.020 ;
        RECT 112.150 142.960 112.470 143.020 ;
        RECT 109.390 142.820 112.470 142.960 ;
        RECT 109.390 142.760 109.710 142.820 ;
        RECT 112.150 142.760 112.470 142.820 ;
        RECT 113.045 142.960 113.335 143.005 ;
        RECT 114.235 142.960 114.525 143.005 ;
        RECT 116.755 142.960 117.045 143.005 ;
        RECT 113.045 142.820 117.045 142.960 ;
        RECT 113.045 142.775 113.335 142.820 ;
        RECT 114.235 142.775 114.525 142.820 ;
        RECT 116.755 142.775 117.045 142.820 ;
        RECT 120.430 142.960 120.750 143.020 ;
        RECT 121.900 142.960 122.040 143.115 ;
        RECT 122.270 143.100 122.590 143.360 ;
        RECT 122.745 143.300 123.035 143.345 ;
        RECT 123.650 143.300 123.970 143.360 ;
        RECT 124.200 143.345 124.340 143.500 ;
        RECT 133.770 143.440 134.090 143.500 ;
        RECT 139.840 143.500 142.280 143.640 ;
        RECT 125.490 143.345 125.810 143.360 ;
        RECT 122.745 143.160 123.970 143.300 ;
        RECT 122.745 143.115 123.035 143.160 ;
        RECT 123.650 143.100 123.970 143.160 ;
        RECT 124.125 143.115 124.415 143.345 ;
        RECT 125.460 143.300 125.810 143.345 ;
        RECT 125.295 143.160 125.810 143.300 ;
        RECT 125.460 143.115 125.810 143.160 ;
        RECT 125.490 143.100 125.810 143.115 ;
        RECT 137.450 143.100 137.770 143.360 ;
        RECT 139.840 143.345 139.980 143.500 ;
        RECT 142.140 143.360 142.280 143.500 ;
        RECT 139.765 143.115 140.055 143.345 ;
        RECT 140.210 143.100 140.530 143.360 ;
        RECT 142.050 143.100 142.370 143.360 ;
        RECT 120.430 142.820 122.040 142.960 ;
        RECT 125.005 142.960 125.295 143.005 ;
        RECT 126.195 142.960 126.485 143.005 ;
        RECT 128.715 142.960 129.005 143.005 ;
        RECT 143.890 142.960 144.210 143.020 ;
        RECT 125.005 142.820 129.005 142.960 ;
        RECT 120.430 142.760 120.750 142.820 ;
        RECT 125.005 142.775 125.295 142.820 ;
        RECT 126.195 142.775 126.485 142.820 ;
        RECT 128.715 142.775 129.005 142.820 ;
        RECT 138.460 142.820 144.210 142.960 ;
        RECT 79.580 142.620 79.720 142.760 ;
        RECT 75.900 142.480 79.720 142.620 ;
        RECT 84.550 142.620 84.840 142.665 ;
        RECT 86.120 142.620 86.410 142.665 ;
        RECT 88.220 142.620 88.510 142.665 ;
        RECT 84.550 142.480 88.510 142.620 ;
        RECT 60.670 142.435 60.960 142.480 ;
        RECT 62.770 142.435 63.060 142.480 ;
        RECT 64.340 142.435 64.630 142.480 ;
        RECT 84.550 142.435 84.840 142.480 ;
        RECT 86.120 142.435 86.410 142.480 ;
        RECT 88.220 142.435 88.510 142.480 ;
        RECT 91.925 142.620 92.215 142.665 ;
        RECT 94.670 142.620 94.990 142.680 ;
        RECT 138.460 142.665 138.600 142.820 ;
        RECT 143.890 142.760 144.210 142.820 ;
        RECT 91.925 142.480 94.990 142.620 ;
        RECT 91.925 142.435 92.215 142.480 ;
        RECT 32.110 142.280 32.430 142.340 ;
        RECT 34.040 142.280 34.180 142.435 ;
        RECT 94.670 142.420 94.990 142.480 ;
        RECT 112.650 142.620 112.940 142.665 ;
        RECT 114.750 142.620 115.040 142.665 ;
        RECT 116.320 142.620 116.610 142.665 ;
        RECT 112.650 142.480 116.610 142.620 ;
        RECT 112.650 142.435 112.940 142.480 ;
        RECT 114.750 142.435 115.040 142.480 ;
        RECT 116.320 142.435 116.610 142.480 ;
        RECT 124.610 142.620 124.900 142.665 ;
        RECT 126.710 142.620 127.000 142.665 ;
        RECT 128.280 142.620 128.570 142.665 ;
        RECT 124.610 142.480 128.570 142.620 ;
        RECT 124.610 142.435 124.900 142.480 ;
        RECT 126.710 142.435 127.000 142.480 ;
        RECT 128.280 142.435 128.570 142.480 ;
        RECT 138.385 142.435 138.675 142.665 ;
        RECT 32.110 142.140 34.180 142.280 ;
        RECT 34.425 142.280 34.715 142.325 ;
        RECT 35.330 142.280 35.650 142.340 ;
        RECT 34.425 142.140 35.650 142.280 ;
        RECT 32.110 142.080 32.430 142.140 ;
        RECT 34.425 142.095 34.715 142.140 ;
        RECT 35.330 142.080 35.650 142.140 ;
        RECT 38.550 142.080 38.870 142.340 ;
        RECT 54.650 142.280 54.970 142.340 ;
        RECT 55.125 142.280 55.415 142.325 ;
        RECT 54.650 142.140 55.415 142.280 ;
        RECT 54.650 142.080 54.970 142.140 ;
        RECT 55.125 142.095 55.415 142.140 ;
        RECT 58.330 142.080 58.650 142.340 ;
        RECT 73.510 142.080 73.830 142.340 ;
        RECT 76.730 142.080 77.050 142.340 ;
        RECT 81.805 142.280 82.095 142.325 ;
        RECT 83.630 142.280 83.950 142.340 ;
        RECT 81.805 142.140 83.950 142.280 ;
        RECT 81.805 142.095 82.095 142.140 ;
        RECT 83.630 142.080 83.950 142.140 ;
        RECT 94.210 142.280 94.530 142.340 ;
        RECT 103.885 142.280 104.175 142.325 ;
        RECT 94.210 142.140 104.175 142.280 ;
        RECT 94.210 142.080 94.530 142.140 ;
        RECT 103.885 142.095 104.175 142.140 ;
        RECT 17.320 141.460 147.040 141.940 ;
        RECT 34.425 141.260 34.715 141.305 ;
        RECT 35.790 141.260 36.110 141.320 ;
        RECT 34.425 141.120 36.110 141.260 ;
        RECT 34.425 141.075 34.715 141.120 ;
        RECT 35.790 141.060 36.110 141.120 ;
        RECT 40.850 141.260 41.170 141.320 ;
        RECT 42.705 141.260 42.995 141.305 ;
        RECT 40.850 141.120 42.995 141.260 ;
        RECT 40.850 141.060 41.170 141.120 ;
        RECT 42.705 141.075 42.995 141.120 ;
        RECT 52.825 141.260 53.115 141.305 ;
        RECT 58.330 141.260 58.650 141.320 ;
        RECT 52.825 141.120 58.650 141.260 ;
        RECT 52.825 141.075 53.115 141.120 ;
        RECT 58.330 141.060 58.650 141.120 ;
        RECT 64.770 141.260 65.090 141.320 ;
        RECT 67.085 141.260 67.375 141.305 ;
        RECT 64.770 141.120 67.375 141.260 ;
        RECT 64.770 141.060 65.090 141.120 ;
        RECT 67.085 141.075 67.375 141.120 ;
        RECT 68.005 141.075 68.295 141.305 ;
        RECT 76.730 141.260 77.050 141.320 ;
        RECT 70.840 141.120 77.050 141.260 ;
        RECT 36.290 140.920 36.580 140.965 ;
        RECT 38.390 140.920 38.680 140.965 ;
        RECT 39.960 140.920 40.250 140.965 ;
        RECT 36.290 140.780 40.250 140.920 ;
        RECT 36.290 140.735 36.580 140.780 ;
        RECT 38.390 140.735 38.680 140.780 ;
        RECT 39.960 140.735 40.250 140.780 ;
        RECT 53.730 140.920 54.050 140.980 ;
        RECT 56.490 140.920 56.810 140.980 ;
        RECT 66.150 140.920 66.470 140.980 ;
        RECT 68.080 140.920 68.220 141.075 ;
        RECT 53.730 140.780 54.880 140.920 ;
        RECT 53.730 140.720 54.050 140.780 ;
        RECT 34.870 140.580 35.190 140.640 ;
        RECT 35.790 140.580 36.110 140.640 ;
        RECT 34.870 140.440 36.110 140.580 ;
        RECT 34.870 140.380 35.190 140.440 ;
        RECT 35.790 140.380 36.110 140.440 ;
        RECT 36.685 140.580 36.975 140.625 ;
        RECT 37.875 140.580 38.165 140.625 ;
        RECT 40.395 140.580 40.685 140.625 ;
        RECT 36.685 140.440 40.685 140.580 ;
        RECT 36.685 140.395 36.975 140.440 ;
        RECT 37.875 140.395 38.165 140.440 ;
        RECT 40.395 140.395 40.685 140.440 ;
        RECT 52.810 140.580 53.130 140.640 ;
        RECT 54.740 140.625 54.880 140.780 ;
        RECT 55.200 140.780 64.080 140.920 ;
        RECT 55.200 140.640 55.340 140.780 ;
        RECT 56.490 140.720 56.810 140.780 ;
        RECT 54.205 140.580 54.495 140.625 ;
        RECT 52.810 140.440 54.495 140.580 ;
        RECT 52.810 140.380 53.130 140.440 ;
        RECT 54.205 140.395 54.495 140.440 ;
        RECT 54.665 140.395 54.955 140.625 ;
        RECT 32.585 140.240 32.875 140.285 ;
        RECT 38.550 140.240 38.870 140.300 ;
        RECT 32.585 140.100 38.870 140.240 ;
        RECT 32.585 140.055 32.875 140.100 ;
        RECT 38.550 140.040 38.870 140.100 ;
        RECT 50.050 140.240 50.370 140.300 ;
        RECT 53.745 140.240 54.035 140.285 ;
        RECT 50.050 140.100 54.035 140.240 ;
        RECT 54.740 140.240 54.880 140.395 ;
        RECT 55.110 140.380 55.430 140.640 ;
        RECT 60.170 140.580 60.490 140.640 ;
        RECT 61.565 140.580 61.855 140.625 ;
        RECT 62.470 140.580 62.790 140.640 ;
        RECT 60.170 140.440 63.620 140.580 ;
        RECT 60.170 140.380 60.490 140.440 ;
        RECT 61.565 140.395 61.855 140.440 ;
        RECT 62.470 140.380 62.790 140.440 ;
        RECT 62.930 140.240 63.250 140.300 ;
        RECT 63.480 140.285 63.620 140.440 ;
        RECT 54.740 140.100 63.250 140.240 ;
        RECT 50.050 140.040 50.370 140.100 ;
        RECT 53.745 140.055 54.035 140.100 ;
        RECT 62.930 140.040 63.250 140.100 ;
        RECT 63.405 140.055 63.695 140.285 ;
        RECT 63.940 140.240 64.080 140.780 ;
        RECT 66.150 140.780 68.220 140.920 ;
        RECT 66.150 140.720 66.470 140.780 ;
        RECT 68.910 140.580 69.230 140.640 ;
        RECT 70.840 140.625 70.980 141.120 ;
        RECT 76.730 141.060 77.050 141.120 ;
        RECT 85.930 141.060 86.250 141.320 ;
        RECT 86.390 141.260 86.710 141.320 ;
        RECT 88.705 141.260 88.995 141.305 ;
        RECT 86.390 141.120 88.995 141.260 ;
        RECT 86.390 141.060 86.710 141.120 ;
        RECT 88.705 141.075 88.995 141.120 ;
        RECT 97.445 141.260 97.735 141.305 ;
        RECT 101.110 141.260 101.430 141.320 ;
        RECT 97.445 141.120 101.430 141.260 ;
        RECT 97.445 141.075 97.735 141.120 ;
        RECT 101.110 141.060 101.430 141.120 ;
        RECT 123.205 141.260 123.495 141.305 ;
        RECT 126.870 141.260 127.190 141.320 ;
        RECT 123.205 141.120 127.190 141.260 ;
        RECT 123.205 141.075 123.495 141.120 ;
        RECT 126.870 141.060 127.190 141.120 ;
        RECT 134.230 141.260 134.550 141.320 ;
        RECT 142.525 141.260 142.815 141.305 ;
        RECT 134.230 141.120 142.815 141.260 ;
        RECT 134.230 141.060 134.550 141.120 ;
        RECT 142.525 141.075 142.815 141.120 ;
        RECT 144.810 141.060 145.130 141.320 ;
        RECT 71.710 140.920 72.000 140.965 ;
        RECT 73.810 140.920 74.100 140.965 ;
        RECT 75.380 140.920 75.670 140.965 ;
        RECT 71.710 140.780 75.670 140.920 ;
        RECT 71.710 140.735 72.000 140.780 ;
        RECT 73.810 140.735 74.100 140.780 ;
        RECT 75.380 140.735 75.670 140.780 ;
        RECT 78.110 140.920 78.430 140.980 ;
        RECT 91.030 140.920 91.320 140.965 ;
        RECT 93.130 140.920 93.420 140.965 ;
        RECT 94.700 140.920 94.990 140.965 ;
        RECT 78.110 140.780 82.940 140.920 ;
        RECT 78.110 140.720 78.430 140.780 ;
        RECT 68.910 140.440 69.600 140.580 ;
        RECT 68.910 140.380 69.230 140.440 ;
        RECT 69.460 140.285 69.600 140.440 ;
        RECT 70.765 140.395 71.055 140.625 ;
        RECT 72.105 140.580 72.395 140.625 ;
        RECT 73.295 140.580 73.585 140.625 ;
        RECT 75.815 140.580 76.105 140.625 ;
        RECT 72.105 140.440 76.105 140.580 ;
        RECT 72.105 140.395 72.395 140.440 ;
        RECT 73.295 140.395 73.585 140.440 ;
        RECT 75.815 140.395 76.105 140.440 ;
        RECT 77.190 140.580 77.510 140.640 ;
        RECT 82.800 140.625 82.940 140.780 ;
        RECT 91.030 140.780 94.990 140.920 ;
        RECT 91.030 140.735 91.320 140.780 ;
        RECT 93.130 140.735 93.420 140.780 ;
        RECT 94.700 140.735 94.990 140.780 ;
        RECT 102.490 140.720 102.810 140.980 ;
        RECT 106.170 140.720 106.490 140.980 ;
        RECT 118.590 140.920 118.910 140.980 ;
        RECT 124.125 140.920 124.415 140.965 ;
        RECT 129.630 140.920 129.950 140.980 ;
        RECT 118.590 140.780 123.420 140.920 ;
        RECT 118.590 140.720 118.910 140.780 ;
        RECT 81.345 140.580 81.635 140.625 ;
        RECT 77.190 140.440 81.635 140.580 ;
        RECT 77.190 140.380 77.510 140.440 ;
        RECT 81.345 140.395 81.635 140.440 ;
        RECT 82.725 140.395 83.015 140.625 ;
        RECT 83.630 140.380 83.950 140.640 ;
        RECT 90.530 140.380 90.850 140.640 ;
        RECT 91.425 140.580 91.715 140.625 ;
        RECT 92.615 140.580 92.905 140.625 ;
        RECT 95.135 140.580 95.425 140.625 ;
        RECT 122.730 140.580 123.050 140.640 ;
        RECT 91.425 140.440 95.425 140.580 ;
        RECT 91.425 140.395 91.715 140.440 ;
        RECT 92.615 140.395 92.905 140.440 ;
        RECT 95.135 140.395 95.425 140.440 ;
        RECT 120.520 140.440 123.050 140.580 ;
        RECT 123.280 140.580 123.420 140.780 ;
        RECT 124.125 140.780 129.950 140.920 ;
        RECT 124.125 140.735 124.415 140.780 ;
        RECT 129.630 140.720 129.950 140.780 ;
        RECT 128.710 140.580 129.030 140.640 ;
        RECT 136.070 140.580 136.390 140.640 ;
        RECT 137.465 140.580 137.755 140.625 ;
        RECT 123.280 140.440 123.880 140.580 ;
        RECT 63.940 140.100 69.140 140.240 ;
        RECT 32.110 139.900 32.430 139.960 ;
        RECT 34.425 139.900 34.715 139.945 ;
        RECT 34.870 139.900 35.190 139.960 ;
        RECT 37.030 139.900 37.320 139.945 ;
        RECT 32.110 139.760 35.190 139.900 ;
        RECT 32.110 139.700 32.430 139.760 ;
        RECT 34.425 139.715 34.715 139.760 ;
        RECT 34.870 139.700 35.190 139.760 ;
        RECT 35.420 139.760 37.320 139.900 ;
        RECT 35.420 139.605 35.560 139.760 ;
        RECT 37.030 139.715 37.320 139.760 ;
        RECT 44.990 139.700 45.310 139.960 ;
        RECT 49.145 139.900 49.435 139.945 ;
        RECT 57.885 139.900 58.175 139.945 ;
        RECT 66.610 139.900 66.930 139.960 ;
        RECT 69.000 139.945 69.140 140.100 ;
        RECT 69.385 140.055 69.675 140.285 ;
        RECT 69.845 140.055 70.135 140.285 ;
        RECT 70.290 140.240 70.610 140.300 ;
        RECT 71.225 140.240 71.515 140.285 ;
        RECT 70.290 140.100 71.515 140.240 ;
        RECT 49.145 139.760 66.930 139.900 ;
        RECT 49.145 139.715 49.435 139.760 ;
        RECT 57.885 139.715 58.175 139.760 ;
        RECT 66.610 139.700 66.930 139.760 ;
        RECT 68.925 139.715 69.215 139.945 ;
        RECT 35.345 139.375 35.635 139.605 ;
        RECT 55.570 139.560 55.890 139.620 ;
        RECT 64.770 139.560 65.090 139.620 ;
        RECT 67.875 139.560 68.165 139.605 ;
        RECT 55.570 139.420 68.165 139.560 ;
        RECT 69.920 139.560 70.060 140.055 ;
        RECT 70.290 140.040 70.610 140.100 ;
        RECT 71.225 140.055 71.515 140.100 ;
        RECT 79.490 140.040 79.810 140.300 ;
        RECT 80.410 140.240 80.730 140.300 ;
        RECT 86.405 140.240 86.695 140.285 ;
        RECT 80.410 140.100 86.695 140.240 ;
        RECT 80.410 140.040 80.730 140.100 ;
        RECT 86.405 140.055 86.695 140.100 ;
        RECT 87.770 140.040 88.090 140.300 ;
        RECT 91.880 140.240 92.170 140.285 ;
        RECT 94.210 140.240 94.530 140.300 ;
        RECT 91.880 140.100 94.530 140.240 ;
        RECT 91.880 140.055 92.170 140.100 ;
        RECT 94.210 140.040 94.530 140.100 ;
        RECT 98.810 140.240 99.130 140.300 ;
        RECT 100.205 140.240 100.495 140.285 ;
        RECT 102.950 140.240 103.270 140.300 ;
        RECT 119.510 140.240 119.830 140.300 ;
        RECT 120.520 140.285 120.660 140.440 ;
        RECT 122.730 140.380 123.050 140.440 ;
        RECT 98.810 140.100 103.270 140.240 ;
        RECT 98.810 140.040 99.130 140.100 ;
        RECT 100.205 140.055 100.495 140.100 ;
        RECT 102.950 140.040 103.270 140.100 ;
        RECT 103.500 140.100 119.830 140.240 ;
        RECT 70.765 139.900 71.055 139.945 ;
        RECT 72.450 139.900 72.740 139.945 ;
        RECT 70.765 139.760 72.740 139.900 ;
        RECT 70.765 139.715 71.055 139.760 ;
        RECT 72.450 139.715 72.740 139.760 ;
        RECT 78.570 139.700 78.890 139.960 ;
        RECT 79.030 139.900 79.350 139.960 ;
        RECT 79.965 139.900 80.255 139.945 ;
        RECT 79.030 139.760 80.255 139.900 ;
        RECT 79.030 139.700 79.350 139.760 ;
        RECT 79.965 139.715 80.255 139.760 ;
        RECT 81.790 139.900 82.110 139.960 ;
        RECT 84.105 139.900 84.395 139.945 ;
        RECT 81.790 139.760 84.395 139.900 ;
        RECT 81.790 139.700 82.110 139.760 ;
        RECT 84.105 139.715 84.395 139.760 ;
        RECT 88.230 139.900 88.550 139.960 ;
        RECT 98.365 139.900 98.655 139.945 ;
        RECT 103.500 139.900 103.640 140.100 ;
        RECT 119.510 140.040 119.830 140.100 ;
        RECT 120.445 140.055 120.735 140.285 ;
        RECT 121.350 140.040 121.670 140.300 ;
        RECT 121.810 140.040 122.130 140.300 ;
        RECT 122.285 140.240 122.575 140.285 ;
        RECT 123.190 140.240 123.510 140.300 ;
        RECT 123.740 140.285 123.880 140.440 ;
        RECT 124.200 140.440 132.160 140.580 ;
        RECT 124.200 140.300 124.340 140.440 ;
        RECT 128.710 140.380 129.030 140.440 ;
        RECT 122.285 140.100 123.510 140.240 ;
        RECT 122.285 140.055 122.575 140.100 ;
        RECT 123.190 140.040 123.510 140.100 ;
        RECT 123.665 140.055 123.955 140.285 ;
        RECT 124.110 140.040 124.430 140.300 ;
        RECT 124.585 140.240 124.875 140.285 ;
        RECT 125.950 140.240 126.270 140.300 ;
        RECT 124.585 140.100 126.270 140.240 ;
        RECT 124.585 140.055 124.875 140.100 ;
        RECT 125.950 140.040 126.270 140.100 ;
        RECT 130.090 140.040 130.410 140.300 ;
        RECT 130.550 140.240 130.870 140.300 ;
        RECT 132.020 140.285 132.160 140.440 ;
        RECT 136.070 140.440 137.755 140.580 ;
        RECT 136.070 140.380 136.390 140.440 ;
        RECT 137.465 140.395 137.755 140.440 ;
        RECT 131.025 140.240 131.315 140.285 ;
        RECT 130.550 140.100 131.315 140.240 ;
        RECT 130.550 140.040 130.870 140.100 ;
        RECT 131.025 140.055 131.315 140.100 ;
        RECT 131.945 140.055 132.235 140.285 ;
        RECT 140.210 140.240 140.530 140.300 ;
        RECT 141.605 140.240 141.895 140.285 ;
        RECT 140.210 140.100 141.895 140.240 ;
        RECT 140.210 140.040 140.530 140.100 ;
        RECT 141.605 140.055 141.895 140.100 ;
        RECT 143.430 140.040 143.750 140.300 ;
        RECT 143.890 140.040 144.210 140.300 ;
        RECT 88.230 139.760 103.640 139.900 ;
        RECT 103.885 139.900 104.175 139.945 ;
        RECT 104.345 139.900 104.635 139.945 ;
        RECT 131.485 139.900 131.775 139.945 ;
        RECT 136.545 139.900 136.835 139.945 ;
        RECT 103.885 139.760 130.320 139.900 ;
        RECT 88.230 139.700 88.550 139.760 ;
        RECT 98.365 139.715 98.655 139.760 ;
        RECT 103.885 139.715 104.175 139.760 ;
        RECT 104.345 139.715 104.635 139.760 ;
        RECT 130.180 139.620 130.320 139.760 ;
        RECT 131.485 139.760 132.160 139.900 ;
        RECT 131.485 139.715 131.775 139.760 ;
        RECT 132.020 139.620 132.160 139.760 ;
        RECT 132.940 139.760 136.835 139.900 ;
        RECT 76.270 139.560 76.590 139.620 ;
        RECT 69.920 139.420 76.590 139.560 ;
        RECT 55.570 139.360 55.890 139.420 ;
        RECT 64.770 139.360 65.090 139.420 ;
        RECT 67.875 139.375 68.165 139.420 ;
        RECT 76.270 139.360 76.590 139.420 ;
        RECT 78.125 139.560 78.415 139.605 ;
        RECT 79.490 139.560 79.810 139.620 ;
        RECT 78.125 139.420 79.810 139.560 ;
        RECT 78.125 139.375 78.415 139.420 ;
        RECT 79.490 139.360 79.810 139.420 ;
        RECT 86.390 139.560 86.710 139.620 ;
        RECT 86.865 139.560 87.155 139.605 ;
        RECT 86.390 139.420 87.155 139.560 ;
        RECT 86.390 139.360 86.710 139.420 ;
        RECT 86.865 139.375 87.155 139.420 ;
        RECT 101.570 139.360 101.890 139.620 ;
        RECT 106.630 139.360 106.950 139.620 ;
        RECT 130.090 139.360 130.410 139.620 ;
        RECT 131.930 139.360 132.250 139.620 ;
        RECT 132.940 139.605 133.080 139.760 ;
        RECT 136.545 139.715 136.835 139.760 ;
        RECT 132.865 139.375 133.155 139.605 ;
        RECT 134.690 139.360 135.010 139.620 ;
        RECT 137.005 139.560 137.295 139.605 ;
        RECT 138.845 139.560 139.135 139.605 ;
        RECT 137.005 139.420 139.135 139.560 ;
        RECT 137.005 139.375 137.295 139.420 ;
        RECT 138.845 139.375 139.135 139.420 ;
        RECT 17.320 138.740 147.040 139.220 ;
        RECT 29.350 138.340 29.670 138.600 ;
        RECT 35.330 138.540 35.650 138.600 ;
        RECT 34.960 138.400 35.650 138.540 ;
        RECT 34.960 138.245 35.100 138.400 ;
        RECT 35.330 138.340 35.650 138.400 ;
        RECT 39.470 138.540 39.790 138.600 ;
        RECT 42.230 138.540 42.550 138.600 ;
        RECT 39.470 138.400 42.550 138.540 ;
        RECT 39.470 138.340 39.790 138.400 ;
        RECT 42.230 138.340 42.550 138.400 ;
        RECT 55.110 138.540 55.430 138.600 ;
        RECT 55.585 138.540 55.875 138.585 ;
        RECT 66.150 138.540 66.470 138.600 ;
        RECT 55.110 138.400 55.875 138.540 ;
        RECT 55.110 138.340 55.430 138.400 ;
        RECT 55.585 138.355 55.875 138.400 ;
        RECT 63.940 138.400 66.470 138.540 ;
        RECT 34.930 138.015 35.220 138.245 ;
        RECT 44.990 138.200 45.310 138.260 ;
        RECT 53.285 138.200 53.575 138.245 ;
        RECT 57.410 138.200 57.730 138.260 ;
        RECT 36.340 138.060 45.680 138.200 ;
        RECT 20.165 137.860 20.455 137.905 ;
        RECT 22.910 137.860 23.230 137.920 ;
        RECT 20.165 137.720 23.230 137.860 ;
        RECT 20.165 137.675 20.455 137.720 ;
        RECT 22.910 137.660 23.230 137.720 ;
        RECT 35.790 137.860 36.110 137.920 ;
        RECT 36.340 137.905 36.480 138.060 ;
        RECT 44.990 138.000 45.310 138.060 ;
        RECT 36.265 137.860 36.555 137.905 ;
        RECT 35.790 137.720 36.555 137.860 ;
        RECT 35.790 137.660 36.110 137.720 ;
        RECT 36.265 137.675 36.555 137.720 ;
        RECT 39.025 137.860 39.315 137.905 ;
        RECT 39.470 137.860 39.790 137.920 ;
        RECT 39.025 137.720 39.790 137.860 ;
        RECT 39.025 137.675 39.315 137.720 ;
        RECT 39.470 137.660 39.790 137.720 ;
        RECT 39.945 137.675 40.235 137.905 ;
        RECT 41.325 137.675 41.615 137.905 ;
        RECT 31.675 137.520 31.965 137.565 ;
        RECT 34.195 137.520 34.485 137.565 ;
        RECT 35.385 137.520 35.675 137.565 ;
        RECT 31.675 137.380 35.675 137.520 ;
        RECT 31.675 137.335 31.965 137.380 ;
        RECT 34.195 137.335 34.485 137.380 ;
        RECT 35.385 137.335 35.675 137.380 ;
        RECT 38.550 137.520 38.870 137.580 ;
        RECT 40.020 137.520 40.160 137.675 ;
        RECT 38.550 137.380 40.160 137.520 ;
        RECT 41.400 137.520 41.540 137.675 ;
        RECT 42.230 137.660 42.550 137.920 ;
        RECT 42.690 137.660 43.010 137.920 ;
        RECT 45.540 137.905 45.680 138.060 ;
        RECT 53.285 138.060 57.730 138.200 ;
        RECT 53.285 138.015 53.575 138.060 ;
        RECT 57.410 138.000 57.730 138.060 ;
        RECT 61.090 138.245 61.410 138.260 ;
        RECT 61.090 138.200 61.440 138.245 ;
        RECT 62.930 138.200 63.250 138.260 ;
        RECT 63.940 138.245 64.080 138.400 ;
        RECT 66.150 138.340 66.470 138.400 ;
        RECT 77.205 138.540 77.495 138.585 ;
        RECT 79.030 138.540 79.350 138.600 ;
        RECT 77.205 138.400 79.350 138.540 ;
        RECT 77.205 138.355 77.495 138.400 ;
        RECT 79.030 138.340 79.350 138.400 ;
        RECT 81.805 138.540 82.095 138.585 ;
        RECT 87.770 138.540 88.090 138.600 ;
        RECT 81.805 138.400 88.090 138.540 ;
        RECT 81.805 138.355 82.095 138.400 ;
        RECT 87.770 138.340 88.090 138.400 ;
        RECT 100.665 138.540 100.955 138.585 ;
        RECT 104.790 138.540 105.110 138.600 ;
        RECT 100.665 138.400 105.110 138.540 ;
        RECT 100.665 138.355 100.955 138.400 ;
        RECT 104.790 138.340 105.110 138.400 ;
        RECT 105.710 138.540 106.030 138.600 ;
        RECT 108.945 138.540 109.235 138.585 ;
        RECT 139.750 138.540 140.070 138.600 ;
        RECT 105.710 138.400 140.070 138.540 ;
        RECT 105.710 138.340 106.030 138.400 ;
        RECT 108.945 138.355 109.235 138.400 ;
        RECT 139.750 138.340 140.070 138.400 ;
        RECT 140.210 138.340 140.530 138.600 ;
        RECT 141.605 138.355 141.895 138.585 ;
        RECT 63.865 138.200 64.155 138.245 ;
        RECT 61.090 138.060 61.605 138.200 ;
        RECT 62.930 138.060 64.155 138.200 ;
        RECT 61.090 138.015 61.440 138.060 ;
        RECT 61.090 138.000 61.410 138.015 ;
        RECT 62.930 138.000 63.250 138.060 ;
        RECT 63.865 138.015 64.155 138.060 ;
        RECT 64.770 138.000 65.090 138.260 ;
        RECT 71.640 138.200 71.930 138.245 ;
        RECT 73.510 138.200 73.830 138.260 ;
        RECT 71.640 138.060 73.830 138.200 ;
        RECT 71.640 138.015 71.930 138.060 ;
        RECT 73.510 138.000 73.830 138.060 ;
        RECT 78.570 138.200 78.890 138.260 ;
        RECT 101.570 138.200 101.890 138.260 ;
        RECT 103.270 138.200 103.560 138.245 ;
        RECT 78.570 138.060 86.620 138.200 ;
        RECT 78.570 138.000 78.890 138.060 ;
        RECT 45.465 137.675 45.755 137.905 ;
        RECT 50.050 137.660 50.370 137.920 ;
        RECT 50.985 137.860 51.275 137.905 ;
        RECT 51.445 137.860 51.735 137.905 ;
        RECT 55.570 137.860 55.890 137.920 ;
        RECT 50.985 137.720 55.890 137.860 ;
        RECT 50.985 137.675 51.275 137.720 ;
        RECT 51.445 137.675 51.735 137.720 ;
        RECT 55.570 137.660 55.890 137.720 ;
        RECT 62.470 137.660 62.790 137.920 ;
        RECT 68.910 137.860 69.230 137.920 ;
        RECT 79.950 137.860 80.270 137.920 ;
        RECT 86.480 137.905 86.620 138.060 ;
        RECT 99.360 138.060 100.420 138.200 ;
        RECT 85.945 137.860 86.235 137.905 ;
        RECT 68.910 137.720 79.720 137.860 ;
        RECT 68.910 137.660 69.230 137.720 ;
        RECT 46.830 137.520 47.150 137.580 ;
        RECT 41.400 137.380 47.150 137.520 ;
        RECT 38.550 137.320 38.870 137.380 ;
        RECT 32.110 137.180 32.400 137.225 ;
        RECT 33.680 137.180 33.970 137.225 ;
        RECT 35.780 137.180 36.070 137.225 ;
        RECT 32.110 137.040 36.070 137.180 ;
        RECT 40.020 137.180 40.160 137.380 ;
        RECT 46.830 137.320 47.150 137.380 ;
        RECT 49.145 137.520 49.435 137.565 ;
        RECT 52.810 137.520 53.130 137.580 ;
        RECT 49.145 137.380 53.130 137.520 ;
        RECT 49.145 137.335 49.435 137.380 ;
        RECT 52.810 137.320 53.130 137.380 ;
        RECT 57.895 137.520 58.185 137.565 ;
        RECT 60.415 137.520 60.705 137.565 ;
        RECT 61.605 137.520 61.895 137.565 ;
        RECT 57.895 137.380 61.895 137.520 ;
        RECT 57.895 137.335 58.185 137.380 ;
        RECT 60.415 137.335 60.705 137.380 ;
        RECT 61.605 137.335 61.895 137.380 ;
        RECT 70.290 137.320 70.610 137.580 ;
        RECT 71.185 137.520 71.475 137.565 ;
        RECT 72.375 137.520 72.665 137.565 ;
        RECT 74.895 137.520 75.185 137.565 ;
        RECT 71.185 137.380 75.185 137.520 ;
        RECT 71.185 137.335 71.475 137.380 ;
        RECT 72.375 137.335 72.665 137.380 ;
        RECT 74.895 137.335 75.185 137.380 ;
        RECT 79.030 137.320 79.350 137.580 ;
        RECT 79.580 137.520 79.720 137.720 ;
        RECT 79.950 137.720 86.235 137.860 ;
        RECT 79.950 137.660 80.270 137.720 ;
        RECT 85.945 137.675 86.235 137.720 ;
        RECT 86.405 137.675 86.695 137.905 ;
        RECT 97.430 137.860 97.750 137.920 ;
        RECT 97.905 137.860 98.195 137.905 ;
        RECT 97.430 137.720 98.195 137.860 ;
        RECT 97.430 137.660 97.750 137.720 ;
        RECT 97.905 137.675 98.195 137.720 ;
        RECT 98.365 137.860 98.655 137.905 ;
        RECT 98.810 137.860 99.130 137.920 ;
        RECT 99.360 137.905 99.500 138.060 ;
        RECT 98.365 137.720 99.130 137.860 ;
        RECT 98.365 137.675 98.655 137.720 ;
        RECT 98.810 137.660 99.130 137.720 ;
        RECT 99.285 137.675 99.575 137.905 ;
        RECT 99.730 137.660 100.050 137.920 ;
        RECT 100.280 137.860 100.420 138.060 ;
        RECT 101.570 138.060 103.560 138.200 ;
        RECT 101.570 138.000 101.890 138.060 ;
        RECT 103.270 138.015 103.560 138.060 ;
        RECT 106.630 138.200 106.950 138.260 ;
        RECT 110.630 138.200 110.920 138.245 ;
        RECT 106.630 138.060 110.920 138.200 ;
        RECT 106.630 138.000 106.950 138.060 ;
        RECT 110.630 138.015 110.920 138.060 ;
        RECT 128.710 138.200 129.030 138.260 ;
        RECT 128.710 138.060 130.320 138.200 ;
        RECT 128.710 138.000 129.030 138.060 ;
        RECT 105.710 137.860 106.030 137.920 ;
        RECT 100.280 137.720 106.030 137.860 ;
        RECT 105.710 137.660 106.030 137.720 ;
        RECT 109.390 137.660 109.710 137.920 ;
        RECT 117.670 137.860 117.990 137.920 ;
        RECT 120.430 137.860 120.750 137.920 ;
        RECT 123.665 137.860 123.955 137.905 ;
        RECT 117.670 137.720 123.955 137.860 ;
        RECT 117.670 137.660 117.990 137.720 ;
        RECT 120.430 137.660 120.750 137.720 ;
        RECT 123.665 137.675 123.955 137.720 ;
        RECT 129.170 137.860 129.490 137.920 ;
        RECT 129.645 137.860 129.935 137.905 ;
        RECT 129.170 137.720 129.935 137.860 ;
        RECT 130.180 137.860 130.320 138.060 ;
        RECT 130.550 138.000 130.870 138.260 ;
        RECT 131.025 138.200 131.315 138.245 ;
        RECT 132.850 138.200 133.170 138.260 ;
        RECT 134.690 138.245 135.010 138.260 ;
        RECT 134.660 138.200 135.010 138.245 ;
        RECT 131.025 138.060 133.170 138.200 ;
        RECT 134.495 138.060 135.010 138.200 ;
        RECT 131.025 138.015 131.315 138.060 ;
        RECT 132.850 138.000 133.170 138.060 ;
        RECT 134.660 138.015 135.010 138.060 ;
        RECT 134.690 138.000 135.010 138.015 ;
        RECT 131.485 137.860 131.775 137.905 ;
        RECT 130.180 137.720 131.775 137.860 ;
        RECT 129.170 137.660 129.490 137.720 ;
        RECT 129.645 137.675 129.935 137.720 ;
        RECT 131.485 137.675 131.775 137.720 ;
        RECT 133.325 137.860 133.615 137.905 ;
        RECT 133.770 137.860 134.090 137.920 ;
        RECT 133.325 137.720 134.090 137.860 ;
        RECT 140.300 137.860 140.440 138.340 ;
        RECT 140.685 137.860 140.975 137.905 ;
        RECT 140.300 137.720 140.975 137.860 ;
        RECT 141.680 137.860 141.820 138.355 ;
        RECT 144.810 138.340 145.130 138.600 ;
        RECT 142.065 137.860 142.355 137.905 ;
        RECT 141.680 137.720 142.355 137.860 ;
        RECT 133.325 137.675 133.615 137.720 ;
        RECT 133.770 137.660 134.090 137.720 ;
        RECT 140.685 137.675 140.975 137.720 ;
        RECT 142.065 137.675 142.355 137.720 ;
        RECT 143.905 137.675 144.195 137.905 ;
        RECT 81.790 137.520 82.110 137.580 ;
        RECT 79.580 137.380 82.110 137.520 ;
        RECT 81.790 137.320 82.110 137.380 ;
        RECT 82.250 137.320 82.570 137.580 ;
        RECT 87.770 137.520 88.090 137.580 ;
        RECT 102.045 137.520 102.335 137.565 ;
        RECT 87.770 137.380 102.335 137.520 ;
        RECT 87.770 137.320 88.090 137.380 ;
        RECT 102.045 137.335 102.335 137.380 ;
        RECT 102.925 137.520 103.215 137.565 ;
        RECT 104.115 137.520 104.405 137.565 ;
        RECT 106.635 137.520 106.925 137.565 ;
        RECT 102.925 137.380 106.925 137.520 ;
        RECT 102.925 137.335 103.215 137.380 ;
        RECT 104.115 137.335 104.405 137.380 ;
        RECT 106.635 137.335 106.925 137.380 ;
        RECT 110.285 137.520 110.575 137.565 ;
        RECT 111.475 137.520 111.765 137.565 ;
        RECT 113.995 137.520 114.285 137.565 ;
        RECT 110.285 137.380 114.285 137.520 ;
        RECT 110.285 137.335 110.575 137.380 ;
        RECT 111.475 137.335 111.765 137.380 ;
        RECT 113.995 137.335 114.285 137.380 ;
        RECT 134.205 137.520 134.495 137.565 ;
        RECT 135.395 137.520 135.685 137.565 ;
        RECT 137.915 137.520 138.205 137.565 ;
        RECT 134.205 137.380 138.205 137.520 ;
        RECT 134.205 137.335 134.495 137.380 ;
        RECT 135.395 137.335 135.685 137.380 ;
        RECT 137.915 137.335 138.205 137.380 ;
        RECT 41.770 137.180 42.090 137.240 ;
        RECT 42.690 137.180 43.010 137.240 ;
        RECT 40.020 137.040 43.010 137.180 ;
        RECT 32.110 136.995 32.400 137.040 ;
        RECT 33.680 136.995 33.970 137.040 ;
        RECT 35.780 136.995 36.070 137.040 ;
        RECT 41.770 136.980 42.090 137.040 ;
        RECT 42.690 136.980 43.010 137.040 ;
        RECT 58.330 137.180 58.620 137.225 ;
        RECT 59.900 137.180 60.190 137.225 ;
        RECT 62.000 137.180 62.290 137.225 ;
        RECT 58.330 137.040 62.290 137.180 ;
        RECT 58.330 136.995 58.620 137.040 ;
        RECT 59.900 136.995 60.190 137.040 ;
        RECT 62.000 136.995 62.290 137.040 ;
        RECT 70.790 137.180 71.080 137.225 ;
        RECT 72.890 137.180 73.180 137.225 ;
        RECT 74.460 137.180 74.750 137.225 ;
        RECT 70.790 137.040 74.750 137.180 ;
        RECT 70.790 136.995 71.080 137.040 ;
        RECT 72.890 136.995 73.180 137.040 ;
        RECT 74.460 136.995 74.750 137.040 ;
        RECT 79.490 137.180 79.810 137.240 ;
        RECT 102.530 137.180 102.820 137.225 ;
        RECT 104.630 137.180 104.920 137.225 ;
        RECT 106.200 137.180 106.490 137.225 ;
        RECT 79.490 137.040 86.620 137.180 ;
        RECT 79.490 136.980 79.810 137.040 ;
        RECT 86.480 136.900 86.620 137.040 ;
        RECT 102.530 137.040 106.490 137.180 ;
        RECT 102.530 136.995 102.820 137.040 ;
        RECT 104.630 136.995 104.920 137.040 ;
        RECT 106.200 136.995 106.490 137.040 ;
        RECT 109.890 137.180 110.180 137.225 ;
        RECT 111.990 137.180 112.280 137.225 ;
        RECT 113.560 137.180 113.850 137.225 ;
        RECT 133.810 137.180 134.100 137.225 ;
        RECT 135.910 137.180 136.200 137.225 ;
        RECT 137.480 137.180 137.770 137.225 ;
        RECT 143.980 137.180 144.120 137.675 ;
        RECT 109.890 137.040 113.850 137.180 ;
        RECT 109.890 136.995 110.180 137.040 ;
        RECT 111.990 136.995 112.280 137.040 ;
        RECT 113.560 136.995 113.850 137.040 ;
        RECT 116.380 137.040 133.080 137.180 ;
        RECT 116.380 136.900 116.520 137.040 ;
        RECT 19.230 136.640 19.550 136.900 ;
        RECT 36.710 136.840 37.030 136.900 ;
        RECT 38.105 136.840 38.395 136.885 ;
        RECT 36.710 136.700 38.395 136.840 ;
        RECT 36.710 136.640 37.030 136.700 ;
        RECT 38.105 136.655 38.395 136.700 ;
        RECT 39.470 136.840 39.790 136.900 ;
        RECT 40.405 136.840 40.695 136.885 ;
        RECT 39.470 136.700 40.695 136.840 ;
        RECT 39.470 136.640 39.790 136.700 ;
        RECT 40.405 136.655 40.695 136.700 ;
        RECT 42.230 136.840 42.550 136.900 ;
        RECT 45.910 136.840 46.230 136.900 ;
        RECT 49.130 136.840 49.450 136.900 ;
        RECT 42.230 136.700 49.450 136.840 ;
        RECT 42.230 136.640 42.550 136.700 ;
        RECT 45.910 136.640 46.230 136.700 ;
        RECT 49.130 136.640 49.450 136.700 ;
        RECT 53.270 136.640 53.590 136.900 ;
        RECT 54.190 136.640 54.510 136.900 ;
        RECT 62.930 136.640 63.250 136.900 ;
        RECT 85.470 136.640 85.790 136.900 ;
        RECT 86.390 136.640 86.710 136.900 ;
        RECT 87.310 136.840 87.630 136.900 ;
        RECT 87.785 136.840 88.075 136.885 ;
        RECT 87.310 136.700 88.075 136.840 ;
        RECT 87.310 136.640 87.630 136.700 ;
        RECT 87.785 136.655 88.075 136.700 ;
        RECT 116.290 136.640 116.610 136.900 ;
        RECT 117.670 136.840 117.990 136.900 ;
        RECT 120.905 136.840 121.195 136.885 ;
        RECT 117.670 136.700 121.195 136.840 ;
        RECT 117.670 136.640 117.990 136.700 ;
        RECT 120.905 136.655 121.195 136.700 ;
        RECT 132.390 136.640 132.710 136.900 ;
        RECT 132.940 136.840 133.080 137.040 ;
        RECT 133.810 137.040 137.770 137.180 ;
        RECT 133.810 136.995 134.100 137.040 ;
        RECT 135.910 136.995 136.200 137.040 ;
        RECT 137.480 136.995 137.770 137.040 ;
        RECT 138.000 137.040 144.120 137.180 ;
        RECT 138.000 136.840 138.140 137.040 ;
        RECT 132.940 136.700 138.140 136.840 ;
        RECT 142.970 136.640 143.290 136.900 ;
        RECT 17.320 136.020 147.040 136.500 ;
        RECT 36.265 135.635 36.555 135.865 ;
        RECT 36.340 135.480 36.480 135.635 ;
        RECT 39.470 135.620 39.790 135.880 ;
        RECT 44.070 135.820 44.390 135.880 ;
        RECT 40.940 135.680 44.390 135.820 ;
        RECT 40.940 135.480 41.080 135.680 ;
        RECT 44.070 135.620 44.390 135.680 ;
        RECT 46.830 135.820 47.150 135.880 ;
        RECT 47.765 135.820 48.055 135.865 ;
        RECT 46.830 135.680 48.055 135.820 ;
        RECT 46.830 135.620 47.150 135.680 ;
        RECT 47.765 135.635 48.055 135.680 ;
        RECT 36.340 135.340 41.080 135.480 ;
        RECT 41.350 135.480 41.640 135.525 ;
        RECT 43.450 135.480 43.740 135.525 ;
        RECT 45.020 135.480 45.310 135.525 ;
        RECT 41.350 135.340 45.310 135.480 ;
        RECT 41.350 135.295 41.640 135.340 ;
        RECT 43.450 135.295 43.740 135.340 ;
        RECT 45.020 135.295 45.310 135.340 ;
        RECT 35.790 135.140 36.110 135.200 ;
        RECT 40.865 135.140 41.155 135.185 ;
        RECT 35.790 135.000 41.155 135.140 ;
        RECT 35.790 134.940 36.110 135.000 ;
        RECT 40.865 134.955 41.155 135.000 ;
        RECT 41.745 135.140 42.035 135.185 ;
        RECT 42.935 135.140 43.225 135.185 ;
        RECT 45.455 135.140 45.745 135.185 ;
        RECT 41.745 135.000 45.745 135.140 ;
        RECT 41.745 134.955 42.035 135.000 ;
        RECT 42.935 134.955 43.225 135.000 ;
        RECT 45.455 134.955 45.745 135.000 ;
        RECT 20.165 134.800 20.455 134.845 ;
        RECT 20.610 134.800 20.930 134.860 ;
        RECT 37.645 134.800 37.935 134.845 ;
        RECT 47.290 134.800 47.610 134.860 ;
        RECT 20.165 134.660 20.930 134.800 ;
        RECT 20.165 134.615 20.455 134.660 ;
        RECT 20.610 134.600 20.930 134.660 ;
        RECT 35.420 134.660 37.415 134.800 ;
        RECT 34.870 134.460 35.190 134.520 ;
        RECT 35.420 134.505 35.560 134.660 ;
        RECT 36.250 134.505 36.570 134.520 ;
        RECT 35.345 134.460 35.635 134.505 ;
        RECT 34.870 134.320 35.635 134.460 ;
        RECT 34.870 134.260 35.190 134.320 ;
        RECT 35.345 134.275 35.635 134.320 ;
        RECT 36.250 134.275 36.635 134.505 ;
        RECT 37.275 134.460 37.415 134.660 ;
        RECT 37.645 134.660 47.610 134.800 ;
        RECT 37.645 134.615 37.935 134.660 ;
        RECT 47.290 134.600 47.610 134.660 ;
        RECT 39.485 134.460 39.775 134.505 ;
        RECT 42.090 134.460 42.380 134.505 ;
        RECT 37.275 134.320 39.775 134.460 ;
        RECT 39.485 134.275 39.775 134.320 ;
        RECT 40.480 134.320 42.380 134.460 ;
        RECT 47.840 134.460 47.980 135.635 ;
        RECT 49.130 135.620 49.450 135.880 ;
        RECT 53.270 135.620 53.590 135.880 ;
        RECT 54.650 135.620 54.970 135.880 ;
        RECT 62.930 135.820 63.250 135.880 ;
        RECT 56.580 135.680 63.250 135.820 ;
        RECT 48.210 135.480 48.530 135.540 ;
        RECT 50.050 135.480 50.370 135.540 ;
        RECT 56.580 135.480 56.720 135.680 ;
        RECT 62.930 135.620 63.250 135.680 ;
        RECT 63.390 135.620 63.710 135.880 ;
        RECT 75.350 135.820 75.670 135.880 ;
        RECT 79.950 135.820 80.270 135.880 ;
        RECT 75.350 135.680 80.270 135.820 ;
        RECT 75.350 135.620 75.670 135.680 ;
        RECT 79.950 135.620 80.270 135.680 ;
        RECT 80.425 135.820 80.715 135.865 ;
        RECT 82.250 135.820 82.570 135.880 ;
        RECT 80.425 135.680 82.570 135.820 ;
        RECT 80.425 135.635 80.715 135.680 ;
        RECT 82.250 135.620 82.570 135.680 ;
        RECT 96.970 135.620 97.290 135.880 ;
        RECT 102.490 135.820 102.810 135.880 ;
        RECT 103.425 135.820 103.715 135.865 ;
        RECT 102.490 135.680 103.715 135.820 ;
        RECT 102.490 135.620 102.810 135.680 ;
        RECT 103.425 135.635 103.715 135.680 ;
        RECT 106.170 135.820 106.490 135.880 ;
        RECT 108.025 135.820 108.315 135.865 ;
        RECT 106.170 135.680 108.315 135.820 ;
        RECT 106.170 135.620 106.490 135.680 ;
        RECT 108.025 135.635 108.315 135.680 ;
        RECT 118.605 135.820 118.895 135.865 ;
        RECT 124.570 135.820 124.890 135.880 ;
        RECT 118.605 135.680 124.890 135.820 ;
        RECT 118.605 135.635 118.895 135.680 ;
        RECT 124.570 135.620 124.890 135.680 ;
        RECT 48.210 135.340 50.370 135.480 ;
        RECT 48.210 135.280 48.530 135.340 ;
        RECT 50.050 135.280 50.370 135.340 ;
        RECT 54.740 135.340 56.720 135.480 ;
        RECT 56.990 135.480 57.280 135.525 ;
        RECT 59.090 135.480 59.380 135.525 ;
        RECT 60.660 135.480 60.950 135.525 ;
        RECT 56.990 135.340 60.950 135.480 ;
        RECT 50.140 134.800 50.280 135.280 ;
        RECT 51.445 134.800 51.735 134.845 ;
        RECT 50.140 134.660 51.735 134.800 ;
        RECT 51.445 134.615 51.735 134.660 ;
        RECT 52.365 134.800 52.655 134.845 ;
        RECT 52.810 134.800 53.130 134.860 ;
        RECT 52.365 134.660 53.130 134.800 ;
        RECT 52.365 134.615 52.655 134.660 ;
        RECT 52.810 134.600 53.130 134.660 ;
        RECT 48.225 134.460 48.515 134.505 ;
        RECT 47.840 134.320 48.515 134.460 ;
        RECT 36.250 134.260 36.570 134.275 ;
        RECT 16.010 134.120 16.330 134.180 ;
        RECT 19.245 134.120 19.535 134.165 ;
        RECT 16.010 133.980 19.535 134.120 ;
        RECT 16.010 133.920 16.330 133.980 ;
        RECT 19.245 133.935 19.535 133.980 ;
        RECT 37.185 134.120 37.475 134.165 ;
        RECT 38.090 134.120 38.410 134.180 ;
        RECT 40.480 134.165 40.620 134.320 ;
        RECT 42.090 134.275 42.380 134.320 ;
        RECT 48.225 134.275 48.515 134.320 ;
        RECT 53.730 134.260 54.050 134.520 ;
        RECT 54.740 134.505 54.880 135.340 ;
        RECT 56.990 135.295 57.280 135.340 ;
        RECT 59.090 135.295 59.380 135.340 ;
        RECT 60.660 135.295 60.950 135.340 ;
        RECT 72.630 135.480 72.920 135.525 ;
        RECT 74.730 135.480 75.020 135.525 ;
        RECT 76.300 135.480 76.590 135.525 ;
        RECT 72.630 135.340 76.590 135.480 ;
        RECT 72.630 135.295 72.920 135.340 ;
        RECT 74.730 135.295 75.020 135.340 ;
        RECT 76.300 135.295 76.590 135.340 ;
        RECT 78.570 135.480 78.890 135.540 ;
        RECT 79.045 135.480 79.335 135.525 ;
        RECT 88.730 135.480 89.020 135.525 ;
        RECT 90.830 135.480 91.120 135.525 ;
        RECT 92.400 135.480 92.690 135.525 ;
        RECT 78.570 135.340 85.240 135.480 ;
        RECT 78.570 135.280 78.890 135.340 ;
        RECT 79.045 135.295 79.335 135.340 ;
        RECT 85.100 135.185 85.240 135.340 ;
        RECT 88.730 135.340 92.690 135.480 ;
        RECT 88.730 135.295 89.020 135.340 ;
        RECT 90.830 135.295 91.120 135.340 ;
        RECT 92.400 135.295 92.690 135.340 ;
        RECT 99.730 135.280 100.050 135.540 ;
        RECT 121.350 135.480 121.640 135.525 ;
        RECT 122.920 135.480 123.210 135.525 ;
        RECT 125.020 135.480 125.310 135.525 ;
        RECT 121.350 135.340 125.310 135.480 ;
        RECT 121.350 135.295 121.640 135.340 ;
        RECT 122.920 135.295 123.210 135.340 ;
        RECT 125.020 135.295 125.310 135.340 ;
        RECT 134.270 135.480 134.560 135.525 ;
        RECT 136.370 135.480 136.660 135.525 ;
        RECT 137.940 135.480 138.230 135.525 ;
        RECT 134.270 135.340 138.230 135.480 ;
        RECT 134.270 135.295 134.560 135.340 ;
        RECT 136.370 135.295 136.660 135.340 ;
        RECT 137.940 135.295 138.230 135.340 ;
        RECT 140.685 135.295 140.975 135.525 ;
        RECT 57.385 135.140 57.675 135.185 ;
        RECT 58.575 135.140 58.865 135.185 ;
        RECT 61.095 135.140 61.385 135.185 ;
        RECT 57.385 135.000 61.385 135.140 ;
        RECT 57.385 134.955 57.675 135.000 ;
        RECT 58.575 134.955 58.865 135.000 ;
        RECT 61.095 134.955 61.385 135.000 ;
        RECT 73.025 135.140 73.315 135.185 ;
        RECT 74.215 135.140 74.505 135.185 ;
        RECT 76.735 135.140 77.025 135.185 ;
        RECT 73.025 135.000 77.025 135.140 ;
        RECT 73.025 134.955 73.315 135.000 ;
        RECT 74.215 134.955 74.505 135.000 ;
        RECT 76.735 134.955 77.025 135.000 ;
        RECT 80.885 135.140 81.175 135.185 ;
        RECT 82.265 135.140 82.555 135.185 ;
        RECT 80.885 135.000 82.555 135.140 ;
        RECT 80.885 134.955 81.175 135.000 ;
        RECT 82.265 134.955 82.555 135.000 ;
        RECT 85.025 134.955 85.315 135.185 ;
        RECT 87.770 135.140 88.090 135.200 ;
        RECT 88.245 135.140 88.535 135.185 ;
        RECT 87.770 135.000 88.535 135.140 ;
        RECT 87.770 134.940 88.090 135.000 ;
        RECT 88.245 134.955 88.535 135.000 ;
        RECT 89.125 135.140 89.415 135.185 ;
        RECT 90.315 135.140 90.605 135.185 ;
        RECT 92.835 135.140 93.125 135.185 ;
        RECT 99.820 135.140 99.960 135.280 ;
        RECT 89.125 135.000 93.125 135.140 ;
        RECT 89.125 134.955 89.415 135.000 ;
        RECT 90.315 134.955 90.605 135.000 ;
        RECT 92.835 134.955 93.125 135.000 ;
        RECT 97.980 135.000 99.960 135.140 ;
        RECT 56.505 134.800 56.795 134.845 ;
        RECT 62.470 134.800 62.790 134.860 ;
        RECT 56.505 134.660 62.790 134.800 ;
        RECT 56.505 134.615 56.795 134.660 ;
        RECT 62.470 134.600 62.790 134.660 ;
        RECT 72.130 134.600 72.450 134.860 ;
        RECT 79.490 134.600 79.810 134.860 ;
        RECT 85.470 134.800 85.790 134.860 ;
        RECT 85.945 134.800 86.235 134.845 ;
        RECT 85.470 134.660 86.235 134.800 ;
        RECT 85.470 134.600 85.790 134.660 ;
        RECT 85.945 134.615 86.235 134.660 ;
        RECT 86.865 134.800 87.155 134.845 ;
        RECT 87.310 134.800 87.630 134.860 ;
        RECT 97.980 134.845 98.120 135.000 ;
        RECT 105.710 134.940 106.030 135.200 ;
        RECT 106.645 135.140 106.935 135.185 ;
        RECT 111.245 135.140 111.535 135.185 ;
        RECT 114.910 135.140 115.230 135.200 ;
        RECT 106.645 135.000 115.230 135.140 ;
        RECT 106.645 134.955 106.935 135.000 ;
        RECT 111.245 134.955 111.535 135.000 ;
        RECT 114.910 134.940 115.230 135.000 ;
        RECT 120.915 135.140 121.205 135.185 ;
        RECT 123.435 135.140 123.725 135.185 ;
        RECT 124.625 135.140 124.915 135.185 ;
        RECT 120.915 135.000 124.915 135.140 ;
        RECT 120.915 134.955 121.205 135.000 ;
        RECT 123.435 134.955 123.725 135.000 ;
        RECT 124.625 134.955 124.915 135.000 ;
        RECT 125.505 135.140 125.795 135.185 ;
        RECT 134.665 135.140 134.955 135.185 ;
        RECT 135.855 135.140 136.145 135.185 ;
        RECT 138.375 135.140 138.665 135.185 ;
        RECT 125.505 135.000 134.000 135.140 ;
        RECT 125.505 134.955 125.795 135.000 ;
        RECT 86.865 134.660 87.630 134.800 ;
        RECT 86.865 134.615 87.155 134.660 ;
        RECT 87.310 134.600 87.630 134.660 ;
        RECT 97.905 134.615 98.195 134.845 ;
        RECT 98.365 134.615 98.655 134.845 ;
        RECT 98.810 134.800 99.130 134.860 ;
        RECT 99.285 134.800 99.575 134.845 ;
        RECT 98.810 134.660 99.575 134.800 ;
        RECT 89.610 134.505 89.930 134.520 ;
        RECT 54.740 134.320 55.035 134.505 ;
        RECT 57.730 134.460 58.020 134.505 ;
        RECT 54.745 134.275 55.035 134.320 ;
        RECT 55.660 134.320 58.020 134.460 ;
        RECT 37.185 133.980 38.410 134.120 ;
        RECT 37.185 133.935 37.475 133.980 ;
        RECT 38.090 133.920 38.410 133.980 ;
        RECT 40.405 133.935 40.695 134.165 ;
        RECT 44.530 134.120 44.850 134.180 ;
        RECT 55.660 134.165 55.800 134.320 ;
        RECT 57.730 134.275 58.020 134.320 ;
        RECT 73.480 134.460 73.770 134.505 ;
        RECT 86.405 134.460 86.695 134.505 ;
        RECT 73.480 134.320 86.695 134.460 ;
        RECT 73.480 134.275 73.770 134.320 ;
        RECT 86.405 134.275 86.695 134.320 ;
        RECT 89.580 134.275 89.930 134.505 ;
        RECT 98.440 134.460 98.580 134.615 ;
        RECT 98.810 134.600 99.130 134.660 ;
        RECT 99.285 134.615 99.575 134.660 ;
        RECT 99.730 134.600 100.050 134.860 ;
        RECT 101.570 134.800 101.890 134.860 ;
        RECT 105.265 134.800 105.555 134.845 ;
        RECT 121.810 134.800 122.130 134.860 ;
        RECT 101.570 134.660 122.130 134.800 ;
        RECT 101.570 134.600 101.890 134.660 ;
        RECT 105.265 134.615 105.555 134.660 ;
        RECT 121.810 134.600 122.130 134.660 ;
        RECT 125.030 134.800 125.350 134.860 ;
        RECT 133.860 134.845 134.000 135.000 ;
        RECT 134.665 135.000 138.665 135.140 ;
        RECT 140.760 135.140 140.900 135.295 ;
        RECT 142.050 135.140 142.370 135.200 ;
        RECT 143.905 135.140 144.195 135.185 ;
        RECT 140.760 135.000 144.195 135.140 ;
        RECT 134.665 134.955 134.955 135.000 ;
        RECT 135.855 134.955 136.145 135.000 ;
        RECT 138.375 134.955 138.665 135.000 ;
        RECT 142.050 134.940 142.370 135.000 ;
        RECT 143.905 134.955 144.195 135.000 ;
        RECT 125.965 134.800 126.255 134.845 ;
        RECT 125.030 134.660 126.255 134.800 ;
        RECT 125.030 134.600 125.350 134.660 ;
        RECT 125.965 134.615 126.255 134.660 ;
        RECT 133.785 134.800 134.075 134.845 ;
        RECT 133.785 134.660 136.300 134.800 ;
        RECT 133.785 134.615 134.075 134.660 ;
        RECT 136.160 134.520 136.300 134.660 ;
        RECT 110.325 134.460 110.615 134.505 ;
        RECT 116.290 134.460 116.610 134.520 ;
        RECT 98.440 134.320 116.610 134.460 ;
        RECT 110.325 134.275 110.615 134.320 ;
        RECT 89.610 134.260 89.930 134.275 ;
        RECT 116.290 134.260 116.610 134.320 ;
        RECT 124.280 134.460 124.570 134.505 ;
        RECT 128.250 134.460 128.570 134.520 ;
        RECT 124.280 134.320 128.570 134.460 ;
        RECT 124.280 134.275 124.570 134.320 ;
        RECT 128.250 134.260 128.570 134.320 ;
        RECT 134.230 134.460 134.550 134.520 ;
        RECT 135.010 134.460 135.300 134.505 ;
        RECT 134.230 134.320 135.300 134.460 ;
        RECT 134.230 134.260 134.550 134.320 ;
        RECT 135.010 134.275 135.300 134.320 ;
        RECT 136.070 134.260 136.390 134.520 ;
        RECT 49.225 134.120 49.515 134.165 ;
        RECT 44.530 133.980 49.515 134.120 ;
        RECT 44.530 133.920 44.850 133.980 ;
        RECT 49.225 133.935 49.515 133.980 ;
        RECT 55.585 133.935 55.875 134.165 ;
        RECT 95.130 133.920 95.450 134.180 ;
        RECT 109.865 134.120 110.155 134.165 ;
        RECT 113.990 134.120 114.310 134.180 ;
        RECT 122.270 134.120 122.590 134.180 ;
        RECT 109.865 133.980 122.590 134.120 ;
        RECT 109.865 133.935 110.155 133.980 ;
        RECT 113.990 133.920 114.310 133.980 ;
        RECT 122.270 133.920 122.590 133.980 ;
        RECT 129.185 134.120 129.475 134.165 ;
        RECT 130.550 134.120 130.870 134.180 ;
        RECT 129.185 133.980 130.870 134.120 ;
        RECT 129.185 133.935 129.475 133.980 ;
        RECT 130.550 133.920 130.870 133.980 ;
        RECT 141.130 133.920 141.450 134.180 ;
        RECT 17.320 133.300 147.040 133.780 ;
        RECT 42.230 133.100 42.550 133.160 ;
        RECT 42.705 133.100 42.995 133.145 ;
        RECT 42.230 132.960 42.995 133.100 ;
        RECT 42.230 132.900 42.550 132.960 ;
        RECT 42.705 132.915 42.995 132.960 ;
        RECT 22.910 132.760 23.230 132.820 ;
        RECT 28.445 132.760 28.735 132.805 ;
        RECT 22.910 132.620 28.735 132.760 ;
        RECT 22.910 132.560 23.230 132.620 ;
        RECT 28.445 132.575 28.735 132.620 ;
        RECT 37.140 132.760 37.430 132.805 ;
        RECT 38.090 132.760 38.410 132.820 ;
        RECT 37.140 132.620 38.410 132.760 ;
        RECT 37.140 132.575 37.430 132.620 ;
        RECT 38.090 132.560 38.410 132.620 ;
        RECT 18.770 132.420 19.090 132.480 ;
        RECT 20.525 132.420 20.815 132.465 ;
        RECT 18.770 132.280 20.815 132.420 ;
        RECT 18.770 132.220 19.090 132.280 ;
        RECT 20.525 132.235 20.815 132.280 ;
        RECT 27.525 132.420 27.815 132.465 ;
        RECT 27.970 132.420 28.290 132.480 ;
        RECT 27.525 132.280 28.290 132.420 ;
        RECT 27.525 132.235 27.815 132.280 ;
        RECT 27.970 132.220 28.290 132.280 ;
        RECT 35.790 132.220 36.110 132.480 ;
        RECT 42.780 132.420 42.920 132.915 ;
        RECT 44.070 132.900 44.390 133.160 ;
        RECT 51.445 133.100 51.735 133.145 ;
        RECT 52.810 133.100 53.130 133.160 ;
        RECT 51.445 132.960 53.130 133.100 ;
        RECT 51.445 132.915 51.735 132.960 ;
        RECT 52.810 132.900 53.130 132.960 ;
        RECT 78.110 132.900 78.430 133.160 ;
        RECT 85.485 133.100 85.775 133.145 ;
        RECT 87.405 133.100 87.695 133.145 ;
        RECT 85.485 132.960 87.695 133.100 ;
        RECT 85.485 132.915 85.775 132.960 ;
        RECT 87.405 132.915 87.695 132.960 ;
        RECT 89.165 133.100 89.455 133.145 ;
        RECT 89.610 133.100 89.930 133.160 ;
        RECT 89.165 132.960 89.930 133.100 ;
        RECT 89.165 132.915 89.455 132.960 ;
        RECT 89.610 132.900 89.930 132.960 ;
        RECT 91.005 133.100 91.295 133.145 ;
        RECT 95.130 133.100 95.450 133.160 ;
        RECT 105.250 133.100 105.570 133.160 ;
        RECT 91.005 132.960 105.570 133.100 ;
        RECT 91.005 132.915 91.295 132.960 ;
        RECT 95.130 132.900 95.450 132.960 ;
        RECT 105.250 132.900 105.570 132.960 ;
        RECT 120.430 133.100 120.750 133.160 ;
        RECT 120.905 133.100 121.195 133.145 ;
        RECT 120.430 132.960 121.195 133.100 ;
        RECT 120.430 132.900 120.750 132.960 ;
        RECT 120.905 132.915 121.195 132.960 ;
        RECT 128.250 132.900 128.570 133.160 ;
        RECT 133.785 133.100 134.075 133.145 ;
        RECT 134.230 133.100 134.550 133.160 ;
        RECT 133.785 132.960 134.550 133.100 ;
        RECT 133.785 132.915 134.075 132.960 ;
        RECT 134.230 132.900 134.550 132.960 ;
        RECT 135.625 133.100 135.915 133.145 ;
        RECT 141.130 133.100 141.450 133.160 ;
        RECT 135.625 132.960 141.450 133.100 ;
        RECT 135.625 132.915 135.915 132.960 ;
        RECT 141.130 132.900 141.450 132.960 ;
        RECT 142.985 132.915 143.275 133.145 ;
        RECT 54.190 132.760 54.510 132.820 ;
        RECT 57.010 132.760 57.300 132.805 ;
        RECT 54.190 132.620 57.300 132.760 ;
        RECT 54.190 132.560 54.510 132.620 ;
        RECT 57.010 132.575 57.300 132.620 ;
        RECT 77.190 132.560 77.510 132.820 ;
        RECT 85.930 132.760 86.250 132.820 ;
        RECT 86.405 132.760 86.695 132.805 ;
        RECT 78.660 132.620 86.695 132.760 ;
        RECT 43.625 132.420 43.915 132.465 ;
        RECT 42.780 132.280 43.915 132.420 ;
        RECT 43.625 132.235 43.915 132.280 ;
        RECT 44.530 132.220 44.850 132.480 ;
        RECT 58.345 132.420 58.635 132.465 ;
        RECT 65.705 132.420 65.995 132.465 ;
        RECT 58.345 132.280 65.995 132.420 ;
        RECT 58.345 132.235 58.635 132.280 ;
        RECT 65.705 132.235 65.995 132.280 ;
        RECT 66.610 132.420 66.930 132.480 ;
        RECT 78.660 132.465 78.800 132.620 ;
        RECT 85.930 132.560 86.250 132.620 ;
        RECT 86.405 132.575 86.695 132.620 ;
        RECT 104.330 132.760 104.650 132.820 ;
        RECT 110.785 132.760 111.075 132.805 ;
        RECT 136.070 132.760 136.390 132.820 ;
        RECT 104.330 132.620 111.075 132.760 ;
        RECT 104.330 132.560 104.650 132.620 ;
        RECT 110.785 132.575 111.075 132.620 ;
        RECT 127.880 132.620 136.390 132.760 ;
        RECT 69.385 132.420 69.675 132.465 ;
        RECT 66.610 132.280 69.675 132.420 ;
        RECT 19.230 131.880 19.550 132.140 ;
        RECT 20.125 132.080 20.415 132.125 ;
        RECT 21.315 132.080 21.605 132.125 ;
        RECT 23.835 132.080 24.125 132.125 ;
        RECT 20.125 131.940 24.125 132.080 ;
        RECT 20.125 131.895 20.415 131.940 ;
        RECT 21.315 131.895 21.605 131.940 ;
        RECT 23.835 131.895 24.125 131.940 ;
        RECT 36.685 132.080 36.975 132.125 ;
        RECT 37.875 132.080 38.165 132.125 ;
        RECT 40.395 132.080 40.685 132.125 ;
        RECT 36.685 131.940 40.685 132.080 ;
        RECT 36.685 131.895 36.975 131.940 ;
        RECT 37.875 131.895 38.165 131.940 ;
        RECT 40.395 131.895 40.685 131.940 ;
        RECT 41.770 132.080 42.090 132.140 ;
        RECT 44.620 132.080 44.760 132.220 ;
        RECT 41.770 131.940 44.760 132.080 ;
        RECT 53.755 132.080 54.045 132.125 ;
        RECT 56.275 132.080 56.565 132.125 ;
        RECT 57.465 132.080 57.755 132.125 ;
        RECT 53.755 131.940 57.755 132.080 ;
        RECT 65.780 132.080 65.920 132.235 ;
        RECT 66.610 132.220 66.930 132.280 ;
        RECT 69.385 132.235 69.675 132.280 ;
        RECT 78.125 132.235 78.415 132.465 ;
        RECT 78.585 132.235 78.875 132.465 ;
        RECT 82.710 132.420 83.030 132.480 ;
        RECT 85.025 132.420 85.315 132.465 ;
        RECT 85.470 132.420 85.790 132.480 ;
        RECT 87.310 132.420 87.630 132.480 ;
        RECT 82.710 132.280 87.630 132.420 ;
        RECT 69.830 132.080 70.150 132.140 ;
        RECT 73.065 132.080 73.355 132.125 ;
        RECT 65.780 131.940 73.355 132.080 ;
        RECT 41.770 131.880 42.090 131.940 ;
        RECT 53.755 131.895 54.045 131.940 ;
        RECT 56.275 131.895 56.565 131.940 ;
        RECT 57.465 131.895 57.755 131.940 ;
        RECT 69.830 131.880 70.150 131.940 ;
        RECT 73.065 131.895 73.355 131.940 ;
        RECT 76.270 132.080 76.590 132.140 ;
        RECT 78.200 132.080 78.340 132.235 ;
        RECT 82.710 132.220 83.030 132.280 ;
        RECT 85.025 132.235 85.315 132.280 ;
        RECT 85.470 132.220 85.790 132.280 ;
        RECT 87.310 132.220 87.630 132.280 ;
        RECT 108.945 132.420 109.235 132.465 ;
        RECT 109.390 132.420 109.710 132.480 ;
        RECT 108.945 132.280 109.710 132.420 ;
        RECT 108.945 132.235 109.235 132.280 ;
        RECT 109.390 132.220 109.710 132.280 ;
        RECT 112.625 132.420 112.915 132.465 ;
        RECT 113.530 132.420 113.850 132.480 ;
        RECT 112.625 132.280 113.850 132.420 ;
        RECT 112.625 132.235 112.915 132.280 ;
        RECT 113.530 132.220 113.850 132.280 ;
        RECT 117.670 132.220 117.990 132.480 ;
        RECT 127.880 132.465 128.020 132.620 ;
        RECT 136.070 132.560 136.390 132.620 ;
        RECT 139.290 132.760 139.610 132.820 ;
        RECT 139.765 132.760 140.055 132.805 ;
        RECT 139.290 132.620 140.055 132.760 ;
        RECT 139.290 132.560 139.610 132.620 ;
        RECT 139.765 132.575 140.055 132.620 ;
        RECT 119.065 132.235 119.355 132.465 ;
        RECT 119.985 132.420 120.275 132.465 ;
        RECT 126.470 132.420 126.760 132.465 ;
        RECT 119.985 132.280 126.760 132.420 ;
        RECT 119.985 132.235 120.275 132.280 ;
        RECT 126.470 132.235 126.760 132.280 ;
        RECT 127.805 132.235 128.095 132.465 ;
        RECT 76.270 131.940 78.340 132.080 ;
        RECT 81.790 132.080 82.110 132.140 ;
        RECT 86.390 132.080 86.710 132.140 ;
        RECT 90.070 132.080 90.390 132.140 ;
        RECT 91.465 132.080 91.755 132.125 ;
        RECT 81.790 131.940 91.755 132.080 ;
        RECT 76.270 131.880 76.590 131.940 ;
        RECT 81.790 131.880 82.110 131.940 ;
        RECT 86.390 131.880 86.710 131.940 ;
        RECT 90.070 131.880 90.390 131.940 ;
        RECT 91.465 131.895 91.755 131.940 ;
        RECT 91.925 131.895 92.215 132.125 ;
        RECT 19.730 131.740 20.020 131.785 ;
        RECT 21.830 131.740 22.120 131.785 ;
        RECT 23.400 131.740 23.690 131.785 ;
        RECT 19.730 131.600 23.690 131.740 ;
        RECT 19.730 131.555 20.020 131.600 ;
        RECT 21.830 131.555 22.120 131.600 ;
        RECT 23.400 131.555 23.690 131.600 ;
        RECT 36.290 131.740 36.580 131.785 ;
        RECT 38.390 131.740 38.680 131.785 ;
        RECT 39.960 131.740 40.250 131.785 ;
        RECT 36.290 131.600 40.250 131.740 ;
        RECT 36.290 131.555 36.580 131.600 ;
        RECT 38.390 131.555 38.680 131.600 ;
        RECT 39.960 131.555 40.250 131.600 ;
        RECT 54.190 131.740 54.480 131.785 ;
        RECT 55.760 131.740 56.050 131.785 ;
        RECT 57.860 131.740 58.150 131.785 ;
        RECT 54.190 131.600 58.150 131.740 ;
        RECT 54.190 131.555 54.480 131.600 ;
        RECT 55.760 131.555 56.050 131.600 ;
        RECT 57.860 131.555 58.150 131.600 ;
        RECT 88.245 131.740 88.535 131.785 ;
        RECT 92.000 131.740 92.140 131.895 ;
        RECT 102.490 131.880 102.810 132.140 ;
        RECT 110.310 131.880 110.630 132.140 ;
        RECT 119.140 132.080 119.280 132.235 ;
        RECT 129.170 132.220 129.490 132.480 ;
        RECT 130.550 132.220 130.870 132.480 ;
        RECT 135.610 132.420 135.930 132.480 ;
        RECT 135.610 132.280 139.520 132.420 ;
        RECT 135.610 132.220 135.930 132.280 ;
        RECT 122.270 132.080 122.590 132.140 ;
        RECT 119.140 131.940 122.590 132.080 ;
        RECT 122.270 131.880 122.590 131.940 ;
        RECT 123.215 132.080 123.505 132.125 ;
        RECT 125.735 132.080 126.025 132.125 ;
        RECT 126.925 132.080 127.215 132.125 ;
        RECT 123.215 131.940 127.215 132.080 ;
        RECT 123.215 131.895 123.505 131.940 ;
        RECT 125.735 131.895 126.025 131.940 ;
        RECT 126.925 131.895 127.215 131.940 ;
        RECT 132.390 132.080 132.710 132.140 ;
        RECT 136.085 132.080 136.375 132.125 ;
        RECT 132.390 131.940 136.375 132.080 ;
        RECT 132.390 131.880 132.710 131.940 ;
        RECT 136.085 131.895 136.375 131.940 ;
        RECT 136.545 131.895 136.835 132.125 ;
        RECT 139.380 132.080 139.520 132.280 ;
        RECT 142.050 132.220 142.370 132.480 ;
        RECT 143.060 132.420 143.200 132.915 ;
        RECT 143.905 132.420 144.195 132.465 ;
        RECT 143.060 132.280 144.195 132.420 ;
        RECT 143.905 132.235 144.195 132.280 ;
        RECT 140.225 132.080 140.515 132.125 ;
        RECT 139.380 131.940 140.515 132.080 ;
        RECT 140.225 131.895 140.515 131.940 ;
        RECT 88.245 131.600 92.140 131.740 ;
        RECT 103.870 131.740 104.190 131.800 ;
        RECT 109.865 131.740 110.155 131.785 ;
        RECT 118.145 131.740 118.435 131.785 ;
        RECT 118.590 131.740 118.910 131.800 ;
        RECT 103.870 131.600 118.910 131.740 ;
        RECT 88.245 131.555 88.535 131.600 ;
        RECT 103.870 131.540 104.190 131.600 ;
        RECT 109.865 131.555 110.155 131.600 ;
        RECT 118.145 131.555 118.435 131.600 ;
        RECT 118.590 131.540 118.910 131.600 ;
        RECT 123.650 131.740 123.940 131.785 ;
        RECT 125.220 131.740 125.510 131.785 ;
        RECT 127.320 131.740 127.610 131.785 ;
        RECT 130.105 131.740 130.395 131.785 ;
        RECT 123.650 131.600 127.610 131.740 ;
        RECT 123.650 131.555 123.940 131.600 ;
        RECT 125.220 131.555 125.510 131.600 ;
        RECT 127.320 131.555 127.610 131.600 ;
        RECT 127.880 131.600 130.395 131.740 ;
        RECT 20.610 131.400 20.930 131.460 ;
        RECT 26.145 131.400 26.435 131.445 ;
        RECT 20.610 131.260 26.435 131.400 ;
        RECT 20.610 131.200 20.930 131.260 ;
        RECT 26.145 131.215 26.435 131.260 ;
        RECT 29.365 131.400 29.655 131.445 ;
        RECT 31.190 131.400 31.510 131.460 ;
        RECT 29.365 131.260 31.510 131.400 ;
        RECT 29.365 131.215 29.655 131.260 ;
        RECT 31.190 131.200 31.510 131.260 ;
        RECT 87.310 131.200 87.630 131.460 ;
        RECT 105.725 131.400 106.015 131.445 ;
        RECT 107.090 131.400 107.410 131.460 ;
        RECT 105.725 131.260 107.410 131.400 ;
        RECT 105.725 131.215 106.015 131.260 ;
        RECT 107.090 131.200 107.410 131.260 ;
        RECT 108.025 131.400 108.315 131.445 ;
        RECT 108.470 131.400 108.790 131.460 ;
        RECT 108.025 131.260 108.790 131.400 ;
        RECT 118.680 131.400 118.820 131.540 ;
        RECT 127.880 131.400 128.020 131.600 ;
        RECT 130.105 131.555 130.395 131.600 ;
        RECT 135.150 131.740 135.470 131.800 ;
        RECT 136.620 131.740 136.760 131.895 ;
        RECT 135.150 131.600 136.760 131.740 ;
        RECT 140.300 131.740 140.440 131.895 ;
        RECT 140.670 131.880 140.990 132.140 ;
        RECT 144.350 131.740 144.670 131.800 ;
        RECT 140.300 131.600 144.670 131.740 ;
        RECT 135.150 131.540 135.470 131.600 ;
        RECT 144.350 131.540 144.670 131.600 ;
        RECT 144.810 131.540 145.130 131.800 ;
        RECT 118.680 131.260 128.020 131.400 ;
        RECT 132.390 131.400 132.710 131.460 ;
        RECT 137.925 131.400 138.215 131.445 ;
        RECT 132.390 131.260 138.215 131.400 ;
        RECT 108.025 131.215 108.315 131.260 ;
        RECT 108.470 131.200 108.790 131.260 ;
        RECT 132.390 131.200 132.710 131.260 ;
        RECT 137.925 131.215 138.215 131.260 ;
        RECT 17.320 130.580 147.040 131.060 ;
        RECT 18.770 130.180 19.090 130.440 ;
        RECT 22.910 130.180 23.230 130.440 ;
        RECT 27.970 130.380 28.290 130.440 ;
        RECT 31.650 130.380 31.970 130.440 ;
        RECT 24.840 130.240 31.970 130.380 ;
        RECT 22.005 129.700 22.295 129.745 ;
        RECT 24.840 129.700 24.980 130.240 ;
        RECT 27.970 130.180 28.290 130.240 ;
        RECT 31.650 130.180 31.970 130.240 ;
        RECT 72.145 130.380 72.435 130.425 ;
        RECT 72.590 130.380 72.910 130.440 ;
        RECT 72.145 130.240 72.910 130.380 ;
        RECT 72.145 130.195 72.435 130.240 ;
        RECT 72.590 130.180 72.910 130.240 ;
        RECT 73.065 130.380 73.355 130.425 ;
        RECT 76.270 130.380 76.590 130.440 ;
        RECT 82.725 130.380 83.015 130.425 ;
        RECT 73.065 130.240 83.015 130.380 ;
        RECT 73.065 130.195 73.355 130.240 ;
        RECT 76.270 130.180 76.590 130.240 ;
        RECT 82.725 130.195 83.015 130.240 ;
        RECT 25.670 130.040 25.960 130.085 ;
        RECT 27.240 130.040 27.530 130.085 ;
        RECT 29.340 130.040 29.630 130.085 ;
        RECT 25.670 129.900 29.630 130.040 ;
        RECT 25.670 129.855 25.960 129.900 ;
        RECT 27.240 129.855 27.530 129.900 ;
        RECT 29.340 129.855 29.630 129.900 ;
        RECT 32.125 130.040 32.415 130.085 ;
        RECT 32.570 130.040 32.890 130.100 ;
        RECT 73.510 130.040 73.830 130.100 ;
        RECT 32.125 129.900 32.890 130.040 ;
        RECT 32.125 129.855 32.415 129.900 ;
        RECT 32.570 129.840 32.890 129.900 ;
        RECT 69.920 129.900 73.830 130.040 ;
        RECT 22.005 129.560 24.980 129.700 ;
        RECT 25.235 129.700 25.525 129.745 ;
        RECT 27.755 129.700 28.045 129.745 ;
        RECT 28.945 129.700 29.235 129.745 ;
        RECT 25.235 129.560 29.235 129.700 ;
        RECT 22.005 129.515 22.295 129.560 ;
        RECT 25.235 129.515 25.525 129.560 ;
        RECT 27.755 129.515 28.045 129.560 ;
        RECT 28.945 129.515 29.235 129.560 ;
        RECT 31.190 129.700 31.510 129.760 ;
        RECT 31.190 129.560 33.260 129.700 ;
        RECT 31.190 129.500 31.510 129.560 ;
        RECT 20.610 129.160 20.930 129.420 ;
        RECT 24.750 129.360 25.070 129.420 ;
        RECT 29.825 129.360 30.115 129.405 ;
        RECT 24.750 129.220 30.115 129.360 ;
        RECT 24.750 129.160 25.070 129.220 ;
        RECT 29.825 129.175 30.115 129.220 ;
        RECT 30.270 129.360 30.590 129.420 ;
        RECT 33.120 129.405 33.260 129.560 ;
        RECT 69.920 129.405 70.060 129.900 ;
        RECT 73.510 129.840 73.830 129.900 ;
        RECT 70.290 129.500 70.610 129.760 ;
        RECT 71.685 129.700 71.975 129.745 ;
        RECT 73.970 129.700 74.290 129.760 ;
        RECT 71.685 129.560 74.290 129.700 ;
        RECT 82.800 129.700 82.940 130.195 ;
        RECT 85.470 130.180 85.790 130.440 ;
        RECT 103.870 130.380 104.190 130.440 ;
        RECT 106.645 130.380 106.935 130.425 ;
        RECT 87.400 130.240 91.680 130.380 ;
        RECT 84.565 130.040 84.855 130.085 ;
        RECT 87.400 130.040 87.540 130.240 ;
        RECT 84.565 129.900 87.540 130.040 ;
        RECT 87.785 130.040 88.075 130.085 ;
        RECT 87.785 129.900 91.220 130.040 ;
        RECT 84.565 129.855 84.855 129.900 ;
        RECT 87.785 129.855 88.075 129.900 ;
        RECT 86.405 129.700 86.695 129.745 ;
        RECT 87.310 129.700 87.630 129.760 ;
        RECT 91.080 129.745 91.220 129.900 ;
        RECT 82.800 129.560 87.630 129.700 ;
        RECT 71.685 129.515 71.975 129.560 ;
        RECT 73.970 129.500 74.290 129.560 ;
        RECT 86.405 129.515 86.695 129.560 ;
        RECT 87.310 129.500 87.630 129.560 ;
        RECT 91.005 129.515 91.295 129.745 ;
        RECT 91.540 129.700 91.680 130.240 ;
        RECT 103.870 130.240 106.935 130.380 ;
        RECT 103.870 130.180 104.190 130.240 ;
        RECT 106.645 130.195 106.935 130.240 ;
        RECT 110.310 130.180 110.630 130.440 ;
        RECT 119.970 130.380 120.290 130.440 ;
        RECT 127.330 130.380 127.650 130.440 ;
        RECT 128.265 130.380 128.555 130.425 ;
        RECT 119.970 130.240 128.555 130.380 ;
        RECT 119.970 130.180 120.290 130.240 ;
        RECT 127.330 130.180 127.650 130.240 ;
        RECT 128.265 130.195 128.555 130.240 ;
        RECT 129.170 130.380 129.490 130.440 ;
        RECT 133.785 130.380 134.075 130.425 ;
        RECT 129.170 130.240 134.075 130.380 ;
        RECT 129.170 130.180 129.490 130.240 ;
        RECT 133.785 130.195 134.075 130.240 ;
        RECT 135.700 130.240 137.680 130.380 ;
        RECT 98.810 130.040 99.130 130.100 ;
        RECT 103.410 130.040 103.730 130.100 ;
        RECT 98.810 129.900 103.730 130.040 ;
        RECT 98.810 129.840 99.130 129.900 ;
        RECT 103.410 129.840 103.730 129.900 ;
        RECT 114.490 130.040 114.780 130.085 ;
        RECT 116.590 130.040 116.880 130.085 ;
        RECT 118.160 130.040 118.450 130.085 ;
        RECT 114.490 129.900 118.450 130.040 ;
        RECT 114.490 129.855 114.780 129.900 ;
        RECT 116.590 129.855 116.880 129.900 ;
        RECT 118.160 129.855 118.450 129.900 ;
        RECT 120.890 129.840 121.210 130.100 ;
        RECT 121.850 130.040 122.140 130.085 ;
        RECT 123.950 130.040 124.240 130.085 ;
        RECT 125.520 130.040 125.810 130.085 ;
        RECT 121.850 129.900 125.810 130.040 ;
        RECT 121.850 129.855 122.140 129.900 ;
        RECT 123.950 129.855 124.240 129.900 ;
        RECT 125.520 129.855 125.810 129.900 ;
        RECT 132.390 129.840 132.710 130.100 ;
        RECT 132.865 130.040 133.155 130.085 ;
        RECT 135.700 130.040 135.840 130.240 ;
        RECT 132.865 129.900 135.840 130.040 ;
        RECT 132.865 129.855 133.155 129.900 ;
        RECT 136.530 129.840 136.850 130.100 ;
        RECT 95.145 129.700 95.435 129.745 ;
        RECT 91.540 129.560 95.435 129.700 ;
        RECT 95.145 129.515 95.435 129.560 ;
        RECT 100.190 129.700 100.510 129.760 ;
        RECT 100.190 129.560 103.640 129.700 ;
        RECT 100.190 129.500 100.510 129.560 ;
        RECT 31.665 129.360 31.955 129.405 ;
        RECT 30.270 129.220 31.955 129.360 ;
        RECT 30.270 129.160 30.590 129.220 ;
        RECT 31.665 129.175 31.955 129.220 ;
        RECT 32.585 129.175 32.875 129.405 ;
        RECT 33.045 129.175 33.335 129.405 ;
        RECT 69.845 129.175 70.135 129.405 ;
        RECT 74.905 129.360 75.195 129.405 ;
        RECT 77.190 129.360 77.510 129.420 ;
        RECT 74.905 129.220 77.510 129.360 ;
        RECT 74.905 129.175 75.195 129.220 ;
        RECT 21.085 129.020 21.375 129.065 ;
        RECT 24.290 129.020 24.610 129.080 ;
        RECT 21.085 128.880 24.610 129.020 ;
        RECT 21.085 128.835 21.375 128.880 ;
        RECT 24.290 128.820 24.610 128.880 ;
        RECT 28.600 129.020 28.890 129.065 ;
        RECT 30.745 129.020 31.035 129.065 ;
        RECT 28.600 128.880 31.035 129.020 ;
        RECT 28.600 128.835 28.890 128.880 ;
        RECT 30.745 128.835 31.035 128.880 ;
        RECT 31.190 129.020 31.510 129.080 ;
        RECT 32.660 129.020 32.800 129.175 ;
        RECT 77.190 129.160 77.510 129.220 ;
        RECT 82.710 129.160 83.030 129.420 ;
        RECT 83.645 129.360 83.935 129.405 ;
        RECT 85.025 129.360 85.315 129.405 ;
        RECT 85.930 129.360 86.250 129.420 ;
        RECT 83.645 129.220 86.250 129.360 ;
        RECT 83.645 129.175 83.935 129.220 ;
        RECT 85.025 129.175 85.315 129.220 ;
        RECT 85.930 129.160 86.250 129.220 ;
        RECT 90.070 129.160 90.390 129.420 ;
        RECT 93.290 129.360 93.610 129.420 ;
        RECT 103.500 129.405 103.640 129.560 ;
        RECT 107.090 129.500 107.410 129.760 ;
        RECT 112.610 129.700 112.930 129.760 ;
        RECT 113.085 129.700 113.375 129.745 ;
        RECT 112.610 129.560 113.375 129.700 ;
        RECT 112.610 129.500 112.930 129.560 ;
        RECT 113.085 129.515 113.375 129.560 ;
        RECT 114.885 129.700 115.175 129.745 ;
        RECT 116.075 129.700 116.365 129.745 ;
        RECT 118.595 129.700 118.885 129.745 ;
        RECT 114.885 129.560 118.885 129.700 ;
        RECT 114.885 129.515 115.175 129.560 ;
        RECT 116.075 129.515 116.365 129.560 ;
        RECT 118.595 129.515 118.885 129.560 ;
        RECT 122.245 129.700 122.535 129.745 ;
        RECT 123.435 129.700 123.725 129.745 ;
        RECT 125.955 129.700 126.245 129.745 ;
        RECT 122.245 129.560 126.245 129.700 ;
        RECT 122.245 129.515 122.535 129.560 ;
        RECT 123.435 129.515 123.725 129.560 ;
        RECT 125.955 129.515 126.245 129.560 ;
        RECT 130.090 129.700 130.410 129.760 ;
        RECT 130.565 129.700 130.855 129.745 ;
        RECT 136.620 129.700 136.760 129.840 ;
        RECT 130.090 129.560 130.855 129.700 ;
        RECT 130.090 129.500 130.410 129.560 ;
        RECT 130.565 129.515 130.855 129.560 ;
        RECT 136.160 129.560 136.760 129.700 ;
        RECT 137.540 129.700 137.680 130.240 ;
        RECT 144.350 130.180 144.670 130.440 ;
        RECT 137.950 130.040 138.240 130.085 ;
        RECT 140.050 130.040 140.340 130.085 ;
        RECT 141.620 130.040 141.910 130.085 ;
        RECT 137.950 129.900 141.910 130.040 ;
        RECT 137.950 129.855 138.240 129.900 ;
        RECT 140.050 129.855 140.340 129.900 ;
        RECT 141.620 129.855 141.910 129.900 ;
        RECT 138.345 129.700 138.635 129.745 ;
        RECT 139.535 129.700 139.825 129.745 ;
        RECT 142.055 129.700 142.345 129.745 ;
        RECT 137.540 129.560 138.140 129.700 ;
        RECT 101.585 129.360 101.875 129.405 ;
        RECT 93.290 129.220 101.875 129.360 ;
        RECT 93.290 129.160 93.610 129.220 ;
        RECT 101.585 129.175 101.875 129.220 ;
        RECT 102.505 129.175 102.795 129.405 ;
        RECT 103.425 129.360 103.715 129.405 ;
        RECT 104.330 129.360 104.650 129.420 ;
        RECT 103.425 129.220 104.650 129.360 ;
        RECT 103.425 129.175 103.715 129.220 ;
        RECT 31.190 128.880 32.800 129.020 ;
        RECT 66.610 129.020 66.930 129.080 ;
        RECT 86.850 129.020 87.170 129.080 ;
        RECT 89.610 129.020 89.930 129.080 ;
        RECT 66.610 128.880 89.930 129.020 ;
        RECT 90.160 129.020 90.300 129.160 ;
        RECT 94.225 129.020 94.515 129.065 ;
        RECT 90.160 128.880 94.515 129.020 ;
        RECT 102.580 129.020 102.720 129.175 ;
        RECT 104.330 129.160 104.650 129.220 ;
        RECT 105.710 129.160 106.030 129.420 ;
        RECT 111.690 129.360 112.010 129.420 ;
        RECT 114.005 129.360 114.295 129.405 ;
        RECT 120.890 129.360 121.210 129.420 ;
        RECT 121.365 129.360 121.655 129.405 ;
        RECT 111.690 129.220 131.700 129.360 ;
        RECT 111.690 129.160 112.010 129.220 ;
        RECT 114.005 129.175 114.295 129.220 ;
        RECT 120.890 129.160 121.210 129.220 ;
        RECT 121.365 129.175 121.655 129.220 ;
        RECT 114.450 129.020 114.770 129.080 ;
        RECT 102.580 128.880 114.770 129.020 ;
        RECT 31.190 128.820 31.510 128.880 ;
        RECT 66.610 128.820 66.930 128.880 ;
        RECT 86.850 128.820 87.170 128.880 ;
        RECT 89.610 128.820 89.930 128.880 ;
        RECT 94.225 128.835 94.515 128.880 ;
        RECT 114.450 128.820 114.770 128.880 ;
        RECT 115.340 129.020 115.630 129.065 ;
        RECT 116.750 129.020 117.070 129.080 ;
        RECT 122.730 129.065 123.050 129.080 ;
        RECT 115.340 128.880 117.070 129.020 ;
        RECT 115.340 128.835 115.630 128.880 ;
        RECT 116.750 128.820 117.070 128.880 ;
        RECT 122.700 128.835 123.050 129.065 ;
        RECT 131.560 129.020 131.700 129.220 ;
        RECT 134.690 129.160 135.010 129.420 ;
        RECT 135.165 129.360 135.455 129.405 ;
        RECT 135.610 129.360 135.930 129.420 ;
        RECT 136.160 129.405 136.300 129.560 ;
        RECT 135.165 129.220 135.930 129.360 ;
        RECT 135.165 129.175 135.455 129.220 ;
        RECT 135.610 129.160 135.930 129.220 ;
        RECT 136.085 129.175 136.375 129.405 ;
        RECT 136.545 129.360 136.835 129.405 ;
        RECT 136.990 129.360 137.310 129.420 ;
        RECT 136.545 129.220 137.310 129.360 ;
        RECT 136.545 129.175 136.835 129.220 ;
        RECT 136.990 129.160 137.310 129.220 ;
        RECT 137.465 129.175 137.755 129.405 ;
        RECT 138.000 129.360 138.140 129.560 ;
        RECT 138.345 129.560 142.345 129.700 ;
        RECT 138.345 129.515 138.635 129.560 ;
        RECT 139.535 129.515 139.825 129.560 ;
        RECT 142.055 129.515 142.345 129.560 ;
        RECT 138.745 129.360 139.035 129.405 ;
        RECT 138.000 129.220 139.035 129.360 ;
        RECT 138.745 129.175 139.035 129.220 ;
        RECT 137.540 129.020 137.680 129.175 ;
        RECT 131.560 128.880 137.680 129.020 ;
        RECT 122.730 128.820 123.050 128.835 ;
        RECT 136.160 128.740 136.300 128.880 ;
        RECT 70.290 128.680 70.610 128.740 ;
        RECT 73.065 128.680 73.355 128.725 ;
        RECT 77.650 128.680 77.970 128.740 ;
        RECT 70.290 128.540 77.970 128.680 ;
        RECT 70.290 128.480 70.610 128.540 ;
        RECT 73.065 128.495 73.355 128.540 ;
        RECT 77.650 128.480 77.970 128.540 ;
        RECT 88.230 128.480 88.550 128.740 ;
        RECT 90.530 128.480 90.850 128.740 ;
        RECT 90.990 128.680 91.310 128.740 ;
        RECT 92.385 128.680 92.675 128.725 ;
        RECT 90.990 128.540 92.675 128.680 ;
        RECT 90.990 128.480 91.310 128.540 ;
        RECT 92.385 128.495 92.675 128.540 ;
        RECT 94.670 128.480 94.990 128.740 ;
        RECT 104.790 128.480 105.110 128.740 ;
        RECT 136.070 128.480 136.390 128.740 ;
        RECT 17.320 127.860 147.040 128.340 ;
        RECT 21.545 127.660 21.835 127.705 ;
        RECT 30.270 127.660 30.590 127.720 ;
        RECT 21.545 127.520 30.590 127.660 ;
        RECT 21.545 127.475 21.835 127.520 ;
        RECT 30.270 127.460 30.590 127.520 ;
        RECT 32.570 127.460 32.890 127.720 ;
        RECT 73.510 127.660 73.830 127.720 ;
        RECT 99.745 127.660 100.035 127.705 ;
        RECT 102.490 127.660 102.810 127.720 ;
        RECT 73.510 127.520 76.960 127.660 ;
        RECT 73.510 127.460 73.830 127.520 ;
        RECT 16.470 127.320 16.790 127.380 ;
        RECT 66.625 127.320 66.915 127.365 ;
        RECT 70.610 127.320 70.900 127.365 ;
        RECT 16.470 127.180 20.840 127.320 ;
        RECT 16.470 127.120 16.790 127.180 ;
        RECT 20.700 127.025 20.840 127.180 ;
        RECT 66.625 127.180 70.900 127.320 ;
        RECT 66.625 127.135 66.915 127.180 ;
        RECT 70.610 127.135 70.900 127.180 ;
        RECT 26.130 127.025 26.450 127.040 ;
        RECT 20.165 126.795 20.455 127.025 ;
        RECT 20.625 126.795 20.915 127.025 ;
        RECT 26.100 126.795 26.450 127.025 ;
        RECT 20.240 126.300 20.380 126.795 ;
        RECT 26.130 126.780 26.450 126.795 ;
        RECT 32.110 126.780 32.430 127.040 ;
        RECT 65.230 126.780 65.550 127.040 ;
        RECT 66.165 126.980 66.455 127.025 ;
        RECT 67.070 126.980 67.390 127.040 ;
        RECT 66.165 126.840 67.390 126.980 ;
        RECT 66.165 126.795 66.455 126.840 ;
        RECT 67.070 126.780 67.390 126.840 ;
        RECT 67.545 126.795 67.835 127.025 ;
        RECT 21.070 126.640 21.390 126.700 ;
        RECT 24.750 126.640 25.070 126.700 ;
        RECT 21.070 126.500 25.070 126.640 ;
        RECT 21.070 126.440 21.390 126.500 ;
        RECT 24.750 126.440 25.070 126.500 ;
        RECT 25.645 126.640 25.935 126.685 ;
        RECT 26.835 126.640 27.125 126.685 ;
        RECT 29.355 126.640 29.645 126.685 ;
        RECT 67.620 126.640 67.760 126.795 ;
        RECT 68.450 126.780 68.770 127.040 ;
        RECT 69.385 126.980 69.675 127.025 ;
        RECT 69.830 126.980 70.150 127.040 ;
        RECT 76.820 127.025 76.960 127.520 ;
        RECT 99.745 127.520 102.810 127.660 ;
        RECT 99.745 127.475 100.035 127.520 ;
        RECT 102.490 127.460 102.810 127.520 ;
        RECT 112.610 127.660 112.930 127.720 ;
        RECT 114.005 127.660 114.295 127.705 ;
        RECT 112.610 127.520 114.295 127.660 ;
        RECT 112.610 127.460 112.930 127.520 ;
        RECT 114.005 127.475 114.295 127.520 ;
        RECT 116.750 127.460 117.070 127.720 ;
        RECT 122.270 127.660 122.590 127.720 ;
        RECT 128.725 127.660 129.015 127.705 ;
        RECT 134.690 127.660 135.010 127.720 ;
        RECT 122.270 127.520 129.015 127.660 ;
        RECT 122.270 127.460 122.590 127.520 ;
        RECT 128.725 127.475 129.015 127.520 ;
        RECT 129.720 127.520 135.010 127.660 ;
        RECT 88.230 127.365 88.550 127.380 ;
        RECT 88.200 127.320 88.550 127.365 ;
        RECT 79.020 127.180 82.940 127.320 ;
        RECT 88.035 127.180 88.550 127.320 ;
        RECT 69.385 126.840 70.150 126.980 ;
        RECT 69.385 126.795 69.675 126.840 ;
        RECT 69.830 126.780 70.150 126.840 ;
        RECT 76.745 126.980 77.035 127.025 ;
        RECT 77.190 126.980 77.510 127.040 ;
        RECT 76.745 126.840 77.510 126.980 ;
        RECT 76.745 126.795 77.035 126.840 ;
        RECT 77.190 126.780 77.510 126.840 ;
        RECT 77.650 127.025 77.970 127.040 ;
        RECT 77.650 126.980 78.005 127.025 ;
        RECT 79.020 126.980 79.160 127.180 ;
        RECT 77.650 126.840 79.160 126.980 ;
        RECT 77.650 126.795 78.005 126.840 ;
        RECT 79.505 126.795 79.795 127.025 ;
        RECT 81.345 126.980 81.635 127.025 ;
        RECT 82.250 126.980 82.570 127.040 ;
        RECT 82.800 127.025 82.940 127.180 ;
        RECT 88.200 127.135 88.550 127.180 ;
        RECT 88.230 127.120 88.550 127.135 ;
        RECT 104.790 127.320 105.110 127.380 ;
        RECT 108.470 127.365 108.790 127.380 ;
        RECT 105.310 127.320 105.600 127.365 ;
        RECT 108.440 127.320 108.790 127.365 ;
        RECT 104.790 127.180 105.600 127.320 ;
        RECT 108.275 127.180 108.790 127.320 ;
        RECT 104.790 127.120 105.110 127.180 ;
        RECT 105.310 127.135 105.600 127.180 ;
        RECT 108.440 127.135 108.790 127.180 ;
        RECT 108.470 127.120 108.790 127.135 ;
        RECT 111.690 127.120 112.010 127.380 ;
        RECT 121.350 127.320 121.670 127.380 ;
        RECT 121.350 127.180 123.880 127.320 ;
        RECT 121.350 127.120 121.670 127.180 ;
        RECT 81.345 126.840 82.570 126.980 ;
        RECT 81.345 126.795 81.635 126.840 ;
        RECT 77.650 126.780 77.970 126.795 ;
        RECT 25.645 126.500 29.645 126.640 ;
        RECT 25.645 126.455 25.935 126.500 ;
        RECT 26.835 126.455 27.125 126.500 ;
        RECT 29.355 126.455 29.645 126.500 ;
        RECT 66.240 126.500 67.760 126.640 ;
        RECT 70.265 126.640 70.555 126.685 ;
        RECT 71.455 126.640 71.745 126.685 ;
        RECT 73.975 126.640 74.265 126.685 ;
        RECT 70.265 126.500 74.265 126.640 ;
        RECT 25.250 126.300 25.540 126.345 ;
        RECT 27.350 126.300 27.640 126.345 ;
        RECT 28.920 126.300 29.210 126.345 ;
        RECT 20.240 126.160 24.980 126.300 ;
        RECT 16.010 125.960 16.330 126.020 ;
        RECT 19.245 125.960 19.535 126.005 ;
        RECT 16.010 125.820 19.535 125.960 ;
        RECT 24.840 125.960 24.980 126.160 ;
        RECT 25.250 126.160 29.210 126.300 ;
        RECT 25.250 126.115 25.540 126.160 ;
        RECT 27.350 126.115 27.640 126.160 ;
        RECT 28.920 126.115 29.210 126.160 ;
        RECT 66.240 126.020 66.380 126.500 ;
        RECT 70.265 126.455 70.555 126.500 ;
        RECT 71.455 126.455 71.745 126.500 ;
        RECT 73.975 126.455 74.265 126.500 ;
        RECT 79.580 126.640 79.720 126.795 ;
        RECT 82.250 126.780 82.570 126.840 ;
        RECT 82.725 126.795 83.015 127.025 ;
        RECT 84.565 126.980 84.855 127.025 ;
        RECT 85.930 126.980 86.250 127.040 ;
        RECT 84.565 126.840 86.250 126.980 ;
        RECT 84.565 126.795 84.855 126.840 ;
        RECT 80.410 126.640 80.730 126.700 ;
        RECT 84.640 126.640 84.780 126.795 ;
        RECT 85.930 126.780 86.250 126.840 ;
        RECT 86.865 126.980 87.155 127.025 ;
        RECT 87.310 126.980 87.630 127.040 ;
        RECT 86.865 126.840 87.630 126.980 ;
        RECT 86.865 126.795 87.155 126.840 ;
        RECT 87.310 126.780 87.630 126.840 ;
        RECT 106.645 126.980 106.935 127.025 ;
        RECT 107.105 126.980 107.395 127.025 ;
        RECT 111.780 126.980 111.920 127.120 ;
        RECT 106.645 126.840 111.920 126.980 ;
        RECT 106.645 126.795 106.935 126.840 ;
        RECT 107.105 126.795 107.395 126.840 ;
        RECT 117.670 126.780 117.990 127.040 ;
        RECT 118.590 126.780 118.910 127.040 ;
        RECT 123.740 127.025 123.880 127.180 ;
        RECT 123.665 126.795 123.955 127.025 ;
        RECT 127.330 126.780 127.650 127.040 ;
        RECT 129.720 127.025 129.860 127.520 ;
        RECT 134.690 127.460 135.010 127.520 ;
        RECT 144.810 127.460 145.130 127.720 ;
        RECT 133.325 127.320 133.615 127.365 ;
        RECT 130.180 127.180 140.900 127.320 ;
        RECT 130.180 127.025 130.320 127.180 ;
        RECT 133.325 127.135 133.615 127.180 ;
        RECT 129.645 126.795 129.935 127.025 ;
        RECT 130.105 126.795 130.395 127.025 ;
        RECT 131.025 126.795 131.315 127.025 ;
        RECT 79.580 126.500 80.730 126.640 ;
        RECT 69.870 126.300 70.160 126.345 ;
        RECT 71.970 126.300 72.260 126.345 ;
        RECT 73.540 126.300 73.830 126.345 ;
        RECT 77.205 126.300 77.495 126.345 ;
        RECT 69.870 126.160 73.830 126.300 ;
        RECT 69.870 126.115 70.160 126.160 ;
        RECT 71.970 126.115 72.260 126.160 ;
        RECT 73.540 126.115 73.830 126.160 ;
        RECT 75.440 126.160 77.495 126.300 ;
        RECT 31.650 125.960 31.970 126.020 ;
        RECT 24.840 125.820 31.970 125.960 ;
        RECT 16.010 125.760 16.330 125.820 ;
        RECT 19.245 125.775 19.535 125.820 ;
        RECT 31.650 125.760 31.970 125.820 ;
        RECT 66.150 125.760 66.470 126.020 ;
        RECT 67.070 125.960 67.390 126.020 ;
        RECT 75.440 125.960 75.580 126.160 ;
        RECT 77.205 126.115 77.495 126.160 ;
        RECT 67.070 125.820 75.580 125.960 ;
        RECT 76.270 125.960 76.590 126.020 ;
        RECT 79.580 125.960 79.720 126.500 ;
        RECT 80.410 126.440 80.730 126.500 ;
        RECT 81.420 126.500 84.780 126.640 ;
        RECT 87.745 126.640 88.035 126.685 ;
        RECT 88.935 126.640 89.225 126.685 ;
        RECT 91.455 126.640 91.745 126.685 ;
        RECT 87.745 126.500 91.745 126.640 ;
        RECT 76.270 125.820 79.720 125.960 ;
        RECT 79.950 125.960 80.270 126.020 ;
        RECT 81.420 126.005 81.560 126.500 ;
        RECT 87.745 126.455 88.035 126.500 ;
        RECT 88.935 126.455 89.225 126.500 ;
        RECT 91.455 126.455 91.745 126.500 ;
        RECT 102.055 126.640 102.345 126.685 ;
        RECT 104.575 126.640 104.865 126.685 ;
        RECT 105.765 126.640 106.055 126.685 ;
        RECT 102.055 126.500 106.055 126.640 ;
        RECT 102.055 126.455 102.345 126.500 ;
        RECT 104.575 126.455 104.865 126.500 ;
        RECT 105.765 126.455 106.055 126.500 ;
        RECT 107.985 126.640 108.275 126.685 ;
        RECT 109.175 126.640 109.465 126.685 ;
        RECT 111.695 126.640 111.985 126.685 ;
        RECT 107.985 126.500 111.985 126.640 ;
        RECT 107.985 126.455 108.275 126.500 ;
        RECT 109.175 126.455 109.465 126.500 ;
        RECT 111.695 126.455 111.985 126.500 ;
        RECT 119.065 126.640 119.355 126.685 ;
        RECT 120.905 126.640 121.195 126.685 ;
        RECT 129.720 126.640 129.860 126.795 ;
        RECT 119.065 126.500 121.195 126.640 ;
        RECT 119.065 126.455 119.355 126.500 ;
        RECT 120.905 126.455 121.195 126.500 ;
        RECT 122.360 126.500 129.860 126.640 ;
        RECT 81.790 126.300 82.110 126.360 ;
        RECT 87.350 126.300 87.640 126.345 ;
        RECT 89.450 126.300 89.740 126.345 ;
        RECT 91.020 126.300 91.310 126.345 ;
        RECT 81.790 126.160 83.400 126.300 ;
        RECT 81.790 126.100 82.110 126.160 ;
        RECT 81.345 125.960 81.635 126.005 ;
        RECT 79.950 125.820 81.635 125.960 ;
        RECT 67.070 125.760 67.390 125.820 ;
        RECT 76.270 125.760 76.590 125.820 ;
        RECT 79.950 125.760 80.270 125.820 ;
        RECT 81.345 125.775 81.635 125.820 ;
        RECT 82.250 125.760 82.570 126.020 ;
        RECT 83.260 126.005 83.400 126.160 ;
        RECT 87.350 126.160 91.310 126.300 ;
        RECT 87.350 126.115 87.640 126.160 ;
        RECT 89.450 126.115 89.740 126.160 ;
        RECT 91.020 126.115 91.310 126.160 ;
        RECT 102.490 126.300 102.780 126.345 ;
        RECT 104.060 126.300 104.350 126.345 ;
        RECT 106.160 126.300 106.450 126.345 ;
        RECT 102.490 126.160 106.450 126.300 ;
        RECT 102.490 126.115 102.780 126.160 ;
        RECT 104.060 126.115 104.350 126.160 ;
        RECT 106.160 126.115 106.450 126.160 ;
        RECT 107.590 126.300 107.880 126.345 ;
        RECT 109.690 126.300 109.980 126.345 ;
        RECT 111.260 126.300 111.550 126.345 ;
        RECT 107.590 126.160 111.550 126.300 ;
        RECT 107.590 126.115 107.880 126.160 ;
        RECT 109.690 126.115 109.980 126.160 ;
        RECT 111.260 126.115 111.550 126.160 ;
        RECT 115.370 126.300 115.690 126.360 ;
        RECT 122.360 126.300 122.500 126.500 ;
        RECT 131.100 126.300 131.240 126.795 ;
        RECT 131.470 126.780 131.790 127.040 ;
        RECT 133.770 126.780 134.090 127.040 ;
        RECT 136.530 126.980 136.850 127.040 ;
        RECT 137.365 126.980 137.655 127.025 ;
        RECT 136.530 126.840 137.655 126.980 ;
        RECT 140.760 126.980 140.900 127.180 ;
        RECT 143.905 126.980 144.195 127.025 ;
        RECT 144.350 126.980 144.670 127.040 ;
        RECT 140.760 126.840 143.200 126.980 ;
        RECT 136.530 126.780 136.850 126.840 ;
        RECT 137.365 126.795 137.655 126.840 ;
        RECT 132.865 126.455 133.155 126.685 ;
        RECT 115.370 126.160 122.500 126.300 ;
        RECT 122.820 126.160 131.240 126.300 ;
        RECT 132.940 126.300 133.080 126.455 ;
        RECT 136.070 126.440 136.390 126.700 ;
        RECT 136.965 126.640 137.255 126.685 ;
        RECT 138.155 126.640 138.445 126.685 ;
        RECT 140.675 126.640 140.965 126.685 ;
        RECT 136.965 126.500 140.965 126.640 ;
        RECT 136.965 126.455 137.255 126.500 ;
        RECT 138.155 126.455 138.445 126.500 ;
        RECT 140.675 126.455 140.965 126.500 ;
        RECT 143.060 126.345 143.200 126.840 ;
        RECT 143.905 126.840 144.670 126.980 ;
        RECT 143.905 126.795 144.195 126.840 ;
        RECT 144.350 126.780 144.670 126.840 ;
        RECT 136.570 126.300 136.860 126.345 ;
        RECT 138.670 126.300 138.960 126.345 ;
        RECT 140.240 126.300 140.530 126.345 ;
        RECT 132.940 126.160 136.300 126.300 ;
        RECT 115.370 126.100 115.690 126.160 ;
        RECT 83.185 125.775 83.475 126.005 ;
        RECT 84.550 125.960 84.870 126.020 ;
        RECT 85.485 125.960 85.775 126.005 ;
        RECT 84.550 125.820 85.775 125.960 ;
        RECT 84.550 125.760 84.870 125.820 ;
        RECT 85.485 125.775 85.775 125.820 ;
        RECT 90.530 125.960 90.850 126.020 ;
        RECT 93.750 125.960 94.070 126.020 ;
        RECT 90.530 125.820 94.070 125.960 ;
        RECT 90.530 125.760 90.850 125.820 ;
        RECT 93.750 125.760 94.070 125.820 ;
        RECT 119.510 125.960 119.830 126.020 ;
        RECT 122.820 125.960 122.960 126.160 ;
        RECT 119.510 125.820 122.960 125.960 ;
        RECT 123.190 125.960 123.510 126.020 ;
        RECT 124.585 125.960 124.875 126.005 ;
        RECT 123.190 125.820 124.875 125.960 ;
        RECT 119.510 125.760 119.830 125.820 ;
        RECT 123.190 125.760 123.510 125.820 ;
        RECT 124.585 125.775 124.875 125.820 ;
        RECT 135.610 125.760 135.930 126.020 ;
        RECT 136.160 125.960 136.300 126.160 ;
        RECT 136.570 126.160 140.530 126.300 ;
        RECT 136.570 126.115 136.860 126.160 ;
        RECT 138.670 126.115 138.960 126.160 ;
        RECT 140.240 126.115 140.530 126.160 ;
        RECT 142.985 126.300 143.275 126.345 ;
        RECT 143.890 126.300 144.210 126.360 ;
        RECT 142.985 126.160 144.210 126.300 ;
        RECT 142.985 126.115 143.275 126.160 ;
        RECT 143.890 126.100 144.210 126.160 ;
        RECT 140.670 125.960 140.990 126.020 ;
        RECT 136.160 125.820 140.990 125.960 ;
        RECT 140.670 125.760 140.990 125.820 ;
        RECT 17.320 125.140 147.040 125.620 ;
        RECT 26.130 124.940 26.450 125.000 ;
        RECT 27.065 124.940 27.355 124.985 ;
        RECT 26.130 124.800 27.355 124.940 ;
        RECT 26.130 124.740 26.450 124.800 ;
        RECT 27.065 124.755 27.355 124.800 ;
        RECT 65.230 124.940 65.550 125.000 ;
        RECT 68.450 124.940 68.770 125.000 ;
        RECT 69.845 124.940 70.135 124.985 ;
        RECT 76.270 124.940 76.590 125.000 ;
        RECT 65.230 124.800 68.220 124.940 ;
        RECT 65.230 124.740 65.550 124.800 ;
        RECT 19.730 124.600 20.020 124.645 ;
        RECT 21.830 124.600 22.120 124.645 ;
        RECT 23.400 124.600 23.690 124.645 ;
        RECT 19.730 124.460 23.690 124.600 ;
        RECT 19.730 124.415 20.020 124.460 ;
        RECT 21.830 124.415 22.120 124.460 ;
        RECT 23.400 124.415 23.690 124.460 ;
        RECT 28.445 124.600 28.735 124.645 ;
        RECT 31.190 124.600 31.510 124.660 ;
        RECT 28.445 124.460 31.510 124.600 ;
        RECT 28.445 124.415 28.735 124.460 ;
        RECT 31.190 124.400 31.510 124.460 ;
        RECT 62.510 124.600 62.800 124.645 ;
        RECT 64.610 124.600 64.900 124.645 ;
        RECT 66.180 124.600 66.470 124.645 ;
        RECT 62.510 124.460 66.470 124.600 ;
        RECT 62.510 124.415 62.800 124.460 ;
        RECT 64.610 124.415 64.900 124.460 ;
        RECT 66.180 124.415 66.470 124.460 ;
        RECT 20.125 124.260 20.415 124.305 ;
        RECT 21.315 124.260 21.605 124.305 ;
        RECT 23.835 124.260 24.125 124.305 ;
        RECT 20.125 124.120 24.125 124.260 ;
        RECT 20.125 124.075 20.415 124.120 ;
        RECT 21.315 124.075 21.605 124.120 ;
        RECT 23.835 124.075 24.125 124.120 ;
        RECT 28.905 124.260 29.195 124.305 ;
        RECT 33.505 124.260 33.795 124.305 ;
        RECT 28.905 124.120 33.795 124.260 ;
        RECT 28.905 124.075 29.195 124.120 ;
        RECT 33.505 124.075 33.795 124.120 ;
        RECT 62.905 124.260 63.195 124.305 ;
        RECT 64.095 124.260 64.385 124.305 ;
        RECT 66.615 124.260 66.905 124.305 ;
        RECT 62.905 124.120 66.905 124.260 ;
        RECT 68.080 124.260 68.220 124.800 ;
        RECT 68.450 124.800 70.135 124.940 ;
        RECT 68.450 124.740 68.770 124.800 ;
        RECT 69.845 124.755 70.135 124.800 ;
        RECT 71.760 124.800 76.590 124.940 ;
        RECT 71.760 124.305 71.900 124.800 ;
        RECT 76.270 124.740 76.590 124.800 ;
        RECT 77.190 124.940 77.510 125.000 ;
        RECT 79.505 124.940 79.795 124.985 ;
        RECT 79.950 124.940 80.270 125.000 ;
        RECT 113.530 124.940 113.850 125.000 ;
        RECT 114.925 124.940 115.215 124.985 ;
        RECT 115.370 124.940 115.690 125.000 ;
        RECT 77.190 124.800 80.270 124.940 ;
        RECT 77.190 124.740 77.510 124.800 ;
        RECT 79.505 124.755 79.795 124.800 ;
        RECT 79.950 124.740 80.270 124.800 ;
        RECT 101.660 124.800 112.840 124.940 ;
        RECT 73.090 124.600 73.380 124.645 ;
        RECT 75.190 124.600 75.480 124.645 ;
        RECT 76.760 124.600 77.050 124.645 ;
        RECT 73.090 124.460 77.050 124.600 ;
        RECT 73.090 124.415 73.380 124.460 ;
        RECT 75.190 124.415 75.480 124.460 ;
        RECT 76.760 124.415 77.050 124.460 ;
        RECT 88.270 124.600 88.560 124.645 ;
        RECT 90.370 124.600 90.660 124.645 ;
        RECT 91.940 124.600 92.230 124.645 ;
        RECT 88.270 124.460 92.230 124.600 ;
        RECT 88.270 124.415 88.560 124.460 ;
        RECT 90.370 124.415 90.660 124.460 ;
        RECT 91.940 124.415 92.230 124.460 ;
        RECT 71.685 124.260 71.975 124.305 ;
        RECT 68.080 124.120 71.975 124.260 ;
        RECT 62.905 124.075 63.195 124.120 ;
        RECT 64.095 124.075 64.385 124.120 ;
        RECT 66.615 124.075 66.905 124.120 ;
        RECT 71.685 124.075 71.975 124.120 ;
        RECT 72.130 124.260 72.450 124.320 ;
        RECT 72.605 124.260 72.895 124.305 ;
        RECT 72.130 124.120 72.895 124.260 ;
        RECT 72.130 124.060 72.450 124.120 ;
        RECT 72.605 124.075 72.895 124.120 ;
        RECT 73.485 124.260 73.775 124.305 ;
        RECT 74.675 124.260 74.965 124.305 ;
        RECT 77.195 124.260 77.485 124.305 ;
        RECT 73.485 124.120 77.485 124.260 ;
        RECT 73.485 124.075 73.775 124.120 ;
        RECT 74.675 124.075 74.965 124.120 ;
        RECT 77.195 124.075 77.485 124.120 ;
        RECT 84.550 124.060 84.870 124.320 ;
        RECT 87.770 124.060 88.090 124.320 ;
        RECT 88.665 124.260 88.955 124.305 ;
        RECT 89.855 124.260 90.145 124.305 ;
        RECT 92.375 124.260 92.665 124.305 ;
        RECT 88.665 124.120 92.665 124.260 ;
        RECT 88.665 124.075 88.955 124.120 ;
        RECT 89.855 124.075 90.145 124.120 ;
        RECT 92.375 124.075 92.665 124.120 ;
        RECT 93.750 124.260 94.070 124.320 ;
        RECT 100.205 124.260 100.495 124.305 ;
        RECT 101.660 124.260 101.800 124.800 ;
        RECT 107.105 124.415 107.395 124.645 ;
        RECT 108.510 124.600 108.800 124.645 ;
        RECT 110.610 124.600 110.900 124.645 ;
        RECT 112.180 124.600 112.470 124.645 ;
        RECT 108.510 124.460 112.470 124.600 ;
        RECT 112.700 124.600 112.840 124.800 ;
        RECT 113.530 124.800 115.690 124.940 ;
        RECT 113.530 124.740 113.850 124.800 ;
        RECT 114.925 124.755 115.215 124.800 ;
        RECT 115.370 124.740 115.690 124.800 ;
        RECT 120.905 124.940 121.195 124.985 ;
        RECT 122.730 124.940 123.050 125.000 ;
        RECT 120.905 124.800 123.050 124.940 ;
        RECT 120.905 124.755 121.195 124.800 ;
        RECT 122.730 124.740 123.050 124.800 ;
        RECT 136.085 124.940 136.375 124.985 ;
        RECT 136.530 124.940 136.850 125.000 ;
        RECT 136.085 124.800 136.850 124.940 ;
        RECT 136.085 124.755 136.375 124.800 ;
        RECT 136.530 124.740 136.850 124.800 ;
        RECT 144.810 124.740 145.130 125.000 ;
        RECT 128.250 124.600 128.570 124.660 ;
        RECT 131.010 124.600 131.330 124.660 ;
        RECT 112.700 124.460 131.330 124.600 ;
        RECT 108.510 124.415 108.800 124.460 ;
        RECT 110.610 124.415 110.900 124.460 ;
        RECT 112.180 124.415 112.470 124.460 ;
        RECT 93.750 124.120 101.800 124.260 ;
        RECT 103.410 124.260 103.730 124.320 ;
        RECT 103.885 124.260 104.175 124.305 ;
        RECT 103.410 124.120 104.175 124.260 ;
        RECT 93.750 124.060 94.070 124.120 ;
        RECT 100.205 124.075 100.495 124.120 ;
        RECT 103.410 124.060 103.730 124.120 ;
        RECT 103.885 124.075 104.175 124.120 ;
        RECT 104.330 124.260 104.650 124.320 ;
        RECT 104.805 124.260 105.095 124.305 ;
        RECT 104.330 124.120 105.095 124.260 ;
        RECT 104.330 124.060 104.650 124.120 ;
        RECT 104.805 124.075 105.095 124.120 ;
        RECT 19.245 123.920 19.535 123.965 ;
        RECT 19.690 123.920 20.010 123.980 ;
        RECT 19.245 123.780 20.010 123.920 ;
        RECT 19.245 123.735 19.535 123.780 ;
        RECT 19.690 123.720 20.010 123.780 ;
        RECT 27.985 123.735 28.275 123.965 ;
        RECT 29.365 123.920 29.655 123.965 ;
        RECT 30.745 123.920 31.035 123.965 ;
        RECT 29.365 123.780 31.035 123.920 ;
        RECT 29.365 123.735 29.655 123.780 ;
        RECT 30.745 123.735 31.035 123.780 ;
        RECT 20.580 123.580 20.870 123.625 ;
        RECT 21.990 123.580 22.310 123.640 ;
        RECT 20.580 123.440 22.310 123.580 ;
        RECT 20.580 123.395 20.870 123.440 ;
        RECT 21.990 123.380 22.310 123.440 ;
        RECT 26.130 123.040 26.450 123.300 ;
        RECT 28.060 123.240 28.200 123.735 ;
        RECT 31.650 123.720 31.970 123.980 ;
        RECT 33.965 123.920 34.255 123.965 ;
        RECT 33.965 123.780 34.365 123.920 ;
        RECT 33.965 123.735 34.255 123.780 ;
        RECT 32.570 123.580 32.890 123.640 ;
        RECT 34.040 123.580 34.180 123.735 ;
        RECT 62.010 123.720 62.330 123.980 ;
        RECT 67.070 123.920 67.390 123.980 ;
        RECT 73.970 123.965 74.290 123.980 ;
        RECT 70.765 123.920 71.055 123.965 ;
        RECT 67.070 123.780 71.055 123.920 ;
        RECT 67.070 123.720 67.390 123.780 ;
        RECT 70.765 123.735 71.055 123.780 ;
        RECT 73.940 123.735 74.290 123.965 ;
        RECT 85.485 123.920 85.775 123.965 ;
        RECT 86.390 123.920 86.710 123.980 ;
        RECT 85.485 123.780 86.710 123.920 ;
        RECT 85.485 123.735 85.775 123.780 ;
        RECT 73.970 123.720 74.290 123.735 ;
        RECT 86.390 123.720 86.710 123.780 ;
        RECT 89.120 123.920 89.410 123.965 ;
        RECT 90.990 123.920 91.310 123.980 ;
        RECT 89.120 123.780 91.310 123.920 ;
        RECT 89.120 123.735 89.410 123.780 ;
        RECT 90.990 123.720 91.310 123.780 ;
        RECT 98.810 123.720 99.130 123.980 ;
        RECT 107.180 123.920 107.320 124.415 ;
        RECT 128.250 124.400 128.570 124.460 ;
        RECT 131.010 124.400 131.330 124.460 ;
        RECT 135.610 124.400 135.930 124.660 ;
        RECT 108.905 124.260 109.195 124.305 ;
        RECT 110.095 124.260 110.385 124.305 ;
        RECT 112.615 124.260 112.905 124.305 ;
        RECT 108.905 124.120 112.905 124.260 ;
        RECT 108.905 124.075 109.195 124.120 ;
        RECT 110.095 124.075 110.385 124.120 ;
        RECT 112.615 124.075 112.905 124.120 ;
        RECT 118.590 124.260 118.910 124.320 ;
        RECT 122.745 124.260 123.035 124.305 ;
        RECT 118.590 124.120 123.035 124.260 ;
        RECT 118.590 124.060 118.910 124.120 ;
        RECT 122.745 124.075 123.035 124.120 ;
        RECT 123.190 124.060 123.510 124.320 ;
        RECT 108.025 123.920 108.315 123.965 ;
        RECT 111.690 123.920 112.010 123.980 ;
        RECT 107.180 123.780 107.780 123.920 ;
        RECT 35.790 123.580 36.110 123.640 ;
        RECT 32.570 123.440 36.110 123.580 ;
        RECT 32.570 123.380 32.890 123.440 ;
        RECT 35.790 123.380 36.110 123.440 ;
        RECT 63.360 123.580 63.650 123.625 ;
        RECT 64.770 123.580 65.090 123.640 ;
        RECT 63.360 123.440 65.090 123.580 ;
        RECT 63.360 123.395 63.650 123.440 ;
        RECT 64.770 123.380 65.090 123.440 ;
        RECT 85.025 123.580 85.315 123.625 ;
        RECT 95.605 123.580 95.895 123.625 ;
        RECT 85.025 123.440 95.895 123.580 ;
        RECT 85.025 123.395 85.315 123.440 ;
        RECT 95.605 123.395 95.895 123.440 ;
        RECT 102.965 123.580 103.255 123.625 ;
        RECT 105.265 123.580 105.555 123.625 ;
        RECT 102.965 123.440 105.555 123.580 ;
        RECT 107.640 123.580 107.780 123.780 ;
        RECT 108.025 123.780 112.010 123.920 ;
        RECT 108.025 123.735 108.315 123.780 ;
        RECT 111.690 123.720 112.010 123.780 ;
        RECT 121.825 123.920 122.115 123.965 ;
        RECT 128.710 123.920 129.030 123.980 ;
        RECT 121.825 123.780 129.030 123.920 ;
        RECT 121.825 123.735 122.115 123.780 ;
        RECT 128.710 123.720 129.030 123.780 ;
        RECT 142.050 123.720 142.370 123.980 ;
        RECT 143.890 123.720 144.210 123.980 ;
        RECT 109.250 123.580 109.540 123.625 ;
        RECT 107.640 123.440 109.540 123.580 ;
        RECT 102.965 123.395 103.255 123.440 ;
        RECT 105.265 123.395 105.555 123.440 ;
        RECT 109.250 123.395 109.540 123.440 ;
        RECT 130.550 123.580 130.870 123.640 ;
        RECT 133.785 123.580 134.075 123.625 ;
        RECT 130.550 123.440 134.075 123.580 ;
        RECT 130.550 123.380 130.870 123.440 ;
        RECT 133.785 123.395 134.075 123.440 ;
        RECT 30.270 123.240 30.590 123.300 ;
        RECT 34.870 123.240 35.190 123.300 ;
        RECT 28.060 123.100 35.190 123.240 ;
        RECT 30.270 123.040 30.590 123.100 ;
        RECT 34.870 123.040 35.190 123.100 ;
        RECT 68.450 123.240 68.770 123.300 ;
        RECT 68.925 123.240 69.215 123.285 ;
        RECT 68.450 123.100 69.215 123.240 ;
        RECT 68.450 123.040 68.770 123.100 ;
        RECT 68.925 123.055 69.215 123.100 ;
        RECT 86.850 123.240 87.170 123.300 ;
        RECT 87.325 123.240 87.615 123.285 ;
        RECT 86.850 123.100 87.615 123.240 ;
        RECT 86.850 123.040 87.170 123.100 ;
        RECT 87.325 123.055 87.615 123.100 ;
        RECT 94.670 123.240 94.990 123.300 ;
        RECT 98.350 123.240 98.670 123.300 ;
        RECT 136.530 123.240 136.850 123.300 ;
        RECT 139.290 123.240 139.610 123.300 ;
        RECT 94.670 123.100 139.610 123.240 ;
        RECT 94.670 123.040 94.990 123.100 ;
        RECT 98.350 123.040 98.670 123.100 ;
        RECT 136.530 123.040 136.850 123.100 ;
        RECT 139.290 123.040 139.610 123.100 ;
        RECT 142.970 123.040 143.290 123.300 ;
        RECT 17.320 122.420 147.040 122.900 ;
        RECT 21.990 122.020 22.310 122.280 ;
        RECT 72.130 122.220 72.450 122.280 ;
        RECT 103.410 122.220 103.730 122.280 ;
        RECT 107.090 122.220 107.410 122.280 ;
        RECT 72.130 122.080 84.320 122.220 ;
        RECT 72.130 122.020 72.450 122.080 ;
        RECT 23.845 121.880 24.135 121.925 ;
        RECT 26.130 121.880 26.450 121.940 ;
        RECT 20.240 121.740 26.450 121.880 ;
        RECT 20.240 121.585 20.380 121.740 ;
        RECT 23.845 121.695 24.135 121.740 ;
        RECT 26.130 121.680 26.450 121.740 ;
        RECT 63.865 121.880 64.155 121.925 ;
        RECT 66.610 121.880 66.930 121.940 ;
        RECT 63.865 121.740 66.930 121.880 ;
        RECT 63.865 121.695 64.155 121.740 ;
        RECT 66.610 121.680 66.930 121.740 ;
        RECT 20.165 121.355 20.455 121.585 ;
        RECT 24.290 121.340 24.610 121.600 ;
        RECT 62.010 121.540 62.330 121.600 ;
        RECT 70.750 121.585 71.070 121.600 ;
        RECT 62.945 121.540 63.235 121.585 ;
        RECT 62.010 121.400 63.235 121.540 ;
        RECT 62.010 121.340 62.330 121.400 ;
        RECT 62.945 121.355 63.235 121.400 ;
        RECT 70.720 121.355 71.070 121.585 ;
        RECT 25.225 121.200 25.515 121.245 ;
        RECT 32.570 121.200 32.890 121.260 ;
        RECT 25.225 121.060 32.890 121.200 ;
        RECT 63.020 121.200 63.160 121.355 ;
        RECT 70.750 121.340 71.070 121.355 ;
        RECT 82.710 121.585 83.030 121.600 ;
        RECT 84.180 121.585 84.320 122.080 ;
        RECT 103.410 122.080 107.410 122.220 ;
        RECT 103.410 122.020 103.730 122.080 ;
        RECT 107.090 122.020 107.410 122.080 ;
        RECT 129.170 122.220 129.490 122.280 ;
        RECT 131.930 122.220 132.250 122.280 ;
        RECT 137.450 122.220 137.770 122.280 ;
        RECT 129.170 122.080 137.770 122.220 ;
        RECT 129.170 122.020 129.490 122.080 ;
        RECT 131.930 122.020 132.250 122.080 ;
        RECT 137.450 122.020 137.770 122.080 ;
        RECT 87.770 121.880 88.090 121.940 ;
        RECT 85.560 121.740 88.090 121.880 ;
        RECT 85.560 121.585 85.700 121.740 ;
        RECT 87.770 121.680 88.090 121.740 ;
        RECT 104.330 121.880 104.650 121.940 ;
        RECT 104.330 121.740 108.700 121.880 ;
        RECT 104.330 121.680 104.650 121.740 ;
        RECT 86.850 121.585 87.170 121.600 ;
        RECT 82.710 121.355 83.060 121.585 ;
        RECT 84.105 121.540 84.395 121.585 ;
        RECT 85.485 121.540 85.775 121.585 ;
        RECT 86.820 121.540 87.170 121.585 ;
        RECT 84.105 121.400 85.775 121.540 ;
        RECT 86.655 121.400 87.170 121.540 ;
        RECT 84.105 121.355 84.395 121.400 ;
        RECT 85.485 121.355 85.775 121.400 ;
        RECT 86.820 121.355 87.170 121.400 ;
        RECT 82.710 121.340 83.030 121.355 ;
        RECT 86.850 121.340 87.170 121.355 ;
        RECT 106.630 121.340 106.950 121.600 ;
        RECT 107.090 121.340 107.410 121.600 ;
        RECT 108.010 121.340 108.330 121.600 ;
        RECT 108.560 121.585 108.700 121.740 ;
        RECT 109.390 121.680 109.710 121.940 ;
        RECT 142.050 121.880 142.370 121.940 ;
        RECT 121.440 121.740 142.370 121.880 ;
        RECT 108.485 121.355 108.775 121.585 ;
        RECT 111.690 121.340 112.010 121.600 ;
        RECT 112.150 121.540 112.470 121.600 ;
        RECT 112.985 121.540 113.275 121.585 ;
        RECT 112.150 121.400 113.275 121.540 ;
        RECT 112.150 121.340 112.470 121.400 ;
        RECT 112.985 121.355 113.275 121.400 ;
        RECT 66.610 121.200 66.930 121.260 ;
        RECT 68.005 121.200 68.295 121.245 ;
        RECT 69.385 121.200 69.675 121.245 ;
        RECT 63.020 121.060 69.675 121.200 ;
        RECT 25.225 121.015 25.515 121.060 ;
        RECT 32.570 121.000 32.890 121.060 ;
        RECT 66.610 121.000 66.930 121.060 ;
        RECT 68.005 121.015 68.295 121.060 ;
        RECT 69.385 121.015 69.675 121.060 ;
        RECT 70.265 121.200 70.555 121.245 ;
        RECT 71.455 121.200 71.745 121.245 ;
        RECT 73.975 121.200 74.265 121.245 ;
        RECT 70.265 121.060 74.265 121.200 ;
        RECT 70.265 121.015 70.555 121.060 ;
        RECT 71.455 121.015 71.745 121.060 ;
        RECT 73.975 121.015 74.265 121.060 ;
        RECT 79.515 121.200 79.805 121.245 ;
        RECT 82.035 121.200 82.325 121.245 ;
        RECT 83.225 121.200 83.515 121.245 ;
        RECT 79.515 121.060 83.515 121.200 ;
        RECT 79.515 121.015 79.805 121.060 ;
        RECT 82.035 121.015 82.325 121.060 ;
        RECT 83.225 121.015 83.515 121.060 ;
        RECT 86.365 121.200 86.655 121.245 ;
        RECT 87.555 121.200 87.845 121.245 ;
        RECT 90.075 121.200 90.365 121.245 ;
        RECT 98.365 121.200 98.655 121.245 ;
        RECT 98.810 121.200 99.130 121.260 ;
        RECT 111.230 121.200 111.550 121.260 ;
        RECT 86.365 121.060 90.365 121.200 ;
        RECT 86.365 121.015 86.655 121.060 ;
        RECT 87.555 121.015 87.845 121.060 ;
        RECT 90.075 121.015 90.365 121.060 ;
        RECT 92.460 121.060 111.550 121.200 ;
        RECT 16.010 120.860 16.330 120.920 ;
        RECT 92.460 120.905 92.600 121.060 ;
        RECT 98.365 121.015 98.655 121.060 ;
        RECT 98.810 121.000 99.130 121.060 ;
        RECT 111.230 121.000 111.550 121.060 ;
        RECT 112.585 121.200 112.875 121.245 ;
        RECT 113.775 121.200 114.065 121.245 ;
        RECT 116.295 121.200 116.585 121.245 ;
        RECT 112.585 121.060 116.585 121.200 ;
        RECT 112.585 121.015 112.875 121.060 ;
        RECT 113.775 121.015 114.065 121.060 ;
        RECT 116.295 121.015 116.585 121.060 ;
        RECT 19.245 120.860 19.535 120.905 ;
        RECT 16.010 120.720 19.535 120.860 ;
        RECT 16.010 120.660 16.330 120.720 ;
        RECT 19.245 120.675 19.535 120.720 ;
        RECT 69.870 120.860 70.160 120.905 ;
        RECT 71.970 120.860 72.260 120.905 ;
        RECT 73.540 120.860 73.830 120.905 ;
        RECT 69.870 120.720 73.830 120.860 ;
        RECT 69.870 120.675 70.160 120.720 ;
        RECT 71.970 120.675 72.260 120.720 ;
        RECT 73.540 120.675 73.830 120.720 ;
        RECT 79.950 120.860 80.240 120.905 ;
        RECT 81.520 120.860 81.810 120.905 ;
        RECT 83.620 120.860 83.910 120.905 ;
        RECT 79.950 120.720 83.910 120.860 ;
        RECT 79.950 120.675 80.240 120.720 ;
        RECT 81.520 120.675 81.810 120.720 ;
        RECT 83.620 120.675 83.910 120.720 ;
        RECT 85.970 120.860 86.260 120.905 ;
        RECT 88.070 120.860 88.360 120.905 ;
        RECT 89.640 120.860 89.930 120.905 ;
        RECT 85.970 120.720 89.930 120.860 ;
        RECT 85.970 120.675 86.260 120.720 ;
        RECT 88.070 120.675 88.360 120.720 ;
        RECT 89.640 120.675 89.930 120.720 ;
        RECT 92.385 120.675 92.675 120.905 ;
        RECT 112.190 120.860 112.480 120.905 ;
        RECT 114.290 120.860 114.580 120.905 ;
        RECT 115.860 120.860 116.150 120.905 ;
        RECT 112.190 120.720 116.150 120.860 ;
        RECT 112.190 120.675 112.480 120.720 ;
        RECT 114.290 120.675 114.580 120.720 ;
        RECT 115.860 120.675 116.150 120.720 ;
        RECT 118.605 120.860 118.895 120.905 ;
        RECT 121.440 120.860 121.580 121.740 ;
        RECT 142.050 121.680 142.370 121.740 ;
        RECT 129.645 121.540 129.935 121.585 ;
        RECT 130.090 121.540 130.410 121.600 ;
        RECT 134.230 121.540 134.550 121.600 ;
        RECT 129.645 121.400 134.550 121.540 ;
        RECT 129.645 121.355 129.935 121.400 ;
        RECT 130.090 121.340 130.410 121.400 ;
        RECT 134.230 121.340 134.550 121.400 ;
        RECT 123.205 121.200 123.495 121.245 ;
        RECT 126.410 121.200 126.730 121.260 ;
        RECT 130.550 121.200 130.870 121.260 ;
        RECT 123.205 121.060 130.870 121.200 ;
        RECT 123.205 121.015 123.495 121.060 ;
        RECT 126.410 121.000 126.730 121.060 ;
        RECT 130.550 121.000 130.870 121.060 ;
        RECT 137.925 121.015 138.215 121.245 ;
        RECT 138.370 121.200 138.690 121.260 ;
        RECT 138.845 121.200 139.135 121.245 ;
        RECT 140.670 121.200 140.990 121.260 ;
        RECT 138.370 121.060 140.990 121.200 ;
        RECT 118.605 120.720 121.580 120.860 ;
        RECT 121.825 120.860 122.115 120.905 ;
        RECT 126.870 120.860 127.190 120.920 ;
        RECT 121.825 120.720 127.190 120.860 ;
        RECT 118.605 120.675 118.895 120.720 ;
        RECT 121.825 120.675 122.115 120.720 ;
        RECT 73.050 120.520 73.370 120.580 ;
        RECT 76.285 120.520 76.575 120.565 ;
        RECT 73.050 120.380 76.575 120.520 ;
        RECT 73.050 120.320 73.370 120.380 ;
        RECT 76.285 120.335 76.575 120.380 ;
        RECT 77.190 120.320 77.510 120.580 ;
        RECT 101.125 120.520 101.415 120.565 ;
        RECT 102.490 120.520 102.810 120.580 ;
        RECT 101.125 120.380 102.810 120.520 ;
        RECT 101.125 120.335 101.415 120.380 ;
        RECT 102.490 120.320 102.810 120.380 ;
        RECT 108.010 120.520 108.330 120.580 ;
        RECT 118.680 120.520 118.820 120.675 ;
        RECT 126.870 120.660 127.190 120.720 ;
        RECT 131.485 120.860 131.775 120.905 ;
        RECT 133.770 120.860 134.090 120.920 ;
        RECT 131.485 120.720 134.090 120.860 ;
        RECT 131.485 120.675 131.775 120.720 ;
        RECT 133.770 120.660 134.090 120.720 ;
        RECT 135.150 120.860 135.470 120.920 ;
        RECT 138.000 120.860 138.140 121.015 ;
        RECT 138.370 121.000 138.690 121.060 ;
        RECT 138.845 121.015 139.135 121.060 ;
        RECT 140.670 121.000 140.990 121.060 ;
        RECT 135.150 120.720 138.140 120.860 ;
        RECT 135.150 120.660 135.470 120.720 ;
        RECT 108.010 120.380 118.820 120.520 ;
        RECT 120.905 120.520 121.195 120.565 ;
        RECT 121.350 120.520 121.670 120.580 ;
        RECT 120.905 120.380 121.670 120.520 ;
        RECT 108.010 120.320 108.330 120.380 ;
        RECT 120.905 120.335 121.195 120.380 ;
        RECT 121.350 120.320 121.670 120.380 ;
        RECT 131.930 120.320 132.250 120.580 ;
        RECT 132.390 120.520 132.710 120.580 ;
        RECT 135.625 120.520 135.915 120.565 ;
        RECT 132.390 120.380 135.915 120.520 ;
        RECT 132.390 120.320 132.710 120.380 ;
        RECT 135.625 120.335 135.915 120.380 ;
        RECT 17.320 119.700 147.040 120.180 ;
        RECT 64.770 119.300 65.090 119.560 ;
        RECT 70.750 119.500 71.070 119.560 ;
        RECT 71.685 119.500 71.975 119.545 ;
        RECT 70.750 119.360 71.975 119.500 ;
        RECT 70.750 119.300 71.070 119.360 ;
        RECT 71.685 119.315 71.975 119.360 ;
        RECT 82.265 119.500 82.555 119.545 ;
        RECT 82.710 119.500 83.030 119.560 ;
        RECT 82.265 119.360 83.030 119.500 ;
        RECT 82.265 119.315 82.555 119.360 ;
        RECT 82.710 119.300 83.030 119.360 ;
        RECT 111.245 119.500 111.535 119.545 ;
        RECT 112.150 119.500 112.470 119.560 ;
        RECT 111.245 119.360 112.470 119.500 ;
        RECT 111.245 119.315 111.535 119.360 ;
        RECT 112.150 119.300 112.470 119.360 ;
        RECT 117.670 119.300 117.990 119.560 ;
        RECT 128.710 119.500 129.030 119.560 ;
        RECT 133.785 119.500 134.075 119.545 ;
        RECT 128.710 119.360 134.075 119.500 ;
        RECT 128.710 119.300 129.030 119.360 ;
        RECT 133.785 119.315 134.075 119.360 ;
        RECT 16.010 119.160 16.330 119.220 ;
        RECT 19.245 119.160 19.535 119.205 ;
        RECT 101.570 119.160 101.890 119.220 ;
        RECT 16.010 119.020 19.535 119.160 ;
        RECT 16.010 118.960 16.330 119.020 ;
        RECT 19.245 118.975 19.535 119.020 ;
        RECT 91.080 119.020 101.890 119.160 ;
        RECT 66.150 118.820 66.470 118.880 ;
        RECT 67.545 118.820 67.835 118.865 ;
        RECT 20.240 118.680 25.670 118.820 ;
        RECT 20.240 118.525 20.380 118.680 ;
        RECT 25.530 118.540 25.670 118.680 ;
        RECT 66.150 118.680 67.835 118.820 ;
        RECT 66.150 118.620 66.470 118.680 ;
        RECT 67.545 118.635 67.835 118.680 ;
        RECT 72.590 118.820 72.910 118.880 ;
        RECT 74.445 118.820 74.735 118.865 ;
        RECT 72.590 118.680 74.735 118.820 ;
        RECT 72.590 118.620 72.910 118.680 ;
        RECT 74.445 118.635 74.735 118.680 ;
        RECT 82.250 118.820 82.570 118.880 ;
        RECT 85.025 118.820 85.315 118.865 ;
        RECT 91.080 118.820 91.220 119.020 ;
        RECT 101.570 118.960 101.890 119.020 ;
        RECT 110.785 119.160 111.075 119.205 ;
        RECT 111.705 119.160 111.995 119.205 ;
        RECT 110.785 119.020 111.995 119.160 ;
        RECT 110.785 118.975 111.075 119.020 ;
        RECT 111.705 118.975 111.995 119.020 ;
        RECT 121.390 119.160 121.680 119.205 ;
        RECT 123.490 119.160 123.780 119.205 ;
        RECT 125.060 119.160 125.350 119.205 ;
        RECT 121.390 119.020 125.350 119.160 ;
        RECT 121.390 118.975 121.680 119.020 ;
        RECT 123.490 118.975 123.780 119.020 ;
        RECT 125.060 118.975 125.350 119.020 ;
        RECT 132.390 118.960 132.710 119.220 ;
        RECT 136.070 119.160 136.390 119.220 ;
        RECT 137.950 119.160 138.240 119.205 ;
        RECT 140.050 119.160 140.340 119.205 ;
        RECT 141.620 119.160 141.910 119.205 ;
        RECT 136.070 119.020 137.680 119.160 ;
        RECT 136.070 118.960 136.390 119.020 ;
        RECT 82.250 118.680 85.315 118.820 ;
        RECT 82.250 118.620 82.570 118.680 ;
        RECT 85.025 118.635 85.315 118.680 ;
        RECT 89.240 118.680 91.220 118.820 ;
        RECT 99.745 118.820 100.035 118.865 ;
        RECT 103.410 118.820 103.730 118.880 ;
        RECT 99.745 118.680 103.730 118.820 ;
        RECT 20.165 118.295 20.455 118.525 ;
        RECT 21.990 118.280 22.310 118.540 ;
        RECT 25.530 118.480 25.990 118.540 ;
        RECT 27.065 118.480 27.355 118.525 ;
        RECT 25.530 118.340 27.355 118.480 ;
        RECT 25.670 118.280 25.990 118.340 ;
        RECT 27.065 118.295 27.355 118.340 ;
        RECT 67.085 118.480 67.375 118.525 ;
        RECT 68.910 118.480 69.230 118.540 ;
        RECT 73.985 118.480 74.275 118.525 ;
        RECT 67.085 118.340 74.275 118.480 ;
        RECT 67.085 118.295 67.375 118.340 ;
        RECT 68.910 118.280 69.230 118.340 ;
        RECT 73.985 118.295 74.275 118.340 ;
        RECT 84.105 118.480 84.395 118.525 ;
        RECT 86.390 118.480 86.710 118.540 ;
        RECT 89.240 118.480 89.380 118.680 ;
        RECT 99.745 118.635 100.035 118.680 ;
        RECT 103.410 118.620 103.730 118.680 ;
        RECT 108.010 118.820 108.330 118.880 ;
        RECT 114.005 118.820 114.295 118.865 ;
        RECT 108.010 118.680 114.295 118.820 ;
        RECT 108.010 118.620 108.330 118.680 ;
        RECT 114.005 118.635 114.295 118.680 ;
        RECT 114.910 118.620 115.230 118.880 ;
        RECT 115.370 118.820 115.690 118.880 ;
        RECT 121.785 118.820 122.075 118.865 ;
        RECT 122.975 118.820 123.265 118.865 ;
        RECT 125.495 118.820 125.785 118.865 ;
        RECT 115.370 118.680 118.820 118.820 ;
        RECT 115.370 118.620 115.690 118.680 ;
        RECT 84.105 118.340 86.710 118.480 ;
        RECT 84.105 118.295 84.395 118.340 ;
        RECT 86.390 118.280 86.710 118.340 ;
        RECT 88.320 118.340 89.380 118.480 ;
        RECT 89.610 118.480 89.930 118.540 ;
        RECT 96.065 118.480 96.355 118.525 ;
        RECT 118.130 118.480 118.450 118.540 ;
        RECT 118.680 118.525 118.820 118.680 ;
        RECT 121.785 118.680 125.785 118.820 ;
        RECT 121.785 118.635 122.075 118.680 ;
        RECT 122.975 118.635 123.265 118.680 ;
        RECT 125.495 118.635 125.785 118.680 ;
        RECT 130.550 118.620 130.870 118.880 ;
        RECT 136.990 118.820 137.310 118.880 ;
        RECT 137.540 118.865 137.680 119.020 ;
        RECT 137.950 119.020 141.910 119.160 ;
        RECT 137.950 118.975 138.240 119.020 ;
        RECT 140.050 118.975 140.340 119.020 ;
        RECT 141.620 118.975 141.910 119.020 ;
        RECT 136.160 118.680 137.310 118.820 ;
        RECT 89.610 118.340 118.450 118.480 ;
        RECT 26.145 118.140 26.435 118.185 ;
        RECT 26.590 118.140 26.910 118.200 ;
        RECT 26.145 118.000 26.910 118.140 ;
        RECT 26.145 117.955 26.435 118.000 ;
        RECT 26.590 117.940 26.910 118.000 ;
        RECT 73.050 118.140 73.370 118.200 ;
        RECT 73.525 118.140 73.815 118.185 ;
        RECT 73.050 118.000 73.815 118.140 ;
        RECT 73.050 117.940 73.370 118.000 ;
        RECT 73.525 117.955 73.815 118.000 ;
        RECT 77.190 118.140 77.510 118.200 ;
        RECT 84.565 118.140 84.855 118.185 ;
        RECT 88.320 118.140 88.460 118.340 ;
        RECT 89.610 118.280 89.930 118.340 ;
        RECT 96.065 118.295 96.355 118.340 ;
        RECT 118.130 118.280 118.450 118.340 ;
        RECT 118.605 118.295 118.895 118.525 ;
        RECT 119.065 118.295 119.355 118.525 ;
        RECT 77.190 118.000 88.460 118.140 ;
        RECT 88.690 118.140 89.010 118.200 ;
        RECT 91.925 118.140 92.215 118.185 ;
        RECT 88.690 118.000 92.215 118.140 ;
        RECT 77.190 117.940 77.510 118.000 ;
        RECT 84.565 117.955 84.855 118.000 ;
        RECT 86.480 117.860 86.620 118.000 ;
        RECT 88.690 117.940 89.010 118.000 ;
        RECT 91.925 117.955 92.215 118.000 ;
        RECT 98.350 117.940 98.670 118.200 ;
        RECT 98.825 118.140 99.115 118.185 ;
        RECT 102.030 118.140 102.350 118.200 ;
        RECT 98.825 118.000 102.350 118.140 ;
        RECT 98.825 117.955 99.115 118.000 ;
        RECT 102.030 117.940 102.350 118.000 ;
        RECT 102.490 117.940 102.810 118.200 ;
        RECT 108.930 117.940 109.250 118.200 ;
        RECT 113.530 117.940 113.850 118.200 ;
        RECT 21.070 117.600 21.390 117.860 ;
        RECT 27.985 117.800 28.275 117.845 ;
        RECT 31.650 117.800 31.970 117.860 ;
        RECT 27.985 117.660 31.970 117.800 ;
        RECT 27.985 117.615 28.275 117.660 ;
        RECT 31.650 117.600 31.970 117.660 ;
        RECT 66.625 117.800 66.915 117.845 ;
        RECT 68.450 117.800 68.770 117.860 ;
        RECT 71.670 117.800 71.990 117.860 ;
        RECT 66.625 117.660 71.990 117.800 ;
        RECT 66.625 117.615 66.915 117.660 ;
        RECT 68.450 117.600 68.770 117.660 ;
        RECT 71.670 117.600 71.990 117.660 ;
        RECT 86.390 117.600 86.710 117.860 ;
        RECT 96.510 117.600 96.830 117.860 ;
        RECT 99.270 117.800 99.590 117.860 ;
        RECT 100.665 117.800 100.955 117.845 ;
        RECT 99.270 117.660 100.955 117.800 ;
        RECT 99.270 117.600 99.590 117.660 ;
        RECT 100.665 117.615 100.955 117.660 ;
        RECT 102.965 117.800 103.255 117.845 ;
        RECT 103.870 117.800 104.190 117.860 ;
        RECT 102.965 117.660 104.190 117.800 ;
        RECT 119.140 117.800 119.280 118.295 ;
        RECT 119.970 118.280 120.290 118.540 ;
        RECT 120.445 118.295 120.735 118.525 ;
        RECT 120.890 118.480 121.210 118.540 ;
        RECT 125.030 118.480 125.350 118.540 ;
        RECT 120.890 118.340 125.350 118.480 ;
        RECT 119.510 118.140 119.830 118.200 ;
        RECT 120.520 118.140 120.660 118.295 ;
        RECT 120.890 118.280 121.210 118.340 ;
        RECT 125.030 118.280 125.350 118.340 ;
        RECT 134.690 118.280 135.010 118.540 ;
        RECT 135.150 118.280 135.470 118.540 ;
        RECT 136.160 118.525 136.300 118.680 ;
        RECT 136.990 118.620 137.310 118.680 ;
        RECT 137.465 118.635 137.755 118.865 ;
        RECT 138.345 118.820 138.635 118.865 ;
        RECT 139.535 118.820 139.825 118.865 ;
        RECT 142.055 118.820 142.345 118.865 ;
        RECT 138.345 118.680 142.345 118.820 ;
        RECT 138.345 118.635 138.635 118.680 ;
        RECT 139.535 118.635 139.825 118.680 ;
        RECT 142.055 118.635 142.345 118.680 ;
        RECT 136.085 118.295 136.375 118.525 ;
        RECT 136.545 118.480 136.835 118.525 ;
        RECT 140.670 118.480 140.990 118.540 ;
        RECT 136.545 118.340 140.990 118.480 ;
        RECT 136.545 118.295 136.835 118.340 ;
        RECT 140.670 118.280 140.990 118.340 ;
        RECT 119.510 118.000 120.660 118.140 ;
        RECT 121.350 118.140 121.670 118.200 ;
        RECT 122.130 118.140 122.420 118.185 ;
        RECT 138.690 118.140 138.980 118.185 ;
        RECT 121.350 118.000 122.420 118.140 ;
        RECT 119.510 117.940 119.830 118.000 ;
        RECT 121.350 117.940 121.670 118.000 ;
        RECT 122.130 117.955 122.420 118.000 ;
        RECT 132.940 118.000 138.980 118.140 ;
        RECT 127.805 117.800 128.095 117.845 ;
        RECT 129.170 117.800 129.490 117.860 ;
        RECT 132.940 117.845 133.080 118.000 ;
        RECT 138.690 117.955 138.980 118.000 ;
        RECT 119.140 117.660 129.490 117.800 ;
        RECT 102.965 117.615 103.255 117.660 ;
        RECT 103.870 117.600 104.190 117.660 ;
        RECT 127.805 117.615 128.095 117.660 ;
        RECT 129.170 117.600 129.490 117.660 ;
        RECT 132.865 117.615 133.155 117.845 ;
        RECT 135.150 117.800 135.470 117.860 ;
        RECT 143.890 117.800 144.210 117.860 ;
        RECT 144.365 117.800 144.655 117.845 ;
        RECT 135.150 117.660 144.655 117.800 ;
        RECT 135.150 117.600 135.470 117.660 ;
        RECT 143.890 117.600 144.210 117.660 ;
        RECT 144.365 117.615 144.655 117.660 ;
        RECT 17.320 116.980 147.040 117.460 ;
        RECT 22.925 116.780 23.215 116.825 ;
        RECT 25.670 116.780 25.990 116.840 ;
        RECT 22.925 116.640 25.990 116.780 ;
        RECT 22.925 116.595 23.215 116.640 ;
        RECT 25.670 116.580 25.990 116.640 ;
        RECT 102.030 116.580 102.350 116.840 ;
        RECT 115.830 116.580 116.150 116.840 ;
        RECT 126.870 116.580 127.190 116.840 ;
        RECT 128.250 116.780 128.570 116.840 ;
        RECT 128.725 116.780 129.015 116.825 ;
        RECT 128.250 116.640 129.015 116.780 ;
        RECT 128.250 116.580 128.570 116.640 ;
        RECT 128.725 116.595 129.015 116.640 ;
        RECT 131.930 116.780 132.250 116.840 ;
        RECT 131.930 116.640 133.080 116.780 ;
        RECT 131.930 116.580 132.250 116.640 ;
        RECT 96.510 116.485 96.830 116.500 ;
        RECT 28.600 116.440 28.890 116.485 ;
        RECT 30.285 116.440 30.575 116.485 ;
        RECT 96.480 116.440 96.830 116.485 ;
        RECT 28.600 116.300 30.575 116.440 ;
        RECT 96.315 116.300 96.830 116.440 ;
        RECT 28.600 116.255 28.890 116.300 ;
        RECT 30.285 116.255 30.575 116.300 ;
        RECT 96.480 116.255 96.830 116.300 ;
        RECT 96.510 116.240 96.830 116.255 ;
        RECT 20.150 115.900 20.470 116.160 ;
        RECT 26.130 116.100 26.450 116.160 ;
        RECT 29.825 116.100 30.115 116.145 ;
        RECT 26.130 115.960 30.115 116.100 ;
        RECT 26.130 115.900 26.450 115.960 ;
        RECT 29.825 115.915 30.115 115.960 ;
        RECT 31.650 115.900 31.970 116.160 ;
        RECT 33.965 116.100 34.255 116.145 ;
        RECT 35.330 116.100 35.650 116.160 ;
        RECT 33.965 115.960 35.650 116.100 ;
        RECT 33.965 115.915 34.255 115.960 ;
        RECT 35.330 115.900 35.650 115.960 ;
        RECT 86.850 116.100 87.170 116.160 ;
        RECT 88.690 116.100 89.010 116.160 ;
        RECT 86.850 115.960 89.010 116.100 ;
        RECT 86.850 115.900 87.170 115.960 ;
        RECT 88.690 115.900 89.010 115.960 ;
        RECT 89.610 115.900 89.930 116.160 ;
        RECT 102.120 116.100 102.260 116.580 ;
        RECT 102.505 116.440 102.795 116.485 ;
        RECT 104.330 116.440 104.650 116.500 ;
        RECT 102.505 116.300 104.650 116.440 ;
        RECT 102.505 116.255 102.795 116.300 ;
        RECT 104.330 116.240 104.650 116.300 ;
        RECT 118.130 116.440 118.450 116.500 ;
        RECT 120.430 116.440 120.750 116.500 ;
        RECT 121.825 116.440 122.115 116.485 ;
        RECT 118.130 116.300 122.115 116.440 ;
        RECT 118.130 116.240 118.450 116.300 ;
        RECT 120.430 116.240 120.750 116.300 ;
        RECT 121.825 116.255 122.115 116.300 ;
        RECT 125.030 116.440 125.350 116.500 ;
        RECT 125.505 116.440 125.795 116.485 ;
        RECT 132.940 116.440 133.080 116.640 ;
        RECT 144.810 116.580 145.130 116.840 ;
        RECT 133.630 116.440 133.920 116.485 ;
        RECT 125.030 116.300 132.620 116.440 ;
        RECT 132.940 116.300 133.920 116.440 ;
        RECT 125.030 116.240 125.350 116.300 ;
        RECT 125.505 116.255 125.795 116.300 ;
        RECT 103.425 116.100 103.715 116.145 ;
        RECT 102.120 115.960 103.715 116.100 ;
        RECT 103.425 115.915 103.715 115.960 ;
        RECT 103.870 115.900 104.190 116.160 ;
        RECT 114.910 116.100 115.230 116.160 ;
        RECT 129.170 116.100 129.490 116.160 ;
        RECT 132.480 116.145 132.620 116.300 ;
        RECT 133.630 116.255 133.920 116.300 ;
        RECT 134.320 116.300 144.120 116.440 ;
        RECT 114.910 115.960 117.440 116.100 ;
        RECT 114.910 115.900 115.230 115.960 ;
        RECT 25.235 115.760 25.525 115.805 ;
        RECT 27.755 115.760 28.045 115.805 ;
        RECT 28.945 115.760 29.235 115.805 ;
        RECT 25.235 115.620 29.235 115.760 ;
        RECT 25.235 115.575 25.525 115.620 ;
        RECT 27.755 115.575 28.045 115.620 ;
        RECT 28.945 115.575 29.235 115.620 ;
        RECT 31.190 115.760 31.510 115.820 ;
        RECT 32.125 115.760 32.415 115.805 ;
        RECT 31.190 115.620 32.415 115.760 ;
        RECT 31.190 115.560 31.510 115.620 ;
        RECT 32.125 115.575 32.415 115.620 ;
        RECT 32.585 115.760 32.875 115.805 ;
        RECT 34.870 115.760 35.190 115.820 ;
        RECT 32.585 115.620 35.190 115.760 ;
        RECT 32.585 115.575 32.875 115.620 ;
        RECT 34.870 115.560 35.190 115.620 ;
        RECT 87.770 115.760 88.090 115.820 ;
        RECT 93.290 115.760 93.610 115.820 ;
        RECT 95.145 115.760 95.435 115.805 ;
        RECT 87.770 115.620 95.435 115.760 ;
        RECT 87.770 115.560 88.090 115.620 ;
        RECT 93.290 115.560 93.610 115.620 ;
        RECT 95.145 115.575 95.435 115.620 ;
        RECT 96.025 115.760 96.315 115.805 ;
        RECT 97.215 115.760 97.505 115.805 ;
        RECT 99.735 115.760 100.025 115.805 ;
        RECT 96.025 115.620 100.025 115.760 ;
        RECT 96.025 115.575 96.315 115.620 ;
        RECT 97.215 115.575 97.505 115.620 ;
        RECT 99.735 115.575 100.025 115.620 ;
        RECT 116.290 115.560 116.610 115.820 ;
        RECT 117.300 115.805 117.440 115.960 ;
        RECT 129.170 115.960 130.780 116.100 ;
        RECT 129.170 115.900 129.490 115.960 ;
        RECT 117.225 115.760 117.515 115.805 ;
        RECT 130.105 115.760 130.395 115.805 ;
        RECT 117.225 115.620 130.395 115.760 ;
        RECT 130.640 115.760 130.780 115.960 ;
        RECT 132.405 115.915 132.695 116.145 ;
        RECT 134.320 116.100 134.460 116.300 ;
        RECT 143.980 116.145 144.120 116.300 ;
        RECT 142.065 116.100 142.355 116.145 ;
        RECT 132.940 115.960 134.460 116.100 ;
        RECT 139.380 115.960 142.355 116.100 ;
        RECT 132.940 115.760 133.080 115.960 ;
        RECT 130.640 115.620 133.080 115.760 ;
        RECT 133.285 115.760 133.575 115.805 ;
        RECT 134.475 115.760 134.765 115.805 ;
        RECT 136.995 115.760 137.285 115.805 ;
        RECT 133.285 115.620 137.285 115.760 ;
        RECT 117.225 115.575 117.515 115.620 ;
        RECT 130.105 115.575 130.395 115.620 ;
        RECT 133.285 115.575 133.575 115.620 ;
        RECT 134.475 115.575 134.765 115.620 ;
        RECT 136.995 115.575 137.285 115.620 ;
        RECT 25.670 115.420 25.960 115.465 ;
        RECT 27.240 115.420 27.530 115.465 ;
        RECT 29.340 115.420 29.630 115.465 ;
        RECT 33.045 115.420 33.335 115.465 ;
        RECT 25.670 115.280 29.630 115.420 ;
        RECT 25.670 115.235 25.960 115.280 ;
        RECT 27.240 115.235 27.530 115.280 ;
        RECT 29.340 115.235 29.630 115.280 ;
        RECT 31.740 115.280 33.335 115.420 ;
        RECT 19.230 115.080 19.550 115.140 ;
        RECT 20.625 115.080 20.915 115.125 ;
        RECT 26.130 115.080 26.450 115.140 ;
        RECT 19.230 114.940 26.450 115.080 ;
        RECT 19.230 114.880 19.550 114.940 ;
        RECT 20.625 114.895 20.915 114.940 ;
        RECT 26.130 114.880 26.450 114.940 ;
        RECT 29.810 115.080 30.130 115.140 ;
        RECT 31.740 115.080 31.880 115.280 ;
        RECT 33.045 115.235 33.335 115.280 ;
        RECT 95.630 115.420 95.920 115.465 ;
        RECT 97.730 115.420 98.020 115.465 ;
        RECT 99.300 115.420 99.590 115.465 ;
        RECT 95.630 115.280 99.590 115.420 ;
        RECT 95.630 115.235 95.920 115.280 ;
        RECT 97.730 115.235 98.020 115.280 ;
        RECT 99.300 115.235 99.590 115.280 ;
        RECT 103.885 115.235 104.175 115.465 ;
        RECT 130.180 115.420 130.320 115.575 ;
        RECT 139.380 115.480 139.520 115.960 ;
        RECT 142.065 115.915 142.355 115.960 ;
        RECT 143.905 115.915 144.195 116.145 ;
        RECT 132.890 115.420 133.180 115.465 ;
        RECT 134.990 115.420 135.280 115.465 ;
        RECT 136.560 115.420 136.850 115.465 ;
        RECT 138.370 115.420 138.690 115.480 ;
        RECT 113.620 115.280 114.680 115.420 ;
        RECT 130.180 115.280 132.620 115.420 ;
        RECT 29.810 114.940 31.880 115.080 ;
        RECT 101.570 115.080 101.890 115.140 ;
        RECT 103.960 115.080 104.100 115.235 ;
        RECT 113.620 115.080 113.760 115.280 ;
        RECT 101.570 114.940 113.760 115.080 ;
        RECT 29.810 114.880 30.130 114.940 ;
        RECT 101.570 114.880 101.890 114.940 ;
        RECT 113.990 114.880 114.310 115.140 ;
        RECT 114.540 115.080 114.680 115.280 ;
        RECT 131.010 115.080 131.330 115.140 ;
        RECT 114.540 114.940 131.330 115.080 ;
        RECT 132.480 115.080 132.620 115.280 ;
        RECT 132.890 115.280 136.850 115.420 ;
        RECT 132.890 115.235 133.180 115.280 ;
        RECT 134.990 115.235 135.280 115.280 ;
        RECT 136.560 115.235 136.850 115.280 ;
        RECT 137.080 115.280 138.690 115.420 ;
        RECT 137.080 115.080 137.220 115.280 ;
        RECT 138.370 115.220 138.690 115.280 ;
        RECT 139.290 115.220 139.610 115.480 ;
        RECT 142.970 115.220 143.290 115.480 ;
        RECT 132.480 114.940 137.220 115.080 ;
        RECT 131.010 114.880 131.330 114.940 ;
        RECT 17.320 114.260 147.040 114.740 ;
        RECT 28.890 114.060 29.210 114.120 ;
        RECT 35.330 114.060 35.650 114.120 ;
        RECT 28.520 113.920 35.650 114.060 ;
        RECT 28.520 113.765 28.660 113.920 ;
        RECT 28.890 113.860 29.210 113.920 ;
        RECT 35.330 113.860 35.650 113.920 ;
        RECT 91.910 114.060 92.230 114.120 ;
        RECT 105.710 114.060 106.030 114.120 ;
        RECT 108.025 114.060 108.315 114.105 ;
        RECT 91.910 113.920 105.480 114.060 ;
        RECT 91.910 113.860 92.230 113.920 ;
        RECT 19.730 113.720 20.020 113.765 ;
        RECT 21.830 113.720 22.120 113.765 ;
        RECT 23.400 113.720 23.690 113.765 ;
        RECT 19.730 113.580 23.690 113.720 ;
        RECT 19.730 113.535 20.020 113.580 ;
        RECT 21.830 113.535 22.120 113.580 ;
        RECT 23.400 113.535 23.690 113.580 ;
        RECT 28.445 113.535 28.735 113.765 ;
        RECT 31.230 113.720 31.520 113.765 ;
        RECT 33.330 113.720 33.620 113.765 ;
        RECT 34.900 113.720 35.190 113.765 ;
        RECT 31.230 113.580 35.190 113.720 ;
        RECT 31.230 113.535 31.520 113.580 ;
        RECT 33.330 113.535 33.620 113.580 ;
        RECT 34.900 113.535 35.190 113.580 ;
        RECT 88.690 113.520 89.010 113.780 ;
        RECT 105.340 113.765 105.480 113.920 ;
        RECT 105.710 113.920 108.315 114.060 ;
        RECT 105.710 113.860 106.030 113.920 ;
        RECT 108.025 113.875 108.315 113.920 ;
        RECT 115.370 114.060 115.690 114.120 ;
        RECT 131.470 114.060 131.790 114.120 ;
        RECT 132.865 114.060 133.155 114.105 ;
        RECT 115.370 113.920 120.200 114.060 ;
        RECT 115.370 113.860 115.690 113.920 ;
        RECT 120.060 113.780 120.200 113.920 ;
        RECT 131.470 113.920 133.155 114.060 ;
        RECT 131.470 113.860 131.790 113.920 ;
        RECT 132.865 113.875 133.155 113.920 ;
        RECT 133.770 113.860 134.090 114.120 ;
        RECT 93.790 113.720 94.080 113.765 ;
        RECT 95.890 113.720 96.180 113.765 ;
        RECT 97.460 113.720 97.750 113.765 ;
        RECT 93.790 113.580 97.750 113.720 ;
        RECT 93.790 113.535 94.080 113.580 ;
        RECT 95.890 113.535 96.180 113.580 ;
        RECT 97.460 113.535 97.750 113.580 ;
        RECT 100.205 113.720 100.495 113.765 ;
        RECT 100.205 113.580 103.640 113.720 ;
        RECT 100.205 113.535 100.495 113.580 ;
        RECT 19.230 113.180 19.550 113.440 ;
        RECT 20.125 113.380 20.415 113.425 ;
        RECT 21.315 113.380 21.605 113.425 ;
        RECT 23.835 113.380 24.125 113.425 ;
        RECT 20.125 113.240 24.125 113.380 ;
        RECT 20.125 113.195 20.415 113.240 ;
        RECT 21.315 113.195 21.605 113.240 ;
        RECT 23.835 113.195 24.125 113.240 ;
        RECT 31.625 113.380 31.915 113.425 ;
        RECT 32.815 113.380 33.105 113.425 ;
        RECT 35.335 113.380 35.625 113.425 ;
        RECT 31.625 113.240 35.625 113.380 ;
        RECT 31.625 113.195 31.915 113.240 ;
        RECT 32.815 113.195 33.105 113.240 ;
        RECT 35.335 113.195 35.625 113.240 ;
        RECT 93.290 113.180 93.610 113.440 ;
        RECT 94.185 113.380 94.475 113.425 ;
        RECT 95.375 113.380 95.665 113.425 ;
        RECT 97.895 113.380 98.185 113.425 ;
        RECT 94.185 113.240 98.185 113.380 ;
        RECT 94.185 113.195 94.475 113.240 ;
        RECT 95.375 113.195 95.665 113.240 ;
        RECT 97.895 113.195 98.185 113.240 ;
        RECT 26.130 113.040 26.450 113.100 ;
        RECT 30.745 113.040 31.035 113.085 ;
        RECT 26.130 112.900 31.035 113.040 ;
        RECT 26.130 112.840 26.450 112.900 ;
        RECT 30.745 112.855 31.035 112.900 ;
        RECT 92.385 113.040 92.675 113.085 ;
        RECT 93.380 113.040 93.520 113.180 ;
        RECT 92.385 112.900 93.520 113.040 ;
        RECT 94.640 113.040 94.930 113.085 ;
        RECT 99.270 113.040 99.590 113.100 ;
        RECT 94.640 112.900 99.590 113.040 ;
        RECT 92.385 112.855 92.675 112.900 ;
        RECT 94.640 112.855 94.930 112.900 ;
        RECT 99.270 112.840 99.590 112.900 ;
        RECT 100.665 113.040 100.955 113.085 ;
        RECT 102.030 113.040 102.350 113.100 ;
        RECT 103.500 113.085 103.640 113.580 ;
        RECT 105.265 113.535 105.555 113.765 ;
        RECT 114.030 113.720 114.320 113.765 ;
        RECT 116.130 113.720 116.420 113.765 ;
        RECT 117.700 113.720 117.990 113.765 ;
        RECT 114.030 113.580 117.990 113.720 ;
        RECT 114.030 113.535 114.320 113.580 ;
        RECT 116.130 113.535 116.420 113.580 ;
        RECT 117.700 113.535 117.990 113.580 ;
        RECT 119.970 113.720 120.290 113.780 ;
        RECT 141.590 113.720 141.910 113.780 ;
        RECT 119.970 113.580 141.910 113.720 ;
        RECT 119.970 113.520 120.290 113.580 ;
        RECT 108.470 113.380 108.790 113.440 ;
        RECT 114.425 113.380 114.715 113.425 ;
        RECT 115.615 113.380 115.905 113.425 ;
        RECT 118.135 113.380 118.425 113.425 ;
        RECT 108.470 113.240 110.540 113.380 ;
        RECT 108.470 113.180 108.790 113.240 ;
        RECT 100.665 112.900 102.350 113.040 ;
        RECT 100.665 112.855 100.955 112.900 ;
        RECT 102.030 112.840 102.350 112.900 ;
        RECT 103.425 113.040 103.715 113.085 ;
        RECT 103.870 113.040 104.190 113.100 ;
        RECT 103.425 112.900 104.190 113.040 ;
        RECT 103.425 112.855 103.715 112.900 ;
        RECT 103.870 112.840 104.190 112.900 ;
        RECT 104.330 113.040 104.650 113.100 ;
        RECT 110.400 113.085 110.540 113.240 ;
        RECT 114.425 113.240 118.425 113.380 ;
        RECT 114.425 113.195 114.715 113.240 ;
        RECT 115.615 113.195 115.905 113.240 ;
        RECT 118.135 113.195 118.425 113.240 ;
        RECT 108.945 113.040 109.235 113.085 ;
        RECT 104.330 112.900 109.235 113.040 ;
        RECT 104.330 112.840 104.650 112.900 ;
        RECT 108.945 112.855 109.235 112.900 ;
        RECT 109.405 112.855 109.695 113.085 ;
        RECT 110.325 112.855 110.615 113.085 ;
        RECT 20.580 112.700 20.870 112.745 ;
        RECT 21.530 112.700 21.850 112.760 ;
        RECT 20.580 112.560 21.850 112.700 ;
        RECT 20.580 112.515 20.870 112.560 ;
        RECT 21.530 112.500 21.850 112.560 ;
        RECT 29.810 112.500 30.130 112.760 ;
        RECT 32.110 112.745 32.430 112.760 ;
        RECT 31.970 112.700 32.430 112.745 ;
        RECT 30.360 112.560 32.430 112.700 ;
        RECT 21.990 112.360 22.310 112.420 ;
        RECT 26.145 112.360 26.435 112.405 ;
        RECT 21.990 112.220 26.435 112.360 ;
        RECT 21.990 112.160 22.310 112.220 ;
        RECT 26.145 112.175 26.435 112.220 ;
        RECT 27.510 112.360 27.830 112.420 ;
        RECT 30.360 112.360 30.500 112.560 ;
        RECT 31.970 112.515 32.430 112.560 ;
        RECT 32.110 112.500 32.430 112.515 ;
        RECT 85.930 112.700 86.250 112.760 ;
        RECT 86.865 112.700 87.155 112.745 ;
        RECT 106.185 112.700 106.475 112.745 ;
        RECT 85.930 112.560 87.155 112.700 ;
        RECT 85.930 112.500 86.250 112.560 ;
        RECT 86.865 112.515 87.155 112.560 ;
        RECT 104.420 112.560 106.475 112.700 ;
        RECT 109.480 112.700 109.620 112.855 ;
        RECT 110.770 112.840 111.090 113.100 ;
        RECT 113.530 112.840 113.850 113.100 ;
        RECT 116.290 113.040 116.610 113.100 ;
        RECT 114.540 112.900 116.610 113.040 ;
        RECT 114.540 112.700 114.680 112.900 ;
        RECT 116.290 112.840 116.610 112.900 ;
        RECT 120.430 113.040 120.750 113.100 ;
        RECT 120.905 113.040 121.195 113.085 ;
        RECT 120.430 112.900 121.195 113.040 ;
        RECT 120.430 112.840 120.750 112.900 ;
        RECT 120.905 112.855 121.195 112.900 ;
        RECT 129.170 113.040 129.490 113.100 ;
        RECT 130.550 113.085 130.870 113.100 ;
        RECT 129.645 113.040 129.935 113.085 ;
        RECT 129.170 112.900 129.935 113.040 ;
        RECT 129.170 112.840 129.490 112.900 ;
        RECT 129.645 112.855 129.935 112.900 ;
        RECT 130.385 112.855 130.870 113.085 ;
        RECT 131.970 113.040 132.260 113.085 ;
        RECT 132.480 113.040 132.620 113.580 ;
        RECT 141.590 113.520 141.910 113.580 ;
        RECT 133.310 113.380 133.630 113.440 ;
        RECT 133.310 113.240 135.840 113.380 ;
        RECT 133.310 113.180 133.630 113.240 ;
        RECT 135.700 113.085 135.840 113.240 ;
        RECT 136.070 113.180 136.390 113.440 ;
        RECT 137.005 113.380 137.295 113.425 ;
        RECT 139.750 113.380 140.070 113.440 ;
        RECT 137.005 113.240 140.070 113.380 ;
        RECT 137.005 113.195 137.295 113.240 ;
        RECT 139.750 113.180 140.070 113.240 ;
        RECT 131.970 112.900 132.620 113.040 ;
        RECT 131.970 112.855 132.260 112.900 ;
        RECT 135.625 112.855 135.915 113.085 ;
        RECT 136.160 113.040 136.300 113.180 ;
        RECT 142.065 113.040 142.355 113.085 ;
        RECT 136.160 112.900 142.355 113.040 ;
        RECT 142.065 112.855 142.355 112.900 ;
        RECT 130.550 112.840 130.870 112.855 ;
        RECT 143.890 112.840 144.210 113.100 ;
        RECT 114.910 112.745 115.230 112.760 ;
        RECT 109.480 112.560 114.680 112.700 ;
        RECT 27.510 112.220 30.500 112.360 ;
        RECT 34.870 112.360 35.190 112.420 ;
        RECT 37.645 112.360 37.935 112.405 ;
        RECT 34.870 112.220 37.935 112.360 ;
        RECT 27.510 112.160 27.830 112.220 ;
        RECT 34.870 112.160 35.190 112.220 ;
        RECT 37.645 112.175 37.935 112.220 ;
        RECT 88.230 112.360 88.550 112.420 ;
        RECT 104.420 112.405 104.560 112.560 ;
        RECT 106.185 112.515 106.475 112.560 ;
        RECT 114.880 112.515 115.230 112.745 ;
        RECT 89.165 112.360 89.455 112.405 ;
        RECT 88.230 112.220 89.455 112.360 ;
        RECT 88.230 112.160 88.550 112.220 ;
        RECT 89.165 112.175 89.455 112.220 ;
        RECT 104.345 112.175 104.635 112.405 ;
        RECT 106.260 112.360 106.400 112.515 ;
        RECT 114.910 112.500 115.230 112.515 ;
        RECT 115.370 112.360 115.690 112.420 ;
        RECT 106.260 112.220 115.690 112.360 ;
        RECT 116.380 112.360 116.520 112.840 ;
        RECT 124.570 112.500 124.890 112.760 ;
        RECT 131.010 112.500 131.330 112.760 ;
        RECT 131.485 112.700 131.775 112.745 ;
        RECT 136.085 112.700 136.375 112.745 ;
        RECT 139.290 112.700 139.610 112.760 ;
        RECT 131.485 112.560 139.610 112.700 ;
        RECT 131.485 112.515 131.775 112.560 ;
        RECT 136.085 112.515 136.375 112.560 ;
        RECT 139.290 112.500 139.610 112.560 ;
        RECT 120.445 112.360 120.735 112.405 ;
        RECT 129.630 112.360 129.950 112.420 ;
        RECT 116.380 112.220 129.950 112.360 ;
        RECT 131.100 112.360 131.240 112.500 ;
        RECT 142.510 112.360 142.830 112.420 ;
        RECT 131.100 112.220 142.830 112.360 ;
        RECT 115.370 112.160 115.690 112.220 ;
        RECT 120.445 112.175 120.735 112.220 ;
        RECT 129.630 112.160 129.950 112.220 ;
        RECT 142.510 112.160 142.830 112.220 ;
        RECT 142.970 112.160 143.290 112.420 ;
        RECT 144.810 112.160 145.130 112.420 ;
        RECT 17.320 111.540 147.040 112.020 ;
        RECT 20.150 111.340 20.470 111.400 ;
        RECT 21.085 111.340 21.375 111.385 ;
        RECT 20.150 111.200 21.375 111.340 ;
        RECT 20.150 111.140 20.470 111.200 ;
        RECT 21.085 111.155 21.375 111.200 ;
        RECT 21.530 111.140 21.850 111.400 ;
        RECT 21.990 111.340 22.310 111.400 ;
        RECT 23.385 111.340 23.675 111.385 ;
        RECT 21.990 111.200 23.675 111.340 ;
        RECT 21.990 111.140 22.310 111.200 ;
        RECT 23.385 111.155 23.675 111.200 ;
        RECT 23.845 111.340 24.135 111.385 ;
        RECT 24.290 111.340 24.610 111.400 ;
        RECT 23.845 111.200 24.610 111.340 ;
        RECT 23.845 111.155 24.135 111.200 ;
        RECT 24.290 111.140 24.610 111.200 ;
        RECT 33.045 111.155 33.335 111.385 ;
        RECT 33.120 111.000 33.260 111.155 ;
        RECT 35.790 111.140 36.110 111.400 ;
        RECT 79.965 111.340 80.255 111.385 ;
        RECT 80.410 111.340 80.730 111.400 ;
        RECT 86.390 111.340 86.710 111.400 ;
        RECT 90.070 111.340 90.390 111.400 ;
        RECT 101.570 111.340 101.890 111.400 ;
        RECT 79.965 111.200 90.390 111.340 ;
        RECT 79.965 111.155 80.255 111.200 ;
        RECT 80.410 111.140 80.730 111.200 ;
        RECT 86.390 111.140 86.710 111.200 ;
        RECT 90.070 111.140 90.390 111.200 ;
        RECT 97.520 111.200 101.890 111.340 ;
        RECT 33.505 111.000 33.795 111.045 ;
        RECT 35.330 111.000 35.650 111.060 ;
        RECT 33.120 110.860 35.650 111.000 ;
        RECT 33.505 110.815 33.795 110.860 ;
        RECT 35.330 110.800 35.650 110.860 ;
        RECT 16.010 110.660 16.330 110.720 ;
        RECT 18.785 110.660 19.075 110.705 ;
        RECT 16.010 110.520 19.075 110.660 ;
        RECT 16.010 110.460 16.330 110.520 ;
        RECT 18.785 110.475 19.075 110.520 ;
        RECT 20.150 110.460 20.470 110.720 ;
        RECT 26.590 110.660 26.910 110.720 ;
        RECT 27.480 110.660 27.770 110.705 ;
        RECT 29.350 110.660 29.670 110.720 ;
        RECT 24.840 110.520 29.670 110.660 ;
        RECT 24.840 110.365 24.980 110.520 ;
        RECT 26.590 110.460 26.910 110.520 ;
        RECT 27.480 110.475 27.770 110.520 ;
        RECT 29.350 110.460 29.670 110.520 ;
        RECT 30.270 110.660 30.590 110.720 ;
        RECT 35.880 110.660 36.020 111.140 ;
        RECT 83.630 111.000 83.950 111.060 ;
        RECT 83.630 110.860 92.140 111.000 ;
        RECT 83.630 110.800 83.950 110.860 ;
        RECT 92.000 110.720 92.140 110.860 ;
        RECT 30.270 110.520 36.020 110.660 ;
        RECT 79.030 110.660 79.350 110.720 ;
        RECT 86.865 110.660 87.155 110.705 ;
        RECT 89.150 110.660 89.470 110.720 ;
        RECT 79.030 110.520 81.100 110.660 ;
        RECT 30.270 110.460 30.590 110.520 ;
        RECT 79.030 110.460 79.350 110.520 ;
        RECT 24.765 110.135 25.055 110.365 ;
        RECT 26.130 110.120 26.450 110.380 ;
        RECT 27.025 110.320 27.315 110.365 ;
        RECT 28.215 110.320 28.505 110.365 ;
        RECT 30.735 110.320 31.025 110.365 ;
        RECT 27.025 110.180 31.025 110.320 ;
        RECT 27.025 110.135 27.315 110.180 ;
        RECT 28.215 110.135 28.505 110.180 ;
        RECT 30.735 110.135 31.025 110.180 ;
        RECT 34.410 110.320 34.730 110.380 ;
        RECT 35.330 110.320 35.650 110.380 ;
        RECT 34.410 110.180 35.650 110.320 ;
        RECT 34.410 110.120 34.730 110.180 ;
        RECT 35.330 110.120 35.650 110.180 ;
        RECT 73.970 110.120 74.290 110.380 ;
        RECT 80.960 110.365 81.100 110.520 ;
        RECT 86.865 110.520 89.470 110.660 ;
        RECT 86.865 110.475 87.155 110.520 ;
        RECT 89.150 110.460 89.470 110.520 ;
        RECT 91.910 110.460 92.230 110.720 ;
        RECT 93.750 110.460 94.070 110.720 ;
        RECT 97.520 110.705 97.660 111.200 ;
        RECT 101.570 111.140 101.890 111.200 ;
        RECT 105.250 111.340 105.570 111.400 ;
        RECT 109.405 111.340 109.695 111.385 ;
        RECT 105.250 111.200 114.680 111.340 ;
        RECT 105.250 111.140 105.570 111.200 ;
        RECT 109.405 111.155 109.695 111.200 ;
        RECT 100.665 110.815 100.955 111.045 ;
        RECT 104.330 111.000 104.650 111.060 ;
        RECT 106.185 111.000 106.475 111.045 ;
        RECT 102.120 110.860 104.100 111.000 ;
        RECT 97.445 110.475 97.735 110.705 ;
        RECT 98.365 110.475 98.655 110.705 ;
        RECT 100.205 110.475 100.495 110.705 ;
        RECT 100.740 110.660 100.880 110.815 ;
        RECT 101.570 110.660 101.890 110.720 ;
        RECT 102.120 110.705 102.260 110.860 ;
        RECT 103.960 110.720 104.100 110.860 ;
        RECT 104.330 110.860 106.475 111.000 ;
        RECT 104.330 110.800 104.650 110.860 ;
        RECT 106.185 110.815 106.475 110.860 ;
        RECT 108.930 111.000 109.250 111.060 ;
        RECT 112.625 111.000 112.915 111.045 ;
        RECT 108.930 110.860 112.915 111.000 ;
        RECT 114.540 111.000 114.680 111.200 ;
        RECT 114.910 111.140 115.230 111.400 ;
        RECT 128.265 111.340 128.555 111.385 ;
        RECT 130.550 111.340 130.870 111.400 ;
        RECT 131.025 111.340 131.315 111.385 ;
        RECT 136.070 111.340 136.390 111.400 ;
        RECT 128.265 111.200 136.390 111.340 ;
        RECT 128.265 111.155 128.555 111.200 ;
        RECT 130.550 111.140 130.870 111.200 ;
        RECT 131.025 111.155 131.315 111.200 ;
        RECT 136.070 111.140 136.390 111.200 ;
        RECT 137.005 111.155 137.295 111.385 ;
        RECT 122.700 111.000 122.990 111.045 ;
        RECT 123.650 111.000 123.970 111.060 ;
        RECT 114.540 110.860 122.270 111.000 ;
        RECT 108.930 110.800 109.250 110.860 ;
        RECT 112.625 110.815 112.915 110.860 ;
        RECT 100.740 110.520 101.890 110.660 ;
        RECT 80.425 110.135 80.715 110.365 ;
        RECT 80.885 110.135 81.175 110.365 ;
        RECT 85.470 110.320 85.790 110.380 ;
        RECT 87.325 110.320 87.615 110.365 ;
        RECT 95.130 110.320 95.450 110.380 ;
        RECT 85.470 110.180 95.450 110.320 ;
        RECT 19.705 109.980 19.995 110.025 ;
        RECT 26.630 109.980 26.920 110.025 ;
        RECT 28.730 109.980 29.020 110.025 ;
        RECT 30.300 109.980 30.590 110.025 ;
        RECT 34.870 109.980 35.190 110.040 ;
        RECT 19.705 109.840 25.670 109.980 ;
        RECT 19.705 109.795 19.995 109.840 ;
        RECT 25.530 109.640 25.670 109.840 ;
        RECT 26.630 109.840 30.590 109.980 ;
        RECT 26.630 109.795 26.920 109.840 ;
        RECT 28.730 109.795 29.020 109.840 ;
        RECT 30.300 109.795 30.590 109.840 ;
        RECT 32.660 109.840 35.190 109.980 ;
        RECT 27.970 109.640 28.290 109.700 ;
        RECT 25.530 109.500 28.290 109.640 ;
        RECT 27.970 109.440 28.290 109.500 ;
        RECT 29.810 109.640 30.130 109.700 ;
        RECT 32.660 109.640 32.800 109.840 ;
        RECT 34.870 109.780 35.190 109.840 ;
        RECT 75.825 109.980 76.115 110.025 ;
        RECT 78.125 109.980 78.415 110.025 ;
        RECT 75.825 109.840 78.415 109.980 ;
        RECT 75.825 109.795 76.115 109.840 ;
        RECT 78.125 109.795 78.415 109.840 ;
        RECT 79.950 109.980 80.270 110.040 ;
        RECT 80.500 109.980 80.640 110.135 ;
        RECT 85.470 110.120 85.790 110.180 ;
        RECT 87.325 110.135 87.615 110.180 ;
        RECT 95.130 110.120 95.450 110.180 ;
        RECT 79.950 109.840 80.640 109.980 ;
        RECT 87.770 109.980 88.090 110.040 ;
        RECT 91.005 109.980 91.295 110.025 ;
        RECT 98.440 109.980 98.580 110.475 ;
        RECT 100.280 110.320 100.420 110.475 ;
        RECT 101.570 110.460 101.890 110.520 ;
        RECT 102.045 110.475 102.335 110.705 ;
        RECT 102.490 110.660 102.810 110.720 ;
        RECT 103.425 110.660 103.715 110.705 ;
        RECT 102.490 110.520 103.715 110.660 ;
        RECT 102.490 110.460 102.810 110.520 ;
        RECT 103.425 110.475 103.715 110.520 ;
        RECT 103.870 110.460 104.190 110.720 ;
        RECT 120.890 110.660 121.210 110.720 ;
        RECT 121.365 110.660 121.655 110.705 ;
        RECT 120.890 110.520 121.655 110.660 ;
        RECT 122.130 110.660 122.270 110.860 ;
        RECT 122.700 110.860 123.970 111.000 ;
        RECT 122.700 110.815 122.990 110.860 ;
        RECT 123.650 110.800 123.970 110.860 ;
        RECT 134.230 111.000 134.550 111.060 ;
        RECT 134.705 111.000 134.995 111.045 ;
        RECT 134.230 110.860 134.995 111.000 ;
        RECT 137.080 111.000 137.220 111.155 ;
        RECT 138.690 111.000 138.980 111.045 ;
        RECT 137.080 110.860 138.980 111.000 ;
        RECT 134.230 110.800 134.550 110.860 ;
        RECT 134.705 110.815 134.995 110.860 ;
        RECT 138.690 110.815 138.980 110.860 ;
        RECT 130.565 110.660 130.855 110.705 ;
        RECT 133.310 110.660 133.630 110.720 ;
        RECT 122.130 110.520 133.630 110.660 ;
        RECT 120.890 110.460 121.210 110.520 ;
        RECT 121.365 110.475 121.655 110.520 ;
        RECT 130.565 110.475 130.855 110.520 ;
        RECT 133.310 110.460 133.630 110.520 ;
        RECT 102.580 110.320 102.720 110.460 ;
        RECT 100.280 110.180 102.720 110.320 ;
        RECT 105.250 110.320 105.570 110.380 ;
        RECT 105.725 110.320 106.015 110.365 ;
        RECT 105.250 110.180 106.015 110.320 ;
        RECT 105.250 110.120 105.570 110.180 ;
        RECT 105.725 110.135 106.015 110.180 ;
        RECT 106.170 110.320 106.490 110.380 ;
        RECT 108.485 110.320 108.775 110.365 ;
        RECT 106.170 110.180 108.775 110.320 ;
        RECT 106.170 110.120 106.490 110.180 ;
        RECT 108.485 110.135 108.775 110.180 ;
        RECT 108.930 110.120 109.250 110.380 ;
        RECT 122.245 110.320 122.535 110.365 ;
        RECT 123.435 110.320 123.725 110.365 ;
        RECT 125.955 110.320 126.245 110.365 ;
        RECT 122.245 110.180 126.245 110.320 ;
        RECT 122.245 110.135 122.535 110.180 ;
        RECT 123.435 110.135 123.725 110.180 ;
        RECT 125.955 110.135 126.245 110.180 ;
        RECT 131.945 110.320 132.235 110.365 ;
        RECT 132.850 110.320 133.170 110.380 ;
        RECT 131.945 110.180 133.170 110.320 ;
        RECT 131.945 110.135 132.235 110.180 ;
        RECT 132.850 110.120 133.170 110.180 ;
        RECT 136.070 110.320 136.390 110.380 ;
        RECT 137.465 110.320 137.755 110.365 ;
        RECT 136.070 110.180 137.755 110.320 ;
        RECT 136.070 110.120 136.390 110.180 ;
        RECT 137.465 110.135 137.755 110.180 ;
        RECT 138.345 110.320 138.635 110.365 ;
        RECT 139.535 110.320 139.825 110.365 ;
        RECT 142.055 110.320 142.345 110.365 ;
        RECT 138.345 110.180 142.345 110.320 ;
        RECT 138.345 110.135 138.635 110.180 ;
        RECT 139.535 110.135 139.825 110.180 ;
        RECT 142.055 110.135 142.345 110.180 ;
        RECT 104.330 109.980 104.650 110.040 ;
        RECT 87.770 109.840 97.200 109.980 ;
        RECT 98.440 109.840 104.650 109.980 ;
        RECT 79.950 109.780 80.270 109.840 ;
        RECT 87.770 109.780 88.090 109.840 ;
        RECT 91.005 109.795 91.295 109.840 ;
        RECT 29.810 109.500 32.800 109.640 ;
        RECT 29.810 109.440 30.130 109.500 ;
        RECT 76.270 109.440 76.590 109.700 ;
        RECT 84.090 109.640 84.410 109.700 ;
        RECT 84.565 109.640 84.855 109.685 ;
        RECT 84.090 109.500 84.855 109.640 ;
        RECT 84.090 109.440 84.410 109.500 ;
        RECT 84.565 109.455 84.855 109.500 ;
        RECT 96.510 109.440 96.830 109.700 ;
        RECT 97.060 109.640 97.200 109.840 ;
        RECT 104.330 109.780 104.650 109.840 ;
        RECT 104.880 109.840 111.920 109.980 ;
        RECT 104.880 109.640 105.020 109.840 ;
        RECT 97.060 109.500 105.020 109.640 ;
        RECT 109.850 109.640 110.170 109.700 ;
        RECT 111.245 109.640 111.535 109.685 ;
        RECT 109.850 109.500 111.535 109.640 ;
        RECT 111.780 109.640 111.920 109.840 ;
        RECT 113.990 109.780 114.310 110.040 ;
        RECT 121.850 109.980 122.140 110.025 ;
        RECT 123.950 109.980 124.240 110.025 ;
        RECT 125.520 109.980 125.810 110.025 ;
        RECT 121.850 109.840 125.810 109.980 ;
        RECT 121.850 109.795 122.140 109.840 ;
        RECT 123.950 109.795 124.240 109.840 ;
        RECT 125.520 109.795 125.810 109.840 ;
        RECT 128.340 109.840 129.400 109.980 ;
        RECT 119.050 109.640 119.370 109.700 ;
        RECT 128.340 109.640 128.480 109.840 ;
        RECT 111.780 109.500 128.480 109.640 ;
        RECT 109.850 109.440 110.170 109.500 ;
        RECT 111.245 109.455 111.535 109.500 ;
        RECT 119.050 109.440 119.370 109.500 ;
        RECT 128.710 109.440 129.030 109.700 ;
        RECT 129.260 109.640 129.400 109.840 ;
        RECT 136.530 109.780 136.850 110.040 ;
        RECT 137.950 109.980 138.240 110.025 ;
        RECT 140.050 109.980 140.340 110.025 ;
        RECT 141.620 109.980 141.910 110.025 ;
        RECT 137.950 109.840 141.910 109.980 ;
        RECT 137.950 109.795 138.240 109.840 ;
        RECT 140.050 109.795 140.340 109.840 ;
        RECT 141.620 109.795 141.910 109.840 ;
        RECT 139.290 109.640 139.610 109.700 ;
        RECT 129.260 109.500 139.610 109.640 ;
        RECT 139.290 109.440 139.610 109.500 ;
        RECT 144.350 109.440 144.670 109.700 ;
        RECT 17.320 108.820 147.040 109.300 ;
        RECT 88.690 108.620 89.010 108.680 ;
        RECT 90.545 108.620 90.835 108.665 ;
        RECT 88.690 108.480 90.835 108.620 ;
        RECT 88.690 108.420 89.010 108.480 ;
        RECT 90.545 108.435 90.835 108.480 ;
        RECT 95.130 108.620 95.450 108.680 ;
        RECT 106.170 108.620 106.490 108.680 ;
        RECT 95.130 108.480 106.490 108.620 ;
        RECT 95.130 108.420 95.450 108.480 ;
        RECT 106.170 108.420 106.490 108.480 ;
        RECT 113.530 108.620 113.850 108.680 ;
        RECT 113.530 108.480 115.140 108.620 ;
        RECT 113.530 108.420 113.850 108.480 ;
        RECT 72.605 108.095 72.895 108.325 ;
        RECT 74.470 108.280 74.760 108.325 ;
        RECT 76.570 108.280 76.860 108.325 ;
        RECT 78.140 108.280 78.430 108.325 ;
        RECT 74.470 108.140 78.430 108.280 ;
        RECT 74.470 108.095 74.760 108.140 ;
        RECT 76.570 108.095 76.860 108.140 ;
        RECT 78.140 108.095 78.430 108.140 ;
        RECT 82.750 108.280 83.040 108.325 ;
        RECT 84.850 108.280 85.140 108.325 ;
        RECT 86.420 108.280 86.710 108.325 ;
        RECT 82.750 108.140 86.710 108.280 ;
        RECT 82.750 108.095 83.040 108.140 ;
        RECT 84.850 108.095 85.140 108.140 ;
        RECT 86.420 108.095 86.710 108.140 ;
        RECT 93.750 108.280 94.070 108.340 ;
        RECT 95.590 108.280 95.910 108.340 ;
        RECT 110.770 108.280 111.060 108.325 ;
        RECT 112.340 108.280 112.630 108.325 ;
        RECT 114.440 108.280 114.730 108.325 ;
        RECT 93.750 108.140 97.200 108.280 ;
        RECT 72.680 107.940 72.820 108.095 ;
        RECT 93.750 108.080 94.070 108.140 ;
        RECT 95.590 108.080 95.910 108.140 ;
        RECT 73.050 107.940 73.370 108.000 ;
        RECT 72.680 107.800 73.370 107.940 ;
        RECT 73.050 107.740 73.370 107.800 ;
        RECT 74.865 107.940 75.155 107.985 ;
        RECT 76.055 107.940 76.345 107.985 ;
        RECT 78.575 107.940 78.865 107.985 ;
        RECT 74.865 107.800 78.865 107.940 ;
        RECT 74.865 107.755 75.155 107.800 ;
        RECT 76.055 107.755 76.345 107.800 ;
        RECT 78.575 107.755 78.865 107.800 ;
        RECT 83.145 107.940 83.435 107.985 ;
        RECT 84.335 107.940 84.625 107.985 ;
        RECT 86.855 107.940 87.145 107.985 ;
        RECT 83.145 107.800 87.145 107.940 ;
        RECT 83.145 107.755 83.435 107.800 ;
        RECT 84.335 107.755 84.625 107.800 ;
        RECT 86.855 107.755 87.145 107.800 ;
        RECT 93.305 107.940 93.595 107.985 ;
        RECT 95.130 107.940 95.450 108.000 ;
        RECT 93.305 107.800 95.450 107.940 ;
        RECT 93.305 107.755 93.595 107.800 ;
        RECT 95.130 107.740 95.450 107.800 ;
        RECT 28.890 107.400 29.210 107.660 ;
        RECT 29.810 107.400 30.130 107.660 ;
        RECT 73.985 107.600 74.275 107.645 ;
        RECT 80.870 107.600 81.190 107.660 ;
        RECT 82.265 107.600 82.555 107.645 ;
        RECT 86.390 107.600 86.710 107.660 ;
        RECT 73.985 107.460 86.710 107.600 ;
        RECT 73.985 107.415 74.275 107.460 ;
        RECT 80.870 107.400 81.190 107.460 ;
        RECT 82.265 107.415 82.555 107.460 ;
        RECT 86.390 107.400 86.710 107.460 ;
        RECT 89.610 107.600 89.930 107.660 ;
        RECT 94.685 107.600 94.975 107.645 ;
        RECT 89.610 107.460 94.975 107.600 ;
        RECT 97.060 107.600 97.200 108.140 ;
        RECT 110.770 108.140 114.730 108.280 ;
        RECT 110.770 108.095 111.060 108.140 ;
        RECT 112.340 108.095 112.630 108.140 ;
        RECT 114.440 108.095 114.730 108.140 ;
        RECT 106.185 107.940 106.475 107.985 ;
        RECT 108.470 107.940 108.790 108.000 ;
        RECT 115.000 107.985 115.140 108.480 ;
        RECT 123.650 108.420 123.970 108.680 ;
        RECT 128.710 108.620 129.030 108.680 ;
        RECT 124.200 108.480 129.030 108.620 ;
        RECT 123.205 108.280 123.495 108.325 ;
        RECT 124.200 108.280 124.340 108.480 ;
        RECT 128.710 108.420 129.030 108.480 ;
        RECT 136.530 108.420 136.850 108.680 ;
        RECT 123.205 108.140 124.340 108.280 ;
        RECT 123.205 108.095 123.495 108.140 ;
        RECT 125.030 108.080 125.350 108.340 ;
        RECT 136.070 108.280 136.390 108.340 ;
        RECT 125.580 108.140 136.390 108.280 ;
        RECT 100.740 107.800 108.790 107.940 ;
        RECT 100.740 107.660 100.880 107.800 ;
        RECT 106.185 107.755 106.475 107.800 ;
        RECT 108.470 107.740 108.790 107.800 ;
        RECT 110.335 107.940 110.625 107.985 ;
        RECT 112.855 107.940 113.145 107.985 ;
        RECT 114.045 107.940 114.335 107.985 ;
        RECT 110.335 107.800 114.335 107.940 ;
        RECT 110.335 107.755 110.625 107.800 ;
        RECT 112.855 107.755 113.145 107.800 ;
        RECT 114.045 107.755 114.335 107.800 ;
        RECT 114.925 107.940 115.215 107.985 ;
        RECT 122.270 107.940 122.590 108.000 ;
        RECT 124.570 107.940 124.890 108.000 ;
        RECT 125.580 107.940 125.720 108.140 ;
        RECT 136.070 108.080 136.390 108.140 ;
        RECT 114.925 107.800 125.720 107.940 ;
        RECT 114.925 107.755 115.215 107.800 ;
        RECT 122.270 107.740 122.590 107.800 ;
        RECT 124.570 107.740 124.890 107.800 ;
        RECT 126.410 107.740 126.730 108.000 ;
        RECT 139.750 107.740 140.070 108.000 ;
        RECT 144.350 107.940 144.670 108.000 ;
        RECT 142.140 107.800 144.670 107.940 ;
        RECT 97.445 107.600 97.735 107.645 ;
        RECT 98.825 107.600 99.115 107.645 ;
        RECT 97.060 107.460 99.115 107.600 ;
        RECT 89.610 107.400 89.930 107.460 ;
        RECT 94.685 107.415 94.975 107.460 ;
        RECT 97.445 107.415 97.735 107.460 ;
        RECT 98.825 107.415 99.115 107.460 ;
        RECT 100.650 107.400 100.970 107.660 ;
        RECT 101.110 107.400 101.430 107.660 ;
        RECT 104.790 107.600 105.110 107.660 ;
        RECT 105.265 107.600 105.555 107.645 ;
        RECT 104.790 107.460 105.555 107.600 ;
        RECT 104.790 107.400 105.110 107.460 ;
        RECT 105.265 107.415 105.555 107.460 ;
        RECT 105.725 107.600 106.015 107.645 ;
        RECT 108.010 107.600 108.330 107.660 ;
        RECT 105.725 107.460 108.330 107.600 ;
        RECT 105.725 107.415 106.015 107.460 ;
        RECT 108.010 107.400 108.330 107.460 ;
        RECT 121.365 107.600 121.655 107.645 ;
        RECT 131.470 107.600 131.790 107.660 ;
        RECT 134.230 107.600 134.550 107.660 ;
        RECT 121.365 107.460 134.550 107.600 ;
        RECT 121.365 107.415 121.655 107.460 ;
        RECT 131.470 107.400 131.790 107.460 ;
        RECT 134.230 107.400 134.550 107.460 ;
        RECT 137.450 107.600 137.770 107.660 ;
        RECT 141.590 107.645 141.910 107.660 ;
        RECT 142.140 107.645 142.280 107.800 ;
        RECT 144.350 107.740 144.670 107.800 ;
        RECT 138.385 107.600 138.675 107.645 ;
        RECT 141.580 107.600 141.910 107.645 ;
        RECT 137.450 107.460 138.675 107.600 ;
        RECT 141.395 107.460 141.910 107.600 ;
        RECT 137.450 107.400 137.770 107.460 ;
        RECT 138.385 107.415 138.675 107.460 ;
        RECT 141.580 107.415 141.910 107.460 ;
        RECT 142.065 107.415 142.355 107.645 ;
        RECT 141.590 107.400 141.910 107.415 ;
        RECT 71.225 107.260 71.515 107.305 ;
        RECT 75.320 107.260 75.610 107.305 ;
        RECT 76.270 107.260 76.590 107.320 ;
        RECT 71.225 107.120 74.200 107.260 ;
        RECT 71.225 107.075 71.515 107.120 ;
        RECT 74.060 106.980 74.200 107.120 ;
        RECT 75.320 107.120 76.590 107.260 ;
        RECT 75.320 107.075 75.610 107.120 ;
        RECT 76.270 107.060 76.590 107.120 ;
        RECT 83.600 107.260 83.890 107.305 ;
        RECT 84.550 107.260 84.870 107.320 ;
        RECT 101.200 107.260 101.340 107.400 ;
        RECT 83.600 107.120 84.870 107.260 ;
        RECT 83.600 107.075 83.890 107.120 ;
        RECT 84.550 107.060 84.870 107.120 ;
        RECT 87.400 107.120 101.340 107.260 ;
        RECT 110.310 107.260 110.630 107.320 ;
        RECT 113.590 107.260 113.880 107.305 ;
        RECT 110.310 107.120 113.880 107.260 ;
        RECT 28.890 106.920 29.210 106.980 ;
        RECT 29.365 106.920 29.655 106.965 ;
        RECT 28.890 106.780 29.655 106.920 ;
        RECT 28.890 106.720 29.210 106.780 ;
        RECT 29.365 106.735 29.655 106.780 ;
        RECT 73.510 106.720 73.830 106.980 ;
        RECT 73.970 106.720 74.290 106.980 ;
        RECT 79.950 106.920 80.270 106.980 ;
        RECT 80.885 106.920 81.175 106.965 ;
        RECT 79.950 106.780 81.175 106.920 ;
        RECT 79.950 106.720 80.270 106.780 ;
        RECT 80.885 106.735 81.175 106.780 ;
        RECT 85.010 106.920 85.330 106.980 ;
        RECT 87.400 106.920 87.540 107.120 ;
        RECT 110.310 107.060 110.630 107.120 ;
        RECT 113.590 107.075 113.880 107.120 ;
        RECT 138.845 107.260 139.135 107.305 ;
        RECT 142.140 107.260 142.280 107.415 ;
        RECT 142.510 107.400 142.830 107.660 ;
        RECT 143.430 107.600 143.750 107.660 ;
        RECT 143.235 107.460 143.750 107.600 ;
        RECT 143.430 107.400 143.750 107.460 ;
        RECT 143.905 107.415 144.195 107.645 ;
        RECT 138.845 107.120 142.280 107.260 ;
        RECT 138.845 107.075 139.135 107.120 ;
        RECT 85.010 106.780 87.540 106.920 ;
        RECT 85.010 106.720 85.330 106.780 ;
        RECT 89.150 106.720 89.470 106.980 ;
        RECT 90.070 106.920 90.390 106.980 ;
        RECT 92.385 106.920 92.675 106.965 ;
        RECT 90.070 106.780 92.675 106.920 ;
        RECT 90.070 106.720 90.390 106.780 ;
        RECT 92.385 106.735 92.675 106.780 ;
        RECT 92.845 106.920 93.135 106.965 ;
        RECT 93.750 106.920 94.070 106.980 ;
        RECT 92.845 106.780 94.070 106.920 ;
        RECT 92.845 106.735 93.135 106.780 ;
        RECT 93.750 106.720 94.070 106.780 ;
        RECT 103.410 106.720 103.730 106.980 ;
        RECT 108.025 106.920 108.315 106.965 ;
        RECT 108.930 106.920 109.250 106.980 ;
        RECT 111.230 106.920 111.550 106.980 ;
        RECT 108.025 106.780 111.550 106.920 ;
        RECT 108.025 106.735 108.315 106.780 ;
        RECT 108.930 106.720 109.250 106.780 ;
        RECT 111.230 106.720 111.550 106.780 ;
        RECT 124.110 106.720 124.430 106.980 ;
        RECT 140.670 106.720 140.990 106.980 ;
        RECT 141.130 106.920 141.450 106.980 ;
        RECT 143.980 106.920 144.120 107.415 ;
        RECT 141.130 106.780 144.120 106.920 ;
        RECT 141.130 106.720 141.450 106.780 ;
        RECT 17.320 106.100 147.040 106.580 ;
        RECT 32.110 105.900 32.430 105.960 ;
        RECT 33.965 105.900 34.255 105.945 ;
        RECT 20.240 105.760 34.255 105.900 ;
        RECT 20.240 105.265 20.380 105.760 ;
        RECT 32.110 105.700 32.430 105.760 ;
        RECT 33.965 105.715 34.255 105.760 ;
        RECT 73.050 105.900 73.370 105.960 ;
        RECT 78.585 105.900 78.875 105.945 ;
        RECT 73.050 105.760 78.875 105.900 ;
        RECT 73.050 105.700 73.370 105.760 ;
        RECT 78.585 105.715 78.875 105.760 ;
        RECT 79.950 105.900 80.270 105.960 ;
        RECT 85.945 105.900 86.235 105.945 ;
        RECT 97.430 105.900 97.750 105.960 ;
        RECT 79.950 105.760 84.780 105.900 ;
        RECT 79.950 105.700 80.270 105.760 ;
        RECT 27.510 105.560 27.830 105.620 ;
        RECT 23.460 105.420 27.830 105.560 ;
        RECT 20.165 105.035 20.455 105.265 ;
        RECT 23.460 104.925 23.600 105.420 ;
        RECT 27.510 105.360 27.830 105.420 ;
        RECT 72.560 105.560 72.850 105.605 ;
        RECT 73.510 105.560 73.830 105.620 ;
        RECT 72.560 105.420 73.830 105.560 ;
        RECT 72.560 105.375 72.850 105.420 ;
        RECT 73.510 105.360 73.830 105.420 ;
        RECT 80.410 105.360 80.730 105.620 ;
        RECT 83.630 105.560 83.950 105.620 ;
        RECT 84.640 105.605 84.780 105.760 ;
        RECT 85.945 105.760 97.750 105.900 ;
        RECT 85.945 105.715 86.235 105.760 ;
        RECT 97.430 105.700 97.750 105.760 ;
        RECT 101.110 105.700 101.430 105.960 ;
        RECT 101.570 105.900 101.890 105.960 ;
        RECT 112.625 105.900 112.915 105.945 ;
        RECT 125.030 105.900 125.350 105.960 ;
        RECT 129.645 105.900 129.935 105.945 ;
        RECT 101.570 105.760 111.000 105.900 ;
        RECT 101.570 105.700 101.890 105.760 ;
        RECT 84.105 105.560 84.395 105.605 ;
        RECT 80.960 105.420 83.400 105.560 ;
        RECT 24.290 105.020 24.610 105.280 ;
        RECT 28.400 105.220 28.690 105.265 ;
        RECT 30.730 105.220 31.050 105.280 ;
        RECT 28.400 105.080 31.050 105.220 ;
        RECT 28.400 105.035 28.690 105.080 ;
        RECT 30.730 105.020 31.050 105.080 ;
        RECT 66.610 105.220 66.930 105.280 ;
        RECT 71.225 105.220 71.515 105.265 ;
        RECT 66.610 105.080 71.515 105.220 ;
        RECT 66.610 105.020 66.930 105.080 ;
        RECT 71.225 105.035 71.515 105.080 ;
        RECT 23.385 104.695 23.675 104.925 ;
        RECT 23.830 104.680 24.150 104.940 ;
        RECT 27.050 104.680 27.370 104.940 ;
        RECT 80.960 104.925 81.100 105.420 ;
        RECT 83.260 105.265 83.400 105.420 ;
        RECT 83.630 105.420 84.395 105.560 ;
        RECT 83.630 105.360 83.950 105.420 ;
        RECT 84.105 105.375 84.395 105.420 ;
        RECT 84.565 105.375 84.855 105.605 ;
        RECT 94.670 105.560 94.990 105.620 ;
        RECT 108.010 105.560 108.330 105.620 ;
        RECT 110.860 105.605 111.000 105.760 ;
        RECT 112.625 105.760 124.800 105.900 ;
        RECT 112.625 105.715 112.915 105.760 ;
        RECT 110.785 105.560 111.075 105.605 ;
        RECT 114.910 105.560 115.230 105.620 ;
        RECT 86.940 105.420 102.720 105.560 ;
        RECT 86.940 105.280 87.080 105.420 ;
        RECT 94.670 105.360 94.990 105.420 ;
        RECT 85.010 105.265 85.330 105.280 ;
        RECT 82.725 105.035 83.015 105.265 ;
        RECT 83.190 105.035 83.480 105.265 ;
        RECT 85.010 105.220 85.340 105.265 ;
        RECT 85.010 105.080 85.525 105.220 ;
        RECT 85.010 105.035 85.340 105.080 ;
        RECT 27.945 104.880 28.235 104.925 ;
        RECT 29.135 104.880 29.425 104.925 ;
        RECT 31.655 104.880 31.945 104.925 ;
        RECT 27.945 104.740 31.945 104.880 ;
        RECT 27.945 104.695 28.235 104.740 ;
        RECT 29.135 104.695 29.425 104.740 ;
        RECT 31.655 104.695 31.945 104.740 ;
        RECT 72.105 104.880 72.395 104.925 ;
        RECT 73.295 104.880 73.585 104.925 ;
        RECT 75.815 104.880 76.105 104.925 ;
        RECT 80.885 104.880 81.175 104.925 ;
        RECT 72.105 104.740 76.105 104.880 ;
        RECT 72.105 104.695 72.395 104.740 ;
        RECT 73.295 104.695 73.585 104.740 ;
        RECT 75.815 104.695 76.105 104.740 ;
        RECT 78.200 104.740 81.175 104.880 ;
        RECT 27.550 104.540 27.840 104.585 ;
        RECT 29.650 104.540 29.940 104.585 ;
        RECT 31.220 104.540 31.510 104.585 ;
        RECT 27.550 104.400 31.510 104.540 ;
        RECT 27.550 104.355 27.840 104.400 ;
        RECT 29.650 104.355 29.940 104.400 ;
        RECT 31.220 104.355 31.510 104.400 ;
        RECT 71.710 104.540 72.000 104.585 ;
        RECT 73.810 104.540 74.100 104.585 ;
        RECT 75.380 104.540 75.670 104.585 ;
        RECT 71.710 104.400 75.670 104.540 ;
        RECT 71.710 104.355 72.000 104.400 ;
        RECT 73.810 104.355 74.100 104.400 ;
        RECT 75.380 104.355 75.670 104.400 ;
        RECT 16.010 104.200 16.330 104.260 ;
        RECT 19.245 104.200 19.535 104.245 ;
        RECT 16.010 104.060 19.535 104.200 ;
        RECT 16.010 104.000 16.330 104.060 ;
        RECT 19.245 104.015 19.535 104.060 ;
        RECT 25.670 104.200 25.990 104.260 ;
        RECT 26.145 104.200 26.435 104.245 ;
        RECT 25.670 104.060 26.435 104.200 ;
        RECT 25.670 104.000 25.990 104.060 ;
        RECT 26.145 104.015 26.435 104.060 ;
        RECT 77.650 104.200 77.970 104.260 ;
        RECT 78.200 104.245 78.340 104.740 ;
        RECT 80.885 104.695 81.175 104.740 ;
        RECT 81.805 104.695 82.095 104.925 ;
        RECT 82.800 104.880 82.940 105.035 ;
        RECT 85.010 105.020 85.330 105.035 ;
        RECT 86.850 105.020 87.170 105.280 ;
        RECT 88.230 105.265 88.550 105.280 ;
        RECT 88.200 105.220 88.550 105.265 ;
        RECT 88.035 105.080 88.550 105.220 ;
        RECT 88.200 105.035 88.550 105.080 ;
        RECT 88.230 105.020 88.550 105.035 ;
        RECT 95.590 105.020 95.910 105.280 ;
        RECT 97.430 105.020 97.750 105.280 ;
        RECT 101.570 105.020 101.890 105.280 ;
        RECT 102.580 105.265 102.720 105.420 ;
        RECT 108.010 105.420 110.080 105.560 ;
        RECT 108.010 105.360 108.330 105.420 ;
        RECT 102.505 105.035 102.795 105.265 ;
        RECT 102.950 105.220 103.270 105.280 ;
        RECT 103.785 105.220 104.075 105.265 ;
        RECT 102.950 105.080 104.075 105.220 ;
        RECT 102.950 105.020 103.270 105.080 ;
        RECT 103.785 105.035 104.075 105.080 ;
        RECT 105.250 105.220 105.570 105.280 ;
        RECT 109.940 105.265 110.080 105.420 ;
        RECT 110.785 105.420 115.230 105.560 ;
        RECT 110.785 105.375 111.075 105.420 ;
        RECT 114.910 105.360 115.230 105.420 ;
        RECT 123.620 105.560 123.910 105.605 ;
        RECT 124.110 105.560 124.430 105.620 ;
        RECT 123.620 105.420 124.430 105.560 ;
        RECT 124.660 105.560 124.800 105.760 ;
        RECT 125.030 105.760 129.935 105.900 ;
        RECT 125.030 105.700 125.350 105.760 ;
        RECT 129.645 105.715 129.935 105.760 ;
        RECT 131.485 105.900 131.775 105.945 ;
        RECT 137.450 105.900 137.770 105.960 ;
        RECT 131.485 105.760 137.770 105.900 ;
        RECT 131.485 105.715 131.775 105.760 ;
        RECT 137.450 105.700 137.770 105.760 ;
        RECT 139.750 105.900 140.070 105.960 ;
        RECT 145.270 105.900 145.590 105.960 ;
        RECT 139.750 105.760 145.590 105.900 ;
        RECT 139.750 105.700 140.070 105.760 ;
        RECT 145.270 105.700 145.590 105.760 ;
        RECT 129.170 105.560 129.490 105.620 ;
        RECT 124.660 105.420 129.490 105.560 ;
        RECT 123.620 105.375 123.910 105.420 ;
        RECT 124.110 105.360 124.430 105.420 ;
        RECT 129.170 105.360 129.490 105.420 ;
        RECT 131.945 105.560 132.235 105.605 ;
        RECT 143.430 105.560 143.750 105.620 ;
        RECT 131.945 105.420 143.750 105.560 ;
        RECT 131.945 105.375 132.235 105.420 ;
        RECT 105.250 105.080 109.160 105.220 ;
        RECT 105.250 105.020 105.570 105.080 ;
        RECT 86.390 104.880 86.710 104.940 ;
        RECT 82.800 104.740 86.710 104.880 ;
        RECT 81.880 104.540 82.020 104.695 ;
        RECT 86.390 104.680 86.710 104.740 ;
        RECT 87.745 104.880 88.035 104.925 ;
        RECT 88.935 104.880 89.225 104.925 ;
        RECT 91.455 104.880 91.745 104.925 ;
        RECT 87.745 104.740 91.745 104.880 ;
        RECT 87.745 104.695 88.035 104.740 ;
        RECT 88.935 104.695 89.225 104.740 ;
        RECT 91.455 104.695 91.745 104.740 ;
        RECT 103.385 104.880 103.675 104.925 ;
        RECT 104.575 104.880 104.865 104.925 ;
        RECT 107.095 104.880 107.385 104.925 ;
        RECT 103.385 104.740 107.385 104.880 ;
        RECT 109.020 104.880 109.160 105.080 ;
        RECT 109.865 105.035 110.155 105.265 ;
        RECT 111.230 105.020 111.550 105.280 ;
        RECT 111.705 105.035 111.995 105.265 ;
        RECT 111.780 104.880 111.920 105.035 ;
        RECT 116.750 104.880 117.070 104.940 ;
        RECT 109.020 104.740 117.070 104.880 ;
        RECT 103.385 104.695 103.675 104.740 ;
        RECT 104.575 104.695 104.865 104.740 ;
        RECT 107.095 104.695 107.385 104.740 ;
        RECT 116.750 104.680 117.070 104.740 ;
        RECT 122.270 104.680 122.590 104.940 ;
        RECT 123.165 104.880 123.455 104.925 ;
        RECT 124.355 104.880 124.645 104.925 ;
        RECT 126.875 104.880 127.165 104.925 ;
        RECT 123.165 104.740 127.165 104.880 ;
        RECT 123.165 104.695 123.455 104.740 ;
        RECT 124.355 104.695 124.645 104.740 ;
        RECT 126.875 104.695 127.165 104.740 ;
        RECT 86.850 104.540 87.170 104.600 ;
        RECT 81.880 104.400 87.170 104.540 ;
        RECT 86.850 104.340 87.170 104.400 ;
        RECT 87.350 104.540 87.640 104.585 ;
        RECT 89.450 104.540 89.740 104.585 ;
        RECT 91.020 104.540 91.310 104.585 ;
        RECT 100.650 104.540 100.970 104.600 ;
        RECT 87.350 104.400 91.310 104.540 ;
        RECT 87.350 104.355 87.640 104.400 ;
        RECT 89.450 104.355 89.740 104.400 ;
        RECT 91.020 104.355 91.310 104.400 ;
        RECT 93.380 104.400 100.970 104.540 ;
        RECT 78.125 104.200 78.415 104.245 ;
        RECT 77.650 104.060 78.415 104.200 ;
        RECT 77.650 104.000 77.970 104.060 ;
        RECT 78.125 104.015 78.415 104.060 ;
        RECT 79.030 104.200 79.350 104.260 ;
        RECT 93.380 104.200 93.520 104.400 ;
        RECT 100.650 104.340 100.970 104.400 ;
        RECT 102.990 104.540 103.280 104.585 ;
        RECT 105.090 104.540 105.380 104.585 ;
        RECT 106.660 104.540 106.950 104.585 ;
        RECT 102.990 104.400 106.950 104.540 ;
        RECT 102.990 104.355 103.280 104.400 ;
        RECT 105.090 104.355 105.380 104.400 ;
        RECT 106.660 104.355 106.950 104.400 ;
        RECT 108.470 104.540 108.790 104.600 ;
        RECT 122.770 104.540 123.060 104.585 ;
        RECT 124.870 104.540 125.160 104.585 ;
        RECT 126.440 104.540 126.730 104.585 ;
        RECT 108.470 104.400 122.270 104.540 ;
        RECT 108.470 104.340 108.790 104.400 ;
        RECT 79.030 104.060 93.520 104.200 ;
        RECT 79.030 104.000 79.350 104.060 ;
        RECT 93.750 104.000 94.070 104.260 ;
        RECT 95.130 104.200 95.450 104.260 ;
        RECT 98.350 104.200 98.670 104.260 ;
        RECT 95.130 104.060 98.670 104.200 ;
        RECT 95.130 104.000 95.450 104.060 ;
        RECT 98.350 104.000 98.670 104.060 ;
        RECT 108.010 104.200 108.330 104.260 ;
        RECT 109.405 104.200 109.695 104.245 ;
        RECT 108.010 104.060 109.695 104.200 ;
        RECT 122.130 104.200 122.270 104.400 ;
        RECT 122.770 104.400 126.730 104.540 ;
        RECT 122.770 104.355 123.060 104.400 ;
        RECT 124.870 104.355 125.160 104.400 ;
        RECT 126.440 104.355 126.730 104.400 ;
        RECT 129.185 104.540 129.475 104.585 ;
        RECT 132.020 104.540 132.160 105.375 ;
        RECT 143.430 105.360 143.750 105.420 ;
        RECT 137.450 105.220 137.770 105.280 ;
        RECT 141.605 105.220 141.895 105.265 ;
        RECT 137.450 105.080 141.895 105.220 ;
        RECT 137.450 105.020 137.770 105.080 ;
        RECT 141.605 105.035 141.895 105.080 ;
        RECT 143.905 105.220 144.195 105.265 ;
        RECT 144.350 105.220 144.670 105.280 ;
        RECT 143.905 105.080 144.670 105.220 ;
        RECT 143.905 105.035 144.195 105.080 ;
        RECT 144.350 105.020 144.670 105.080 ;
        RECT 132.850 104.680 133.170 104.940 ;
        RECT 137.910 104.680 138.230 104.940 ;
        RECT 138.845 104.880 139.135 104.925 ;
        RECT 139.750 104.880 140.070 104.940 ;
        RECT 138.845 104.740 140.070 104.880 ;
        RECT 138.845 104.695 139.135 104.740 ;
        RECT 139.750 104.680 140.070 104.740 ;
        RECT 142.050 104.680 142.370 104.940 ;
        RECT 142.525 104.695 142.815 104.925 ;
        RECT 139.290 104.540 139.610 104.600 ;
        RECT 142.600 104.540 142.740 104.695 ;
        RECT 129.185 104.400 132.160 104.540 ;
        RECT 132.480 104.400 142.740 104.540 ;
        RECT 129.185 104.355 129.475 104.400 ;
        RECT 132.480 104.200 132.620 104.400 ;
        RECT 139.290 104.340 139.610 104.400 ;
        RECT 144.810 104.340 145.130 104.600 ;
        RECT 122.130 104.060 132.620 104.200 ;
        RECT 133.310 104.200 133.630 104.260 ;
        RECT 135.625 104.200 135.915 104.245 ;
        RECT 133.310 104.060 135.915 104.200 ;
        RECT 108.010 104.000 108.330 104.060 ;
        RECT 109.405 104.015 109.695 104.060 ;
        RECT 133.310 104.000 133.630 104.060 ;
        RECT 135.625 104.015 135.915 104.060 ;
        RECT 136.530 104.200 136.850 104.260 ;
        RECT 139.765 104.200 140.055 104.245 ;
        RECT 136.530 104.060 140.055 104.200 ;
        RECT 136.530 104.000 136.850 104.060 ;
        RECT 139.765 104.015 140.055 104.060 ;
        RECT 17.320 103.380 147.040 103.860 ;
        RECT 19.245 103.180 19.535 103.225 ;
        RECT 20.150 103.180 20.470 103.240 ;
        RECT 24.290 103.180 24.610 103.240 ;
        RECT 19.245 103.040 24.610 103.180 ;
        RECT 19.245 102.995 19.535 103.040 ;
        RECT 20.150 102.980 20.470 103.040 ;
        RECT 24.290 102.980 24.610 103.040 ;
        RECT 30.730 102.980 31.050 103.240 ;
        RECT 84.550 102.980 84.870 103.240 ;
        RECT 86.390 103.180 86.710 103.240 ;
        RECT 88.705 103.180 88.995 103.225 ;
        RECT 86.390 103.040 88.995 103.180 ;
        RECT 86.390 102.980 86.710 103.040 ;
        RECT 88.705 102.995 88.995 103.040 ;
        RECT 102.950 102.980 103.270 103.240 ;
        RECT 110.310 102.980 110.630 103.240 ;
        RECT 124.570 103.180 124.890 103.240 ;
        RECT 132.850 103.180 133.170 103.240 ;
        RECT 114.540 103.040 133.170 103.180 ;
        RECT 21.990 102.840 22.280 102.885 ;
        RECT 23.560 102.840 23.850 102.885 ;
        RECT 25.660 102.840 25.950 102.885 ;
        RECT 21.990 102.700 25.950 102.840 ;
        RECT 21.990 102.655 22.280 102.700 ;
        RECT 23.560 102.655 23.850 102.700 ;
        RECT 25.660 102.655 25.950 102.700 ;
        RECT 63.890 102.840 64.180 102.885 ;
        RECT 65.990 102.840 66.280 102.885 ;
        RECT 67.560 102.840 67.850 102.885 ;
        RECT 63.890 102.700 67.850 102.840 ;
        RECT 63.890 102.655 64.180 102.700 ;
        RECT 65.990 102.655 66.280 102.700 ;
        RECT 67.560 102.655 67.850 102.700 ;
        RECT 68.450 102.840 68.770 102.900 ;
        RECT 73.970 102.840 74.290 102.900 ;
        RECT 68.450 102.700 82.480 102.840 ;
        RECT 68.450 102.640 68.770 102.700 ;
        RECT 73.970 102.640 74.290 102.700 ;
        RECT 21.555 102.500 21.845 102.545 ;
        RECT 24.075 102.500 24.365 102.545 ;
        RECT 25.265 102.500 25.555 102.545 ;
        RECT 21.555 102.360 25.555 102.500 ;
        RECT 21.555 102.315 21.845 102.360 ;
        RECT 24.075 102.315 24.365 102.360 ;
        RECT 25.265 102.315 25.555 102.360 ;
        RECT 27.510 102.500 27.830 102.560 ;
        RECT 33.505 102.500 33.795 102.545 ;
        RECT 27.510 102.360 33.795 102.500 ;
        RECT 27.510 102.300 27.830 102.360 ;
        RECT 33.505 102.315 33.795 102.360 ;
        RECT 64.285 102.500 64.575 102.545 ;
        RECT 65.475 102.500 65.765 102.545 ;
        RECT 67.995 102.500 68.285 102.545 ;
        RECT 64.285 102.360 68.285 102.500 ;
        RECT 64.285 102.315 64.575 102.360 ;
        RECT 65.475 102.315 65.765 102.360 ;
        RECT 67.995 102.315 68.285 102.360 ;
        RECT 71.210 102.500 71.530 102.560 ;
        RECT 73.525 102.500 73.815 102.545 ;
        RECT 79.030 102.500 79.350 102.560 ;
        RECT 82.340 102.545 82.480 102.700 ;
        RECT 84.090 102.640 84.410 102.900 ;
        RECT 103.410 102.640 103.730 102.900 ;
        RECT 109.850 102.640 110.170 102.900 ;
        RECT 71.210 102.360 79.350 102.500 ;
        RECT 71.210 102.300 71.530 102.360 ;
        RECT 73.525 102.315 73.815 102.360 ;
        RECT 79.030 102.300 79.350 102.360 ;
        RECT 82.265 102.500 82.555 102.545 ;
        RECT 96.510 102.500 96.830 102.560 ;
        RECT 82.265 102.360 96.830 102.500 ;
        RECT 82.265 102.315 82.555 102.360 ;
        RECT 96.510 102.300 96.830 102.360 ;
        RECT 98.350 102.500 98.670 102.560 ;
        RECT 101.110 102.500 101.430 102.560 ;
        RECT 114.005 102.500 114.295 102.545 ;
        RECT 114.540 102.500 114.680 103.040 ;
        RECT 124.570 102.980 124.890 103.040 ;
        RECT 132.850 102.980 133.170 103.040 ;
        RECT 117.710 102.840 118.000 102.885 ;
        RECT 119.810 102.840 120.100 102.885 ;
        RECT 121.380 102.840 121.670 102.885 ;
        RECT 117.710 102.700 121.670 102.840 ;
        RECT 117.710 102.655 118.000 102.700 ;
        RECT 119.810 102.655 120.100 102.700 ;
        RECT 121.380 102.655 121.670 102.700 ;
        RECT 132.405 102.840 132.695 102.885 ;
        RECT 133.310 102.840 133.630 102.900 ;
        RECT 132.405 102.700 133.630 102.840 ;
        RECT 132.405 102.655 132.695 102.700 ;
        RECT 133.310 102.640 133.630 102.700 ;
        RECT 136.570 102.840 136.860 102.885 ;
        RECT 138.670 102.840 138.960 102.885 ;
        RECT 140.240 102.840 140.530 102.885 ;
        RECT 136.570 102.700 140.530 102.840 ;
        RECT 136.570 102.655 136.860 102.700 ;
        RECT 138.670 102.655 138.960 102.700 ;
        RECT 140.240 102.655 140.530 102.700 ;
        RECT 98.350 102.360 114.680 102.500 ;
        RECT 118.105 102.500 118.395 102.545 ;
        RECT 119.295 102.500 119.585 102.545 ;
        RECT 121.815 102.500 122.105 102.545 ;
        RECT 118.105 102.360 122.105 102.500 ;
        RECT 98.350 102.300 98.670 102.360 ;
        RECT 101.110 102.300 101.430 102.360 ;
        RECT 114.005 102.315 114.295 102.360 ;
        RECT 118.105 102.315 118.395 102.360 ;
        RECT 119.295 102.315 119.585 102.360 ;
        RECT 121.815 102.315 122.105 102.360 ;
        RECT 126.410 102.500 126.730 102.560 ;
        RECT 130.565 102.500 130.855 102.545 ;
        RECT 126.410 102.360 130.855 102.500 ;
        RECT 126.410 102.300 126.730 102.360 ;
        RECT 130.565 102.315 130.855 102.360 ;
        RECT 136.070 102.300 136.390 102.560 ;
        RECT 136.965 102.500 137.255 102.545 ;
        RECT 138.155 102.500 138.445 102.545 ;
        RECT 140.675 102.500 140.965 102.545 ;
        RECT 136.965 102.360 140.965 102.500 ;
        RECT 136.965 102.315 137.255 102.360 ;
        RECT 138.155 102.315 138.445 102.360 ;
        RECT 140.675 102.315 140.965 102.360 ;
        RECT 24.865 102.160 25.155 102.205 ;
        RECT 25.670 102.160 25.990 102.220 ;
        RECT 24.865 102.020 25.990 102.160 ;
        RECT 24.865 101.975 25.155 102.020 ;
        RECT 25.670 101.960 25.990 102.020 ;
        RECT 26.145 102.160 26.435 102.205 ;
        RECT 27.050 102.160 27.370 102.220 ;
        RECT 26.145 102.020 27.370 102.160 ;
        RECT 26.145 101.975 26.435 102.020 ;
        RECT 27.050 101.960 27.370 102.020 ;
        RECT 32.110 102.160 32.430 102.220 ;
        RECT 32.585 102.160 32.875 102.205 ;
        RECT 32.110 102.020 32.875 102.160 ;
        RECT 32.110 101.960 32.430 102.020 ;
        RECT 32.585 101.975 32.875 102.020 ;
        RECT 61.550 102.160 61.870 102.220 ;
        RECT 63.405 102.160 63.695 102.205 ;
        RECT 66.610 102.160 66.930 102.220 ;
        RECT 72.590 102.160 72.910 102.220 ;
        RECT 78.110 102.160 78.430 102.220 ;
        RECT 61.550 102.020 66.930 102.160 ;
        RECT 72.395 102.020 78.430 102.160 ;
        RECT 61.550 101.960 61.870 102.020 ;
        RECT 63.405 101.975 63.695 102.020 ;
        RECT 66.610 101.960 66.930 102.020 ;
        RECT 72.590 101.960 72.910 102.020 ;
        RECT 78.110 101.960 78.430 102.020 ;
        RECT 89.610 101.960 89.930 102.220 ;
        RECT 91.465 102.160 91.755 102.205 ;
        RECT 93.750 102.160 94.070 102.220 ;
        RECT 91.465 102.020 94.070 102.160 ;
        RECT 91.465 101.975 91.755 102.020 ;
        RECT 93.750 101.960 94.070 102.020 ;
        RECT 105.265 102.160 105.555 102.205 ;
        RECT 108.025 102.160 108.315 102.205 ;
        RECT 109.390 102.160 109.710 102.220 ;
        RECT 105.265 102.020 109.710 102.160 ;
        RECT 105.265 101.975 105.555 102.020 ;
        RECT 108.025 101.975 108.315 102.020 ;
        RECT 109.390 101.960 109.710 102.020 ;
        RECT 114.450 102.160 114.770 102.220 ;
        RECT 114.925 102.160 115.215 102.205 ;
        RECT 114.450 102.020 115.215 102.160 ;
        RECT 114.450 101.960 114.770 102.020 ;
        RECT 114.925 101.975 115.215 102.020 ;
        RECT 117.225 102.160 117.515 102.205 ;
        RECT 122.270 102.160 122.590 102.220 ;
        RECT 142.510 102.160 142.830 102.220 ;
        RECT 143.905 102.160 144.195 102.205 ;
        RECT 117.225 102.020 122.590 102.160 ;
        RECT 117.225 101.975 117.515 102.020 ;
        RECT 122.270 101.960 122.590 102.020 ;
        RECT 129.720 102.020 142.830 102.160 ;
        RECT 64.770 101.865 65.090 101.880 ;
        RECT 64.740 101.635 65.090 101.865 ;
        RECT 73.065 101.820 73.355 101.865 ;
        RECT 64.770 101.620 65.090 101.635 ;
        RECT 70.380 101.680 73.355 101.820 ;
        RECT 70.380 101.540 70.520 101.680 ;
        RECT 73.065 101.635 73.355 101.680 ;
        RECT 89.150 101.820 89.470 101.880 ;
        RECT 90.085 101.820 90.375 101.865 ;
        RECT 89.150 101.680 90.375 101.820 ;
        RECT 89.150 101.620 89.470 101.680 ;
        RECT 90.085 101.635 90.375 101.680 ;
        RECT 90.530 101.820 90.850 101.880 ;
        RECT 97.430 101.820 97.750 101.880 ;
        RECT 118.590 101.865 118.910 101.880 ;
        RECT 90.530 101.680 97.750 101.820 ;
        RECT 30.730 101.480 31.050 101.540 ;
        RECT 33.045 101.480 33.335 101.525 ;
        RECT 30.730 101.340 33.335 101.480 ;
        RECT 30.730 101.280 31.050 101.340 ;
        RECT 33.045 101.295 33.335 101.340 ;
        RECT 70.290 101.280 70.610 101.540 ;
        RECT 70.750 101.280 71.070 101.540 ;
        RECT 90.160 101.480 90.300 101.635 ;
        RECT 90.530 101.620 90.850 101.680 ;
        RECT 97.430 101.620 97.750 101.680 ;
        RECT 114.540 101.680 118.360 101.820 ;
        RECT 114.540 101.540 114.680 101.680 ;
        RECT 91.910 101.480 92.230 101.540 ;
        RECT 90.160 101.340 92.230 101.480 ;
        RECT 91.910 101.280 92.230 101.340 ;
        RECT 114.450 101.280 114.770 101.540 ;
        RECT 116.765 101.480 117.055 101.525 ;
        RECT 117.670 101.480 117.990 101.540 ;
        RECT 116.765 101.340 117.990 101.480 ;
        RECT 118.220 101.480 118.360 101.680 ;
        RECT 118.560 101.635 118.910 101.865 ;
        RECT 118.590 101.620 118.910 101.635 ;
        RECT 124.125 101.480 124.415 101.525 ;
        RECT 129.720 101.480 129.860 102.020 ;
        RECT 142.510 101.960 142.830 102.020 ;
        RECT 143.060 102.020 144.195 102.160 ;
        RECT 137.310 101.820 137.600 101.865 ;
        RECT 132.940 101.680 137.600 101.820 ;
        RECT 132.940 101.525 133.080 101.680 ;
        RECT 137.310 101.635 137.600 101.680 ;
        RECT 118.220 101.340 129.860 101.480 ;
        RECT 116.765 101.295 117.055 101.340 ;
        RECT 117.670 101.280 117.990 101.340 ;
        RECT 124.125 101.295 124.415 101.340 ;
        RECT 132.865 101.295 133.155 101.525 ;
        RECT 137.910 101.480 138.230 101.540 ;
        RECT 143.060 101.525 143.200 102.020 ;
        RECT 143.905 101.975 144.195 102.020 ;
        RECT 142.985 101.480 143.275 101.525 ;
        RECT 137.910 101.340 143.275 101.480 ;
        RECT 137.910 101.280 138.230 101.340 ;
        RECT 142.985 101.295 143.275 101.340 ;
        RECT 144.810 101.280 145.130 101.540 ;
        RECT 17.320 100.660 147.040 101.140 ;
        RECT 18.310 100.460 18.630 100.520 ;
        RECT 19.245 100.460 19.535 100.505 ;
        RECT 18.310 100.320 19.535 100.460 ;
        RECT 18.310 100.260 18.630 100.320 ;
        RECT 19.245 100.275 19.535 100.320 ;
        RECT 30.730 100.260 31.050 100.520 ;
        RECT 64.325 100.460 64.615 100.505 ;
        RECT 64.770 100.460 65.090 100.520 ;
        RECT 64.325 100.320 65.090 100.460 ;
        RECT 64.325 100.275 64.615 100.320 ;
        RECT 64.770 100.260 65.090 100.320 ;
        RECT 93.750 100.460 94.070 100.520 ;
        RECT 118.130 100.460 118.450 100.520 ;
        RECT 93.750 100.320 118.450 100.460 ;
        RECT 93.750 100.260 94.070 100.320 ;
        RECT 118.130 100.260 118.450 100.320 ;
        RECT 118.590 100.260 118.910 100.520 ;
        RECT 136.085 100.275 136.375 100.505 ;
        RECT 142.050 100.460 142.370 100.520 ;
        RECT 143.445 100.460 143.735 100.505 ;
        RECT 142.050 100.320 143.735 100.460 ;
        RECT 30.285 100.120 30.575 100.165 ;
        RECT 25.530 99.980 30.575 100.120 ;
        RECT 20.150 99.580 20.470 99.840 ;
        RECT 21.990 99.780 22.310 99.840 ;
        RECT 25.530 99.780 25.670 99.980 ;
        RECT 30.285 99.935 30.575 99.980 ;
        RECT 66.625 100.120 66.915 100.165 ;
        RECT 67.070 100.120 67.390 100.180 ;
        RECT 68.450 100.120 68.770 100.180 ;
        RECT 66.625 99.980 68.770 100.120 ;
        RECT 66.625 99.935 66.915 99.980 ;
        RECT 67.070 99.920 67.390 99.980 ;
        RECT 68.450 99.920 68.770 99.980 ;
        RECT 107.105 100.120 107.395 100.165 ;
        RECT 109.390 100.120 109.710 100.180 ;
        RECT 112.610 100.120 112.930 100.180 ;
        RECT 116.305 100.120 116.595 100.165 ;
        RECT 107.105 99.980 116.595 100.120 ;
        RECT 136.160 100.120 136.300 100.275 ;
        RECT 142.050 100.260 142.370 100.320 ;
        RECT 143.445 100.275 143.735 100.320 ;
        RECT 137.770 100.120 138.060 100.165 ;
        RECT 136.160 99.980 138.060 100.120 ;
        RECT 107.105 99.935 107.395 99.980 ;
        RECT 109.390 99.920 109.710 99.980 ;
        RECT 112.610 99.920 112.930 99.980 ;
        RECT 116.305 99.935 116.595 99.980 ;
        RECT 137.770 99.935 138.060 99.980 ;
        RECT 21.160 99.640 25.670 99.780 ;
        RECT 26.705 99.780 26.995 99.825 ;
        RECT 26.705 99.640 28.660 99.780 ;
        RECT 21.160 99.145 21.300 99.640 ;
        RECT 21.990 99.580 22.310 99.640 ;
        RECT 26.705 99.595 26.995 99.640 ;
        RECT 23.395 99.440 23.685 99.485 ;
        RECT 25.915 99.440 26.205 99.485 ;
        RECT 27.105 99.440 27.395 99.485 ;
        RECT 23.395 99.300 27.395 99.440 ;
        RECT 23.395 99.255 23.685 99.300 ;
        RECT 25.915 99.255 26.205 99.300 ;
        RECT 27.105 99.255 27.395 99.300 ;
        RECT 27.985 99.255 28.275 99.485 ;
        RECT 21.085 98.915 21.375 99.145 ;
        RECT 23.830 99.100 24.120 99.145 ;
        RECT 25.400 99.100 25.690 99.145 ;
        RECT 27.500 99.100 27.790 99.145 ;
        RECT 23.830 98.960 27.790 99.100 ;
        RECT 23.830 98.915 24.120 98.960 ;
        RECT 25.400 98.915 25.690 98.960 ;
        RECT 27.500 98.915 27.790 98.960 ;
        RECT 27.050 98.760 27.370 98.820 ;
        RECT 28.060 98.760 28.200 99.255 ;
        RECT 28.520 99.145 28.660 99.640 ;
        RECT 28.890 99.440 29.210 99.500 ;
        RECT 31.205 99.440 31.495 99.485 ;
        RECT 28.890 99.300 31.495 99.440 ;
        RECT 28.890 99.240 29.210 99.300 ;
        RECT 31.205 99.255 31.495 99.300 ;
        RECT 71.670 99.440 71.990 99.500 ;
        RECT 103.870 99.440 104.190 99.500 ;
        RECT 113.990 99.440 114.310 99.500 ;
        RECT 71.670 99.300 104.190 99.440 ;
        RECT 71.670 99.240 71.990 99.300 ;
        RECT 103.870 99.240 104.190 99.300 ;
        RECT 104.420 99.300 114.310 99.440 ;
        RECT 116.380 99.440 116.520 99.935 ;
        RECT 116.750 99.780 117.070 99.840 ;
        RECT 132.390 99.780 132.710 99.840 ;
        RECT 135.610 99.780 135.930 99.840 ;
        RECT 116.750 99.640 135.930 99.780 ;
        RECT 116.750 99.580 117.070 99.640 ;
        RECT 132.390 99.580 132.710 99.640 ;
        RECT 135.610 99.580 135.930 99.640 ;
        RECT 136.070 99.780 136.390 99.840 ;
        RECT 136.545 99.780 136.835 99.825 ;
        RECT 136.070 99.640 136.835 99.780 ;
        RECT 136.070 99.580 136.390 99.640 ;
        RECT 136.545 99.595 136.835 99.640 ;
        RECT 143.430 99.780 143.750 99.840 ;
        RECT 143.905 99.780 144.195 99.825 ;
        RECT 143.430 99.640 144.195 99.780 ;
        RECT 143.430 99.580 143.750 99.640 ;
        RECT 143.905 99.595 144.195 99.640 ;
        RECT 116.380 99.300 118.360 99.440 ;
        RECT 28.445 98.915 28.735 99.145 ;
        RECT 65.245 99.100 65.535 99.145 ;
        RECT 70.750 99.100 71.070 99.160 ;
        RECT 65.245 98.960 71.070 99.100 ;
        RECT 65.245 98.915 65.535 98.960 ;
        RECT 70.750 98.900 71.070 98.960 ;
        RECT 78.110 99.100 78.430 99.160 ;
        RECT 86.390 99.100 86.710 99.160 ;
        RECT 104.420 99.100 104.560 99.300 ;
        RECT 113.990 99.240 114.310 99.300 ;
        RECT 78.110 98.960 104.560 99.100 ;
        RECT 78.110 98.900 78.430 98.960 ;
        RECT 86.390 98.900 86.710 98.960 ;
        RECT 108.930 98.900 109.250 99.160 ;
        RECT 117.670 98.900 117.990 99.160 ;
        RECT 118.220 99.100 118.360 99.300 ;
        RECT 133.770 99.240 134.090 99.500 ;
        RECT 137.425 99.440 137.715 99.485 ;
        RECT 138.615 99.440 138.905 99.485 ;
        RECT 141.135 99.440 141.425 99.485 ;
        RECT 137.425 99.300 141.425 99.440 ;
        RECT 137.425 99.255 137.715 99.300 ;
        RECT 138.615 99.255 138.905 99.300 ;
        RECT 141.135 99.255 141.425 99.300 ;
        RECT 131.010 99.100 131.330 99.160 ;
        RECT 118.220 98.960 131.330 99.100 ;
        RECT 131.010 98.900 131.330 98.960 ;
        RECT 135.625 99.100 135.915 99.145 ;
        RECT 136.530 99.100 136.850 99.160 ;
        RECT 135.625 98.960 136.850 99.100 ;
        RECT 135.625 98.915 135.915 98.960 ;
        RECT 136.530 98.900 136.850 98.960 ;
        RECT 137.030 99.100 137.320 99.145 ;
        RECT 139.130 99.100 139.420 99.145 ;
        RECT 140.700 99.100 140.990 99.145 ;
        RECT 137.030 98.960 140.990 99.100 ;
        RECT 137.030 98.915 137.320 98.960 ;
        RECT 139.130 98.915 139.420 98.960 ;
        RECT 140.700 98.915 140.990 98.960 ;
        RECT 27.050 98.620 28.200 98.760 ;
        RECT 79.490 98.760 79.810 98.820 ;
        RECT 83.170 98.760 83.490 98.820 ;
        RECT 89.610 98.760 89.930 98.820 ;
        RECT 94.670 98.760 94.990 98.820 ;
        RECT 79.490 98.620 94.990 98.760 ;
        RECT 27.050 98.560 27.370 98.620 ;
        RECT 79.490 98.560 79.810 98.620 ;
        RECT 83.170 98.560 83.490 98.620 ;
        RECT 89.610 98.560 89.930 98.620 ;
        RECT 94.670 98.560 94.990 98.620 ;
        RECT 109.390 98.560 109.710 98.820 ;
        RECT 111.690 98.760 112.010 98.820 ;
        RECT 129.630 98.760 129.950 98.820 ;
        RECT 111.690 98.620 129.950 98.760 ;
        RECT 111.690 98.560 112.010 98.620 ;
        RECT 129.630 98.560 129.950 98.620 ;
        RECT 144.810 98.560 145.130 98.820 ;
        RECT 17.320 97.940 147.040 98.420 ;
        RECT 24.750 97.740 25.070 97.800 ;
        RECT 27.985 97.740 28.275 97.785 ;
        RECT 24.750 97.600 28.275 97.740 ;
        RECT 24.750 97.540 25.070 97.600 ;
        RECT 27.985 97.555 28.275 97.600 ;
        RECT 29.825 97.555 30.115 97.785 ;
        RECT 30.745 97.740 31.035 97.785 ;
        RECT 31.190 97.740 31.510 97.800 ;
        RECT 30.745 97.600 31.510 97.740 ;
        RECT 30.745 97.555 31.035 97.600 ;
        RECT 21.990 97.400 22.280 97.445 ;
        RECT 23.560 97.400 23.850 97.445 ;
        RECT 25.660 97.400 25.950 97.445 ;
        RECT 21.990 97.260 25.950 97.400 ;
        RECT 29.900 97.400 30.040 97.555 ;
        RECT 31.190 97.540 31.510 97.600 ;
        RECT 35.805 97.740 36.095 97.785 ;
        RECT 74.445 97.740 74.735 97.785 ;
        RECT 94.210 97.740 94.530 97.800 ;
        RECT 114.450 97.740 114.770 97.800 ;
        RECT 35.805 97.600 36.480 97.740 ;
        RECT 35.805 97.555 36.095 97.600 ;
        RECT 35.330 97.400 35.650 97.460 ;
        RECT 29.900 97.260 35.650 97.400 ;
        RECT 21.990 97.215 22.280 97.260 ;
        RECT 23.560 97.215 23.850 97.260 ;
        RECT 25.660 97.215 25.950 97.260 ;
        RECT 35.330 97.200 35.650 97.260 ;
        RECT 21.555 97.060 21.845 97.105 ;
        RECT 24.075 97.060 24.365 97.105 ;
        RECT 25.265 97.060 25.555 97.105 ;
        RECT 34.885 97.060 35.175 97.105 ;
        RECT 21.555 96.920 25.555 97.060 ;
        RECT 21.555 96.875 21.845 96.920 ;
        RECT 24.075 96.875 24.365 96.920 ;
        RECT 25.265 96.875 25.555 96.920 ;
        RECT 28.980 96.920 35.175 97.060 ;
        RECT 26.145 96.720 26.435 96.765 ;
        RECT 27.050 96.720 27.370 96.780 ;
        RECT 26.145 96.580 27.370 96.720 ;
        RECT 26.145 96.535 26.435 96.580 ;
        RECT 27.050 96.520 27.370 96.580 ;
        RECT 27.970 96.720 28.290 96.780 ;
        RECT 28.980 96.765 29.120 96.920 ;
        RECT 28.905 96.720 29.195 96.765 ;
        RECT 27.970 96.580 29.195 96.720 ;
        RECT 27.970 96.520 28.290 96.580 ;
        RECT 28.905 96.535 29.195 96.580 ;
        RECT 29.810 96.520 30.130 96.780 ;
        RECT 31.740 96.765 31.880 96.920 ;
        RECT 34.885 96.875 35.175 96.920 ;
        RECT 31.665 96.535 31.955 96.765 ;
        RECT 32.570 96.720 32.890 96.780 ;
        RECT 33.045 96.720 33.335 96.765 ;
        RECT 32.570 96.580 33.335 96.720 ;
        RECT 32.570 96.520 32.890 96.580 ;
        RECT 33.045 96.535 33.335 96.580 ;
        RECT 33.965 96.535 34.255 96.765 ;
        RECT 24.920 96.380 25.210 96.425 ;
        RECT 25.670 96.380 25.990 96.440 ;
        RECT 24.920 96.240 25.990 96.380 ;
        RECT 24.920 96.195 25.210 96.240 ;
        RECT 25.670 96.180 25.990 96.240 ;
        RECT 31.190 96.380 31.510 96.440 ;
        RECT 34.040 96.380 34.180 96.535 ;
        RECT 34.410 96.520 34.730 96.780 ;
        RECT 35.330 96.720 35.650 96.780 ;
        RECT 35.805 96.720 36.095 96.765 ;
        RECT 35.330 96.580 36.095 96.720 ;
        RECT 35.330 96.520 35.650 96.580 ;
        RECT 35.805 96.535 36.095 96.580 ;
        RECT 36.340 96.380 36.480 97.600 ;
        RECT 74.445 97.600 94.530 97.740 ;
        RECT 74.445 97.555 74.735 97.600 ;
        RECT 94.210 97.540 94.530 97.600 ;
        RECT 99.820 97.600 114.770 97.740 ;
        RECT 63.865 97.400 64.155 97.445 ;
        RECT 69.370 97.400 69.690 97.460 ;
        RECT 63.865 97.260 69.690 97.400 ;
        RECT 63.865 97.215 64.155 97.260 ;
        RECT 69.370 97.200 69.690 97.260 ;
        RECT 80.885 97.400 81.175 97.445 ;
        RECT 84.105 97.400 84.395 97.445 ;
        RECT 99.820 97.400 99.960 97.600 ;
        RECT 114.450 97.540 114.770 97.600 ;
        RECT 117.685 97.740 117.975 97.785 ;
        RECT 119.510 97.740 119.830 97.800 ;
        RECT 117.685 97.600 119.830 97.740 ;
        RECT 117.685 97.555 117.975 97.600 ;
        RECT 119.510 97.540 119.830 97.600 ;
        RECT 122.130 97.600 144.120 97.740 ;
        RECT 111.690 97.400 112.010 97.460 ;
        RECT 80.885 97.260 84.395 97.400 ;
        RECT 80.885 97.215 81.175 97.260 ;
        RECT 84.105 97.215 84.395 97.260 ;
        RECT 92.460 97.260 99.960 97.400 ;
        RECT 101.660 97.260 112.010 97.400 ;
        RECT 61.090 97.060 61.410 97.120 ;
        RECT 62.025 97.060 62.315 97.105 ;
        RECT 67.070 97.060 67.390 97.120 ;
        RECT 61.090 96.920 67.390 97.060 ;
        RECT 61.090 96.860 61.410 96.920 ;
        RECT 62.025 96.875 62.315 96.920 ;
        RECT 67.070 96.860 67.390 96.920 ;
        RECT 70.765 97.060 71.055 97.105 ;
        RECT 71.210 97.060 71.530 97.120 ;
        RECT 74.430 97.060 74.750 97.120 ;
        RECT 83.630 97.060 83.950 97.120 ;
        RECT 70.765 96.920 71.530 97.060 ;
        RECT 70.765 96.875 71.055 96.920 ;
        RECT 71.210 96.860 71.530 96.920 ;
        RECT 72.680 96.920 83.950 97.060 ;
        RECT 68.450 96.720 68.770 96.780 ;
        RECT 72.680 96.765 72.820 96.920 ;
        RECT 74.430 96.860 74.750 96.920 ;
        RECT 83.630 96.860 83.950 96.920 ;
        RECT 87.325 97.060 87.615 97.105 ;
        RECT 87.770 97.060 88.090 97.120 ;
        RECT 87.325 96.920 88.090 97.060 ;
        RECT 87.325 96.875 87.615 96.920 ;
        RECT 87.770 96.860 88.090 96.920 ;
        RECT 71.685 96.720 71.975 96.765 ;
        RECT 68.450 96.580 71.975 96.720 ;
        RECT 68.450 96.520 68.770 96.580 ;
        RECT 71.685 96.535 71.975 96.580 ;
        RECT 72.605 96.535 72.895 96.765 ;
        RECT 73.525 96.535 73.815 96.765 ;
        RECT 79.045 96.720 79.335 96.765 ;
        RECT 85.930 96.720 86.250 96.780 ;
        RECT 79.045 96.580 86.250 96.720 ;
        RECT 79.045 96.535 79.335 96.580 ;
        RECT 31.190 96.240 36.480 96.380 ;
        RECT 69.385 96.380 69.675 96.425 ;
        RECT 72.130 96.380 72.450 96.440 ;
        RECT 69.385 96.240 72.450 96.380 ;
        RECT 31.190 96.180 31.510 96.240 ;
        RECT 69.385 96.195 69.675 96.240 ;
        RECT 72.130 96.180 72.450 96.240 ;
        RECT 73.050 96.180 73.370 96.440 ;
        RECT 73.600 96.380 73.740 96.535 ;
        RECT 85.930 96.520 86.250 96.580 ;
        RECT 86.390 96.520 86.710 96.780 ;
        RECT 90.530 96.520 90.850 96.780 ;
        RECT 91.285 96.720 91.575 96.765 ;
        RECT 92.460 96.720 92.600 97.260 ;
        RECT 101.660 97.105 101.800 97.260 ;
        RECT 111.690 97.200 112.010 97.260 ;
        RECT 114.910 97.400 115.230 97.460 ;
        RECT 117.210 97.400 117.530 97.460 ;
        RECT 114.910 97.260 117.530 97.400 ;
        RECT 114.910 97.200 115.230 97.260 ;
        RECT 101.585 96.875 101.875 97.105 ;
        RECT 103.410 97.060 103.730 97.120 ;
        RECT 104.805 97.060 105.095 97.105 ;
        RECT 105.710 97.060 106.030 97.120 ;
        RECT 103.410 96.920 106.030 97.060 ;
        RECT 103.410 96.860 103.730 96.920 ;
        RECT 104.805 96.875 105.095 96.920 ;
        RECT 105.710 96.860 106.030 96.920 ;
        RECT 108.470 97.060 108.790 97.120 ;
        RECT 111.245 97.060 111.535 97.105 ;
        RECT 108.470 96.920 111.535 97.060 ;
        RECT 108.470 96.860 108.790 96.920 ;
        RECT 111.245 96.875 111.535 96.920 ;
        RECT 113.620 96.920 115.140 97.060 ;
        RECT 91.285 96.580 92.600 96.720 ;
        RECT 92.830 96.765 93.150 96.780 ;
        RECT 92.830 96.720 93.160 96.765 ;
        RECT 96.050 96.720 96.370 96.780 ;
        RECT 100.205 96.720 100.495 96.765 ;
        RECT 92.830 96.580 93.345 96.720 ;
        RECT 96.050 96.580 100.495 96.720 ;
        RECT 91.285 96.535 91.575 96.580 ;
        RECT 92.830 96.535 93.160 96.580 ;
        RECT 92.830 96.520 93.150 96.535 ;
        RECT 96.050 96.520 96.370 96.580 ;
        RECT 100.205 96.535 100.495 96.580 ;
        RECT 110.785 96.720 111.075 96.765 ;
        RECT 113.620 96.720 113.760 96.920 ;
        RECT 115.000 96.780 115.140 96.920 ;
        RECT 110.785 96.580 113.760 96.720 ;
        RECT 110.785 96.535 111.075 96.580 ;
        RECT 114.465 96.535 114.755 96.765 ;
        RECT 114.910 96.720 115.230 96.780 ;
        RECT 115.920 96.765 116.060 97.260 ;
        RECT 117.210 97.200 117.530 97.260 ;
        RECT 118.130 97.060 118.450 97.120 ;
        RECT 122.130 97.060 122.270 97.600 ;
        RECT 128.265 97.400 128.555 97.445 ;
        RECT 130.550 97.400 130.870 97.460 ;
        RECT 128.265 97.260 130.870 97.400 ;
        RECT 128.265 97.215 128.555 97.260 ;
        RECT 130.550 97.200 130.870 97.260 ;
        RECT 131.010 97.200 131.330 97.460 ;
        RECT 135.625 97.400 135.915 97.445 ;
        RECT 136.530 97.400 136.850 97.460 ;
        RECT 135.625 97.260 136.850 97.400 ;
        RECT 135.625 97.215 135.915 97.260 ;
        RECT 136.530 97.200 136.850 97.260 ;
        RECT 118.130 96.920 122.270 97.060 ;
        RECT 126.410 97.060 126.730 97.120 ;
        RECT 133.770 97.060 134.090 97.120 ;
        RECT 126.410 96.920 134.090 97.060 ;
        RECT 118.130 96.860 118.450 96.920 ;
        RECT 126.410 96.860 126.730 96.920 ;
        RECT 133.770 96.860 134.090 96.920 ;
        RECT 136.085 97.060 136.375 97.105 ;
        RECT 136.990 97.060 137.310 97.120 ;
        RECT 136.085 96.920 137.310 97.060 ;
        RECT 136.085 96.875 136.375 96.920 ;
        RECT 136.990 96.860 137.310 96.920 ;
        RECT 116.750 96.765 117.070 96.780 ;
        RECT 114.910 96.580 115.425 96.720 ;
        RECT 75.350 96.380 75.670 96.440 ;
        RECT 85.010 96.380 85.330 96.440 ;
        RECT 86.480 96.380 86.620 96.520 ;
        RECT 73.600 96.240 85.330 96.380 ;
        RECT 75.350 96.180 75.670 96.240 ;
        RECT 85.010 96.180 85.330 96.240 ;
        RECT 86.020 96.240 86.620 96.380 ;
        RECT 90.070 96.380 90.390 96.440 ;
        RECT 91.925 96.380 92.215 96.425 ;
        RECT 90.070 96.240 92.215 96.380 ;
        RECT 19.230 95.840 19.550 96.100 ;
        RECT 33.950 96.040 34.270 96.100 ;
        RECT 35.790 96.040 36.110 96.100 ;
        RECT 36.725 96.040 37.015 96.085 ;
        RECT 33.950 95.900 37.015 96.040 ;
        RECT 33.950 95.840 34.270 95.900 ;
        RECT 35.790 95.840 36.110 95.900 ;
        RECT 36.725 95.855 37.015 95.900 ;
        RECT 64.310 95.840 64.630 96.100 ;
        RECT 67.070 96.040 67.390 96.100 ;
        RECT 67.545 96.040 67.835 96.085 ;
        RECT 67.070 95.900 67.835 96.040 ;
        RECT 67.070 95.840 67.390 95.900 ;
        RECT 67.545 95.855 67.835 95.900 ;
        RECT 68.910 96.040 69.230 96.100 ;
        RECT 69.845 96.040 70.135 96.085 ;
        RECT 68.910 95.900 70.135 96.040 ;
        RECT 68.910 95.840 69.230 95.900 ;
        RECT 69.845 95.855 70.135 95.900 ;
        RECT 81.345 96.040 81.635 96.085 ;
        RECT 81.790 96.040 82.110 96.100 ;
        RECT 86.020 96.085 86.160 96.240 ;
        RECT 90.070 96.180 90.390 96.240 ;
        RECT 91.925 96.195 92.215 96.240 ;
        RECT 92.385 96.195 92.675 96.425 ;
        RECT 99.730 96.380 100.050 96.440 ;
        RECT 93.840 96.240 100.050 96.380 ;
        RECT 81.345 95.900 82.110 96.040 ;
        RECT 81.345 95.855 81.635 95.900 ;
        RECT 81.790 95.840 82.110 95.900 ;
        RECT 85.945 95.855 86.235 96.085 ;
        RECT 86.405 96.040 86.695 96.085 ;
        RECT 87.310 96.040 87.630 96.100 ;
        RECT 92.460 96.040 92.600 96.195 ;
        RECT 93.840 96.085 93.980 96.240 ;
        RECT 99.730 96.180 100.050 96.240 ;
        RECT 103.870 96.380 104.190 96.440 ;
        RECT 113.070 96.380 113.390 96.440 ;
        RECT 103.870 96.240 113.390 96.380 ;
        RECT 103.870 96.180 104.190 96.240 ;
        RECT 113.070 96.180 113.390 96.240 ;
        RECT 86.405 95.900 92.600 96.040 ;
        RECT 86.405 95.855 86.695 95.900 ;
        RECT 87.310 95.840 87.630 95.900 ;
        RECT 93.765 95.855 94.055 96.085 ;
        RECT 96.510 96.040 96.830 96.100 ;
        RECT 99.270 96.040 99.590 96.100 ;
        RECT 96.510 95.900 99.590 96.040 ;
        RECT 96.510 95.840 96.830 95.900 ;
        RECT 99.270 95.840 99.590 95.900 ;
        RECT 102.030 95.840 102.350 96.100 ;
        RECT 104.330 95.840 104.650 96.100 ;
        RECT 108.470 95.840 108.790 96.100 ;
        RECT 110.310 95.840 110.630 96.100 ;
        RECT 114.540 96.040 114.680 96.535 ;
        RECT 114.910 96.520 115.230 96.580 ;
        RECT 115.845 96.535 116.135 96.765 ;
        RECT 116.750 96.720 117.080 96.765 ;
        RECT 130.565 96.720 130.855 96.765 ;
        RECT 131.470 96.720 131.790 96.780 ;
        RECT 131.945 96.720 132.235 96.765 ;
        RECT 116.750 96.580 117.265 96.720 ;
        RECT 130.565 96.580 132.235 96.720 ;
        RECT 116.750 96.535 117.080 96.580 ;
        RECT 130.565 96.535 130.855 96.580 ;
        RECT 116.750 96.520 117.070 96.535 ;
        RECT 131.470 96.520 131.790 96.580 ;
        RECT 131.945 96.535 132.235 96.580 ;
        RECT 135.610 96.720 135.930 96.780 ;
        RECT 137.465 96.720 137.755 96.765 ;
        RECT 135.610 96.580 137.755 96.720 ;
        RECT 135.610 96.520 135.930 96.580 ;
        RECT 137.465 96.535 137.755 96.580 ;
        RECT 137.910 96.520 138.230 96.780 ;
        RECT 139.305 96.720 139.595 96.765 ;
        RECT 142.050 96.720 142.370 96.780 ;
        RECT 143.980 96.765 144.120 97.600 ;
        RECT 139.305 96.580 142.370 96.720 ;
        RECT 139.305 96.535 139.595 96.580 ;
        RECT 142.050 96.520 142.370 96.580 ;
        RECT 143.905 96.535 144.195 96.765 ;
        RECT 116.305 96.195 116.595 96.425 ;
        RECT 115.370 96.040 115.690 96.100 ;
        RECT 114.540 95.900 115.690 96.040 ;
        RECT 116.380 96.040 116.520 96.195 ;
        RECT 129.630 96.180 129.950 96.440 ;
        RECT 138.370 96.180 138.690 96.440 ;
        RECT 147.110 96.380 147.430 96.440 ;
        RECT 143.060 96.240 147.430 96.380 ;
        RECT 116.750 96.040 117.070 96.100 ;
        RECT 116.380 95.900 117.070 96.040 ;
        RECT 115.370 95.840 115.690 95.900 ;
        RECT 116.750 95.840 117.070 95.900 ;
        RECT 128.710 95.840 129.030 96.100 ;
        RECT 136.545 96.040 136.835 96.085 ;
        RECT 141.130 96.040 141.450 96.100 ;
        RECT 143.060 96.085 143.200 96.240 ;
        RECT 147.110 96.180 147.430 96.240 ;
        RECT 136.545 95.900 141.450 96.040 ;
        RECT 136.545 95.855 136.835 95.900 ;
        RECT 141.130 95.840 141.450 95.900 ;
        RECT 142.985 95.855 143.275 96.085 ;
        RECT 144.825 96.040 145.115 96.085 ;
        RECT 150.330 96.040 150.650 96.100 ;
        RECT 144.825 95.900 150.650 96.040 ;
        RECT 144.825 95.855 145.115 95.900 ;
        RECT 150.330 95.840 150.650 95.900 ;
        RECT 17.320 95.220 147.040 95.700 ;
        RECT 25.670 95.020 25.990 95.080 ;
        RECT 26.145 95.020 26.435 95.065 ;
        RECT 25.670 94.880 26.435 95.020 ;
        RECT 25.670 94.820 25.990 94.880 ;
        RECT 26.145 94.835 26.435 94.880 ;
        RECT 68.465 94.835 68.755 95.065 ;
        RECT 24.305 94.680 24.595 94.725 ;
        RECT 20.240 94.540 24.595 94.680 ;
        RECT 19.230 94.340 19.550 94.400 ;
        RECT 20.240 94.385 20.380 94.540 ;
        RECT 24.305 94.495 24.595 94.540 ;
        RECT 28.890 94.480 29.210 94.740 ;
        RECT 35.330 94.680 35.650 94.740 ;
        RECT 33.120 94.540 35.650 94.680 ;
        RECT 20.165 94.340 20.455 94.385 ;
        RECT 19.230 94.200 20.455 94.340 ;
        RECT 19.230 94.140 19.550 94.200 ;
        RECT 20.165 94.155 20.455 94.200 ;
        RECT 21.990 94.140 22.310 94.400 ;
        RECT 23.830 94.140 24.150 94.400 ;
        RECT 25.670 94.340 25.990 94.400 ;
        RECT 28.445 94.340 28.735 94.385 ;
        RECT 25.670 94.200 28.735 94.340 ;
        RECT 28.980 94.340 29.120 94.480 ;
        RECT 31.190 94.340 31.510 94.400 ;
        RECT 28.980 94.200 31.510 94.340 ;
        RECT 25.670 94.140 25.990 94.200 ;
        RECT 28.445 94.155 28.735 94.200 ;
        RECT 31.190 94.140 31.510 94.200 ;
        RECT 32.110 94.340 32.430 94.400 ;
        RECT 33.120 94.340 33.260 94.540 ;
        RECT 35.330 94.480 35.650 94.540 ;
        RECT 35.805 94.680 36.095 94.725 ;
        RECT 36.710 94.680 37.030 94.740 ;
        RECT 61.090 94.680 61.410 94.740 ;
        RECT 62.900 94.680 63.190 94.725 ;
        RECT 64.310 94.680 64.630 94.740 ;
        RECT 35.805 94.540 42.000 94.680 ;
        RECT 35.805 94.495 36.095 94.540 ;
        RECT 36.710 94.480 37.030 94.540 ;
        RECT 32.110 94.200 33.260 94.340 ;
        RECT 32.110 94.140 32.430 94.200 ;
        RECT 33.490 94.140 33.810 94.400 ;
        RECT 37.645 94.340 37.935 94.385 ;
        RECT 38.550 94.340 38.870 94.400 ;
        RECT 37.645 94.200 38.870 94.340 ;
        RECT 37.645 94.155 37.935 94.200 ;
        RECT 38.550 94.140 38.870 94.200 ;
        RECT 39.025 94.340 39.315 94.385 ;
        RECT 39.560 94.340 39.700 94.540 ;
        RECT 41.860 94.400 42.000 94.540 ;
        RECT 61.090 94.540 62.700 94.680 ;
        RECT 61.090 94.480 61.410 94.540 ;
        RECT 39.025 94.200 39.700 94.340 ;
        RECT 39.930 94.340 40.250 94.400 ;
        RECT 40.405 94.340 40.695 94.385 ;
        RECT 39.930 94.200 40.695 94.340 ;
        RECT 39.025 94.155 39.315 94.200 ;
        RECT 39.930 94.140 40.250 94.200 ;
        RECT 40.405 94.155 40.695 94.200 ;
        RECT 41.310 94.140 41.630 94.400 ;
        RECT 41.770 94.140 42.090 94.400 ;
        RECT 61.550 94.140 61.870 94.400 ;
        RECT 62.560 94.340 62.700 94.540 ;
        RECT 62.900 94.540 64.630 94.680 ;
        RECT 68.540 94.680 68.680 94.835 ;
        RECT 69.370 94.820 69.690 95.080 ;
        RECT 70.750 95.020 71.070 95.080 ;
        RECT 71.225 95.020 71.515 95.065 ;
        RECT 70.750 94.880 71.515 95.020 ;
        RECT 70.750 94.820 71.070 94.880 ;
        RECT 71.225 94.835 71.515 94.880 ;
        RECT 71.685 95.020 71.975 95.065 ;
        RECT 73.050 95.020 73.370 95.080 ;
        RECT 71.685 94.880 73.370 95.020 ;
        RECT 71.685 94.835 71.975 94.880 ;
        RECT 71.760 94.680 71.900 94.835 ;
        RECT 73.050 94.820 73.370 94.880 ;
        RECT 73.970 95.020 74.290 95.080 ;
        RECT 87.770 95.020 88.090 95.080 ;
        RECT 73.970 94.880 88.090 95.020 ;
        RECT 73.970 94.820 74.290 94.880 ;
        RECT 87.770 94.820 88.090 94.880 ;
        RECT 89.610 94.820 89.930 95.080 ;
        RECT 90.070 94.820 90.390 95.080 ;
        RECT 92.830 95.020 93.150 95.080 ;
        RECT 103.410 95.020 103.730 95.080 ;
        RECT 92.830 94.880 103.730 95.020 ;
        RECT 92.830 94.820 93.150 94.880 ;
        RECT 103.410 94.820 103.730 94.880 ;
        RECT 103.870 95.020 104.190 95.080 ;
        RECT 104.345 95.020 104.635 95.065 ;
        RECT 103.870 94.880 104.635 95.020 ;
        RECT 103.870 94.820 104.190 94.880 ;
        RECT 104.345 94.835 104.635 94.880 ;
        RECT 108.930 95.020 109.250 95.080 ;
        RECT 114.465 95.020 114.755 95.065 ;
        RECT 117.670 95.020 117.990 95.080 ;
        RECT 122.745 95.020 123.035 95.065 ;
        RECT 126.870 95.020 127.190 95.080 ;
        RECT 136.085 95.020 136.375 95.065 ;
        RECT 136.530 95.020 136.850 95.080 ;
        RECT 108.930 94.880 114.755 95.020 ;
        RECT 108.930 94.820 109.250 94.880 ;
        RECT 114.465 94.835 114.755 94.880 ;
        RECT 116.380 94.880 127.190 95.020 ;
        RECT 68.540 94.540 71.900 94.680 ;
        RECT 72.130 94.680 72.450 94.740 ;
        RECT 79.490 94.680 79.810 94.740 ;
        RECT 72.130 94.540 79.810 94.680 ;
        RECT 62.900 94.495 63.190 94.540 ;
        RECT 64.310 94.480 64.630 94.540 ;
        RECT 72.130 94.480 72.450 94.540 ;
        RECT 79.490 94.480 79.810 94.540 ;
        RECT 85.930 94.680 86.250 94.740 ;
        RECT 108.440 94.680 108.730 94.725 ;
        RECT 109.390 94.680 109.710 94.740 ;
        RECT 85.930 94.540 91.220 94.680 ;
        RECT 85.930 94.480 86.250 94.540 ;
        RECT 64.770 94.340 65.090 94.400 ;
        RECT 62.560 94.200 65.090 94.340 ;
        RECT 64.770 94.140 65.090 94.200 ;
        RECT 73.510 94.140 73.830 94.400 ;
        RECT 78.110 94.140 78.430 94.400 ;
        RECT 80.425 94.340 80.715 94.385 ;
        RECT 80.870 94.340 81.190 94.400 ;
        RECT 81.790 94.385 82.110 94.400 ;
        RECT 81.760 94.340 82.110 94.385 ;
        RECT 80.425 94.200 81.190 94.340 ;
        RECT 81.595 94.200 82.110 94.340 ;
        RECT 91.080 94.340 91.220 94.540 ;
        RECT 103.960 94.540 105.020 94.680 ;
        RECT 91.925 94.340 92.215 94.385 ;
        RECT 93.750 94.340 94.070 94.400 ;
        RECT 96.425 94.340 96.715 94.385 ;
        RECT 91.080 94.200 94.070 94.340 ;
        RECT 80.425 94.155 80.715 94.200 ;
        RECT 80.870 94.140 81.190 94.200 ;
        RECT 81.760 94.155 82.110 94.200 ;
        RECT 91.925 94.155 92.215 94.200 ;
        RECT 81.790 94.140 82.110 94.155 ;
        RECT 93.750 94.140 94.070 94.200 ;
        RECT 94.300 94.200 96.715 94.340 ;
        RECT 23.385 93.815 23.675 94.045 ;
        RECT 23.920 94.000 24.060 94.140 ;
        RECT 28.905 94.000 29.195 94.045 ;
        RECT 23.920 93.860 29.195 94.000 ;
        RECT 28.905 93.815 29.195 93.860 ;
        RECT 16.930 93.660 17.250 93.720 ;
        RECT 21.085 93.660 21.375 93.705 ;
        RECT 16.930 93.520 21.375 93.660 ;
        RECT 23.460 93.660 23.600 93.815 ;
        RECT 28.430 93.660 28.750 93.720 ;
        RECT 23.460 93.520 28.750 93.660 ;
        RECT 28.980 93.660 29.120 93.815 ;
        RECT 29.350 93.800 29.670 94.060 ;
        RECT 31.665 94.000 31.955 94.045 ;
        RECT 34.425 94.000 34.715 94.045 ;
        RECT 35.330 94.000 35.650 94.060 ;
        RECT 31.665 93.860 34.180 94.000 ;
        RECT 31.665 93.815 31.955 93.860 ;
        RECT 32.585 93.660 32.875 93.705 ;
        RECT 28.980 93.520 32.875 93.660 ;
        RECT 34.040 93.660 34.180 93.860 ;
        RECT 34.425 93.860 35.650 94.000 ;
        RECT 34.425 93.815 34.715 93.860 ;
        RECT 35.330 93.800 35.650 93.860 ;
        RECT 38.105 94.000 38.395 94.045 ;
        RECT 40.850 94.000 41.170 94.060 ;
        RECT 38.105 93.860 41.170 94.000 ;
        RECT 38.105 93.815 38.395 93.860 ;
        RECT 40.850 93.800 41.170 93.860 ;
        RECT 62.445 94.000 62.735 94.045 ;
        RECT 63.635 94.000 63.925 94.045 ;
        RECT 66.155 94.000 66.445 94.045 ;
        RECT 62.445 93.860 66.445 94.000 ;
        RECT 62.445 93.815 62.735 93.860 ;
        RECT 63.635 93.815 63.925 93.860 ;
        RECT 66.155 93.815 66.445 93.860 ;
        RECT 71.670 94.000 71.990 94.060 ;
        RECT 72.145 94.000 72.435 94.045 ;
        RECT 71.670 93.860 72.435 94.000 ;
        RECT 71.670 93.800 71.990 93.860 ;
        RECT 72.145 93.815 72.435 93.860 ;
        RECT 78.585 93.815 78.875 94.045 ;
        RECT 79.505 93.815 79.795 94.045 ;
        RECT 81.305 94.000 81.595 94.045 ;
        RECT 82.495 94.000 82.785 94.045 ;
        RECT 85.015 94.000 85.305 94.045 ;
        RECT 90.545 94.000 90.835 94.045 ;
        RECT 92.830 94.000 93.150 94.060 ;
        RECT 94.300 94.045 94.440 94.200 ;
        RECT 96.425 94.155 96.715 94.200 ;
        RECT 101.110 94.340 101.430 94.400 ;
        RECT 103.960 94.340 104.100 94.540 ;
        RECT 101.110 94.200 104.100 94.340 ;
        RECT 104.880 94.340 105.020 94.540 ;
        RECT 108.440 94.540 109.710 94.680 ;
        RECT 108.440 94.495 108.730 94.540 ;
        RECT 109.390 94.480 109.710 94.540 ;
        RECT 110.310 94.680 110.630 94.740 ;
        RECT 116.380 94.725 116.520 94.880 ;
        RECT 117.670 94.820 117.990 94.880 ;
        RECT 122.745 94.835 123.035 94.880 ;
        RECT 126.870 94.820 127.190 94.880 ;
        RECT 127.420 94.880 135.840 95.020 ;
        RECT 116.305 94.680 116.595 94.725 ;
        RECT 110.310 94.540 116.595 94.680 ;
        RECT 110.310 94.480 110.630 94.540 ;
        RECT 116.305 94.495 116.595 94.540 ;
        RECT 117.210 94.680 117.530 94.740 ;
        RECT 127.420 94.680 127.560 94.880 ;
        RECT 117.210 94.540 127.560 94.680 ;
        RECT 127.760 94.680 128.050 94.725 ;
        RECT 128.710 94.680 129.030 94.740 ;
        RECT 127.760 94.540 129.030 94.680 ;
        RECT 117.210 94.480 117.530 94.540 ;
        RECT 127.760 94.495 128.050 94.540 ;
        RECT 128.710 94.480 129.030 94.540 ;
        RECT 131.010 94.680 131.330 94.740 ;
        RECT 134.245 94.680 134.535 94.725 ;
        RECT 131.010 94.540 134.535 94.680 ;
        RECT 135.700 94.680 135.840 94.880 ;
        RECT 136.085 94.880 136.850 95.020 ;
        RECT 136.085 94.835 136.375 94.880 ;
        RECT 136.530 94.820 136.850 94.880 ;
        RECT 137.450 95.020 137.770 95.080 ;
        RECT 137.925 95.020 138.215 95.065 ;
        RECT 137.450 94.880 138.215 95.020 ;
        RECT 137.450 94.820 137.770 94.880 ;
        RECT 137.925 94.835 138.215 94.880 ;
        RECT 138.370 94.820 138.690 95.080 ;
        RECT 138.460 94.680 138.600 94.820 ;
        RECT 135.700 94.540 141.360 94.680 ;
        RECT 131.010 94.480 131.330 94.540 ;
        RECT 134.245 94.495 134.535 94.540 ;
        RECT 105.710 94.340 106.030 94.400 ;
        RECT 116.750 94.340 117.070 94.400 ;
        RECT 120.890 94.340 121.210 94.400 ;
        RECT 141.220 94.385 141.360 94.540 ;
        RECT 138.385 94.340 138.675 94.385 ;
        RECT 104.880 94.200 105.480 94.340 ;
        RECT 101.110 94.140 101.430 94.200 ;
        RECT 81.305 93.860 85.305 94.000 ;
        RECT 81.305 93.815 81.595 93.860 ;
        RECT 82.495 93.815 82.785 93.860 ;
        RECT 85.015 93.815 85.305 93.860 ;
        RECT 86.940 93.860 93.150 94.000 ;
        RECT 38.565 93.660 38.855 93.705 ;
        RECT 43.610 93.660 43.930 93.720 ;
        RECT 34.040 93.520 38.320 93.660 ;
        RECT 16.930 93.460 17.250 93.520 ;
        RECT 21.085 93.475 21.375 93.520 ;
        RECT 28.430 93.460 28.750 93.520 ;
        RECT 32.585 93.475 32.875 93.520 ;
        RECT 38.180 93.380 38.320 93.520 ;
        RECT 38.565 93.520 43.930 93.660 ;
        RECT 38.565 93.475 38.855 93.520 ;
        RECT 43.610 93.460 43.930 93.520 ;
        RECT 59.725 93.475 60.015 93.705 ;
        RECT 62.050 93.660 62.340 93.705 ;
        RECT 64.150 93.660 64.440 93.705 ;
        RECT 65.720 93.660 66.010 93.705 ;
        RECT 62.050 93.520 66.010 93.660 ;
        RECT 62.050 93.475 62.340 93.520 ;
        RECT 64.150 93.475 64.440 93.520 ;
        RECT 65.720 93.475 66.010 93.520 ;
        RECT 75.365 93.660 75.655 93.705 ;
        RECT 76.285 93.660 76.575 93.705 ;
        RECT 75.365 93.520 76.575 93.660 ;
        RECT 75.365 93.475 75.655 93.520 ;
        RECT 76.285 93.475 76.575 93.520 ;
        RECT 78.110 93.660 78.430 93.720 ;
        RECT 78.660 93.660 78.800 93.815 ;
        RECT 78.110 93.520 78.800 93.660 ;
        RECT 18.310 93.320 18.630 93.380 ;
        RECT 19.245 93.320 19.535 93.365 ;
        RECT 18.310 93.180 19.535 93.320 ;
        RECT 18.310 93.120 18.630 93.180 ;
        RECT 19.245 93.135 19.535 93.180 ;
        RECT 26.130 93.320 26.450 93.380 ;
        RECT 26.605 93.320 26.895 93.365 ;
        RECT 26.130 93.180 26.895 93.320 ;
        RECT 26.130 93.120 26.450 93.180 ;
        RECT 26.605 93.135 26.895 93.180 ;
        RECT 27.510 93.320 27.830 93.380 ;
        RECT 33.490 93.320 33.810 93.380 ;
        RECT 27.510 93.180 33.810 93.320 ;
        RECT 27.510 93.120 27.830 93.180 ;
        RECT 33.490 93.120 33.810 93.180 ;
        RECT 33.950 93.120 34.270 93.380 ;
        RECT 34.870 93.320 35.190 93.380 ;
        RECT 36.725 93.320 37.015 93.365 ;
        RECT 34.870 93.180 37.015 93.320 ;
        RECT 34.870 93.120 35.190 93.180 ;
        RECT 36.725 93.135 37.015 93.180 ;
        RECT 38.090 93.120 38.410 93.380 ;
        RECT 41.325 93.320 41.615 93.365 ;
        RECT 44.530 93.320 44.850 93.380 ;
        RECT 41.325 93.180 44.850 93.320 ;
        RECT 41.325 93.135 41.615 93.180 ;
        RECT 44.530 93.120 44.850 93.180 ;
        RECT 58.790 93.120 59.110 93.380 ;
        RECT 59.800 93.320 59.940 93.475 ;
        RECT 78.110 93.460 78.430 93.520 ;
        RECT 66.150 93.320 66.470 93.380 ;
        RECT 59.800 93.180 66.470 93.320 ;
        RECT 66.150 93.120 66.470 93.180 ;
        RECT 75.810 93.120 76.130 93.380 ;
        RECT 79.580 93.320 79.720 93.815 ;
        RECT 80.910 93.660 81.200 93.705 ;
        RECT 83.010 93.660 83.300 93.705 ;
        RECT 84.580 93.660 84.870 93.705 ;
        RECT 80.910 93.520 84.870 93.660 ;
        RECT 80.910 93.475 81.200 93.520 ;
        RECT 83.010 93.475 83.300 93.520 ;
        RECT 84.580 93.475 84.870 93.520 ;
        RECT 85.470 93.320 85.790 93.380 ;
        RECT 86.940 93.320 87.080 93.860 ;
        RECT 90.545 93.815 90.835 93.860 ;
        RECT 92.830 93.800 93.150 93.860 ;
        RECT 94.225 93.815 94.515 94.045 ;
        RECT 95.130 93.800 95.450 94.060 ;
        RECT 105.340 94.045 105.480 94.200 ;
        RECT 105.710 94.200 112.380 94.340 ;
        RECT 105.710 94.140 106.030 94.200 ;
        RECT 96.025 94.000 96.315 94.045 ;
        RECT 97.215 94.000 97.505 94.045 ;
        RECT 99.735 94.000 100.025 94.045 ;
        RECT 96.025 93.860 100.025 94.000 ;
        RECT 96.025 93.815 96.315 93.860 ;
        RECT 97.215 93.815 97.505 93.860 ;
        RECT 99.735 93.815 100.025 93.860 ;
        RECT 104.805 93.815 105.095 94.045 ;
        RECT 105.265 93.815 105.555 94.045 ;
        RECT 93.305 93.475 93.595 93.705 ;
        RECT 95.630 93.660 95.920 93.705 ;
        RECT 97.730 93.660 98.020 93.705 ;
        RECT 99.300 93.660 99.590 93.705 ;
        RECT 102.505 93.660 102.795 93.705 ;
        RECT 95.630 93.520 99.590 93.660 ;
        RECT 95.630 93.475 95.920 93.520 ;
        RECT 97.730 93.475 98.020 93.520 ;
        RECT 99.300 93.475 99.590 93.520 ;
        RECT 99.820 93.520 102.795 93.660 ;
        RECT 79.580 93.180 87.080 93.320 ;
        RECT 85.470 93.120 85.790 93.180 ;
        RECT 87.310 93.120 87.630 93.380 ;
        RECT 87.770 93.120 88.090 93.380 ;
        RECT 93.380 93.320 93.520 93.475 ;
        RECT 99.820 93.320 99.960 93.520 ;
        RECT 102.505 93.475 102.795 93.520 ;
        RECT 93.380 93.180 99.960 93.320 ;
        RECT 102.045 93.320 102.335 93.365 ;
        RECT 102.950 93.320 103.270 93.380 ;
        RECT 104.880 93.320 105.020 93.815 ;
        RECT 107.090 93.800 107.410 94.060 ;
        RECT 107.985 94.000 108.275 94.045 ;
        RECT 109.175 94.000 109.465 94.045 ;
        RECT 111.695 94.000 111.985 94.045 ;
        RECT 107.985 93.860 111.985 94.000 ;
        RECT 112.240 94.000 112.380 94.200 ;
        RECT 116.750 94.200 121.210 94.340 ;
        RECT 116.750 94.140 117.070 94.200 ;
        RECT 120.890 94.140 121.210 94.200 ;
        RECT 126.040 94.200 136.755 94.340 ;
        RECT 117.685 94.000 117.975 94.045 ;
        RECT 112.240 93.860 117.975 94.000 ;
        RECT 107.985 93.815 108.275 93.860 ;
        RECT 109.175 93.815 109.465 93.860 ;
        RECT 111.695 93.815 111.985 93.860 ;
        RECT 117.685 93.815 117.975 93.860 ;
        RECT 123.205 94.000 123.495 94.045 ;
        RECT 123.650 94.000 123.970 94.060 ;
        RECT 123.205 93.860 123.970 94.000 ;
        RECT 123.205 93.815 123.495 93.860 ;
        RECT 107.590 93.660 107.880 93.705 ;
        RECT 109.690 93.660 109.980 93.705 ;
        RECT 111.260 93.660 111.550 93.705 ;
        RECT 107.590 93.520 111.550 93.660 ;
        RECT 107.590 93.475 107.880 93.520 ;
        RECT 109.690 93.475 109.980 93.520 ;
        RECT 111.260 93.475 111.550 93.520 ;
        RECT 114.005 93.660 114.295 93.705 ;
        RECT 116.750 93.660 117.070 93.720 ;
        RECT 114.005 93.520 117.070 93.660 ;
        RECT 117.760 93.660 117.900 93.815 ;
        RECT 123.650 93.800 123.970 93.860 ;
        RECT 124.125 94.000 124.415 94.045 ;
        RECT 124.570 94.000 124.890 94.060 ;
        RECT 124.125 93.860 124.890 94.000 ;
        RECT 124.125 93.815 124.415 93.860 ;
        RECT 124.570 93.800 124.890 93.860 ;
        RECT 126.040 93.660 126.180 94.200 ;
        RECT 126.425 93.815 126.715 94.045 ;
        RECT 127.305 94.000 127.595 94.045 ;
        RECT 128.495 94.000 128.785 94.045 ;
        RECT 131.015 94.000 131.305 94.045 ;
        RECT 127.305 93.860 131.305 94.000 ;
        RECT 127.305 93.815 127.595 93.860 ;
        RECT 128.495 93.815 128.785 93.860 ;
        RECT 131.015 93.815 131.305 93.860 ;
        RECT 133.770 94.000 134.090 94.060 ;
        RECT 135.165 94.000 135.455 94.045 ;
        RECT 133.770 93.860 135.455 94.000 ;
        RECT 117.760 93.520 126.180 93.660 ;
        RECT 114.005 93.475 114.295 93.520 ;
        RECT 116.750 93.460 117.070 93.520 ;
        RECT 102.045 93.180 105.020 93.320 ;
        RECT 116.290 93.320 116.610 93.380 ;
        RECT 120.905 93.320 121.195 93.365 ;
        RECT 116.290 93.180 121.195 93.320 ;
        RECT 126.500 93.320 126.640 93.815 ;
        RECT 133.770 93.800 134.090 93.860 ;
        RECT 135.165 93.815 135.455 93.860 ;
        RECT 126.910 93.660 127.200 93.705 ;
        RECT 129.010 93.660 129.300 93.705 ;
        RECT 130.580 93.660 130.870 93.705 ;
        RECT 136.070 93.660 136.390 93.720 ;
        RECT 126.910 93.520 130.870 93.660 ;
        RECT 126.910 93.475 127.200 93.520 ;
        RECT 129.010 93.475 129.300 93.520 ;
        RECT 130.580 93.475 130.870 93.520 ;
        RECT 131.100 93.520 136.390 93.660 ;
        RECT 136.615 93.660 136.755 94.200 ;
        RECT 138.385 94.200 140.900 94.340 ;
        RECT 138.385 94.155 138.675 94.200 ;
        RECT 139.290 93.800 139.610 94.060 ;
        RECT 140.760 94.000 140.900 94.200 ;
        RECT 141.145 94.155 141.435 94.385 ;
        RECT 141.605 94.155 141.895 94.385 ;
        RECT 141.680 94.000 141.820 94.155 ;
        RECT 142.050 94.140 142.370 94.400 ;
        RECT 142.985 94.340 143.275 94.385 ;
        RECT 143.890 94.340 144.210 94.400 ;
        RECT 142.985 94.200 144.210 94.340 ;
        RECT 142.985 94.155 143.275 94.200 ;
        RECT 143.890 94.140 144.210 94.200 ;
        RECT 140.760 93.860 141.820 94.000 ;
        RECT 141.220 93.720 141.360 93.860 ;
        RECT 139.750 93.660 140.070 93.720 ;
        RECT 136.615 93.520 140.070 93.660 ;
        RECT 131.100 93.320 131.240 93.520 ;
        RECT 136.070 93.460 136.390 93.520 ;
        RECT 139.750 93.460 140.070 93.520 ;
        RECT 141.130 93.460 141.450 93.720 ;
        RECT 126.500 93.180 131.240 93.320 ;
        RECT 102.045 93.135 102.335 93.180 ;
        RECT 102.950 93.120 103.270 93.180 ;
        RECT 116.290 93.120 116.610 93.180 ;
        RECT 120.905 93.135 121.195 93.180 ;
        RECT 133.310 93.120 133.630 93.380 ;
        RECT 137.450 93.320 137.770 93.380 ;
        RECT 140.225 93.320 140.515 93.365 ;
        RECT 137.450 93.180 140.515 93.320 ;
        RECT 137.450 93.120 137.770 93.180 ;
        RECT 140.225 93.135 140.515 93.180 ;
        RECT 144.350 93.320 144.670 93.380 ;
        RECT 144.825 93.320 145.115 93.365 ;
        RECT 144.350 93.180 145.115 93.320 ;
        RECT 144.350 93.120 144.670 93.180 ;
        RECT 144.825 93.135 145.115 93.180 ;
        RECT 17.320 92.500 147.040 92.980 ;
        RECT 31.665 92.300 31.955 92.345 ;
        RECT 32.110 92.300 32.430 92.360 ;
        RECT 42.230 92.300 42.550 92.360 ;
        RECT 61.550 92.300 61.870 92.360 ;
        RECT 31.665 92.160 32.430 92.300 ;
        RECT 31.665 92.115 31.955 92.160 ;
        RECT 32.110 92.100 32.430 92.160 ;
        RECT 36.340 92.160 42.550 92.300 ;
        RECT 22.030 91.960 22.320 92.005 ;
        RECT 24.130 91.960 24.420 92.005 ;
        RECT 25.700 91.960 25.990 92.005 ;
        RECT 22.030 91.820 25.990 91.960 ;
        RECT 22.030 91.775 22.320 91.820 ;
        RECT 24.130 91.775 24.420 91.820 ;
        RECT 25.700 91.775 25.990 91.820 ;
        RECT 22.425 91.620 22.715 91.665 ;
        RECT 23.615 91.620 23.905 91.665 ;
        RECT 26.135 91.620 26.425 91.665 ;
        RECT 35.330 91.620 35.650 91.680 ;
        RECT 22.425 91.480 26.425 91.620 ;
        RECT 22.425 91.435 22.715 91.480 ;
        RECT 23.615 91.435 23.905 91.480 ;
        RECT 26.135 91.435 26.425 91.480 ;
        RECT 32.200 91.480 35.650 91.620 ;
        RECT 32.200 91.340 32.340 91.480 ;
        RECT 21.545 91.280 21.835 91.325 ;
        RECT 27.050 91.280 27.370 91.340 ;
        RECT 21.545 91.140 27.370 91.280 ;
        RECT 21.545 91.095 21.835 91.140 ;
        RECT 27.050 91.080 27.370 91.140 ;
        RECT 27.510 91.280 27.830 91.340 ;
        RECT 28.905 91.280 29.195 91.325 ;
        RECT 27.510 91.140 29.195 91.280 ;
        RECT 27.510 91.080 27.830 91.140 ;
        RECT 28.905 91.095 29.195 91.140 ;
        RECT 29.825 91.280 30.115 91.325 ;
        RECT 32.110 91.280 32.430 91.340 ;
        RECT 29.825 91.140 32.430 91.280 ;
        RECT 29.825 91.095 30.115 91.140 ;
        RECT 32.110 91.080 32.430 91.140 ;
        RECT 32.570 91.080 32.890 91.340 ;
        RECT 33.950 91.080 34.270 91.340 ;
        RECT 34.960 91.325 35.100 91.480 ;
        RECT 35.330 91.420 35.650 91.480 ;
        RECT 36.340 91.325 36.480 92.160 ;
        RECT 42.230 92.100 42.550 92.160 ;
        RECT 57.960 92.160 61.870 92.300 ;
        RECT 41.310 91.760 41.630 92.020 ;
        RECT 48.210 91.760 48.530 92.020 ;
        RECT 39.025 91.620 39.315 91.665 ;
        RECT 37.720 91.480 39.315 91.620 ;
        RECT 37.720 91.325 37.860 91.480 ;
        RECT 39.025 91.435 39.315 91.480 ;
        RECT 39.470 91.620 39.790 91.680 ;
        RECT 41.400 91.620 41.540 91.760 ;
        RECT 57.960 91.665 58.100 92.160 ;
        RECT 61.550 92.100 61.870 92.160 ;
        RECT 64.785 92.300 65.075 92.345 ;
        RECT 68.450 92.300 68.770 92.360 ;
        RECT 71.210 92.300 71.530 92.360 ;
        RECT 85.025 92.300 85.315 92.345 ;
        RECT 90.530 92.300 90.850 92.360 ;
        RECT 64.785 92.160 71.530 92.300 ;
        RECT 64.785 92.115 65.075 92.160 ;
        RECT 68.450 92.100 68.770 92.160 ;
        RECT 71.210 92.100 71.530 92.160 ;
        RECT 71.760 92.160 82.480 92.300 ;
        RECT 58.370 91.960 58.660 92.005 ;
        RECT 60.470 91.960 60.760 92.005 ;
        RECT 62.040 91.960 62.330 92.005 ;
        RECT 58.370 91.820 62.330 91.960 ;
        RECT 58.370 91.775 58.660 91.820 ;
        RECT 60.470 91.775 60.760 91.820 ;
        RECT 62.040 91.775 62.330 91.820 ;
        RECT 65.730 91.960 66.020 92.005 ;
        RECT 67.830 91.960 68.120 92.005 ;
        RECT 69.400 91.960 69.690 92.005 ;
        RECT 65.730 91.820 69.690 91.960 ;
        RECT 65.730 91.775 66.020 91.820 ;
        RECT 67.830 91.775 68.120 91.820 ;
        RECT 69.400 91.775 69.690 91.820 ;
        RECT 48.685 91.620 48.975 91.665 ;
        RECT 39.470 91.480 42.460 91.620 ;
        RECT 39.470 91.420 39.790 91.480 ;
        RECT 34.885 91.095 35.175 91.325 ;
        RECT 36.265 91.095 36.555 91.325 ;
        RECT 37.645 91.095 37.935 91.325 ;
        RECT 38.565 91.095 38.855 91.325 ;
        RECT 39.945 91.280 40.235 91.325 ;
        RECT 40.390 91.280 40.710 91.340 ;
        RECT 42.320 91.325 42.460 91.480 ;
        RECT 45.080 91.480 48.975 91.620 ;
        RECT 45.080 91.325 45.220 91.480 ;
        RECT 48.685 91.435 48.975 91.480 ;
        RECT 57.885 91.435 58.175 91.665 ;
        RECT 58.765 91.620 59.055 91.665 ;
        RECT 59.955 91.620 60.245 91.665 ;
        RECT 62.475 91.620 62.765 91.665 ;
        RECT 58.765 91.480 62.765 91.620 ;
        RECT 58.765 91.435 59.055 91.480 ;
        RECT 59.955 91.435 60.245 91.480 ;
        RECT 62.475 91.435 62.765 91.480 ;
        RECT 66.125 91.620 66.415 91.665 ;
        RECT 67.315 91.620 67.605 91.665 ;
        RECT 69.835 91.620 70.125 91.665 ;
        RECT 66.125 91.480 70.125 91.620 ;
        RECT 66.125 91.435 66.415 91.480 ;
        RECT 67.315 91.435 67.605 91.480 ;
        RECT 69.835 91.435 70.125 91.480 ;
        RECT 39.945 91.140 40.710 91.280 ;
        RECT 39.945 91.095 40.235 91.140 ;
        RECT 22.880 90.940 23.170 90.985 ;
        RECT 26.590 90.940 26.910 91.000 ;
        RECT 22.880 90.800 26.910 90.940 ;
        RECT 22.880 90.755 23.170 90.800 ;
        RECT 26.590 90.740 26.910 90.800 ;
        RECT 33.490 90.940 33.810 91.000 ;
        RECT 36.710 90.940 37.030 91.000 ;
        RECT 33.490 90.800 37.030 90.940 ;
        RECT 38.640 90.940 38.780 91.095 ;
        RECT 40.390 91.080 40.710 91.140 ;
        RECT 41.325 91.095 41.615 91.325 ;
        RECT 42.245 91.095 42.535 91.325 ;
        RECT 43.625 91.095 43.915 91.325 ;
        RECT 45.005 91.095 45.295 91.325 ;
        RECT 45.925 91.280 46.215 91.325 ;
        RECT 46.830 91.280 47.150 91.340 ;
        RECT 45.925 91.140 47.150 91.280 ;
        RECT 45.925 91.095 46.215 91.140 ;
        RECT 40.850 90.940 41.170 91.000 ;
        RECT 38.640 90.800 41.170 90.940 ;
        RECT 41.400 90.940 41.540 91.095 ;
        RECT 42.705 90.940 42.995 90.985 ;
        RECT 41.400 90.800 42.995 90.940 ;
        RECT 33.490 90.740 33.810 90.800 ;
        RECT 36.710 90.740 37.030 90.800 ;
        RECT 40.850 90.740 41.170 90.800 ;
        RECT 42.705 90.755 42.995 90.800 ;
        RECT 28.430 90.400 28.750 90.660 ;
        RECT 29.365 90.600 29.655 90.645 ;
        RECT 31.190 90.600 31.510 90.660 ;
        RECT 29.365 90.460 31.510 90.600 ;
        RECT 29.365 90.415 29.655 90.460 ;
        RECT 31.190 90.400 31.510 90.460 ;
        RECT 35.330 90.400 35.650 90.660 ;
        RECT 39.930 90.600 40.250 90.660 ;
        RECT 43.700 90.600 43.840 91.095 ;
        RECT 46.830 91.080 47.150 91.140 ;
        RECT 59.220 91.095 59.510 91.325 ;
        RECT 61.550 91.280 61.870 91.340 ;
        RECT 65.245 91.280 65.535 91.325 ;
        RECT 61.550 91.140 65.535 91.280 ;
        RECT 46.385 90.755 46.675 90.985 ;
        RECT 58.790 90.940 59.110 91.000 ;
        RECT 59.340 90.940 59.480 91.095 ;
        RECT 61.550 91.080 61.870 91.140 ;
        RECT 65.245 91.095 65.535 91.140 ;
        RECT 68.450 91.280 68.770 91.340 ;
        RECT 70.290 91.280 70.610 91.340 ;
        RECT 71.760 91.280 71.900 92.160 ;
        RECT 74.930 91.960 75.220 92.005 ;
        RECT 77.030 91.960 77.320 92.005 ;
        RECT 78.600 91.960 78.890 92.005 ;
        RECT 74.930 91.820 78.890 91.960 ;
        RECT 74.930 91.775 75.220 91.820 ;
        RECT 77.030 91.775 77.320 91.820 ;
        RECT 78.600 91.775 78.890 91.820 ;
        RECT 75.325 91.620 75.615 91.665 ;
        RECT 76.515 91.620 76.805 91.665 ;
        RECT 79.035 91.620 79.325 91.665 ;
        RECT 75.325 91.480 79.325 91.620 ;
        RECT 75.325 91.435 75.615 91.480 ;
        RECT 76.515 91.435 76.805 91.480 ;
        RECT 79.035 91.435 79.325 91.480 ;
        RECT 68.450 91.140 71.900 91.280 ;
        RECT 72.605 91.280 72.895 91.325 ;
        RECT 73.050 91.280 73.370 91.340 ;
        RECT 72.605 91.140 73.370 91.280 ;
        RECT 68.450 91.080 68.770 91.140 ;
        RECT 70.290 91.080 70.610 91.140 ;
        RECT 72.605 91.095 72.895 91.140 ;
        RECT 73.050 91.080 73.370 91.140 ;
        RECT 74.445 91.280 74.735 91.325 ;
        RECT 80.870 91.280 81.190 91.340 ;
        RECT 82.340 91.325 82.480 92.160 ;
        RECT 85.025 92.160 90.850 92.300 ;
        RECT 85.025 92.115 85.315 92.160 ;
        RECT 90.530 92.100 90.850 92.160 ;
        RECT 92.370 92.300 92.690 92.360 ;
        RECT 94.225 92.300 94.515 92.345 ;
        RECT 92.370 92.160 94.515 92.300 ;
        RECT 92.370 92.100 92.690 92.160 ;
        RECT 94.225 92.115 94.515 92.160 ;
        RECT 102.965 92.300 103.255 92.345 ;
        RECT 104.330 92.300 104.650 92.360 ;
        RECT 102.965 92.160 104.650 92.300 ;
        RECT 102.965 92.115 103.255 92.160 ;
        RECT 104.330 92.100 104.650 92.160 ;
        RECT 106.630 92.100 106.950 92.360 ;
        RECT 123.650 92.300 123.970 92.360 ;
        RECT 125.950 92.300 126.270 92.360 ;
        RECT 129.645 92.300 129.935 92.345 ;
        RECT 136.070 92.300 136.390 92.360 ;
        RECT 123.650 92.160 129.935 92.300 ;
        RECT 123.650 92.100 123.970 92.160 ;
        RECT 125.950 92.100 126.270 92.160 ;
        RECT 129.645 92.115 129.935 92.160 ;
        RECT 134.320 92.160 136.390 92.300 ;
        RECT 87.810 91.960 88.100 92.005 ;
        RECT 89.910 91.960 90.200 92.005 ;
        RECT 91.480 91.960 91.770 92.005 ;
        RECT 82.845 91.820 87.540 91.960 ;
        RECT 74.445 91.140 81.190 91.280 ;
        RECT 74.445 91.095 74.735 91.140 ;
        RECT 80.870 91.080 81.190 91.140 ;
        RECT 82.265 91.095 82.555 91.325 ;
        RECT 58.790 90.800 59.480 90.940 ;
        RECT 66.580 90.940 66.870 90.985 ;
        RECT 67.990 90.940 68.310 91.000 ;
        RECT 66.580 90.800 68.310 90.940 ;
        RECT 39.930 90.460 43.840 90.600 ;
        RECT 45.910 90.600 46.230 90.660 ;
        RECT 46.460 90.600 46.600 90.755 ;
        RECT 58.790 90.740 59.110 90.800 ;
        RECT 66.580 90.755 66.870 90.800 ;
        RECT 67.990 90.740 68.310 90.800 ;
        RECT 69.830 90.940 70.150 91.000 ;
        RECT 75.810 90.985 76.130 91.000 ;
        RECT 75.780 90.940 76.130 90.985 ;
        RECT 69.830 90.800 73.740 90.940 ;
        RECT 75.615 90.800 76.130 90.940 ;
        RECT 80.960 90.940 81.100 91.080 ;
        RECT 82.845 91.000 82.985 91.820 ;
        RECT 85.010 91.620 85.330 91.680 ;
        RECT 87.400 91.665 87.540 91.820 ;
        RECT 87.810 91.820 91.770 91.960 ;
        RECT 87.810 91.775 88.100 91.820 ;
        RECT 89.910 91.775 90.200 91.820 ;
        RECT 91.480 91.775 91.770 91.820 ;
        RECT 93.750 91.960 94.070 92.020 ;
        RECT 94.685 91.960 94.975 92.005 ;
        RECT 93.750 91.820 94.975 91.960 ;
        RECT 93.750 91.760 94.070 91.820 ;
        RECT 94.685 91.775 94.975 91.820 ;
        RECT 96.550 91.960 96.840 92.005 ;
        RECT 98.650 91.960 98.940 92.005 ;
        RECT 100.220 91.960 100.510 92.005 ;
        RECT 105.250 91.960 105.570 92.020 ;
        RECT 108.510 91.960 108.800 92.005 ;
        RECT 110.610 91.960 110.900 92.005 ;
        RECT 112.180 91.960 112.470 92.005 ;
        RECT 96.550 91.820 100.510 91.960 ;
        RECT 96.550 91.775 96.840 91.820 ;
        RECT 98.650 91.775 98.940 91.820 ;
        RECT 100.220 91.775 100.510 91.820 ;
        RECT 102.580 91.820 105.940 91.960 ;
        RECT 83.260 91.480 85.330 91.620 ;
        RECT 83.260 91.325 83.400 91.480 ;
        RECT 85.010 91.420 85.330 91.480 ;
        RECT 87.325 91.435 87.615 91.665 ;
        RECT 88.205 91.620 88.495 91.665 ;
        RECT 89.395 91.620 89.685 91.665 ;
        RECT 91.915 91.620 92.205 91.665 ;
        RECT 88.205 91.480 92.205 91.620 ;
        RECT 88.205 91.435 88.495 91.480 ;
        RECT 89.395 91.435 89.685 91.480 ;
        RECT 91.915 91.435 92.205 91.480 ;
        RECT 95.130 91.620 95.450 91.680 ;
        RECT 96.065 91.620 96.355 91.665 ;
        RECT 95.130 91.480 96.355 91.620 ;
        RECT 95.130 91.420 95.450 91.480 ;
        RECT 96.065 91.435 96.355 91.480 ;
        RECT 96.945 91.620 97.235 91.665 ;
        RECT 98.135 91.620 98.425 91.665 ;
        RECT 100.655 91.620 100.945 91.665 ;
        RECT 96.945 91.480 100.945 91.620 ;
        RECT 96.945 91.435 97.235 91.480 ;
        RECT 98.135 91.435 98.425 91.480 ;
        RECT 100.655 91.435 100.945 91.480 ;
        RECT 83.185 91.095 83.475 91.325 ;
        RECT 84.105 91.095 84.395 91.325 ;
        RECT 82.710 90.940 83.030 91.000 ;
        RECT 80.960 90.800 83.030 90.940 ;
        RECT 69.830 90.740 70.150 90.800 ;
        RECT 45.910 90.460 46.600 90.600 ;
        RECT 39.930 90.400 40.250 90.460 ;
        RECT 45.910 90.400 46.230 90.460 ;
        RECT 72.130 90.400 72.450 90.660 ;
        RECT 73.600 90.645 73.740 90.800 ;
        RECT 75.780 90.755 76.130 90.800 ;
        RECT 75.810 90.740 76.130 90.755 ;
        RECT 82.710 90.740 83.030 90.800 ;
        RECT 83.645 90.755 83.935 90.985 ;
        RECT 73.525 90.415 73.815 90.645 ;
        RECT 78.110 90.600 78.430 90.660 ;
        RECT 81.345 90.600 81.635 90.645 ;
        RECT 83.720 90.600 83.860 90.755 ;
        RECT 78.110 90.460 83.860 90.600 ;
        RECT 84.180 90.600 84.320 91.095 ;
        RECT 95.590 91.080 95.910 91.340 ;
        RECT 102.580 91.280 102.720 91.820 ;
        RECT 105.250 91.760 105.570 91.820 ;
        RECT 102.950 91.620 103.270 91.680 ;
        RECT 102.950 91.480 104.100 91.620 ;
        RECT 102.950 91.420 103.270 91.480 ;
        RECT 103.960 91.325 104.100 91.480 ;
        RECT 103.425 91.280 103.715 91.325 ;
        RECT 97.060 91.140 102.720 91.280 ;
        RECT 103.040 91.140 103.715 91.280 ;
        RECT 88.660 90.940 88.950 90.985 ;
        RECT 89.610 90.940 89.930 91.000 ;
        RECT 93.290 90.940 93.610 91.000 ;
        RECT 97.060 90.940 97.200 91.140 ;
        RECT 88.660 90.800 89.930 90.940 ;
        RECT 88.660 90.755 88.950 90.800 ;
        RECT 89.610 90.740 89.930 90.800 ;
        RECT 90.620 90.800 97.200 90.940 ;
        RECT 97.400 90.940 97.690 90.985 ;
        RECT 101.570 90.940 101.890 91.000 ;
        RECT 97.400 90.800 101.890 90.940 ;
        RECT 89.150 90.600 89.470 90.660 ;
        RECT 90.620 90.600 90.760 90.800 ;
        RECT 93.290 90.740 93.610 90.800 ;
        RECT 97.400 90.755 97.690 90.800 ;
        RECT 101.570 90.740 101.890 90.800 ;
        RECT 84.180 90.460 90.760 90.600 ;
        RECT 94.210 90.600 94.530 90.660 ;
        RECT 103.040 90.600 103.180 91.140 ;
        RECT 103.425 91.095 103.715 91.140 ;
        RECT 103.890 91.095 104.180 91.325 ;
        RECT 104.330 91.280 104.650 91.340 ;
        RECT 105.800 91.325 105.940 91.820 ;
        RECT 108.510 91.820 112.470 91.960 ;
        RECT 108.510 91.775 108.800 91.820 ;
        RECT 110.610 91.775 110.900 91.820 ;
        RECT 112.180 91.775 112.470 91.820 ;
        RECT 115.870 91.960 116.160 92.005 ;
        RECT 117.970 91.960 118.260 92.005 ;
        RECT 119.540 91.960 119.830 92.005 ;
        RECT 115.870 91.820 119.830 91.960 ;
        RECT 115.870 91.775 116.160 91.820 ;
        RECT 117.970 91.775 118.260 91.820 ;
        RECT 119.540 91.775 119.830 91.820 ;
        RECT 123.230 91.960 123.520 92.005 ;
        RECT 125.330 91.960 125.620 92.005 ;
        RECT 126.900 91.960 127.190 92.005 ;
        RECT 123.230 91.820 127.190 91.960 ;
        RECT 123.230 91.775 123.520 91.820 ;
        RECT 125.330 91.775 125.620 91.820 ;
        RECT 126.900 91.775 127.190 91.820 ;
        RECT 131.010 91.760 131.330 92.020 ;
        RECT 108.905 91.620 109.195 91.665 ;
        RECT 110.095 91.620 110.385 91.665 ;
        RECT 112.615 91.620 112.905 91.665 ;
        RECT 108.905 91.480 112.905 91.620 ;
        RECT 108.905 91.435 109.195 91.480 ;
        RECT 110.095 91.435 110.385 91.480 ;
        RECT 112.615 91.435 112.905 91.480 ;
        RECT 116.265 91.620 116.555 91.665 ;
        RECT 117.455 91.620 117.745 91.665 ;
        RECT 119.975 91.620 120.265 91.665 ;
        RECT 116.265 91.480 120.265 91.620 ;
        RECT 116.265 91.435 116.555 91.480 ;
        RECT 117.455 91.435 117.745 91.480 ;
        RECT 119.975 91.435 120.265 91.480 ;
        RECT 123.625 91.620 123.915 91.665 ;
        RECT 124.815 91.620 125.105 91.665 ;
        RECT 127.335 91.620 127.625 91.665 ;
        RECT 123.625 91.480 127.625 91.620 ;
        RECT 123.625 91.435 123.915 91.480 ;
        RECT 124.815 91.435 125.105 91.480 ;
        RECT 127.335 91.435 127.625 91.480 ;
        RECT 132.405 91.620 132.695 91.665 ;
        RECT 133.770 91.620 134.090 91.680 ;
        RECT 134.320 91.665 134.460 92.160 ;
        RECT 136.070 92.100 136.390 92.160 ;
        RECT 141.130 92.100 141.450 92.360 ;
        RECT 134.730 91.960 135.020 92.005 ;
        RECT 136.830 91.960 137.120 92.005 ;
        RECT 138.400 91.960 138.690 92.005 ;
        RECT 134.730 91.820 138.690 91.960 ;
        RECT 134.730 91.775 135.020 91.820 ;
        RECT 136.830 91.775 137.120 91.820 ;
        RECT 138.400 91.775 138.690 91.820 ;
        RECT 132.405 91.480 134.090 91.620 ;
        RECT 132.405 91.435 132.695 91.480 ;
        RECT 133.770 91.420 134.090 91.480 ;
        RECT 134.245 91.435 134.535 91.665 ;
        RECT 135.125 91.620 135.415 91.665 ;
        RECT 136.315 91.620 136.605 91.665 ;
        RECT 138.835 91.620 139.125 91.665 ;
        RECT 135.125 91.480 139.125 91.620 ;
        RECT 135.125 91.435 135.415 91.480 ;
        RECT 136.315 91.435 136.605 91.480 ;
        RECT 138.835 91.435 139.125 91.480 ;
        RECT 144.825 91.620 145.115 91.665 ;
        RECT 145.270 91.620 145.590 91.680 ;
        RECT 144.825 91.480 145.590 91.620 ;
        RECT 144.825 91.435 145.115 91.480 ;
        RECT 145.270 91.420 145.590 91.480 ;
        RECT 105.265 91.280 105.555 91.325 ;
        RECT 104.330 91.140 105.555 91.280 ;
        RECT 104.330 91.080 104.650 91.140 ;
        RECT 105.265 91.095 105.555 91.140 ;
        RECT 105.750 91.095 106.040 91.325 ;
        RECT 107.090 91.280 107.410 91.340 ;
        RECT 108.025 91.280 108.315 91.325 ;
        RECT 115.385 91.280 115.675 91.325 ;
        RECT 122.730 91.280 123.050 91.340 ;
        RECT 107.090 91.140 123.050 91.280 ;
        RECT 107.090 91.080 107.410 91.140 ;
        RECT 108.025 91.095 108.315 91.140 ;
        RECT 115.385 91.095 115.675 91.140 ;
        RECT 122.730 91.080 123.050 91.140 ;
        RECT 135.580 91.280 135.870 91.325 ;
        RECT 136.990 91.280 137.310 91.340 ;
        RECT 135.580 91.140 137.310 91.280 ;
        RECT 135.580 91.095 135.870 91.140 ;
        RECT 136.990 91.080 137.310 91.140 ;
        RECT 104.790 90.740 105.110 91.000 ;
        RECT 107.550 90.940 107.870 91.000 ;
        RECT 109.250 90.940 109.540 90.985 ;
        RECT 107.550 90.800 109.540 90.940 ;
        RECT 107.550 90.740 107.870 90.800 ;
        RECT 109.250 90.755 109.540 90.800 ;
        RECT 115.830 90.940 116.150 91.000 ;
        RECT 124.110 90.985 124.430 91.000 ;
        RECT 116.610 90.940 116.900 90.985 ;
        RECT 115.830 90.800 116.900 90.940 ;
        RECT 115.830 90.740 116.150 90.800 ;
        RECT 116.610 90.755 116.900 90.800 ;
        RECT 124.080 90.755 124.430 90.985 ;
        RECT 143.445 90.940 143.735 90.985 ;
        RECT 124.110 90.740 124.430 90.755 ;
        RECT 138.000 90.800 143.735 90.940 ;
        RECT 138.000 90.660 138.140 90.800 ;
        RECT 143.445 90.755 143.735 90.800 ;
        RECT 94.210 90.460 103.180 90.600 ;
        RECT 113.070 90.600 113.390 90.660 ;
        RECT 114.910 90.600 115.230 90.660 ;
        RECT 113.070 90.460 115.230 90.600 ;
        RECT 78.110 90.400 78.430 90.460 ;
        RECT 81.345 90.415 81.635 90.460 ;
        RECT 89.150 90.400 89.470 90.460 ;
        RECT 94.210 90.400 94.530 90.460 ;
        RECT 113.070 90.400 113.390 90.460 ;
        RECT 114.910 90.400 115.230 90.460 ;
        RECT 118.130 90.600 118.450 90.660 ;
        RECT 122.285 90.600 122.575 90.645 ;
        RECT 118.130 90.460 122.575 90.600 ;
        RECT 118.130 90.400 118.450 90.460 ;
        RECT 122.285 90.415 122.575 90.460 ;
        RECT 130.090 90.400 130.410 90.660 ;
        RECT 132.850 90.600 133.170 90.660 ;
        RECT 137.910 90.600 138.230 90.660 ;
        RECT 132.850 90.460 138.230 90.600 ;
        RECT 132.850 90.400 133.170 90.460 ;
        RECT 137.910 90.400 138.230 90.460 ;
        RECT 141.590 90.400 141.910 90.660 ;
        RECT 143.890 90.400 144.210 90.660 ;
        RECT 17.320 89.780 147.040 90.260 ;
        RECT 19.245 89.580 19.535 89.625 ;
        RECT 25.670 89.580 25.990 89.640 ;
        RECT 19.245 89.440 25.990 89.580 ;
        RECT 19.245 89.395 19.535 89.440 ;
        RECT 25.670 89.380 25.990 89.440 ;
        RECT 26.590 89.380 26.910 89.640 ;
        RECT 28.430 89.380 28.750 89.640 ;
        RECT 28.905 89.580 29.195 89.625 ;
        RECT 30.730 89.580 31.050 89.640 ;
        RECT 31.665 89.580 31.955 89.625 ;
        RECT 28.905 89.440 31.955 89.580 ;
        RECT 28.905 89.395 29.195 89.440 ;
        RECT 30.730 89.380 31.050 89.440 ;
        RECT 31.665 89.395 31.955 89.440 ;
        RECT 33.950 89.580 34.270 89.640 ;
        RECT 33.950 89.440 34.640 89.580 ;
        RECT 33.950 89.380 34.270 89.440 ;
        RECT 24.920 89.240 25.210 89.285 ;
        RECT 26.130 89.240 26.450 89.300 ;
        RECT 24.920 89.100 26.450 89.240 ;
        RECT 24.920 89.055 25.210 89.100 ;
        RECT 26.130 89.040 26.450 89.100 ;
        RECT 27.510 89.240 27.830 89.300 ;
        RECT 34.500 89.240 34.640 89.440 ;
        RECT 41.770 89.380 42.090 89.640 ;
        RECT 43.610 89.380 43.930 89.640 ;
        RECT 48.210 89.580 48.530 89.640 ;
        RECT 57.425 89.580 57.715 89.625 ;
        RECT 48.210 89.440 57.715 89.580 ;
        RECT 48.210 89.380 48.530 89.440 ;
        RECT 57.425 89.395 57.715 89.440 ;
        RECT 67.530 89.580 67.850 89.640 ;
        RECT 68.910 89.580 69.230 89.640 ;
        RECT 67.530 89.440 69.230 89.580 ;
        RECT 67.530 89.380 67.850 89.440 ;
        RECT 68.910 89.380 69.230 89.440 ;
        RECT 71.685 89.580 71.975 89.625 ;
        RECT 72.130 89.580 72.450 89.640 ;
        RECT 71.685 89.440 72.450 89.580 ;
        RECT 71.685 89.395 71.975 89.440 ;
        RECT 72.130 89.380 72.450 89.440 ;
        RECT 76.285 89.580 76.575 89.625 ;
        RECT 91.450 89.580 91.770 89.640 ;
        RECT 94.225 89.580 94.515 89.625 ;
        RECT 76.285 89.440 91.220 89.580 ;
        RECT 76.285 89.395 76.575 89.440 ;
        RECT 34.885 89.240 35.175 89.285 ;
        RECT 27.510 89.100 34.180 89.240 ;
        RECT 34.500 89.100 35.175 89.240 ;
        RECT 27.510 89.040 27.830 89.100 ;
        RECT 31.190 88.900 31.510 88.960 ;
        RECT 33.045 88.900 33.335 88.945 ;
        RECT 31.190 88.760 33.335 88.900 ;
        RECT 31.190 88.700 31.510 88.760 ;
        RECT 33.045 88.715 33.335 88.760 ;
        RECT 33.490 88.700 33.810 88.960 ;
        RECT 34.040 88.920 34.180 89.100 ;
        RECT 34.885 89.055 35.175 89.100 ;
        RECT 35.330 89.240 35.650 89.300 ;
        RECT 61.550 89.240 61.870 89.300 ;
        RECT 35.330 89.100 37.400 89.240 ;
        RECT 35.330 89.040 35.650 89.100 ;
        RECT 37.260 88.945 37.400 89.100 ;
        RECT 38.180 89.100 41.540 89.240 ;
        RECT 34.040 88.850 34.640 88.920 ;
        RECT 35.805 88.900 36.095 88.945 ;
        RECT 34.960 88.850 36.095 88.900 ;
        RECT 34.040 88.780 36.095 88.850 ;
        RECT 34.500 88.760 36.095 88.780 ;
        RECT 34.500 88.710 35.100 88.760 ;
        RECT 35.805 88.715 36.095 88.760 ;
        RECT 37.185 88.715 37.475 88.945 ;
        RECT 37.630 88.900 37.950 88.960 ;
        RECT 38.180 88.945 38.320 89.100 ;
        RECT 38.105 88.900 38.395 88.945 ;
        RECT 37.630 88.760 38.395 88.900 ;
        RECT 37.630 88.700 37.950 88.760 ;
        RECT 38.105 88.715 38.395 88.760 ;
        RECT 38.550 88.700 38.870 88.960 ;
        RECT 39.470 88.700 39.790 88.960 ;
        RECT 40.850 88.700 41.170 88.960 ;
        RECT 41.400 88.945 41.540 89.100 ;
        RECT 60.720 89.100 61.870 89.240 ;
        RECT 41.325 88.715 41.615 88.945 ;
        RECT 42.230 88.700 42.550 88.960 ;
        RECT 44.530 88.700 44.850 88.960 ;
        RECT 45.910 88.700 46.230 88.960 ;
        RECT 56.950 88.900 57.270 88.960 ;
        RECT 60.720 88.945 60.860 89.100 ;
        RECT 61.550 89.040 61.870 89.100 ;
        RECT 62.010 88.945 62.330 88.960 ;
        RECT 58.345 88.900 58.635 88.945 ;
        RECT 56.950 88.760 58.635 88.900 ;
        RECT 56.950 88.700 57.270 88.760 ;
        RECT 58.345 88.715 58.635 88.760 ;
        RECT 60.645 88.715 60.935 88.945 ;
        RECT 61.980 88.715 62.330 88.945 ;
        RECT 71.225 88.900 71.515 88.945 ;
        RECT 71.670 88.900 71.990 88.960 ;
        RECT 71.225 88.760 71.990 88.900 ;
        RECT 72.220 88.900 72.360 89.380 ;
        RECT 74.430 89.040 74.750 89.300 ;
        RECT 84.980 89.240 85.270 89.285 ;
        RECT 85.930 89.240 86.250 89.300 ;
        RECT 84.980 89.100 86.250 89.240 ;
        RECT 84.980 89.055 85.270 89.100 ;
        RECT 85.930 89.040 86.250 89.100 ;
        RECT 73.510 88.900 73.830 88.960 ;
        RECT 72.220 88.760 73.830 88.900 ;
        RECT 71.225 88.715 71.515 88.760 ;
        RECT 62.010 88.700 62.330 88.715 ;
        RECT 71.670 88.700 71.990 88.760 ;
        RECT 73.510 88.700 73.830 88.760 ;
        RECT 74.905 88.715 75.195 88.945 ;
        RECT 21.555 88.560 21.845 88.605 ;
        RECT 24.075 88.560 24.365 88.605 ;
        RECT 25.265 88.560 25.555 88.605 ;
        RECT 21.555 88.420 25.555 88.560 ;
        RECT 21.555 88.375 21.845 88.420 ;
        RECT 24.075 88.375 24.365 88.420 ;
        RECT 25.265 88.375 25.555 88.420 ;
        RECT 26.145 88.560 26.435 88.605 ;
        RECT 27.050 88.560 27.370 88.620 ;
        RECT 26.145 88.420 27.370 88.560 ;
        RECT 26.145 88.375 26.435 88.420 ;
        RECT 27.050 88.360 27.370 88.420 ;
        RECT 29.350 88.360 29.670 88.620 ;
        RECT 32.585 88.375 32.875 88.605 ;
        RECT 33.965 88.560 34.255 88.605 ;
        RECT 35.330 88.560 35.650 88.620 ;
        RECT 33.965 88.420 35.650 88.560 ;
        RECT 33.965 88.375 34.255 88.420 ;
        RECT 21.990 88.220 22.280 88.265 ;
        RECT 23.560 88.220 23.850 88.265 ;
        RECT 25.660 88.220 25.950 88.265 ;
        RECT 21.990 88.080 25.950 88.220 ;
        RECT 32.660 88.220 32.800 88.375 ;
        RECT 35.330 88.360 35.650 88.420 ;
        RECT 36.250 88.560 36.570 88.620 ;
        RECT 38.640 88.560 38.780 88.700 ;
        RECT 39.945 88.560 40.235 88.605 ;
        RECT 40.390 88.560 40.710 88.620 ;
        RECT 36.250 88.420 40.710 88.560 ;
        RECT 36.250 88.360 36.570 88.420 ;
        RECT 39.945 88.375 40.235 88.420 ;
        RECT 40.390 88.360 40.710 88.420 ;
        RECT 61.525 88.560 61.815 88.605 ;
        RECT 62.715 88.560 63.005 88.605 ;
        RECT 65.235 88.560 65.525 88.605 ;
        RECT 72.590 88.560 72.910 88.620 ;
        RECT 73.970 88.560 74.290 88.620 ;
        RECT 61.525 88.420 65.525 88.560 ;
        RECT 72.395 88.420 74.290 88.560 ;
        RECT 61.525 88.375 61.815 88.420 ;
        RECT 62.715 88.375 63.005 88.420 ;
        RECT 65.235 88.375 65.525 88.420 ;
        RECT 72.590 88.360 72.910 88.420 ;
        RECT 73.970 88.360 74.290 88.420 ;
        RECT 38.565 88.220 38.855 88.265 ;
        RECT 32.660 88.080 38.855 88.220 ;
        RECT 21.990 88.035 22.280 88.080 ;
        RECT 23.560 88.035 23.850 88.080 ;
        RECT 25.660 88.035 25.950 88.080 ;
        RECT 38.565 88.035 38.855 88.080 ;
        RECT 61.130 88.220 61.420 88.265 ;
        RECT 63.230 88.220 63.520 88.265 ;
        RECT 64.800 88.220 65.090 88.265 ;
        RECT 61.130 88.080 65.090 88.220 ;
        RECT 61.130 88.035 61.420 88.080 ;
        RECT 63.230 88.035 63.520 88.080 ;
        RECT 64.800 88.035 65.090 88.080 ;
        RECT 68.910 88.220 69.230 88.280 ;
        RECT 74.980 88.220 75.120 88.715 ;
        RECT 75.350 88.700 75.670 88.960 ;
        RECT 82.710 88.900 83.030 88.960 ;
        RECT 91.080 88.945 91.220 89.440 ;
        RECT 91.450 89.440 92.600 89.580 ;
        RECT 91.450 89.380 91.770 89.440 ;
        RECT 92.460 89.285 92.600 89.440 ;
        RECT 94.225 89.440 101.340 89.580 ;
        RECT 94.225 89.395 94.515 89.440 ;
        RECT 92.385 89.240 92.675 89.285 ;
        RECT 101.200 89.240 101.340 89.440 ;
        RECT 101.570 89.380 101.890 89.640 ;
        RECT 107.105 89.580 107.395 89.625 ;
        RECT 107.550 89.580 107.870 89.640 ;
        RECT 107.105 89.440 107.870 89.580 ;
        RECT 107.105 89.395 107.395 89.440 ;
        RECT 107.550 89.380 107.870 89.440 ;
        RECT 114.925 89.580 115.215 89.625 ;
        RECT 115.830 89.580 116.150 89.640 ;
        RECT 114.925 89.440 116.150 89.580 ;
        RECT 114.925 89.395 115.215 89.440 ;
        RECT 115.830 89.380 116.150 89.440 ;
        RECT 117.670 89.380 117.990 89.640 ;
        RECT 118.130 89.380 118.450 89.640 ;
        RECT 130.550 89.580 130.870 89.640 ;
        RECT 131.025 89.580 131.315 89.625 ;
        RECT 130.550 89.440 131.315 89.580 ;
        RECT 130.550 89.380 130.870 89.440 ;
        RECT 131.025 89.395 131.315 89.440 ;
        RECT 132.850 89.380 133.170 89.640 ;
        RECT 133.310 89.580 133.630 89.640 ;
        RECT 135.150 89.580 135.470 89.640 ;
        RECT 139.750 89.580 140.070 89.640 ;
        RECT 133.310 89.440 135.470 89.580 ;
        RECT 133.310 89.380 133.630 89.440 ;
        RECT 135.150 89.380 135.470 89.440 ;
        RECT 137.080 89.440 140.070 89.580 ;
        RECT 110.770 89.240 111.090 89.300 ;
        RECT 92.385 89.100 98.120 89.240 ;
        RECT 101.200 89.100 111.090 89.240 ;
        RECT 92.385 89.055 92.675 89.100 ;
        RECT 83.645 88.900 83.935 88.945 ;
        RECT 82.710 88.760 83.935 88.900 ;
        RECT 82.710 88.700 83.030 88.760 ;
        RECT 83.645 88.715 83.935 88.760 ;
        RECT 91.005 88.715 91.295 88.945 ;
        RECT 91.745 88.900 92.035 88.945 ;
        RECT 91.745 88.760 92.600 88.900 ;
        RECT 91.745 88.715 92.035 88.760 ;
        RECT 92.460 88.620 92.600 88.760 ;
        RECT 92.830 88.700 93.150 88.960 ;
        RECT 93.290 88.945 93.610 88.960 ;
        RECT 93.290 88.900 93.620 88.945 ;
        RECT 94.670 88.900 94.990 88.960 ;
        RECT 96.985 88.900 97.275 88.945 ;
        RECT 93.290 88.760 93.805 88.900 ;
        RECT 94.670 88.760 97.275 88.900 ;
        RECT 93.290 88.715 93.620 88.760 ;
        RECT 93.290 88.700 93.610 88.715 ;
        RECT 94.670 88.700 94.990 88.760 ;
        RECT 96.985 88.715 97.275 88.760 ;
        RECT 84.525 88.560 84.815 88.605 ;
        RECT 85.715 88.560 86.005 88.605 ;
        RECT 88.235 88.560 88.525 88.605 ;
        RECT 84.525 88.420 88.525 88.560 ;
        RECT 84.525 88.375 84.815 88.420 ;
        RECT 85.715 88.375 86.005 88.420 ;
        RECT 88.235 88.375 88.525 88.420 ;
        RECT 92.370 88.360 92.690 88.620 ;
        RECT 93.750 88.560 94.070 88.620 ;
        RECT 97.430 88.560 97.750 88.620 ;
        RECT 93.750 88.420 97.750 88.560 ;
        RECT 93.750 88.360 94.070 88.420 ;
        RECT 97.430 88.360 97.750 88.420 ;
        RECT 68.910 88.080 75.120 88.220 ;
        RECT 84.130 88.220 84.420 88.265 ;
        RECT 86.230 88.220 86.520 88.265 ;
        RECT 87.800 88.220 88.090 88.265 ;
        RECT 84.130 88.080 88.090 88.220 ;
        RECT 68.910 88.020 69.230 88.080 ;
        RECT 84.130 88.035 84.420 88.080 ;
        RECT 86.230 88.035 86.520 88.080 ;
        RECT 87.800 88.035 88.090 88.080 ;
        RECT 90.070 88.220 90.390 88.280 ;
        RECT 90.545 88.220 90.835 88.265 ;
        RECT 90.070 88.080 90.835 88.220 ;
        RECT 90.070 88.020 90.390 88.080 ;
        RECT 90.545 88.035 90.835 88.080 ;
        RECT 32.570 87.880 32.890 87.940 ;
        RECT 36.710 87.880 37.030 87.940 ;
        RECT 32.570 87.740 37.030 87.880 ;
        RECT 32.570 87.680 32.890 87.740 ;
        RECT 36.710 87.680 37.030 87.740 ;
        RECT 39.010 87.880 39.330 87.940 ;
        RECT 39.485 87.880 39.775 87.925 ;
        RECT 39.010 87.740 39.775 87.880 ;
        RECT 39.010 87.680 39.330 87.740 ;
        RECT 39.485 87.695 39.775 87.740 ;
        RECT 45.465 87.880 45.755 87.925 ;
        RECT 46.830 87.880 47.150 87.940 ;
        RECT 48.670 87.880 48.990 87.940 ;
        RECT 45.465 87.740 48.990 87.880 ;
        RECT 45.465 87.695 45.755 87.740 ;
        RECT 46.830 87.680 47.150 87.740 ;
        RECT 48.670 87.680 48.990 87.740 ;
        RECT 69.370 87.680 69.690 87.940 ;
        RECT 95.130 87.680 95.450 87.940 ;
        RECT 97.980 87.880 98.120 89.100 ;
        RECT 110.770 89.040 111.090 89.100 ;
        RECT 112.610 89.040 112.930 89.300 ;
        RECT 122.730 89.240 123.050 89.300 ;
        RECT 122.730 89.100 136.760 89.240 ;
        RECT 122.730 89.040 123.050 89.100 ;
        RECT 99.270 88.700 99.590 88.960 ;
        RECT 98.365 88.560 98.655 88.605 ;
        RECT 100.650 88.560 100.970 88.620 ;
        RECT 98.365 88.420 100.970 88.560 ;
        RECT 98.365 88.375 98.655 88.420 ;
        RECT 100.650 88.360 100.970 88.420 ;
        RECT 104.805 88.560 105.095 88.605 ;
        RECT 112.700 88.560 112.840 89.040 ;
        RECT 123.740 88.945 123.880 89.100 ;
        RECT 136.620 88.960 136.760 89.100 ;
        RECT 123.665 88.715 123.955 88.945 ;
        RECT 125.000 88.900 125.290 88.945 ;
        RECT 130.090 88.900 130.410 88.960 ;
        RECT 125.000 88.760 130.410 88.900 ;
        RECT 125.000 88.715 125.290 88.760 ;
        RECT 130.090 88.700 130.410 88.760 ;
        RECT 136.070 88.700 136.390 88.960 ;
        RECT 136.530 88.700 136.850 88.960 ;
        RECT 113.530 88.560 113.850 88.620 ;
        RECT 104.805 88.420 113.850 88.560 ;
        RECT 104.805 88.375 105.095 88.420 ;
        RECT 113.530 88.360 113.850 88.420 ;
        RECT 119.050 88.360 119.370 88.620 ;
        RECT 124.545 88.560 124.835 88.605 ;
        RECT 125.735 88.560 126.025 88.605 ;
        RECT 128.255 88.560 128.545 88.605 ;
        RECT 124.545 88.420 128.545 88.560 ;
        RECT 124.545 88.375 124.835 88.420 ;
        RECT 125.735 88.375 126.025 88.420 ;
        RECT 128.255 88.375 128.545 88.420 ;
        RECT 134.245 88.560 134.535 88.605 ;
        RECT 137.080 88.560 137.220 89.440 ;
        RECT 139.750 89.380 140.070 89.440 ;
        RECT 143.445 89.580 143.735 89.625 ;
        RECT 143.890 89.580 144.210 89.640 ;
        RECT 143.445 89.440 144.210 89.580 ;
        RECT 143.445 89.395 143.735 89.440 ;
        RECT 143.890 89.380 144.210 89.440 ;
        RECT 141.130 89.240 141.450 89.300 ;
        RECT 141.130 89.100 144.120 89.240 ;
        RECT 141.130 89.040 141.450 89.100 ;
        RECT 137.880 88.900 138.170 88.945 ;
        RECT 139.750 88.900 140.070 88.960 ;
        RECT 143.980 88.945 144.120 89.100 ;
        RECT 137.880 88.760 140.070 88.900 ;
        RECT 137.880 88.715 138.170 88.760 ;
        RECT 139.750 88.700 140.070 88.760 ;
        RECT 143.905 88.715 144.195 88.945 ;
        RECT 134.245 88.420 137.220 88.560 ;
        RECT 137.425 88.560 137.715 88.605 ;
        RECT 138.615 88.560 138.905 88.605 ;
        RECT 141.135 88.560 141.425 88.605 ;
        RECT 137.425 88.420 141.425 88.560 ;
        RECT 134.245 88.375 134.535 88.420 ;
        RECT 137.425 88.375 137.715 88.420 ;
        RECT 138.615 88.375 138.905 88.420 ;
        RECT 141.135 88.375 141.425 88.420 ;
        RECT 101.125 88.220 101.415 88.265 ;
        RECT 102.030 88.220 102.350 88.280 ;
        RECT 101.125 88.080 102.350 88.220 ;
        RECT 101.125 88.035 101.415 88.080 ;
        RECT 102.030 88.020 102.350 88.080 ;
        RECT 106.645 88.220 106.935 88.265 ;
        RECT 108.470 88.220 108.790 88.280 ;
        RECT 106.645 88.080 108.790 88.220 ;
        RECT 106.645 88.035 106.935 88.080 ;
        RECT 108.470 88.020 108.790 88.080 ;
        RECT 114.465 88.220 114.755 88.265 ;
        RECT 115.845 88.220 116.135 88.265 ;
        RECT 114.465 88.080 116.135 88.220 ;
        RECT 114.465 88.035 114.755 88.080 ;
        RECT 115.845 88.035 116.135 88.080 ;
        RECT 124.150 88.220 124.440 88.265 ;
        RECT 126.250 88.220 126.540 88.265 ;
        RECT 127.820 88.220 128.110 88.265 ;
        RECT 124.150 88.080 128.110 88.220 ;
        RECT 124.150 88.035 124.440 88.080 ;
        RECT 126.250 88.035 126.540 88.080 ;
        RECT 127.820 88.035 128.110 88.080 ;
        RECT 129.170 88.220 129.490 88.280 ;
        RECT 130.090 88.220 130.410 88.280 ;
        RECT 129.170 88.080 130.410 88.220 ;
        RECT 129.170 88.020 129.490 88.080 ;
        RECT 130.090 88.020 130.410 88.080 ;
        RECT 130.565 88.220 130.855 88.265 ;
        RECT 131.470 88.220 131.790 88.280 ;
        RECT 130.565 88.080 131.790 88.220 ;
        RECT 130.565 88.035 130.855 88.080 ;
        RECT 131.470 88.020 131.790 88.080 ;
        RECT 133.770 88.220 134.090 88.280 ;
        RECT 136.530 88.220 136.850 88.280 ;
        RECT 133.770 88.080 136.850 88.220 ;
        RECT 133.770 88.020 134.090 88.080 ;
        RECT 136.530 88.020 136.850 88.080 ;
        RECT 137.030 88.220 137.320 88.265 ;
        RECT 139.130 88.220 139.420 88.265 ;
        RECT 140.700 88.220 140.990 88.265 ;
        RECT 137.030 88.080 140.990 88.220 ;
        RECT 137.030 88.035 137.320 88.080 ;
        RECT 139.130 88.035 139.420 88.080 ;
        RECT 140.700 88.035 140.990 88.080 ;
        RECT 104.790 87.880 105.110 87.940 ;
        RECT 97.980 87.740 105.110 87.880 ;
        RECT 104.790 87.680 105.110 87.740 ;
        RECT 129.630 87.880 129.950 87.940 ;
        RECT 135.165 87.880 135.455 87.925 ;
        RECT 129.630 87.740 135.455 87.880 ;
        RECT 129.630 87.680 129.950 87.740 ;
        RECT 135.165 87.695 135.455 87.740 ;
        RECT 144.810 87.680 145.130 87.940 ;
        RECT 17.320 87.060 147.040 87.540 ;
        RECT 26.145 86.860 26.435 86.905 ;
        RECT 28.890 86.860 29.210 86.920 ;
        RECT 26.145 86.720 29.210 86.860 ;
        RECT 26.145 86.675 26.435 86.720 ;
        RECT 28.890 86.660 29.210 86.720 ;
        RECT 29.810 86.860 30.130 86.920 ;
        RECT 32.125 86.860 32.415 86.905 ;
        RECT 29.810 86.720 32.415 86.860 ;
        RECT 29.810 86.660 30.130 86.720 ;
        RECT 32.125 86.675 32.415 86.720 ;
        RECT 33.580 86.720 36.020 86.860 ;
        RECT 21.085 86.520 21.375 86.565 ;
        RECT 24.765 86.520 25.055 86.565 ;
        RECT 33.580 86.520 33.720 86.720 ;
        RECT 21.085 86.380 24.520 86.520 ;
        RECT 21.085 86.335 21.375 86.380 ;
        RECT 15.090 86.180 15.410 86.240 ;
        RECT 24.380 86.180 24.520 86.380 ;
        RECT 24.765 86.380 33.720 86.520 ;
        RECT 33.965 86.520 34.255 86.565 ;
        RECT 34.870 86.520 35.190 86.580 ;
        RECT 33.965 86.380 35.190 86.520 ;
        RECT 35.880 86.520 36.020 86.720 ;
        RECT 36.250 86.660 36.570 86.920 ;
        RECT 36.710 86.860 37.030 86.920 ;
        RECT 39.025 86.860 39.315 86.905 ;
        RECT 39.470 86.860 39.790 86.920 ;
        RECT 36.710 86.720 38.780 86.860 ;
        RECT 36.710 86.660 37.030 86.720 ;
        RECT 37.630 86.520 37.950 86.580 ;
        RECT 35.880 86.380 37.950 86.520 ;
        RECT 24.765 86.335 25.055 86.380 ;
        RECT 33.965 86.335 34.255 86.380 ;
        RECT 34.870 86.320 35.190 86.380 ;
        RECT 37.630 86.320 37.950 86.380 ;
        RECT 38.090 86.320 38.410 86.580 ;
        RECT 38.640 86.520 38.780 86.720 ;
        RECT 39.025 86.720 39.790 86.860 ;
        RECT 39.025 86.675 39.315 86.720 ;
        RECT 39.470 86.660 39.790 86.720 ;
        RECT 40.850 86.860 41.170 86.920 ;
        RECT 41.325 86.860 41.615 86.905 ;
        RECT 44.545 86.860 44.835 86.905 ;
        RECT 40.850 86.720 41.615 86.860 ;
        RECT 40.850 86.660 41.170 86.720 ;
        RECT 41.325 86.675 41.615 86.720 ;
        RECT 41.860 86.720 44.835 86.860 ;
        RECT 41.860 86.520 42.000 86.720 ;
        RECT 44.545 86.675 44.835 86.720 ;
        RECT 48.670 86.860 48.990 86.920 ;
        RECT 54.205 86.860 54.495 86.905 ;
        RECT 48.670 86.720 54.495 86.860 ;
        RECT 48.670 86.660 48.990 86.720 ;
        RECT 54.205 86.675 54.495 86.720 ;
        RECT 62.010 86.660 62.330 86.920 ;
        RECT 67.990 86.660 68.310 86.920 ;
        RECT 85.930 86.660 86.250 86.920 ;
        RECT 89.610 86.660 89.930 86.920 ;
        RECT 115.370 86.860 115.690 86.920 ;
        RECT 117.225 86.860 117.515 86.905 ;
        RECT 115.370 86.720 117.515 86.860 ;
        RECT 115.370 86.660 115.690 86.720 ;
        RECT 117.225 86.675 117.515 86.720 ;
        RECT 119.970 86.860 120.290 86.920 ;
        RECT 125.950 86.860 126.270 86.920 ;
        RECT 119.970 86.720 126.270 86.860 ;
        RECT 119.970 86.660 120.290 86.720 ;
        RECT 125.950 86.660 126.270 86.720 ;
        RECT 130.105 86.860 130.395 86.905 ;
        RECT 131.010 86.860 131.330 86.920 ;
        RECT 130.105 86.720 131.330 86.860 ;
        RECT 130.105 86.675 130.395 86.720 ;
        RECT 131.010 86.660 131.330 86.720 ;
        RECT 133.785 86.860 134.075 86.905 ;
        RECT 138.830 86.860 139.150 86.920 ;
        RECT 133.785 86.720 139.150 86.860 ;
        RECT 133.785 86.675 134.075 86.720 ;
        RECT 138.830 86.660 139.150 86.720 ;
        RECT 139.750 86.660 140.070 86.920 ;
        RECT 38.640 86.380 42.000 86.520 ;
        RECT 42.230 86.520 42.550 86.580 ;
        RECT 50.985 86.520 51.275 86.565 ;
        RECT 42.230 86.380 51.275 86.520 ;
        RECT 42.230 86.320 42.550 86.380 ;
        RECT 50.985 86.335 51.275 86.380 ;
        RECT 56.965 86.520 57.255 86.565 ;
        RECT 60.170 86.520 60.490 86.580 ;
        RECT 56.965 86.380 60.490 86.520 ;
        RECT 56.965 86.335 57.255 86.380 ;
        RECT 60.170 86.320 60.490 86.380 ;
        RECT 62.945 86.520 63.235 86.565 ;
        RECT 67.070 86.520 67.390 86.580 ;
        RECT 62.945 86.380 67.390 86.520 ;
        RECT 62.945 86.335 63.235 86.380 ;
        RECT 67.070 86.320 67.390 86.380 ;
        RECT 67.545 86.520 67.835 86.565 ;
        RECT 69.370 86.520 69.690 86.580 ;
        RECT 67.545 86.380 69.690 86.520 ;
        RECT 67.545 86.335 67.835 86.380 ;
        RECT 69.370 86.320 69.690 86.380 ;
        RECT 85.485 86.520 85.775 86.565 ;
        RECT 87.770 86.520 88.090 86.580 ;
        RECT 85.485 86.380 88.090 86.520 ;
        RECT 85.485 86.335 85.775 86.380 ;
        RECT 87.770 86.320 88.090 86.380 ;
        RECT 89.165 86.520 89.455 86.565 ;
        RECT 95.130 86.520 95.450 86.580 ;
        RECT 89.165 86.380 95.450 86.520 ;
        RECT 89.165 86.335 89.455 86.380 ;
        RECT 95.130 86.320 95.450 86.380 ;
        RECT 95.590 86.520 95.910 86.580 ;
        RECT 97.905 86.520 98.195 86.565 ;
        RECT 95.590 86.380 98.195 86.520 ;
        RECT 95.590 86.320 95.910 86.380 ;
        RECT 97.905 86.335 98.195 86.380 ;
        RECT 113.530 86.520 113.850 86.580 ;
        RECT 115.845 86.520 116.135 86.565 ;
        RECT 116.290 86.520 116.610 86.580 ;
        RECT 113.530 86.380 114.220 86.520 ;
        RECT 113.530 86.320 113.850 86.380 ;
        RECT 38.180 86.180 38.320 86.320 ;
        RECT 71.670 86.180 71.990 86.240 ;
        RECT 15.090 86.040 24.060 86.180 ;
        RECT 24.380 86.040 34.180 86.180 ;
        RECT 15.090 85.980 15.410 86.040 ;
        RECT 18.310 85.840 18.630 85.900 ;
        RECT 23.920 85.885 24.060 86.040 ;
        RECT 18.785 85.840 19.075 85.885 ;
        RECT 18.310 85.700 19.075 85.840 ;
        RECT 18.310 85.640 18.630 85.700 ;
        RECT 18.785 85.655 19.075 85.700 ;
        RECT 20.165 85.655 20.455 85.885 ;
        RECT 23.385 85.655 23.675 85.885 ;
        RECT 23.845 85.655 24.135 85.885 ;
        RECT 24.750 85.840 25.070 85.900 ;
        RECT 25.225 85.840 25.515 85.885 ;
        RECT 24.750 85.700 25.515 85.840 ;
        RECT 11.870 85.500 12.190 85.560 ;
        RECT 20.240 85.500 20.380 85.655 ;
        RECT 23.460 85.500 23.600 85.655 ;
        RECT 24.750 85.640 25.070 85.700 ;
        RECT 25.225 85.655 25.515 85.700 ;
        RECT 28.430 85.640 28.750 85.900 ;
        RECT 30.745 85.840 31.035 85.885 ;
        RECT 31.190 85.840 31.510 85.900 ;
        RECT 30.745 85.700 31.510 85.840 ;
        RECT 30.745 85.655 31.035 85.700 ;
        RECT 31.190 85.640 31.510 85.700 ;
        RECT 33.045 85.655 33.335 85.885 ;
        RECT 25.670 85.500 25.990 85.560 ;
        RECT 11.870 85.360 20.380 85.500 ;
        RECT 21.160 85.360 23.140 85.500 ;
        RECT 23.460 85.360 25.990 85.500 ;
        RECT 11.870 85.300 12.190 85.360 ;
        RECT 19.705 85.160 19.995 85.205 ;
        RECT 21.160 85.160 21.300 85.360 ;
        RECT 19.705 85.020 21.300 85.160 ;
        RECT 21.530 85.160 21.850 85.220 ;
        RECT 22.465 85.160 22.755 85.205 ;
        RECT 21.530 85.020 22.755 85.160 ;
        RECT 23.000 85.160 23.140 85.360 ;
        RECT 25.670 85.300 25.990 85.360 ;
        RECT 27.510 85.500 27.830 85.560 ;
        RECT 33.120 85.500 33.260 85.655 ;
        RECT 33.490 85.640 33.810 85.900 ;
        RECT 27.510 85.360 33.260 85.500 ;
        RECT 34.040 85.500 34.180 86.040 ;
        RECT 34.500 86.040 38.320 86.180 ;
        RECT 59.800 86.040 71.990 86.180 ;
        RECT 34.500 85.885 34.640 86.040 ;
        RECT 34.425 85.655 34.715 85.885 ;
        RECT 34.870 85.840 35.190 85.900 ;
        RECT 35.345 85.840 35.635 85.885 ;
        RECT 34.870 85.700 35.635 85.840 ;
        RECT 34.870 85.640 35.190 85.700 ;
        RECT 35.345 85.655 35.635 85.700 ;
        RECT 38.090 85.640 38.410 85.900 ;
        RECT 40.850 85.840 41.170 85.900 ;
        RECT 42.245 85.840 42.535 85.885 ;
        RECT 40.850 85.700 42.535 85.840 ;
        RECT 40.850 85.640 41.170 85.700 ;
        RECT 42.245 85.655 42.535 85.700 ;
        RECT 44.070 85.840 44.390 85.900 ;
        RECT 45.465 85.840 45.755 85.885 ;
        RECT 44.070 85.700 45.755 85.840 ;
        RECT 44.070 85.640 44.390 85.700 ;
        RECT 45.465 85.655 45.755 85.700 ;
        RECT 47.290 85.840 47.610 85.900 ;
        RECT 48.685 85.840 48.975 85.885 ;
        RECT 47.290 85.700 48.975 85.840 ;
        RECT 47.290 85.640 47.610 85.700 ;
        RECT 48.685 85.655 48.975 85.700 ;
        RECT 50.510 85.840 50.830 85.900 ;
        RECT 51.905 85.840 52.195 85.885 ;
        RECT 50.510 85.700 52.195 85.840 ;
        RECT 50.510 85.640 50.830 85.700 ;
        RECT 51.905 85.655 52.195 85.700 ;
        RECT 53.730 85.840 54.050 85.900 ;
        RECT 55.125 85.840 55.415 85.885 ;
        RECT 53.730 85.700 55.415 85.840 ;
        RECT 53.730 85.640 54.050 85.700 ;
        RECT 55.125 85.655 55.415 85.700 ;
        RECT 57.870 85.640 58.190 85.900 ;
        RECT 59.800 85.885 59.940 86.040 ;
        RECT 71.670 85.980 71.990 86.040 ;
        RECT 72.590 85.980 72.910 86.240 ;
        RECT 83.645 86.180 83.935 86.225 ;
        RECT 86.850 86.180 87.170 86.240 ;
        RECT 83.645 86.040 87.170 86.180 ;
        RECT 83.645 85.995 83.935 86.040 ;
        RECT 86.850 85.980 87.170 86.040 ;
        RECT 87.310 86.180 87.630 86.240 ;
        RECT 114.080 86.225 114.220 86.380 ;
        RECT 115.845 86.380 116.610 86.520 ;
        RECT 115.845 86.335 116.135 86.380 ;
        RECT 116.290 86.320 116.610 86.380 ;
        RECT 118.130 86.520 118.450 86.580 ;
        RECT 123.665 86.520 123.955 86.565 ;
        RECT 118.130 86.380 123.955 86.520 ;
        RECT 118.130 86.320 118.450 86.380 ;
        RECT 123.665 86.335 123.955 86.380 ;
        RECT 125.030 86.520 125.350 86.580 ;
        RECT 131.485 86.520 131.775 86.565 ;
        RECT 137.450 86.520 137.770 86.580 ;
        RECT 125.030 86.380 131.775 86.520 ;
        RECT 125.030 86.320 125.350 86.380 ;
        RECT 131.485 86.335 131.775 86.380 ;
        RECT 137.135 86.380 137.770 86.520 ;
        RECT 87.310 86.040 91.680 86.180 ;
        RECT 87.310 85.980 87.630 86.040 ;
        RECT 59.725 85.655 60.015 85.885 ;
        RECT 61.565 85.840 61.855 85.885 ;
        RECT 67.530 85.840 67.850 85.900 ;
        RECT 61.565 85.700 67.850 85.840 ;
        RECT 61.565 85.655 61.855 85.700 ;
        RECT 67.530 85.640 67.850 85.700 ;
        RECT 71.210 85.640 71.530 85.900 ;
        RECT 73.510 85.640 73.830 85.900 ;
        RECT 77.650 85.640 77.970 85.900 ;
        RECT 78.110 85.640 78.430 85.900 ;
        RECT 79.950 85.640 80.270 85.900 ;
        RECT 45.910 85.500 46.230 85.560 ;
        RECT 63.390 85.500 63.710 85.560 ;
        RECT 34.040 85.360 46.230 85.500 ;
        RECT 27.510 85.300 27.830 85.360 ;
        RECT 45.910 85.300 46.230 85.360 ;
        RECT 58.880 85.360 63.710 85.500 ;
        RECT 27.600 85.160 27.740 85.300 ;
        RECT 23.000 85.020 27.740 85.160 ;
        RECT 27.970 85.160 28.290 85.220 ;
        RECT 29.365 85.160 29.655 85.205 ;
        RECT 27.970 85.020 29.655 85.160 ;
        RECT 19.705 84.975 19.995 85.020 ;
        RECT 21.530 84.960 21.850 85.020 ;
        RECT 22.465 84.975 22.755 85.020 ;
        RECT 27.970 84.960 28.290 85.020 ;
        RECT 29.365 84.975 29.655 85.020 ;
        RECT 31.665 85.160 31.955 85.205 ;
        RECT 39.010 85.160 39.330 85.220 ;
        RECT 31.665 85.020 39.330 85.160 ;
        RECT 31.665 84.975 31.955 85.020 ;
        RECT 39.010 84.960 39.330 85.020 ;
        RECT 47.750 84.960 48.070 85.220 ;
        RECT 58.880 85.205 59.020 85.360 ;
        RECT 63.390 85.300 63.710 85.360 ;
        RECT 64.325 85.500 64.615 85.545 ;
        RECT 64.770 85.500 65.090 85.560 ;
        RECT 65.705 85.500 65.995 85.545 ;
        RECT 64.325 85.360 65.995 85.500 ;
        RECT 64.325 85.315 64.615 85.360 ;
        RECT 64.770 85.300 65.090 85.360 ;
        RECT 65.705 85.315 65.995 85.360 ;
        RECT 66.150 85.500 66.470 85.560 ;
        RECT 86.940 85.500 87.080 85.980 ;
        RECT 91.540 85.885 91.680 86.040 ;
        RECT 114.005 85.995 114.295 86.225 ;
        RECT 118.590 86.180 118.910 86.240 ;
        RECT 124.570 86.180 124.890 86.240 ;
        RECT 126.885 86.180 127.175 86.225 ;
        RECT 118.590 86.040 122.270 86.180 ;
        RECT 118.590 85.980 118.910 86.040 ;
        RECT 91.465 85.655 91.755 85.885 ;
        RECT 91.910 85.640 92.230 85.900 ;
        RECT 94.210 85.840 94.530 85.900 ;
        RECT 95.145 85.840 95.435 85.885 ;
        RECT 94.210 85.700 95.435 85.840 ;
        RECT 94.210 85.640 94.530 85.700 ;
        RECT 95.145 85.655 95.435 85.700 ;
        RECT 96.985 85.840 97.275 85.885 ;
        RECT 97.430 85.840 97.750 85.900 ;
        RECT 96.985 85.700 97.750 85.840 ;
        RECT 96.985 85.655 97.275 85.700 ;
        RECT 97.430 85.640 97.750 85.700 ;
        RECT 100.665 85.840 100.955 85.885 ;
        RECT 102.950 85.840 103.270 85.900 ;
        RECT 100.665 85.700 103.270 85.840 ;
        RECT 100.665 85.655 100.955 85.700 ;
        RECT 102.950 85.640 103.270 85.700 ;
        RECT 103.885 85.840 104.175 85.885 ;
        RECT 104.330 85.840 104.650 85.900 ;
        RECT 103.885 85.700 104.650 85.840 ;
        RECT 103.885 85.655 104.175 85.700 ;
        RECT 104.330 85.640 104.650 85.700 ;
        RECT 107.105 85.840 107.395 85.885 ;
        RECT 108.010 85.840 108.330 85.900 ;
        RECT 107.105 85.700 108.330 85.840 ;
        RECT 107.105 85.655 107.395 85.700 ;
        RECT 108.010 85.640 108.330 85.700 ;
        RECT 110.325 85.840 110.615 85.885 ;
        RECT 111.230 85.840 111.550 85.900 ;
        RECT 110.325 85.700 111.550 85.840 ;
        RECT 110.325 85.655 110.615 85.700 ;
        RECT 111.230 85.640 111.550 85.700 ;
        RECT 113.070 85.840 113.390 85.900 ;
        RECT 113.545 85.840 113.835 85.885 ;
        RECT 113.070 85.700 113.835 85.840 ;
        RECT 113.070 85.640 113.390 85.700 ;
        RECT 113.545 85.655 113.835 85.700 ;
        RECT 118.145 85.840 118.435 85.885 ;
        RECT 119.510 85.840 119.830 85.900 ;
        RECT 118.145 85.700 119.830 85.840 ;
        RECT 118.145 85.655 118.435 85.700 ;
        RECT 119.510 85.640 119.830 85.700 ;
        RECT 119.970 85.640 120.290 85.900 ;
        RECT 120.890 85.640 121.210 85.900 ;
        RECT 122.130 85.840 122.270 86.040 ;
        RECT 124.570 86.040 127.175 86.180 ;
        RECT 124.570 85.980 124.890 86.040 ;
        RECT 126.885 85.995 127.175 86.040 ;
        RECT 127.805 86.180 128.095 86.225 ;
        RECT 131.010 86.180 131.330 86.240 ;
        RECT 127.805 86.040 131.330 86.180 ;
        RECT 127.805 85.995 128.095 86.040 ;
        RECT 131.010 85.980 131.330 86.040 ;
        RECT 122.745 85.840 123.035 85.885 ;
        RECT 122.130 85.700 123.035 85.840 ;
        RECT 122.745 85.655 123.035 85.700 ;
        RECT 125.950 85.640 126.270 85.900 ;
        RECT 130.550 85.640 130.870 85.900 ;
        RECT 132.390 85.840 132.710 85.900 ;
        RECT 134.475 85.840 134.765 85.885 ;
        RECT 132.390 85.700 134.765 85.840 ;
        RECT 132.390 85.640 132.710 85.700 ;
        RECT 134.475 85.655 134.765 85.700 ;
        RECT 135.150 85.640 135.470 85.900 ;
        RECT 135.610 85.640 135.930 85.900 ;
        RECT 136.530 85.840 136.850 85.900 ;
        RECT 137.135 85.885 137.275 86.380 ;
        RECT 137.450 86.320 137.770 86.380 ;
        RECT 139.305 86.520 139.595 86.565 ;
        RECT 141.590 86.520 141.910 86.580 ;
        RECT 139.305 86.380 141.910 86.520 ;
        RECT 139.305 86.335 139.595 86.380 ;
        RECT 141.590 86.320 141.910 86.380 ;
        RECT 144.825 86.335 145.115 86.565 ;
        RECT 138.370 86.180 138.690 86.240 ;
        RECT 144.900 86.180 145.040 86.335 ;
        RECT 138.370 86.040 145.040 86.180 ;
        RECT 138.370 85.980 138.690 86.040 ;
        RECT 136.335 85.700 136.850 85.840 ;
        RECT 136.530 85.640 136.850 85.700 ;
        RECT 137.005 85.655 137.295 85.885 ;
        RECT 137.450 85.640 137.770 85.900 ;
        RECT 140.210 85.640 140.530 85.900 ;
        RECT 142.050 85.640 142.370 85.900 ;
        RECT 142.970 85.840 143.290 85.900 ;
        RECT 143.905 85.840 144.195 85.885 ;
        RECT 142.970 85.700 144.195 85.840 ;
        RECT 142.970 85.640 143.290 85.700 ;
        RECT 143.905 85.655 144.195 85.700 ;
        RECT 87.325 85.500 87.615 85.545 ;
        RECT 66.150 85.360 69.600 85.500 ;
        RECT 86.940 85.360 87.615 85.500 ;
        RECT 66.150 85.300 66.470 85.360 ;
        RECT 58.805 84.975 59.095 85.205 ;
        RECT 60.645 85.160 60.935 85.205 ;
        RECT 66.610 85.160 66.930 85.220 ;
        RECT 69.460 85.205 69.600 85.360 ;
        RECT 87.325 85.315 87.615 85.360 ;
        RECT 89.150 85.500 89.470 85.560 ;
        RECT 92.370 85.500 92.690 85.560 ;
        RECT 114.910 85.500 115.230 85.560 ;
        RECT 89.150 85.360 91.220 85.500 ;
        RECT 89.150 85.300 89.470 85.360 ;
        RECT 60.645 85.020 66.930 85.160 ;
        RECT 60.645 84.975 60.935 85.020 ;
        RECT 66.610 84.960 66.930 85.020 ;
        RECT 69.385 84.975 69.675 85.205 ;
        RECT 73.050 85.160 73.370 85.220 ;
        RECT 74.445 85.160 74.735 85.205 ;
        RECT 73.050 85.020 74.735 85.160 ;
        RECT 73.050 84.960 73.370 85.020 ;
        RECT 74.445 84.975 74.735 85.020 ;
        RECT 76.270 85.160 76.590 85.220 ;
        RECT 76.745 85.160 77.035 85.205 ;
        RECT 76.270 85.020 77.035 85.160 ;
        RECT 76.270 84.960 76.590 85.020 ;
        RECT 76.745 84.975 77.035 85.020 ;
        RECT 79.045 85.160 79.335 85.205 ;
        RECT 79.490 85.160 79.810 85.220 ;
        RECT 79.045 85.020 79.810 85.160 ;
        RECT 79.045 84.975 79.335 85.020 ;
        RECT 79.490 84.960 79.810 85.020 ;
        RECT 80.885 85.160 81.175 85.205 ;
        RECT 82.710 85.160 83.030 85.220 ;
        RECT 80.885 85.020 83.030 85.160 ;
        RECT 80.885 84.975 81.175 85.020 ;
        RECT 82.710 84.960 83.030 85.020 ;
        RECT 85.930 85.160 86.250 85.220 ;
        RECT 90.545 85.160 90.835 85.205 ;
        RECT 85.930 85.020 90.835 85.160 ;
        RECT 91.080 85.160 91.220 85.360 ;
        RECT 92.370 85.360 94.670 85.500 ;
        RECT 92.370 85.300 92.690 85.360 ;
        RECT 92.845 85.160 93.135 85.205 ;
        RECT 91.080 85.020 93.135 85.160 ;
        RECT 94.530 85.160 94.670 85.360 ;
        RECT 114.910 85.360 117.900 85.500 ;
        RECT 114.910 85.300 115.230 85.360 ;
        RECT 96.065 85.160 96.355 85.205 ;
        RECT 94.530 85.020 96.355 85.160 ;
        RECT 85.930 84.960 86.250 85.020 ;
        RECT 90.545 84.975 90.835 85.020 ;
        RECT 92.845 84.975 93.135 85.020 ;
        RECT 96.065 84.975 96.355 85.020 ;
        RECT 98.810 85.160 99.130 85.220 ;
        RECT 99.745 85.160 100.035 85.205 ;
        RECT 98.810 85.020 100.035 85.160 ;
        RECT 98.810 84.960 99.130 85.020 ;
        RECT 99.745 84.975 100.035 85.020 ;
        RECT 102.030 85.160 102.350 85.220 ;
        RECT 102.965 85.160 103.255 85.205 ;
        RECT 102.030 85.020 103.255 85.160 ;
        RECT 102.030 84.960 102.350 85.020 ;
        RECT 102.965 84.975 103.255 85.020 ;
        RECT 105.250 85.160 105.570 85.220 ;
        RECT 106.185 85.160 106.475 85.205 ;
        RECT 105.250 85.020 106.475 85.160 ;
        RECT 105.250 84.960 105.570 85.020 ;
        RECT 106.185 84.975 106.475 85.020 ;
        RECT 108.470 85.160 108.790 85.220 ;
        RECT 109.405 85.160 109.695 85.205 ;
        RECT 108.470 85.020 109.695 85.160 ;
        RECT 108.470 84.960 108.790 85.020 ;
        RECT 109.405 84.975 109.695 85.020 ;
        RECT 111.690 85.160 112.010 85.220 ;
        RECT 112.625 85.160 112.915 85.205 ;
        RECT 111.690 85.020 112.915 85.160 ;
        RECT 111.690 84.960 112.010 85.020 ;
        RECT 112.625 84.975 112.915 85.020 ;
        RECT 116.290 84.960 116.610 85.220 ;
        RECT 117.760 85.160 117.900 85.360 ;
        RECT 118.590 85.300 118.910 85.560 ;
        RECT 119.050 85.300 119.370 85.560 ;
        RECT 121.350 85.500 121.670 85.560 ;
        RECT 131.010 85.500 131.330 85.560 ;
        RECT 121.350 85.360 125.260 85.500 ;
        RECT 121.350 85.300 121.670 85.360 ;
        RECT 125.120 85.205 125.260 85.360 ;
        RECT 131.010 85.360 134.460 85.500 ;
        RECT 131.010 85.300 131.330 85.360 ;
        RECT 121.825 85.160 122.115 85.205 ;
        RECT 117.760 85.020 122.115 85.160 ;
        RECT 121.825 84.975 122.115 85.020 ;
        RECT 125.045 84.975 125.335 85.205 ;
        RECT 128.265 85.160 128.555 85.205 ;
        RECT 132.850 85.160 133.170 85.220 ;
        RECT 128.265 85.020 133.170 85.160 ;
        RECT 134.320 85.160 134.460 85.360 ;
        RECT 141.145 85.160 141.435 85.205 ;
        RECT 134.320 85.020 141.435 85.160 ;
        RECT 128.265 84.975 128.555 85.020 ;
        RECT 132.850 84.960 133.170 85.020 ;
        RECT 141.145 84.975 141.435 85.020 ;
        RECT 142.970 84.960 143.290 85.220 ;
        RECT 17.320 84.340 147.040 84.820 ;
        RECT 33.490 84.140 33.810 84.200 ;
        RECT 47.750 84.140 48.070 84.200 ;
        RECT 33.490 84.000 48.070 84.140 ;
        RECT 33.490 83.940 33.810 84.000 ;
        RECT 47.750 83.940 48.070 84.000 ;
        RECT 57.870 84.140 58.190 84.200 ;
        RECT 68.910 84.140 69.230 84.200 ;
        RECT 57.870 84.000 69.230 84.140 ;
        RECT 57.870 83.940 58.190 84.000 ;
        RECT 68.910 83.940 69.230 84.000 ;
        RECT 116.290 84.140 116.610 84.200 ;
        RECT 124.110 84.140 124.430 84.200 ;
        RECT 116.290 84.000 124.430 84.140 ;
        RECT 116.290 83.940 116.610 84.000 ;
        RECT 124.110 83.940 124.430 84.000 ;
        RECT 104.790 83.800 105.110 83.860 ;
        RECT 119.050 83.800 119.370 83.860 ;
        RECT 135.610 83.800 135.930 83.860 ;
        RECT 104.790 83.660 135.930 83.800 ;
        RECT 104.790 83.600 105.110 83.660 ;
        RECT 119.050 83.600 119.370 83.660 ;
        RECT 135.610 83.600 135.930 83.660 ;
        RECT 127.790 80.400 128.110 80.460 ;
        RECT 136.070 80.400 136.390 80.460 ;
        RECT 127.790 80.260 136.390 80.400 ;
        RECT 127.790 80.200 128.110 80.260 ;
        RECT 136.070 80.200 136.390 80.260 ;
        RECT 140.670 80.060 140.990 80.120 ;
        RECT 144.810 80.060 145.130 80.120 ;
        RECT 140.670 79.920 145.130 80.060 ;
        RECT 140.670 79.860 140.990 79.920 ;
        RECT 144.810 79.860 145.130 79.920 ;
        RECT 134.230 79.380 134.550 79.440 ;
        RECT 142.970 79.380 143.290 79.440 ;
        RECT 134.230 79.240 143.290 79.380 ;
        RECT 134.230 79.180 134.550 79.240 ;
        RECT 142.970 79.180 143.290 79.240 ;
        RECT 158.295 7.555 160.610 222.955 ;
        RECT 7.615 7.020 160.610 7.555 ;
        RECT 0.510 4.540 160.610 7.020 ;
        RECT 7.615 4.445 160.610 4.540 ;
      LAYER met2 ;
        RECT 60.790 213.440 64.260 213.450 ;
        RECT 60.260 213.170 64.260 213.440 ;
        RECT 80.900 213.370 82.640 213.380 ;
        RECT 83.130 213.370 85.220 213.380 ;
        RECT 79.580 213.290 79.720 213.300 ;
        RECT 32.870 212.235 34.410 212.605 ;
        RECT 60.260 211.050 60.400 213.170 ;
        RECT 75.720 213.010 79.720 213.290 ;
        RECT 79.580 211.730 79.720 213.010 ;
        RECT 80.900 212.920 85.220 213.370 ;
        RECT 96.800 213.310 99.660 213.330 ;
        RECT 86.010 213.030 90.010 213.310 ;
        RECT 95.660 213.050 99.660 213.310 ;
        RECT 82.790 212.750 82.970 212.920 ;
        RECT 79.520 211.410 79.780 211.730 ;
        RECT 82.800 211.050 82.940 212.750 ;
        RECT 86.020 211.390 86.160 213.030 ;
        RECT 95.680 211.730 95.820 213.050 ;
        RECT 87.800 211.410 88.060 211.730 ;
        RECT 95.620 211.410 95.880 211.730 ;
        RECT 85.960 211.070 86.220 211.390 ;
        RECT 60.200 210.730 60.460 211.050 ;
        RECT 82.740 210.730 83.000 211.050 ;
        RECT 87.340 210.730 87.600 211.050 ;
        RECT 51.920 210.390 52.180 210.710 ;
        RECT 84.580 210.390 84.840 210.710 ;
        RECT 36.170 209.515 37.710 209.885 ;
        RECT 32.870 206.795 34.410 207.165 ;
        RECT 51.000 205.970 51.260 206.290 ;
        RECT 49.160 204.610 49.420 204.930 ;
        RECT 36.170 204.075 37.710 204.445 ;
        RECT 49.220 203.910 49.360 204.610 ;
        RECT 49.160 203.590 49.420 203.910 ;
        RECT 45.480 203.250 45.740 203.570 ;
        RECT 32.870 201.355 34.410 201.725 ;
        RECT 45.540 200.510 45.680 203.250 ;
        RECT 50.540 202.910 50.800 203.230 ;
        RECT 45.940 201.890 46.200 202.210 ;
        RECT 43.640 200.190 43.900 200.510 ;
        RECT 45.480 200.190 45.740 200.510 ;
        RECT 36.170 198.635 37.710 199.005 ;
        RECT 32.870 195.915 34.410 196.285 ;
        RECT 42.720 195.090 42.980 195.410 ;
        RECT 21.560 194.410 21.820 194.730 ;
        RECT 26.160 194.410 26.420 194.730 ;
        RECT 32.140 194.410 32.400 194.730 ;
        RECT 21.620 192.690 21.760 194.410 ;
        RECT 21.560 192.370 21.820 192.690 ;
        RECT 18.800 192.030 19.060 192.350 ;
        RECT 18.860 189.825 19.000 192.030 ;
        RECT 18.790 189.455 19.070 189.825 ;
        RECT 21.620 187.590 21.760 192.370 ;
        RECT 25.240 192.030 25.500 192.350 ;
        RECT 25.700 192.030 25.960 192.350 ;
        RECT 24.780 191.350 25.040 191.670 ;
        RECT 23.860 191.010 24.120 191.330 ;
        RECT 22.940 188.630 23.200 188.950 ;
        RECT 21.560 187.270 21.820 187.590 ;
        RECT 23.000 184.870 23.140 188.630 ;
        RECT 23.920 187.250 24.060 191.010 ;
        RECT 23.860 186.930 24.120 187.250 ;
        RECT 22.940 184.550 23.200 184.870 ;
        RECT 24.840 183.510 24.980 191.350 ;
        RECT 25.300 189.290 25.440 192.030 ;
        RECT 25.240 188.970 25.500 189.290 ;
        RECT 25.300 187.590 25.440 188.970 ;
        RECT 25.240 187.270 25.500 187.590 ;
        RECT 24.780 183.190 25.040 183.510 ;
        RECT 24.840 179.090 24.980 183.190 ;
        RECT 25.760 183.170 25.900 192.030 ;
        RECT 26.220 188.950 26.360 194.410 ;
        RECT 28.920 194.070 29.180 194.390 ;
        RECT 27.080 193.730 27.340 194.050 ;
        RECT 26.160 188.630 26.420 188.950 ;
        RECT 26.160 185.570 26.420 185.890 ;
        RECT 26.220 184.190 26.360 185.570 ;
        RECT 27.140 184.870 27.280 193.730 ;
        RECT 28.980 189.290 29.120 194.070 ;
        RECT 32.200 191.670 32.340 194.410 ;
        RECT 39.500 194.070 39.760 194.390 ;
        RECT 36.170 193.195 37.710 193.565 ;
        RECT 39.560 193.030 39.700 194.070 ;
        RECT 39.960 193.730 40.220 194.050 ;
        RECT 39.500 192.710 39.760 193.030 ;
        RECT 35.820 192.030 36.080 192.350 ;
        RECT 32.140 191.580 32.400 191.670 ;
        RECT 31.740 191.440 32.400 191.580 ;
        RECT 31.740 189.290 31.880 191.440 ;
        RECT 32.140 191.350 32.400 191.440 ;
        RECT 32.870 190.475 34.410 190.845 ;
        RECT 35.880 190.310 36.020 192.030 ;
        RECT 40.020 191.750 40.160 193.730 ;
        RECT 40.880 192.030 41.140 192.350 ;
        RECT 39.560 191.610 40.160 191.750 ;
        RECT 39.560 191.580 39.700 191.610 ;
        RECT 39.100 191.440 39.700 191.580 ;
        RECT 39.100 191.185 39.240 191.440 ;
        RECT 40.420 191.350 40.680 191.670 ;
        RECT 39.960 191.240 40.220 191.330 ;
        RECT 39.030 190.815 39.310 191.185 ;
        RECT 39.560 191.100 40.220 191.240 ;
        RECT 35.820 189.990 36.080 190.310 ;
        RECT 39.100 189.290 39.240 190.815 ;
        RECT 28.920 188.970 29.180 189.290 ;
        RECT 31.680 188.970 31.940 189.290 ;
        RECT 32.600 189.030 32.860 189.290 ;
        RECT 33.980 189.030 34.240 189.290 ;
        RECT 32.600 188.970 34.240 189.030 ;
        RECT 39.040 188.970 39.300 189.290 ;
        RECT 28.460 188.290 28.720 188.610 ;
        RECT 28.520 186.910 28.660 188.290 ;
        RECT 28.980 187.590 29.120 188.970 ;
        RECT 30.760 188.290 31.020 188.610 ;
        RECT 28.920 187.270 29.180 187.590 ;
        RECT 28.460 186.590 28.720 186.910 ;
        RECT 28.980 186.570 29.120 187.270 ;
        RECT 28.920 186.250 29.180 186.570 ;
        RECT 27.540 185.570 27.800 185.890 ;
        RECT 27.080 184.550 27.340 184.870 ;
        RECT 26.160 183.870 26.420 184.190 ;
        RECT 25.700 182.850 25.960 183.170 ;
        RECT 25.700 181.150 25.960 181.470 ;
        RECT 24.780 178.770 25.040 179.090 ;
        RECT 25.760 178.070 25.900 181.150 ;
        RECT 26.220 181.130 26.360 183.870 ;
        RECT 27.600 183.850 27.740 185.570 ;
        RECT 27.540 183.530 27.800 183.850 ;
        RECT 30.820 183.170 30.960 188.290 ;
        RECT 31.740 187.250 31.880 188.970 ;
        RECT 32.140 188.630 32.400 188.950 ;
        RECT 32.660 188.890 34.180 188.970 ;
        RECT 31.680 187.160 31.940 187.250 ;
        RECT 31.280 187.020 31.940 187.160 ;
        RECT 31.280 186.570 31.420 187.020 ;
        RECT 31.680 186.930 31.940 187.020 ;
        RECT 31.220 186.250 31.480 186.570 ;
        RECT 31.280 185.890 31.420 186.250 ;
        RECT 31.220 185.570 31.480 185.890 ;
        RECT 32.200 183.510 32.340 188.630 ;
        RECT 32.660 188.610 32.800 188.890 ;
        RECT 32.600 188.290 32.860 188.610 ;
        RECT 32.660 186.230 32.800 188.290 ;
        RECT 36.170 187.755 37.710 188.125 ;
        RECT 35.820 186.590 36.080 186.910 ;
        RECT 37.200 186.590 37.460 186.910 ;
        RECT 38.580 186.590 38.840 186.910 ;
        RECT 32.600 185.910 32.860 186.230 ;
        RECT 34.900 185.910 35.160 186.230 ;
        RECT 32.870 185.035 34.410 185.405 ;
        RECT 32.140 183.190 32.400 183.510 ;
        RECT 30.760 182.850 31.020 183.170 ;
        RECT 26.160 180.810 26.420 181.130 ;
        RECT 26.220 178.410 26.360 180.810 ;
        RECT 34.960 180.790 35.100 185.910 ;
        RECT 35.360 184.550 35.620 184.870 ;
        RECT 35.420 182.150 35.560 184.550 ;
        RECT 35.880 183.850 36.020 186.590 ;
        RECT 37.260 185.890 37.400 186.590 ;
        RECT 37.200 185.570 37.460 185.890 ;
        RECT 35.820 183.530 36.080 183.850 ;
        RECT 35.360 181.830 35.620 182.150 ;
        RECT 35.880 181.810 36.020 183.530 ;
        RECT 37.260 183.510 37.400 185.570 ;
        RECT 38.640 183.850 38.780 186.590 ;
        RECT 39.100 184.870 39.240 188.970 ;
        RECT 39.560 186.910 39.700 191.100 ;
        RECT 39.960 191.010 40.220 191.100 ;
        RECT 40.480 189.970 40.620 191.350 ;
        RECT 40.420 189.650 40.680 189.970 ;
        RECT 40.480 186.910 40.620 189.650 ;
        RECT 40.940 189.290 41.080 192.030 ;
        RECT 42.780 191.330 42.920 195.090 ;
        RECT 43.700 192.690 43.840 200.190 ;
        RECT 46.000 199.830 46.140 201.890 ;
        RECT 45.940 199.510 46.200 199.830 ;
        RECT 50.600 198.470 50.740 202.910 ;
        RECT 50.540 198.150 50.800 198.470 ;
        RECT 51.060 197.790 51.200 205.970 ;
        RECT 51.000 197.470 51.260 197.790 ;
        RECT 50.540 196.790 50.800 197.110 ;
        RECT 43.640 192.370 43.900 192.690 ;
        RECT 46.400 192.370 46.660 192.690 ;
        RECT 43.180 191.690 43.440 192.010 ;
        RECT 42.720 191.010 42.980 191.330 ;
        RECT 40.880 188.970 41.140 189.290 ;
        RECT 41.340 188.630 41.600 188.950 ;
        RECT 41.400 186.910 41.540 188.630 ;
        RECT 42.780 186.990 42.920 191.010 ;
        RECT 43.240 189.290 43.380 191.690 ;
        RECT 43.180 188.970 43.440 189.290 ;
        RECT 43.240 187.590 43.380 188.970 ;
        RECT 43.180 187.270 43.440 187.590 ;
        RECT 39.500 186.590 39.760 186.910 ;
        RECT 40.420 186.590 40.680 186.910 ;
        RECT 41.340 186.590 41.600 186.910 ;
        RECT 42.780 186.850 43.380 186.990 ;
        RECT 43.240 186.570 43.380 186.850 ;
        RECT 39.960 186.250 40.220 186.570 ;
        RECT 43.180 186.250 43.440 186.570 ;
        RECT 39.040 184.550 39.300 184.870 ;
        RECT 38.580 183.530 38.840 183.850 ;
        RECT 39.500 183.530 39.760 183.850 ;
        RECT 37.200 183.190 37.460 183.510 ;
        RECT 36.170 182.315 37.710 182.685 ;
        RECT 36.280 181.830 36.540 182.150 ;
        RECT 35.820 181.490 36.080 181.810 ;
        RECT 35.360 181.150 35.620 181.470 ;
        RECT 34.900 180.470 35.160 180.790 ;
        RECT 29.380 180.130 29.640 180.450 ;
        RECT 28.000 178.770 28.260 179.090 ;
        RECT 26.160 178.090 26.420 178.410 ;
        RECT 27.080 178.090 27.340 178.410 ;
        RECT 25.700 177.750 25.960 178.070 ;
        RECT 22.480 177.410 22.740 177.730 ;
        RECT 22.540 176.370 22.680 177.410 ;
        RECT 22.480 176.050 22.740 176.370 ;
        RECT 25.760 175.010 25.900 177.750 ;
        RECT 26.220 176.030 26.360 178.090 ;
        RECT 27.140 176.370 27.280 178.090 ;
        RECT 27.080 176.050 27.340 176.370 ;
        RECT 26.160 175.710 26.420 176.030 ;
        RECT 26.620 175.030 26.880 175.350 ;
        RECT 25.240 174.690 25.500 175.010 ;
        RECT 25.700 174.690 25.960 175.010 ;
        RECT 25.300 172.970 25.440 174.690 ;
        RECT 25.760 173.990 25.900 174.690 ;
        RECT 25.700 173.670 25.960 173.990 ;
        RECT 25.240 172.650 25.500 172.970 ;
        RECT 21.100 166.530 21.360 166.850 ;
        RECT 19.260 161.770 19.520 162.090 ;
        RECT 19.320 159.710 19.460 161.770 ;
        RECT 20.180 161.090 20.440 161.410 ;
        RECT 20.240 160.390 20.380 161.090 ;
        RECT 20.180 160.070 20.440 160.390 ;
        RECT 19.260 159.390 19.520 159.710 ;
        RECT 21.160 158.690 21.300 166.530 ;
        RECT 22.020 165.170 22.280 165.490 ;
        RECT 21.560 163.810 21.820 164.130 ;
        RECT 21.620 160.390 21.760 163.810 ;
        RECT 22.080 161.410 22.220 165.170 ;
        RECT 23.400 164.040 23.660 164.130 ;
        RECT 23.400 163.900 24.060 164.040 ;
        RECT 23.400 163.810 23.660 163.900 ;
        RECT 22.020 161.090 22.280 161.410 ;
        RECT 21.560 160.070 21.820 160.390 ;
        RECT 22.080 160.050 22.220 161.090 ;
        RECT 23.920 160.050 24.060 163.900 ;
        RECT 25.300 160.390 25.440 172.650 ;
        RECT 26.680 167.530 26.820 175.030 ;
        RECT 26.620 167.210 26.880 167.530 ;
        RECT 26.680 165.490 26.820 167.210 ;
        RECT 27.540 166.870 27.800 167.190 ;
        RECT 26.620 165.170 26.880 165.490 ;
        RECT 27.600 165.150 27.740 166.870 ;
        RECT 27.540 164.830 27.800 165.150 ;
        RECT 26.160 164.150 26.420 164.470 ;
        RECT 26.220 163.110 26.360 164.150 ;
        RECT 27.080 163.810 27.340 164.130 ;
        RECT 27.140 163.110 27.280 163.810 ;
        RECT 26.160 162.790 26.420 163.110 ;
        RECT 27.080 162.790 27.340 163.110 ;
        RECT 27.600 162.090 27.740 164.830 ;
        RECT 27.540 161.770 27.800 162.090 ;
        RECT 27.540 161.150 27.800 161.410 ;
        RECT 28.060 161.150 28.200 178.770 ;
        RECT 29.440 178.410 29.580 180.130 ;
        RECT 32.870 179.595 34.410 179.965 ;
        RECT 32.140 179.110 32.400 179.430 ;
        RECT 31.220 178.770 31.480 179.090 ;
        RECT 30.300 178.430 30.560 178.750 ;
        RECT 29.380 178.090 29.640 178.410 ;
        RECT 29.440 175.430 29.580 178.090 ;
        RECT 30.360 176.710 30.500 178.430 ;
        RECT 30.300 176.390 30.560 176.710 ;
        RECT 31.280 176.370 31.420 178.770 ;
        RECT 32.200 176.710 32.340 179.110 ;
        RECT 35.420 178.410 35.560 181.150 ;
        RECT 35.820 180.810 36.080 181.130 ;
        RECT 35.880 178.410 36.020 180.810 ;
        RECT 35.360 178.090 35.620 178.410 ;
        RECT 35.820 178.090 36.080 178.410 ;
        RECT 36.340 177.640 36.480 181.830 ;
        RECT 39.560 181.130 39.700 183.530 ;
        RECT 40.020 181.470 40.160 186.250 ;
        RECT 40.880 185.910 41.140 186.230 ;
        RECT 40.420 185.570 40.680 185.890 ;
        RECT 40.480 183.850 40.620 185.570 ;
        RECT 40.420 183.530 40.680 183.850 ;
        RECT 40.940 183.510 41.080 185.910 ;
        RECT 42.720 185.570 42.980 185.890 ;
        RECT 42.260 183.590 42.520 183.850 ;
        RECT 42.780 183.590 42.920 185.570 ;
        RECT 43.240 184.530 43.380 186.250 ;
        RECT 43.180 184.210 43.440 184.530 ;
        RECT 42.260 183.530 42.920 183.590 ;
        RECT 40.880 183.190 41.140 183.510 ;
        RECT 42.320 183.450 42.920 183.530 ;
        RECT 41.340 182.850 41.600 183.170 ;
        RECT 41.800 182.850 42.060 183.170 ;
        RECT 41.400 181.470 41.540 182.850 ;
        RECT 41.860 181.810 42.000 182.850 ;
        RECT 41.800 181.490 42.060 181.810 ;
        RECT 39.960 181.150 40.220 181.470 ;
        RECT 41.340 181.150 41.600 181.470 ;
        RECT 39.500 180.810 39.760 181.130 ;
        RECT 36.740 180.470 37.000 180.790 ;
        RECT 36.800 178.410 36.940 180.470 ;
        RECT 39.500 180.130 39.760 180.450 ;
        RECT 36.740 178.090 37.000 178.410 ;
        RECT 37.660 178.090 37.920 178.410 ;
        RECT 38.580 178.090 38.840 178.410 ;
        RECT 37.720 177.730 37.860 178.090 ;
        RECT 35.880 177.500 36.480 177.640 ;
        RECT 32.140 176.390 32.400 176.710 ;
        RECT 31.220 176.050 31.480 176.370 ;
        RECT 29.440 175.290 30.040 175.430 ;
        RECT 34.900 175.370 35.160 175.690 ;
        RECT 29.900 175.010 30.040 175.290 ;
        RECT 29.380 174.690 29.640 175.010 ;
        RECT 29.840 174.690 30.100 175.010 ;
        RECT 29.440 172.630 29.580 174.690 ;
        RECT 32.870 174.155 34.410 174.525 ;
        RECT 29.380 172.310 29.640 172.630 ;
        RECT 34.960 170.590 35.100 175.370 ;
        RECT 34.900 170.270 35.160 170.590 ;
        RECT 32.870 168.715 34.410 169.085 ;
        RECT 29.380 167.890 29.640 168.210 ;
        RECT 28.920 166.530 29.180 166.850 ;
        RECT 28.980 165.150 29.120 166.530 ;
        RECT 29.440 165.150 29.580 167.890 ;
        RECT 33.980 167.210 34.240 167.530 ;
        RECT 31.680 166.870 31.940 167.190 ;
        RECT 28.920 164.830 29.180 165.150 ;
        RECT 29.380 164.830 29.640 165.150 ;
        RECT 28.460 164.490 28.720 164.810 ;
        RECT 28.520 161.410 28.660 164.490 ;
        RECT 28.980 163.110 29.120 164.830 ;
        RECT 31.740 164.810 31.880 166.870 ;
        RECT 34.040 165.830 34.180 167.210 ;
        RECT 33.980 165.510 34.240 165.830 ;
        RECT 32.140 164.830 32.400 165.150 ;
        RECT 31.680 164.490 31.940 164.810 ;
        RECT 30.760 163.810 31.020 164.130 ;
        RECT 31.680 163.810 31.940 164.130 ;
        RECT 28.920 162.790 29.180 163.110 ;
        RECT 27.540 161.090 28.200 161.150 ;
        RECT 28.460 161.090 28.720 161.410 ;
        RECT 27.600 161.010 28.200 161.090 ;
        RECT 25.240 160.070 25.500 160.390 ;
        RECT 28.060 160.050 28.200 161.010 ;
        RECT 22.020 159.730 22.280 160.050 ;
        RECT 23.860 159.730 24.120 160.050 ;
        RECT 28.000 159.730 28.260 160.050 ;
        RECT 28.980 159.030 29.120 162.790 ;
        RECT 30.300 161.770 30.560 162.090 ;
        RECT 29.840 161.430 30.100 161.750 ;
        RECT 29.900 160.050 30.040 161.430 ;
        RECT 30.360 160.390 30.500 161.770 ;
        RECT 30.820 160.390 30.960 163.810 ;
        RECT 30.300 160.070 30.560 160.390 ;
        RECT 30.760 160.070 31.020 160.390 ;
        RECT 29.840 159.730 30.100 160.050 ;
        RECT 28.920 158.710 29.180 159.030 ;
        RECT 31.740 158.690 31.880 163.810 ;
        RECT 32.200 163.110 32.340 164.830 ;
        RECT 34.960 164.470 35.100 170.270 ;
        RECT 35.360 166.870 35.620 167.190 ;
        RECT 35.420 164.810 35.560 166.870 ;
        RECT 35.880 165.830 36.020 177.500 ;
        RECT 37.660 177.410 37.920 177.730 ;
        RECT 38.120 177.410 38.380 177.730 ;
        RECT 36.170 176.875 37.710 177.245 ;
        RECT 38.180 176.110 38.320 177.410 ;
        RECT 38.640 176.370 38.780 178.090 ;
        RECT 39.040 176.390 39.300 176.710 ;
        RECT 37.720 176.030 38.320 176.110 ;
        RECT 38.580 176.050 38.840 176.370 ;
        RECT 37.660 175.970 38.320 176.030 ;
        RECT 37.660 175.710 37.920 175.970 ;
        RECT 38.580 174.690 38.840 175.010 ;
        RECT 38.640 173.650 38.780 174.690 ;
        RECT 38.580 173.330 38.840 173.650 ;
        RECT 38.120 172.650 38.380 172.970 ;
        RECT 36.170 171.435 37.710 171.805 ;
        RECT 38.180 171.270 38.320 172.650 ;
        RECT 37.200 170.950 37.460 171.270 ;
        RECT 38.120 170.950 38.380 171.270 ;
        RECT 36.280 170.270 36.540 170.590 ;
        RECT 36.340 168.550 36.480 170.270 ;
        RECT 37.260 168.550 37.400 170.950 ;
        RECT 38.580 170.270 38.840 170.590 ;
        RECT 36.280 168.230 36.540 168.550 ;
        RECT 37.200 168.230 37.460 168.550 ;
        RECT 38.640 168.210 38.780 170.270 ;
        RECT 39.100 169.570 39.240 176.390 ;
        RECT 39.560 172.970 39.700 180.130 ;
        RECT 42.320 179.430 42.460 183.450 ;
        RECT 42.720 181.150 42.980 181.470 ;
        RECT 42.260 179.110 42.520 179.430 ;
        RECT 39.960 178.090 40.220 178.410 ;
        RECT 40.020 176.710 40.160 178.090 ;
        RECT 40.420 177.750 40.680 178.070 ;
        RECT 39.960 176.390 40.220 176.710 ;
        RECT 40.480 175.690 40.620 177.750 ;
        RECT 42.780 176.030 42.920 181.150 ;
        RECT 42.720 175.710 42.980 176.030 ;
        RECT 40.420 175.370 40.680 175.690 ;
        RECT 39.960 175.030 40.220 175.350 ;
        RECT 40.020 173.650 40.160 175.030 ;
        RECT 39.960 173.330 40.220 173.650 ;
        RECT 39.500 172.650 39.760 172.970 ;
        RECT 40.020 171.270 40.160 173.330 ;
        RECT 43.240 172.970 43.380 184.210 ;
        RECT 43.700 178.750 43.840 192.370 ;
        RECT 45.020 192.030 45.280 192.350 ;
        RECT 45.480 192.030 45.740 192.350 ;
        RECT 45.080 186.910 45.220 192.030 ;
        RECT 45.540 188.950 45.680 192.030 ;
        RECT 46.460 189.970 46.600 192.370 ;
        RECT 46.400 189.650 46.660 189.970 ;
        RECT 45.940 189.310 46.200 189.630 ;
        RECT 45.480 188.630 45.740 188.950 ;
        RECT 45.020 186.590 45.280 186.910 ;
        RECT 45.080 186.310 45.220 186.590 ;
        RECT 44.160 186.170 45.220 186.310 ;
        RECT 44.160 182.150 44.300 186.170 ;
        RECT 45.540 184.170 45.680 188.630 ;
        RECT 46.000 184.530 46.140 189.310 ;
        RECT 46.460 188.950 46.600 189.650 ;
        RECT 50.600 189.630 50.740 196.790 ;
        RECT 51.460 196.450 51.720 196.770 ;
        RECT 51.520 193.030 51.660 196.450 ;
        RECT 51.460 192.710 51.720 193.030 ;
        RECT 51.980 192.690 52.120 210.390 ;
        RECT 55.140 209.030 55.400 209.350 ;
        RECT 55.200 208.670 55.340 209.030 ;
        RECT 64.340 208.690 64.600 209.010 ;
        RECT 53.760 208.350 54.020 208.670 ;
        RECT 55.140 208.350 55.400 208.670 ;
        RECT 60.660 208.350 60.920 208.670 ;
        RECT 52.380 208.010 52.640 208.330 ;
        RECT 52.440 197.790 52.580 208.010 ;
        RECT 53.300 205.630 53.560 205.950 ;
        RECT 53.360 202.210 53.500 205.630 ;
        RECT 53.300 201.890 53.560 202.210 ;
        RECT 53.360 200.170 53.500 201.890 ;
        RECT 53.820 201.190 53.960 208.350 ;
        RECT 54.220 207.330 54.480 207.650 ;
        RECT 54.280 203.230 54.420 207.330 ;
        RECT 54.680 205.290 54.940 205.610 ;
        RECT 54.220 202.910 54.480 203.230 ;
        RECT 53.760 200.870 54.020 201.190 ;
        RECT 53.300 199.850 53.560 200.170 ;
        RECT 54.220 199.850 54.480 200.170 ;
        RECT 52.380 197.470 52.640 197.790 ;
        RECT 52.840 194.750 53.100 195.070 ;
        RECT 52.900 193.030 53.040 194.750 ;
        RECT 54.280 194.730 54.420 199.850 ;
        RECT 54.740 199.830 54.880 205.290 ;
        RECT 55.200 202.210 55.340 208.350 ;
        RECT 56.980 208.010 57.240 208.330 ;
        RECT 55.600 207.330 55.860 207.650 ;
        RECT 55.660 205.610 55.800 207.330 ;
        RECT 57.040 206.630 57.180 208.010 ;
        RECT 60.200 207.670 60.460 207.990 ;
        RECT 56.980 206.310 57.240 206.630 ;
        RECT 55.600 205.290 55.860 205.610 ;
        RECT 55.140 201.890 55.400 202.210 ;
        RECT 57.040 199.830 57.180 206.310 ;
        RECT 59.740 202.230 60.000 202.550 ;
        RECT 59.800 200.850 59.940 202.230 ;
        RECT 59.740 200.760 60.000 200.850 ;
        RECT 59.340 200.620 60.000 200.760 ;
        RECT 59.340 199.830 59.480 200.620 ;
        RECT 59.740 200.530 60.000 200.620 ;
        RECT 60.260 200.510 60.400 207.670 ;
        RECT 60.720 201.190 60.860 208.350 ;
        RECT 64.400 204.930 64.540 208.690 ;
        RECT 68.480 208.350 68.740 208.670 ;
        RECT 68.940 208.350 69.200 208.670 ;
        RECT 70.780 208.350 71.040 208.670 ;
        RECT 65.260 207.330 65.520 207.650 ;
        RECT 64.340 204.610 64.600 204.930 ;
        RECT 61.120 201.890 61.380 202.210 ;
        RECT 60.660 200.870 60.920 201.190 ;
        RECT 60.200 200.190 60.460 200.510 ;
        RECT 61.180 200.170 61.320 201.890 ;
        RECT 62.960 200.190 63.220 200.510 ;
        RECT 61.120 199.850 61.380 200.170 ;
        RECT 61.580 199.850 61.840 200.170 ;
        RECT 54.680 199.510 54.940 199.830 ;
        RECT 56.520 199.510 56.780 199.830 ;
        RECT 56.980 199.510 57.240 199.830 ;
        RECT 59.280 199.510 59.540 199.830 ;
        RECT 59.740 199.510 60.000 199.830 ;
        RECT 56.580 197.790 56.720 199.510 ;
        RECT 56.520 197.470 56.780 197.790 ;
        RECT 57.040 195.150 57.180 199.510 ;
        RECT 58.360 199.170 58.620 199.490 ;
        RECT 56.580 195.010 57.180 195.150 ;
        RECT 54.220 194.410 54.480 194.730 ;
        RECT 56.580 194.470 56.720 195.010 ;
        RECT 53.760 194.070 54.020 194.390 ;
        RECT 52.840 192.710 53.100 193.030 ;
        RECT 51.920 192.370 52.180 192.690 ;
        RECT 51.920 191.690 52.180 192.010 ;
        RECT 50.540 189.310 50.800 189.630 ;
        RECT 46.400 188.630 46.660 188.950 ;
        RECT 46.460 186.570 46.600 188.630 ;
        RECT 46.860 188.290 47.120 188.610 ;
        RECT 46.920 187.250 47.060 188.290 ;
        RECT 46.860 186.930 47.120 187.250 ;
        RECT 46.400 186.250 46.660 186.570 ;
        RECT 45.940 184.210 46.200 184.530 ;
        RECT 45.080 184.030 45.680 184.170 ;
        RECT 45.080 183.170 45.220 184.030 ;
        RECT 46.000 183.510 46.140 184.210 ;
        RECT 46.460 183.850 46.600 186.250 ;
        RECT 50.600 185.890 50.740 189.310 ;
        RECT 51.980 187.590 52.120 191.690 ;
        RECT 52.380 191.185 52.640 191.330 ;
        RECT 52.370 190.815 52.650 191.185 ;
        RECT 53.300 191.010 53.560 191.330 ;
        RECT 52.380 188.970 52.640 189.290 ;
        RECT 51.920 187.270 52.180 187.590 ;
        RECT 52.440 186.910 52.580 188.970 ;
        RECT 53.360 188.610 53.500 191.010 ;
        RECT 53.300 188.290 53.560 188.610 ;
        RECT 53.820 187.250 53.960 194.070 ;
        RECT 54.280 192.350 54.420 194.410 ;
        RECT 56.120 194.390 56.720 194.470 ;
        RECT 56.060 194.330 56.720 194.390 ;
        RECT 56.060 194.070 56.320 194.330 ;
        RECT 55.140 193.730 55.400 194.050 ;
        RECT 55.200 193.030 55.340 193.730 ;
        RECT 55.140 192.710 55.400 193.030 ;
        RECT 54.220 192.030 54.480 192.350 ;
        RECT 54.680 191.350 54.940 191.670 ;
        RECT 54.220 188.970 54.480 189.290 ;
        RECT 54.280 187.590 54.420 188.970 ;
        RECT 54.740 187.590 54.880 191.350 ;
        RECT 55.200 189.710 55.340 192.710 ;
        RECT 55.200 189.630 55.800 189.710 ;
        RECT 55.200 189.570 55.860 189.630 ;
        RECT 55.600 189.310 55.860 189.570 ;
        RECT 55.140 188.970 55.400 189.290 ;
        RECT 55.200 187.590 55.340 188.970 ;
        RECT 54.220 187.270 54.480 187.590 ;
        RECT 54.680 187.270 54.940 187.590 ;
        RECT 55.140 187.270 55.400 187.590 ;
        RECT 53.760 186.930 54.020 187.250 ;
        RECT 51.000 186.590 51.260 186.910 ;
        RECT 52.380 186.590 52.640 186.910 ;
        RECT 50.540 185.570 50.800 185.890 ;
        RECT 51.060 184.530 51.200 186.590 ;
        RECT 51.000 184.210 51.260 184.530 ;
        RECT 52.380 184.210 52.640 184.530 ;
        RECT 46.400 183.530 46.660 183.850 ;
        RECT 45.940 183.190 46.200 183.510 ;
        RECT 45.020 182.850 45.280 183.170 ;
        RECT 44.100 181.830 44.360 182.150 ;
        RECT 43.640 178.430 43.900 178.750 ;
        RECT 43.640 174.690 43.900 175.010 ;
        RECT 43.700 173.310 43.840 174.690 ;
        RECT 43.640 172.990 43.900 173.310 ;
        RECT 43.180 172.650 43.440 172.970 ;
        RECT 43.640 172.310 43.900 172.630 ;
        RECT 40.420 171.970 40.680 172.290 ;
        RECT 41.340 171.970 41.600 172.290 ;
        RECT 39.960 170.950 40.220 171.270 ;
        RECT 40.480 170.590 40.620 171.970 ;
        RECT 40.420 170.270 40.680 170.590 ;
        RECT 39.040 169.250 39.300 169.570 ;
        RECT 39.500 168.230 39.760 168.550 ;
        RECT 38.580 167.890 38.840 168.210 ;
        RECT 36.170 165.995 37.710 166.365 ;
        RECT 35.820 165.510 36.080 165.830 ;
        RECT 39.560 165.150 39.700 168.230 ;
        RECT 39.500 164.830 39.760 165.150 ;
        RECT 40.420 164.830 40.680 165.150 ;
        RECT 35.360 164.490 35.620 164.810 ;
        RECT 39.560 164.550 39.700 164.830 ;
        RECT 34.900 164.150 35.160 164.470 ;
        RECT 39.560 164.410 40.160 164.550 ;
        RECT 32.870 163.275 34.410 163.645 ;
        RECT 32.140 162.790 32.400 163.110 ;
        RECT 32.140 161.430 32.400 161.750 ;
        RECT 32.200 160.390 32.340 161.430 ;
        RECT 34.960 161.410 35.100 164.150 ;
        RECT 38.120 163.810 38.380 164.130 ;
        RECT 39.500 163.810 39.760 164.130 ;
        RECT 34.900 161.090 35.160 161.410 ;
        RECT 36.170 160.555 37.710 160.925 ;
        RECT 32.140 160.070 32.400 160.390 ;
        RECT 36.740 159.390 37.000 159.710 ;
        RECT 21.100 158.370 21.360 158.690 ;
        RECT 31.680 158.370 31.940 158.690 ;
        RECT 32.870 157.835 34.410 158.205 ;
        RECT 36.800 157.670 36.940 159.390 ;
        RECT 36.740 157.350 37.000 157.670 ;
        RECT 38.180 156.310 38.320 163.810 ;
        RECT 38.580 161.090 38.840 161.410 ;
        RECT 38.640 156.310 38.780 161.090 ;
        RECT 39.560 157.670 39.700 163.810 ;
        RECT 40.020 162.090 40.160 164.410 ;
        RECT 40.480 163.110 40.620 164.830 ;
        RECT 40.420 162.790 40.680 163.110 ;
        RECT 40.480 162.090 40.620 162.790 ;
        RECT 39.960 161.770 40.220 162.090 ;
        RECT 40.420 161.770 40.680 162.090 ;
        RECT 40.020 160.390 40.160 161.770 ;
        RECT 41.400 161.750 41.540 171.970 ;
        RECT 43.700 171.270 43.840 172.310 ;
        RECT 43.640 170.950 43.900 171.270 ;
        RECT 43.640 166.870 43.900 167.190 ;
        RECT 43.700 165.830 43.840 166.870 ;
        RECT 41.800 165.510 42.060 165.830 ;
        RECT 43.640 165.510 43.900 165.830 ;
        RECT 41.340 161.430 41.600 161.750 ;
        RECT 39.960 160.070 40.220 160.390 ;
        RECT 39.500 157.350 39.760 157.670 ;
        RECT 38.120 155.990 38.380 156.310 ;
        RECT 38.580 155.990 38.840 156.310 ;
        RECT 36.170 155.115 37.710 155.485 ;
        RECT 16.040 153.950 16.300 154.270 ;
        RECT 16.100 153.105 16.240 153.950 ;
        RECT 16.030 152.735 16.310 153.105 ;
        RECT 32.870 152.395 34.410 152.765 ;
        RECT 35.360 151.910 35.620 152.230 ;
        RECT 32.600 150.890 32.860 151.210 ;
        RECT 15.890 149.110 16.310 149.560 ;
        RECT 32.660 148.830 32.800 150.890 ;
        RECT 33.520 150.550 33.780 150.870 ;
        RECT 29.380 148.510 29.640 148.830 ;
        RECT 32.600 148.510 32.860 148.830 ;
        RECT 29.440 143.050 29.580 148.510 ;
        RECT 32.660 148.230 32.800 148.510 ;
        RECT 33.580 148.490 33.720 150.550 ;
        RECT 33.980 150.210 34.240 150.530 ;
        RECT 34.040 149.170 34.180 150.210 ;
        RECT 35.420 149.420 35.560 151.910 ;
        RECT 35.820 151.570 36.080 151.890 ;
        RECT 34.500 149.280 35.560 149.420 ;
        RECT 33.980 148.850 34.240 149.170 ;
        RECT 32.200 148.090 32.800 148.230 ;
        RECT 33.520 148.170 33.780 148.490 ;
        RECT 34.500 148.150 34.640 149.280 ;
        RECT 34.900 148.510 35.160 148.830 ;
        RECT 32.200 146.790 32.340 148.090 ;
        RECT 34.440 147.830 34.700 148.150 ;
        RECT 32.870 146.955 34.410 147.325 ;
        RECT 32.140 146.470 32.400 146.790 ;
        RECT 34.960 145.770 35.100 148.510 ;
        RECT 34.900 145.450 35.160 145.770 ;
        RECT 29.380 142.730 29.640 143.050 ;
        RECT 29.440 138.630 29.580 142.730 ;
        RECT 32.140 142.050 32.400 142.370 ;
        RECT 32.200 139.990 32.340 142.050 ;
        RECT 32.870 141.515 34.410 141.885 ;
        RECT 34.960 140.670 35.100 145.450 ;
        RECT 35.420 143.050 35.560 149.280 ;
        RECT 35.880 148.830 36.020 151.570 ;
        RECT 39.040 151.230 39.300 151.550 ;
        RECT 38.580 150.890 38.840 151.210 ;
        RECT 38.120 150.550 38.380 150.870 ;
        RECT 36.170 149.675 37.710 150.045 ;
        RECT 35.820 148.510 36.080 148.830 ;
        RECT 36.280 147.490 36.540 147.810 ;
        RECT 36.340 145.430 36.480 147.490 ;
        RECT 38.180 146.450 38.320 150.550 ;
        RECT 38.120 146.130 38.380 146.450 ;
        RECT 36.280 145.110 36.540 145.430 ;
        RECT 35.820 144.770 36.080 145.090 ;
        RECT 35.360 142.730 35.620 143.050 ;
        RECT 35.360 142.050 35.620 142.370 ;
        RECT 34.900 140.350 35.160 140.670 ;
        RECT 32.140 139.670 32.400 139.990 ;
        RECT 34.900 139.670 35.160 139.990 ;
        RECT 29.380 138.310 29.640 138.630 ;
        RECT 22.940 137.630 23.200 137.950 ;
        RECT 19.260 136.610 19.520 136.930 ;
        RECT 19.320 135.425 19.460 136.610 ;
        RECT 19.250 135.055 19.530 135.425 ;
        RECT 20.640 134.570 20.900 134.890 ;
        RECT 16.040 133.890 16.300 134.210 ;
        RECT 16.100 132.705 16.240 133.890 ;
        RECT 16.030 132.335 16.310 132.705 ;
        RECT 18.800 132.190 19.060 132.510 ;
        RECT 18.860 130.470 19.000 132.190 ;
        RECT 19.260 131.850 19.520 132.170 ;
        RECT 18.800 130.150 19.060 130.470 ;
        RECT 16.490 128.255 16.770 128.625 ;
        RECT 16.560 127.410 16.700 128.255 ;
        RECT 16.500 127.090 16.760 127.410 ;
        RECT 16.040 125.905 16.300 126.050 ;
        RECT 16.030 125.535 16.310 125.905 ;
        RECT 19.320 124.430 19.460 131.850 ;
        RECT 20.700 131.490 20.840 134.570 ;
        RECT 23.000 132.850 23.140 137.630 ;
        RECT 32.870 136.075 34.410 136.445 ;
        RECT 34.960 134.550 35.100 139.670 ;
        RECT 35.420 138.630 35.560 142.050 ;
        RECT 35.880 141.350 36.020 144.770 ;
        RECT 36.170 144.235 37.710 144.605 ;
        RECT 38.180 144.070 38.320 146.130 ;
        RECT 38.640 145.770 38.780 150.890 ;
        RECT 39.100 145.770 39.240 151.230 ;
        RECT 41.860 151.210 42.000 165.510 ;
        RECT 44.160 165.150 44.300 181.830 ;
        RECT 44.560 178.090 44.820 178.410 ;
        RECT 44.620 170.250 44.760 178.090 ;
        RECT 45.080 176.370 45.220 182.850 ;
        RECT 46.460 180.790 46.600 183.530 ;
        RECT 47.780 181.150 48.040 181.470 ;
        RECT 46.400 180.470 46.660 180.790 ;
        RECT 47.840 178.410 47.980 181.150 ;
        RECT 47.780 178.090 48.040 178.410 ;
        RECT 45.480 177.410 45.740 177.730 ;
        RECT 45.020 176.050 45.280 176.370 ;
        RECT 45.540 176.030 45.680 177.410 ;
        RECT 45.480 175.710 45.740 176.030 ;
        RECT 45.940 175.710 46.200 176.030 ;
        RECT 46.000 173.990 46.140 175.710 ;
        RECT 45.940 173.670 46.200 173.990 ;
        RECT 48.240 172.650 48.500 172.970 ;
        RECT 48.300 170.590 48.440 172.650 ;
        RECT 48.240 170.270 48.500 170.590 ;
        RECT 44.560 169.930 44.820 170.250 ;
        RECT 45.480 169.930 45.740 170.250 ;
        RECT 46.860 169.930 47.120 170.250 ;
        RECT 48.700 169.930 48.960 170.250 ;
        RECT 50.540 169.930 50.800 170.250 ;
        RECT 44.620 168.550 44.760 169.930 ;
        RECT 44.560 168.230 44.820 168.550 ;
        RECT 45.540 167.870 45.680 169.930 ;
        RECT 45.940 169.250 46.200 169.570 ;
        RECT 45.480 167.550 45.740 167.870 ;
        RECT 45.020 166.530 45.280 166.850 ;
        RECT 45.080 165.150 45.220 166.530 ;
        RECT 45.540 165.830 45.680 167.550 ;
        RECT 45.480 165.510 45.740 165.830 ;
        RECT 46.000 165.150 46.140 169.250 ;
        RECT 46.920 168.210 47.060 169.930 ;
        RECT 48.760 168.550 48.900 169.930 ;
        RECT 47.780 168.230 48.040 168.550 ;
        RECT 48.700 168.230 48.960 168.550 ;
        RECT 46.860 167.890 47.120 168.210 ;
        RECT 47.840 167.530 47.980 168.230 ;
        RECT 50.600 167.530 50.740 169.930 ;
        RECT 47.780 167.210 48.040 167.530 ;
        RECT 50.540 167.210 50.800 167.530 ;
        RECT 47.320 166.530 47.580 166.850 ;
        RECT 47.380 165.150 47.520 166.530 ;
        RECT 44.100 164.830 44.360 165.150 ;
        RECT 45.020 164.830 45.280 165.150 ;
        RECT 45.940 164.830 46.200 165.150 ;
        RECT 46.400 164.830 46.660 165.150 ;
        RECT 47.320 164.830 47.580 165.150 ;
        RECT 43.180 164.490 43.440 164.810 ;
        RECT 43.240 161.750 43.380 164.490 ;
        RECT 46.000 163.190 46.140 164.830 ;
        RECT 46.460 164.130 46.600 164.830 ;
        RECT 47.840 164.130 47.980 167.210 ;
        RECT 46.400 163.810 46.660 164.130 ;
        RECT 47.320 163.810 47.580 164.130 ;
        RECT 47.780 163.810 48.040 164.130 ;
        RECT 46.000 163.050 47.060 163.190 ;
        RECT 47.380 163.110 47.520 163.810 ;
        RECT 43.180 161.430 43.440 161.750 ;
        RECT 43.240 160.390 43.380 161.430 ;
        RECT 46.400 161.090 46.660 161.410 ;
        RECT 43.180 160.070 43.440 160.390 ;
        RECT 46.460 159.710 46.600 161.090 ;
        RECT 46.400 159.390 46.660 159.710 ;
        RECT 41.800 151.120 42.060 151.210 ;
        RECT 41.800 150.980 42.920 151.120 ;
        RECT 41.800 150.890 42.060 150.980 ;
        RECT 39.500 150.550 39.760 150.870 ;
        RECT 39.560 150.270 39.700 150.550 ;
        RECT 39.560 150.130 40.160 150.270 ;
        RECT 40.020 147.810 40.160 150.130 ;
        RECT 39.960 147.490 40.220 147.810 ;
        RECT 40.020 145.770 40.160 147.490 ;
        RECT 42.780 145.770 42.920 150.980 ;
        RECT 46.920 150.870 47.060 163.050 ;
        RECT 47.320 162.790 47.580 163.110 ;
        RECT 47.380 162.430 47.520 162.790 ;
        RECT 47.320 162.110 47.580 162.430 ;
        RECT 47.840 162.090 47.980 163.810 ;
        RECT 50.600 162.090 50.740 167.210 ;
        RECT 47.780 161.770 48.040 162.090 ;
        RECT 50.540 161.770 50.800 162.090 ;
        RECT 47.780 151.910 48.040 152.230 ;
        RECT 46.860 150.550 47.120 150.870 ;
        RECT 46.400 150.210 46.660 150.530 ;
        RECT 47.320 150.210 47.580 150.530 ;
        RECT 46.460 148.830 46.600 150.210 ;
        RECT 47.380 149.170 47.520 150.210 ;
        RECT 47.840 149.170 47.980 151.910 ;
        RECT 50.540 150.210 50.800 150.530 ;
        RECT 47.320 148.850 47.580 149.170 ;
        RECT 47.780 148.850 48.040 149.170 ;
        RECT 46.400 148.510 46.660 148.830 ;
        RECT 46.860 148.510 47.120 148.830 ;
        RECT 46.920 145.770 47.060 148.510 ;
        RECT 47.840 146.450 47.980 148.850 ;
        RECT 50.600 148.830 50.740 150.210 ;
        RECT 50.080 148.510 50.340 148.830 ;
        RECT 50.540 148.510 50.800 148.830 ;
        RECT 50.140 147.810 50.280 148.510 ;
        RECT 51.060 148.490 51.200 184.210 ;
        RECT 51.920 172.310 52.180 172.630 ;
        RECT 51.980 171.270 52.120 172.310 ;
        RECT 51.920 170.950 52.180 171.270 ;
        RECT 52.440 167.870 52.580 184.210 ;
        RECT 54.740 183.510 54.880 187.270 ;
        RECT 55.600 186.590 55.860 186.910 ;
        RECT 55.660 184.530 55.800 186.590 ;
        RECT 56.120 186.230 56.260 194.070 ;
        RECT 58.420 194.050 58.560 199.170 ;
        RECT 59.340 197.110 59.480 199.510 ;
        RECT 59.800 197.790 59.940 199.510 ;
        RECT 59.740 197.470 60.000 197.790 ;
        RECT 59.280 196.790 59.540 197.110 ;
        RECT 58.820 194.750 59.080 195.070 ;
        RECT 58.360 193.730 58.620 194.050 ;
        RECT 58.880 192.350 59.020 194.750 ;
        RECT 58.820 192.030 59.080 192.350 ;
        RECT 59.280 192.030 59.540 192.350 ;
        RECT 57.440 191.920 57.700 192.010 ;
        RECT 57.040 191.780 57.700 191.920 ;
        RECT 57.040 191.330 57.180 191.780 ;
        RECT 57.440 191.690 57.700 191.780 ;
        RECT 56.980 191.010 57.240 191.330 ;
        RECT 57.440 191.010 57.700 191.330 ;
        RECT 57.500 190.310 57.640 191.010 ;
        RECT 57.440 189.990 57.700 190.310 ;
        RECT 57.900 189.650 58.160 189.970 ;
        RECT 57.440 188.970 57.700 189.290 ;
        RECT 56.520 188.290 56.780 188.610 ;
        RECT 56.060 185.910 56.320 186.230 ;
        RECT 55.600 184.210 55.860 184.530 ;
        RECT 56.580 183.850 56.720 188.290 ;
        RECT 57.500 187.500 57.640 188.970 ;
        RECT 57.040 187.360 57.640 187.500 ;
        RECT 57.040 186.910 57.180 187.360 ;
        RECT 56.980 186.590 57.240 186.910 ;
        RECT 57.440 186.590 57.700 186.910 ;
        RECT 57.040 183.850 57.180 186.590 ;
        RECT 57.500 184.190 57.640 186.590 ;
        RECT 57.960 186.230 58.100 189.650 ;
        RECT 59.340 189.290 59.480 192.030 ;
        RECT 59.280 188.970 59.540 189.290 ;
        RECT 59.800 186.910 59.940 197.470 ;
        RECT 61.640 195.750 61.780 199.850 ;
        RECT 63.020 198.470 63.160 200.190 ;
        RECT 64.400 200.170 64.540 204.610 ;
        RECT 64.340 199.850 64.600 200.170 ;
        RECT 62.960 198.150 63.220 198.470 ;
        RECT 65.320 197.790 65.460 207.330 ;
        RECT 65.720 205.290 65.980 205.610 ;
        RECT 65.780 202.890 65.920 205.290 ;
        RECT 68.540 203.910 68.680 208.350 ;
        RECT 68.480 203.590 68.740 203.910 ;
        RECT 66.180 202.910 66.440 203.230 ;
        RECT 65.720 202.570 65.980 202.890 ;
        RECT 65.780 200.510 65.920 202.570 ;
        RECT 65.720 200.190 65.980 200.510 ;
        RECT 66.240 199.490 66.380 202.910 ;
        RECT 69.000 201.190 69.140 208.350 ;
        RECT 69.400 207.330 69.660 207.650 ;
        RECT 69.460 205.270 69.600 207.330 ;
        RECT 69.400 204.950 69.660 205.270 ;
        RECT 69.400 202.910 69.660 203.230 ;
        RECT 69.460 201.190 69.600 202.910 ;
        RECT 68.940 200.870 69.200 201.190 ;
        RECT 69.400 200.870 69.660 201.190 ;
        RECT 67.100 199.510 67.360 199.830 ;
        RECT 66.180 199.170 66.440 199.490 ;
        RECT 65.260 197.470 65.520 197.790 ;
        RECT 61.580 195.430 61.840 195.750 ;
        RECT 60.660 195.090 60.920 195.410 ;
        RECT 60.200 191.010 60.460 191.330 ;
        RECT 60.260 187.250 60.400 191.010 ;
        RECT 60.720 189.630 60.860 195.090 ;
        RECT 61.640 192.350 61.780 195.430 ;
        RECT 62.500 194.410 62.760 194.730 ;
        RECT 61.580 192.030 61.840 192.350 ;
        RECT 61.120 191.010 61.380 191.330 ;
        RECT 60.660 189.310 60.920 189.630 ;
        RECT 61.180 189.030 61.320 191.010 ;
        RECT 60.720 188.890 61.320 189.030 ;
        RECT 60.720 187.590 60.860 188.890 ;
        RECT 61.120 188.290 61.380 188.610 ;
        RECT 61.180 187.590 61.320 188.290 ;
        RECT 60.660 187.270 60.920 187.590 ;
        RECT 61.120 187.270 61.380 187.590 ;
        RECT 60.200 186.930 60.460 187.250 ;
        RECT 59.280 186.590 59.540 186.910 ;
        RECT 59.740 186.590 60.000 186.910 ;
        RECT 61.580 186.590 61.840 186.910 ;
        RECT 57.900 185.910 58.160 186.230 ;
        RECT 57.440 183.870 57.700 184.190 ;
        RECT 56.520 183.530 56.780 183.850 ;
        RECT 56.980 183.530 57.240 183.850 ;
        RECT 54.680 183.190 54.940 183.510 ;
        RECT 54.220 182.850 54.480 183.170 ;
        RECT 52.840 181.150 53.100 181.470 ;
        RECT 52.900 178.750 53.040 181.150 ;
        RECT 54.280 179.090 54.420 182.850 ;
        RECT 57.500 181.470 57.640 183.870 ;
        RECT 55.600 181.150 55.860 181.470 ;
        RECT 57.440 181.150 57.700 181.470 ;
        RECT 54.220 178.770 54.480 179.090 ;
        RECT 52.840 178.430 53.100 178.750 ;
        RECT 52.900 172.970 53.040 178.430 ;
        RECT 53.300 177.750 53.560 178.070 ;
        RECT 52.840 172.650 53.100 172.970 ;
        RECT 53.360 169.570 53.500 177.750 ;
        RECT 53.300 169.250 53.560 169.570 ;
        RECT 55.660 167.870 55.800 181.150 ;
        RECT 57.960 179.090 58.100 185.910 ;
        RECT 59.340 183.170 59.480 186.590 ;
        RECT 61.120 186.250 61.380 186.570 ;
        RECT 61.180 184.170 61.320 186.250 ;
        RECT 61.640 184.870 61.780 186.590 ;
        RECT 61.580 184.550 61.840 184.870 ;
        RECT 61.180 184.030 61.780 184.170 ;
        RECT 60.200 183.530 60.460 183.850 ;
        RECT 59.280 182.850 59.540 183.170 ;
        RECT 60.260 181.810 60.400 183.530 ;
        RECT 61.640 183.170 61.780 184.030 ;
        RECT 62.040 183.530 62.300 183.850 ;
        RECT 61.580 182.850 61.840 183.170 ;
        RECT 60.200 181.490 60.460 181.810 ;
        RECT 59.740 180.810 60.000 181.130 ;
        RECT 58.360 180.130 58.620 180.450 ;
        RECT 57.900 178.770 58.160 179.090 ;
        RECT 58.420 178.070 58.560 180.130 ;
        RECT 59.800 178.410 59.940 180.810 ;
        RECT 60.260 180.450 60.400 181.490 ;
        RECT 60.660 181.150 60.920 181.470 ;
        RECT 60.200 180.130 60.460 180.450 ;
        RECT 60.720 178.410 60.860 181.150 ;
        RECT 61.640 178.410 61.780 182.850 ;
        RECT 62.100 181.470 62.240 183.530 ;
        RECT 62.040 181.150 62.300 181.470 ;
        RECT 62.560 180.870 62.700 194.410 ;
        RECT 66.240 192.010 66.380 199.170 ;
        RECT 67.160 197.110 67.300 199.510 ;
        RECT 68.480 199.170 68.740 199.490 ;
        RECT 68.540 198.130 68.680 199.170 ;
        RECT 68.480 197.810 68.740 198.130 ;
        RECT 68.940 197.130 69.200 197.450 ;
        RECT 67.100 196.790 67.360 197.110 ;
        RECT 67.560 196.450 67.820 196.770 ;
        RECT 67.620 195.750 67.760 196.450 ;
        RECT 67.560 195.430 67.820 195.750 ;
        RECT 69.000 192.350 69.140 197.130 ;
        RECT 66.640 192.030 66.900 192.350 ;
        RECT 68.940 192.030 69.200 192.350 ;
        RECT 62.960 191.690 63.220 192.010 ;
        RECT 66.180 191.690 66.440 192.010 ;
        RECT 63.020 184.190 63.160 191.690 ;
        RECT 65.260 191.350 65.520 191.670 ;
        RECT 63.880 191.010 64.140 191.330 ;
        RECT 63.940 189.970 64.080 191.010 ;
        RECT 63.880 189.650 64.140 189.970 ;
        RECT 65.320 189.290 65.460 191.350 ;
        RECT 65.710 190.815 65.990 191.185 ;
        RECT 65.780 189.290 65.920 190.815 ;
        RECT 66.240 190.310 66.380 191.690 ;
        RECT 66.700 190.310 66.840 192.030 ;
        RECT 67.100 191.690 67.360 192.010 ;
        RECT 66.180 189.990 66.440 190.310 ;
        RECT 66.640 189.990 66.900 190.310 ;
        RECT 67.160 189.630 67.300 191.690 ;
        RECT 67.100 189.310 67.360 189.630 ;
        RECT 65.260 188.970 65.520 189.290 ;
        RECT 65.720 188.970 65.980 189.290 ;
        RECT 67.160 186.230 67.300 189.310 ;
        RECT 69.000 189.290 69.140 192.030 ;
        RECT 69.460 189.970 69.600 200.870 ;
        RECT 70.840 200.850 70.980 208.350 ;
        RECT 82.740 208.010 83.000 208.330 ;
        RECT 71.700 207.330 71.960 207.650 ;
        RECT 71.760 203.230 71.900 207.330 ;
        RECT 82.800 204.930 82.940 208.010 ;
        RECT 80.440 204.610 80.700 204.930 ;
        RECT 82.740 204.610 83.000 204.930 ;
        RECT 80.500 203.230 80.640 204.610 ;
        RECT 71.240 202.910 71.500 203.230 ;
        RECT 71.700 202.910 71.960 203.230 ;
        RECT 80.440 202.910 80.700 203.230 ;
        RECT 81.820 202.910 82.080 203.230 ;
        RECT 71.300 202.630 71.440 202.910 ;
        RECT 71.300 202.490 71.900 202.630 ;
        RECT 70.780 200.530 71.040 200.850 ;
        RECT 70.840 197.790 70.980 200.530 ;
        RECT 71.760 200.170 71.900 202.490 ;
        RECT 71.700 199.850 71.960 200.170 ;
        RECT 70.780 197.470 71.040 197.790 ;
        RECT 69.860 191.010 70.120 191.330 ;
        RECT 69.400 189.650 69.660 189.970 ;
        RECT 69.920 189.290 70.060 191.010 ;
        RECT 68.940 188.970 69.200 189.290 ;
        RECT 69.860 188.970 70.120 189.290 ;
        RECT 71.240 188.630 71.500 188.950 ;
        RECT 69.400 188.290 69.660 188.610 ;
        RECT 69.460 186.910 69.600 188.290 ;
        RECT 71.300 187.590 71.440 188.630 ;
        RECT 71.240 187.270 71.500 187.590 ;
        RECT 69.400 186.590 69.660 186.910 ;
        RECT 67.100 185.910 67.360 186.230 ;
        RECT 63.880 185.570 64.140 185.890 ;
        RECT 69.860 185.570 70.120 185.890 ;
        RECT 62.960 183.870 63.220 184.190 ;
        RECT 63.940 181.810 64.080 185.570 ;
        RECT 69.920 184.530 70.060 185.570 ;
        RECT 69.860 184.210 70.120 184.530 ;
        RECT 69.920 183.850 70.060 184.210 ;
        RECT 69.860 183.530 70.120 183.850 ;
        RECT 71.240 183.530 71.500 183.850 ;
        RECT 66.180 182.850 66.440 183.170 ;
        RECT 65.260 181.830 65.520 182.150 ;
        RECT 63.880 181.490 64.140 181.810 ;
        RECT 65.320 181.470 65.460 181.830 ;
        RECT 65.720 181.490 65.980 181.810 ;
        RECT 63.420 181.150 63.680 181.470 ;
        RECT 65.260 181.150 65.520 181.470 ;
        RECT 62.560 180.730 63.160 180.870 ;
        RECT 62.500 180.130 62.760 180.450 ;
        RECT 62.560 178.410 62.700 180.130 ;
        RECT 63.020 179.090 63.160 180.730 ;
        RECT 63.480 179.090 63.620 181.150 ;
        RECT 62.960 178.770 63.220 179.090 ;
        RECT 63.420 178.770 63.680 179.090 ;
        RECT 59.740 178.090 60.000 178.410 ;
        RECT 60.200 178.090 60.460 178.410 ;
        RECT 60.660 178.090 60.920 178.410 ;
        RECT 61.580 178.090 61.840 178.410 ;
        RECT 62.500 178.090 62.760 178.410 ;
        RECT 58.360 177.750 58.620 178.070 ;
        RECT 60.260 176.710 60.400 178.090 ;
        RECT 60.200 176.390 60.460 176.710 ;
        RECT 60.720 176.370 60.860 178.090 ;
        RECT 62.040 176.390 62.300 176.710 ;
        RECT 60.660 176.050 60.920 176.370 ;
        RECT 62.100 176.030 62.240 176.390 ;
        RECT 63.020 176.110 63.160 178.770 ;
        RECT 63.880 178.090 64.140 178.410 ;
        RECT 63.940 176.710 64.080 178.090 ;
        RECT 63.880 176.390 64.140 176.710 ;
        RECT 63.020 176.030 63.620 176.110 ;
        RECT 62.040 175.710 62.300 176.030 ;
        RECT 63.020 175.970 63.680 176.030 ;
        RECT 63.420 175.710 63.680 175.970 ;
        RECT 65.320 174.750 65.460 181.150 ;
        RECT 64.860 174.610 65.460 174.750 ;
        RECT 58.360 173.330 58.620 173.650 ;
        RECT 56.980 170.950 57.240 171.270 ;
        RECT 57.040 170.250 57.180 170.950 ;
        RECT 58.420 170.590 58.560 173.330 ;
        RECT 61.120 172.310 61.380 172.630 ;
        RECT 58.360 170.270 58.620 170.590 ;
        RECT 61.180 170.250 61.320 172.310 ;
        RECT 63.420 171.970 63.680 172.290 ;
        RECT 63.480 170.250 63.620 171.970 ;
        RECT 56.980 169.930 57.240 170.250 ;
        RECT 61.120 169.930 61.380 170.250 ;
        RECT 63.420 169.930 63.680 170.250 ;
        RECT 52.380 167.550 52.640 167.870 ;
        RECT 55.600 167.550 55.860 167.870 ;
        RECT 52.440 148.830 52.580 167.550 ;
        RECT 54.220 164.830 54.480 165.150 ;
        RECT 54.280 163.110 54.420 164.830 ;
        RECT 55.660 164.810 55.800 167.550 ;
        RECT 57.040 167.530 57.180 169.930 ;
        RECT 58.360 169.250 58.620 169.570 ;
        RECT 58.820 169.250 59.080 169.570 ;
        RECT 56.980 167.210 57.240 167.530 ;
        RECT 58.420 165.490 58.560 169.250 ;
        RECT 58.880 167.530 59.020 169.250 ;
        RECT 58.820 167.210 59.080 167.530 ;
        RECT 58.360 165.170 58.620 165.490 ;
        RECT 55.600 164.490 55.860 164.810 ;
        RECT 54.220 162.790 54.480 163.110 ;
        RECT 55.660 160.050 55.800 164.490 ;
        RECT 55.600 159.730 55.860 160.050 ;
        RECT 62.500 158.370 62.760 158.690 ;
        RECT 56.060 157.010 56.320 157.330 ;
        RECT 56.120 154.270 56.260 157.010 ;
        RECT 57.440 156.330 57.700 156.650 ;
        RECT 57.500 154.950 57.640 156.330 ;
        RECT 61.580 155.990 61.840 156.310 ;
        RECT 57.440 154.630 57.700 154.950 ;
        RECT 57.960 154.270 59.480 154.350 ;
        RECT 56.060 154.180 56.320 154.270 ;
        RECT 57.960 154.210 59.540 154.270 ;
        RECT 56.060 154.040 56.720 154.180 ;
        RECT 56.060 153.950 56.320 154.040 ;
        RECT 56.580 151.890 56.720 154.040 ;
        RECT 57.960 153.590 58.100 154.210 ;
        RECT 59.280 153.950 59.540 154.210 ;
        RECT 58.820 153.610 59.080 153.930 ;
        RECT 57.900 153.270 58.160 153.590 ;
        RECT 56.520 151.570 56.780 151.890 ;
        RECT 58.880 151.630 59.020 153.610 ;
        RECT 60.660 152.930 60.920 153.250 ;
        RECT 60.720 152.230 60.860 152.930 ;
        RECT 60.660 151.910 60.920 152.230 ;
        RECT 55.140 150.890 55.400 151.210 ;
        RECT 56.060 150.890 56.320 151.210 ;
        RECT 56.580 150.950 56.720 151.570 ;
        RECT 58.880 151.550 60.400 151.630 ;
        RECT 58.820 151.490 60.400 151.550 ;
        RECT 58.820 151.230 59.080 151.490 ;
        RECT 54.680 150.210 54.940 150.530 ;
        RECT 54.740 149.170 54.880 150.210 ;
        RECT 52.900 148.830 54.420 148.910 ;
        RECT 54.680 148.850 54.940 149.170 ;
        RECT 51.460 148.510 51.720 148.830 ;
        RECT 52.380 148.510 52.640 148.830 ;
        RECT 52.900 148.770 54.480 148.830 ;
        RECT 51.000 148.170 51.260 148.490 ;
        RECT 50.080 147.490 50.340 147.810 ;
        RECT 51.520 146.790 51.660 148.510 ;
        RECT 52.900 148.490 53.040 148.770 ;
        RECT 54.220 148.510 54.480 148.770 ;
        RECT 52.840 148.170 53.100 148.490 ;
        RECT 51.460 146.470 51.720 146.790 ;
        RECT 47.780 146.130 48.040 146.450 ;
        RECT 38.580 145.450 38.840 145.770 ;
        RECT 39.040 145.450 39.300 145.770 ;
        RECT 39.960 145.450 40.220 145.770 ;
        RECT 40.880 145.450 41.140 145.770 ;
        RECT 42.260 145.450 42.520 145.770 ;
        RECT 42.720 145.450 42.980 145.770 ;
        RECT 46.860 145.450 47.120 145.770 ;
        RECT 38.120 143.750 38.380 144.070 ;
        RECT 38.640 143.390 38.780 145.450 ;
        RECT 39.100 144.070 39.240 145.450 ;
        RECT 39.040 143.750 39.300 144.070 ;
        RECT 38.580 143.070 38.840 143.390 ;
        RECT 39.100 143.050 39.240 143.750 ;
        RECT 40.020 143.730 40.160 145.450 ;
        RECT 40.940 144.070 41.080 145.450 ;
        RECT 42.320 145.090 42.460 145.450 ;
        RECT 42.260 144.770 42.520 145.090 ;
        RECT 45.940 144.770 46.200 145.090 ;
        RECT 40.880 143.750 41.140 144.070 ;
        RECT 39.960 143.410 40.220 143.730 ;
        RECT 39.040 142.730 39.300 143.050 ;
        RECT 38.580 142.050 38.840 142.370 ;
        RECT 35.820 141.030 36.080 141.350 ;
        RECT 35.820 140.350 36.080 140.670 ;
        RECT 35.360 138.310 35.620 138.630 ;
        RECT 35.880 137.950 36.020 140.350 ;
        RECT 38.640 140.330 38.780 142.050 ;
        RECT 40.940 141.350 41.080 143.750 ;
        RECT 40.880 141.030 41.140 141.350 ;
        RECT 38.580 140.010 38.840 140.330 ;
        RECT 36.170 138.795 37.710 139.165 ;
        RECT 35.820 137.630 36.080 137.950 ;
        RECT 35.880 135.230 36.020 137.630 ;
        RECT 38.640 137.610 38.780 140.010 ;
        RECT 45.020 139.670 45.280 139.990 ;
        RECT 39.500 138.310 39.760 138.630 ;
        RECT 42.260 138.310 42.520 138.630 ;
        RECT 39.560 137.950 39.700 138.310 ;
        RECT 42.320 137.950 42.460 138.310 ;
        RECT 45.080 138.290 45.220 139.670 ;
        RECT 45.020 137.970 45.280 138.290 ;
        RECT 39.500 137.630 39.760 137.950 ;
        RECT 42.260 137.630 42.520 137.950 ;
        RECT 42.720 137.630 42.980 137.950 ;
        RECT 38.580 137.290 38.840 137.610 ;
        RECT 41.800 136.950 42.060 137.270 ;
        RECT 36.740 136.610 37.000 136.930 ;
        RECT 39.500 136.610 39.760 136.930 ;
        RECT 36.800 135.870 36.940 136.610 ;
        RECT 39.560 135.910 39.700 136.610 ;
        RECT 36.340 135.730 36.940 135.870 ;
        RECT 35.820 134.910 36.080 135.230 ;
        RECT 34.900 134.230 35.160 134.550 ;
        RECT 22.940 132.530 23.200 132.850 ;
        RECT 20.640 131.170 20.900 131.490 ;
        RECT 20.700 129.450 20.840 131.170 ;
        RECT 23.000 130.470 23.140 132.530 ;
        RECT 35.880 132.510 36.020 134.910 ;
        RECT 36.340 134.550 36.480 135.730 ;
        RECT 39.500 135.590 39.760 135.910 ;
        RECT 36.280 134.230 36.540 134.550 ;
        RECT 38.120 133.890 38.380 134.210 ;
        RECT 36.170 133.355 37.710 133.725 ;
        RECT 38.180 132.850 38.320 133.890 ;
        RECT 38.120 132.530 38.380 132.850 ;
        RECT 28.000 132.190 28.260 132.510 ;
        RECT 35.820 132.190 36.080 132.510 ;
        RECT 28.060 130.470 28.200 132.190 ;
        RECT 41.860 132.170 42.000 136.950 ;
        RECT 42.320 136.930 42.460 137.630 ;
        RECT 42.780 137.270 42.920 137.630 ;
        RECT 42.720 136.950 42.980 137.270 ;
        RECT 46.000 136.930 46.140 144.770 ;
        RECT 46.920 137.610 47.060 145.450 ;
        RECT 52.900 140.670 53.040 148.170 ;
        RECT 55.200 148.150 55.340 150.890 ;
        RECT 56.120 149.170 56.260 150.890 ;
        RECT 56.580 150.870 57.640 150.950 ;
        RECT 56.520 150.810 57.640 150.870 ;
        RECT 56.520 150.550 56.780 150.810 ;
        RECT 56.980 150.210 57.240 150.530 ;
        RECT 56.060 148.850 56.320 149.170 ;
        RECT 57.040 148.830 57.180 150.210 ;
        RECT 56.520 148.510 56.780 148.830 ;
        RECT 56.980 148.510 57.240 148.830 ;
        RECT 55.140 147.830 55.400 148.150 ;
        RECT 54.680 147.490 54.940 147.810 ;
        RECT 54.220 143.410 54.480 143.730 ;
        RECT 53.760 143.070 54.020 143.390 ;
        RECT 53.820 141.010 53.960 143.070 ;
        RECT 53.760 140.690 54.020 141.010 ;
        RECT 52.840 140.350 53.100 140.670 ;
        RECT 50.080 140.010 50.340 140.330 ;
        RECT 50.140 137.950 50.280 140.010 ;
        RECT 50.080 137.630 50.340 137.950 ;
        RECT 46.860 137.290 47.120 137.610 ;
        RECT 42.260 136.610 42.520 136.930 ;
        RECT 45.940 136.610 46.200 136.930 ;
        RECT 42.320 133.190 42.460 136.610 ;
        RECT 46.920 135.910 47.060 137.290 ;
        RECT 49.160 136.610 49.420 136.930 ;
        RECT 49.220 135.910 49.360 136.610 ;
        RECT 44.100 135.590 44.360 135.910 ;
        RECT 46.860 135.590 47.120 135.910 ;
        RECT 49.160 135.590 49.420 135.910 ;
        RECT 44.160 133.190 44.300 135.590 ;
        RECT 50.140 135.570 50.280 137.630 ;
        RECT 52.900 137.610 53.040 140.350 ;
        RECT 54.280 140.070 54.420 143.410 ;
        RECT 54.740 143.390 54.880 147.490 ;
        RECT 54.680 143.070 54.940 143.390 ;
        RECT 55.600 143.070 55.860 143.390 ;
        RECT 54.680 142.050 54.940 142.370 ;
        RECT 53.820 139.930 54.420 140.070 ;
        RECT 52.840 137.290 53.100 137.610 ;
        RECT 48.240 135.310 48.500 135.570 ;
        RECT 47.380 135.250 48.500 135.310 ;
        RECT 50.080 135.250 50.340 135.570 ;
        RECT 47.380 135.170 48.440 135.250 ;
        RECT 47.380 134.890 47.520 135.170 ;
        RECT 52.900 134.890 53.040 137.290 ;
        RECT 53.300 136.610 53.560 136.930 ;
        RECT 53.360 135.910 53.500 136.610 ;
        RECT 53.300 135.590 53.560 135.910 ;
        RECT 47.320 134.570 47.580 134.890 ;
        RECT 52.840 134.570 53.100 134.890 ;
        RECT 44.560 133.890 44.820 134.210 ;
        RECT 42.260 132.870 42.520 133.190 ;
        RECT 44.100 132.870 44.360 133.190 ;
        RECT 44.620 132.510 44.760 133.890 ;
        RECT 52.900 133.190 53.040 134.570 ;
        RECT 53.820 134.550 53.960 139.930 ;
        RECT 54.220 136.610 54.480 136.930 ;
        RECT 53.760 134.230 54.020 134.550 ;
        RECT 52.840 132.870 53.100 133.190 ;
        RECT 54.280 132.850 54.420 136.610 ;
        RECT 54.740 135.910 54.880 142.050 ;
        RECT 55.140 140.350 55.400 140.670 ;
        RECT 55.200 138.630 55.340 140.350 ;
        RECT 55.660 139.650 55.800 143.070 ;
        RECT 56.580 141.010 56.720 148.510 ;
        RECT 57.500 145.090 57.640 150.810 ;
        RECT 58.360 148.510 58.620 148.830 ;
        RECT 58.420 146.450 58.560 148.510 ;
        RECT 58.820 147.490 59.080 147.810 ;
        RECT 58.360 146.130 58.620 146.450 ;
        RECT 57.440 144.770 57.700 145.090 ;
        RECT 56.520 140.690 56.780 141.010 ;
        RECT 55.600 139.330 55.860 139.650 ;
        RECT 55.140 138.310 55.400 138.630 ;
        RECT 55.660 137.950 55.800 139.330 ;
        RECT 57.500 138.290 57.640 144.770 ;
        RECT 58.880 143.730 59.020 147.490 ;
        RECT 58.820 143.410 59.080 143.730 ;
        RECT 60.260 143.390 60.400 151.490 ;
        RECT 60.720 150.530 60.860 151.910 ;
        RECT 61.120 150.550 61.380 150.870 ;
        RECT 60.660 150.210 60.920 150.530 ;
        RECT 61.180 148.830 61.320 150.550 ;
        RECT 61.640 149.170 61.780 155.990 ;
        RECT 62.040 155.650 62.300 155.970 ;
        RECT 62.100 154.610 62.240 155.650 ;
        RECT 62.560 154.950 62.700 158.370 ;
        RECT 62.960 156.670 63.220 156.990 ;
        RECT 62.500 154.630 62.760 154.950 ;
        RECT 62.040 154.290 62.300 154.610 ;
        RECT 61.580 148.850 61.840 149.170 ;
        RECT 63.020 148.830 63.160 156.670 ;
        RECT 64.860 156.650 65.000 174.610 ;
        RECT 65.260 173.670 65.520 173.990 ;
        RECT 65.320 169.570 65.460 173.670 ;
        RECT 65.780 170.250 65.920 181.490 ;
        RECT 66.240 181.130 66.380 182.850 ;
        RECT 71.300 181.550 71.440 183.530 ;
        RECT 71.760 182.150 71.900 199.850 ;
        RECT 72.620 196.790 72.880 197.110 ;
        RECT 72.680 187.250 72.820 196.790 ;
        RECT 80.500 195.410 80.640 202.910 ;
        RECT 81.880 201.190 82.020 202.910 ;
        RECT 81.820 200.870 82.080 201.190 ;
        RECT 82.800 200.170 82.940 204.610 ;
        RECT 82.740 199.850 83.000 200.170 ;
        RECT 80.900 196.450 81.160 196.770 ;
        RECT 80.440 195.090 80.700 195.410 ;
        RECT 79.980 194.410 80.240 194.730 ;
        RECT 80.040 193.030 80.180 194.410 ;
        RECT 79.980 192.710 80.240 193.030 ;
        RECT 80.500 192.690 80.640 195.090 ;
        RECT 80.960 194.730 81.100 196.450 ;
        RECT 81.360 195.430 81.620 195.750 ;
        RECT 81.420 195.070 81.560 195.430 ;
        RECT 81.360 194.750 81.620 195.070 ;
        RECT 80.900 194.410 81.160 194.730 ;
        RECT 82.280 194.070 82.540 194.390 ;
        RECT 78.600 192.370 78.860 192.690 ;
        RECT 80.440 192.370 80.700 192.690 ;
        RECT 75.380 191.690 75.640 192.010 ;
        RECT 73.540 191.010 73.800 191.330 ;
        RECT 72.620 186.930 72.880 187.250 ;
        RECT 71.700 181.830 71.960 182.150 ;
        RECT 72.160 181.830 72.420 182.150 ;
        RECT 70.380 181.470 71.440 181.550 ;
        RECT 66.640 181.150 66.900 181.470 ;
        RECT 70.320 181.410 71.440 181.470 ;
        RECT 70.320 181.150 70.580 181.410 ;
        RECT 66.180 180.810 66.440 181.130 ;
        RECT 66.700 178.750 66.840 181.150 ;
        RECT 71.300 180.450 71.440 181.410 ;
        RECT 72.220 181.130 72.360 181.830 ;
        RECT 72.160 180.810 72.420 181.130 ;
        RECT 72.680 180.870 72.820 186.930 ;
        RECT 73.600 186.910 73.740 191.010 ;
        RECT 75.440 190.310 75.580 191.690 ;
        RECT 75.380 189.990 75.640 190.310 ;
        RECT 78.660 189.290 78.800 192.370 ;
        RECT 82.340 192.350 82.480 194.070 ;
        RECT 82.740 193.730 83.000 194.050 ;
        RECT 82.800 192.350 82.940 193.730 ;
        RECT 80.900 192.030 81.160 192.350 ;
        RECT 82.280 192.030 82.540 192.350 ;
        RECT 82.740 192.030 83.000 192.350 ;
        RECT 78.600 188.970 78.860 189.290 ;
        RECT 78.660 187.590 78.800 188.970 ;
        RECT 78.600 187.270 78.860 187.590 ;
        RECT 73.540 186.590 73.800 186.910 ;
        RECT 73.600 184.530 73.740 186.590 ;
        RECT 73.540 184.210 73.800 184.530 ;
        RECT 73.600 182.150 73.740 184.210 ;
        RECT 80.960 183.510 81.100 192.030 ;
        RECT 84.120 188.290 84.380 188.610 ;
        RECT 84.180 187.250 84.320 188.290 ;
        RECT 84.120 186.930 84.380 187.250 ;
        RECT 82.280 185.570 82.540 185.890 ;
        RECT 81.820 184.210 82.080 184.530 ;
        RECT 81.360 183.870 81.620 184.190 ;
        RECT 80.900 183.190 81.160 183.510 ;
        RECT 73.540 181.830 73.800 182.150 ;
        RECT 72.680 180.790 73.740 180.870 ;
        RECT 74.000 180.810 74.260 181.130 ;
        RECT 72.680 180.730 73.800 180.790 ;
        RECT 73.540 180.470 73.800 180.730 ;
        RECT 70.780 180.130 71.040 180.450 ;
        RECT 71.240 180.130 71.500 180.450 ;
        RECT 72.620 180.130 72.880 180.450 ;
        RECT 66.640 178.430 66.900 178.750 ;
        RECT 70.840 178.410 70.980 180.130 ;
        RECT 72.680 178.750 72.820 180.130 ;
        RECT 72.620 178.430 72.880 178.750 ;
        RECT 70.780 178.090 71.040 178.410 ;
        RECT 66.640 177.750 66.900 178.070 ;
        RECT 66.180 176.050 66.440 176.370 ;
        RECT 66.240 172.630 66.380 176.050 ;
        RECT 66.700 176.030 66.840 177.750 ;
        RECT 72.680 176.030 72.820 178.430 ;
        RECT 73.600 178.070 73.740 180.470 ;
        RECT 73.540 177.750 73.800 178.070 ;
        RECT 66.640 175.710 66.900 176.030 ;
        RECT 72.620 175.710 72.880 176.030 ;
        RECT 66.700 173.990 66.840 175.710 ;
        RECT 66.640 173.670 66.900 173.990 ;
        RECT 72.680 172.970 72.820 175.710 ;
        RECT 73.080 175.370 73.340 175.690 ;
        RECT 73.140 173.990 73.280 175.370 ;
        RECT 73.080 173.670 73.340 173.990 ;
        RECT 66.640 172.650 66.900 172.970 ;
        RECT 68.480 172.650 68.740 172.970 ;
        RECT 72.620 172.650 72.880 172.970 ;
        RECT 66.180 172.310 66.440 172.630 ;
        RECT 66.240 170.930 66.380 172.310 ;
        RECT 66.180 170.610 66.440 170.930 ;
        RECT 65.720 169.930 65.980 170.250 ;
        RECT 65.260 169.250 65.520 169.570 ;
        RECT 65.320 165.830 65.460 169.250 ;
        RECT 65.780 168.550 65.920 169.930 ;
        RECT 65.720 168.230 65.980 168.550 ;
        RECT 66.240 168.210 66.380 170.610 ;
        RECT 66.700 170.590 66.840 172.650 ;
        RECT 68.020 172.310 68.280 172.630 ;
        RECT 67.560 171.970 67.820 172.290 ;
        RECT 67.620 171.270 67.760 171.970 ;
        RECT 68.080 171.270 68.220 172.310 ;
        RECT 67.560 170.950 67.820 171.270 ;
        RECT 68.020 170.950 68.280 171.270 ;
        RECT 66.640 170.270 66.900 170.590 ;
        RECT 68.540 169.910 68.680 172.650 ;
        RECT 68.940 171.970 69.200 172.290 ;
        RECT 68.480 169.590 68.740 169.910 ;
        RECT 66.180 167.890 66.440 168.210 ;
        RECT 69.000 167.530 69.140 171.970 ;
        RECT 73.600 170.930 73.740 177.750 ;
        RECT 74.060 177.730 74.200 180.810 ;
        RECT 80.960 179.430 81.100 183.190 ;
        RECT 81.420 181.130 81.560 183.870 ;
        RECT 81.880 182.150 82.020 184.210 ;
        RECT 81.820 181.830 82.080 182.150 ;
        RECT 82.340 181.810 82.480 185.570 ;
        RECT 84.640 184.170 84.780 210.390 ;
        RECT 85.500 210.050 85.760 210.370 ;
        RECT 85.560 205.270 85.700 210.050 ;
        RECT 85.960 208.010 86.220 208.330 ;
        RECT 85.500 204.950 85.760 205.270 ;
        RECT 86.020 203.910 86.160 208.010 ;
        RECT 87.400 203.910 87.540 210.730 ;
        RECT 85.960 203.590 86.220 203.910 ;
        RECT 87.340 203.590 87.600 203.910 ;
        RECT 86.420 203.250 86.680 203.570 ;
        RECT 86.480 201.190 86.620 203.250 ;
        RECT 86.420 200.870 86.680 201.190 ;
        RECT 86.480 200.170 86.620 200.870 ;
        RECT 86.420 199.850 86.680 200.170 ;
        RECT 85.960 199.170 86.220 199.490 ;
        RECT 85.040 196.450 85.300 196.770 ;
        RECT 85.100 189.290 85.240 196.450 ;
        RECT 86.020 195.750 86.160 199.170 ;
        RECT 85.960 195.430 86.220 195.750 ;
        RECT 85.960 194.070 86.220 194.390 ;
        RECT 86.020 193.030 86.160 194.070 ;
        RECT 85.960 192.710 86.220 193.030 ;
        RECT 85.040 188.970 85.300 189.290 ;
        RECT 85.960 188.290 86.220 188.610 ;
        RECT 86.020 187.590 86.160 188.290 ;
        RECT 85.960 187.270 86.220 187.590 ;
        RECT 84.640 184.030 85.240 184.170 ;
        RECT 82.280 181.490 82.540 181.810 ;
        RECT 81.360 180.810 81.620 181.130 ;
        RECT 80.900 179.110 81.160 179.430 ;
        RECT 81.420 178.410 81.560 180.810 ;
        RECT 81.360 178.090 81.620 178.410 ;
        RECT 74.000 177.410 74.260 177.730 ;
        RECT 78.140 174.690 78.400 175.010 ;
        RECT 74.460 172.310 74.720 172.630 ;
        RECT 73.540 170.610 73.800 170.930 ;
        RECT 74.520 169.910 74.660 172.310 ;
        RECT 78.200 171.270 78.340 174.690 ;
        RECT 83.660 172.650 83.920 172.970 ;
        RECT 78.140 170.950 78.400 171.270 ;
        RECT 83.720 170.930 83.860 172.650 ;
        RECT 83.660 170.610 83.920 170.930 ;
        RECT 78.140 170.270 78.400 170.590 ;
        RECT 74.460 169.590 74.720 169.910 ;
        RECT 68.940 167.210 69.200 167.530 ;
        RECT 78.200 166.850 78.340 170.270 ;
        RECT 83.720 167.870 83.860 170.610 ;
        RECT 84.580 169.250 84.840 169.570 ;
        RECT 83.660 167.550 83.920 167.870 ;
        RECT 78.140 166.530 78.400 166.850 ;
        RECT 65.260 165.510 65.520 165.830 ;
        RECT 83.200 165.060 83.460 165.150 ;
        RECT 82.800 164.920 83.460 165.060 ;
        RECT 82.800 162.090 82.940 164.920 ;
        RECT 83.200 164.830 83.460 164.920 ;
        RECT 83.720 164.810 83.860 167.550 ;
        RECT 83.660 164.490 83.920 164.810 ;
        RECT 83.720 162.430 83.860 164.490 ;
        RECT 84.640 163.110 84.780 169.250 ;
        RECT 85.100 167.870 85.240 184.030 ;
        RECT 86.880 183.190 87.140 183.510 ;
        RECT 85.960 180.130 86.220 180.450 ;
        RECT 86.020 178.070 86.160 180.130 ;
        RECT 85.960 177.750 86.220 178.070 ;
        RECT 86.420 177.750 86.680 178.070 ;
        RECT 86.480 175.690 86.620 177.750 ;
        RECT 86.420 175.370 86.680 175.690 ;
        RECT 86.480 172.970 86.620 175.370 ;
        RECT 86.420 172.650 86.680 172.970 ;
        RECT 85.040 167.550 85.300 167.870 ;
        RECT 85.100 164.130 85.240 167.550 ;
        RECT 85.960 164.490 86.220 164.810 ;
        RECT 85.040 163.810 85.300 164.130 ;
        RECT 84.580 162.790 84.840 163.110 ;
        RECT 86.020 162.770 86.160 164.490 ;
        RECT 85.960 162.450 86.220 162.770 ;
        RECT 83.660 162.110 83.920 162.430 ;
        RECT 82.740 161.770 83.000 162.090 ;
        RECT 84.120 161.770 84.380 162.090 ;
        RECT 82.800 160.050 82.940 161.770 ;
        RECT 82.740 159.730 83.000 160.050 ;
        RECT 84.180 159.710 84.320 161.770 ;
        RECT 86.940 161.750 87.080 183.190 ;
        RECT 87.340 166.530 87.600 166.850 ;
        RECT 87.400 165.490 87.540 166.530 ;
        RECT 87.860 165.490 88.000 211.410 ;
        RECT 89.180 210.730 89.440 211.050 ;
        RECT 103.440 210.730 103.700 211.050 ;
        RECT 88.260 210.050 88.520 210.370 ;
        RECT 87.340 165.170 87.600 165.490 ;
        RECT 87.800 165.170 88.060 165.490 ;
        RECT 87.860 162.770 88.000 165.170 ;
        RECT 88.320 165.150 88.460 210.050 ;
        RECT 89.240 209.350 89.380 210.730 ;
        RECT 89.640 210.390 89.900 210.710 ;
        RECT 89.700 209.350 89.840 210.390 ;
        RECT 91.020 210.050 91.280 210.370 ;
        RECT 89.180 209.030 89.440 209.350 ;
        RECT 89.640 209.030 89.900 209.350 ;
        RECT 90.560 208.690 90.820 209.010 ;
        RECT 89.640 206.310 89.900 206.630 ;
        RECT 89.700 203.230 89.840 206.310 ;
        RECT 90.620 203.230 90.760 208.690 ;
        RECT 91.080 203.230 91.220 210.050 ;
        RECT 93.320 209.030 93.580 209.350 ;
        RECT 93.380 208.670 93.520 209.030 ;
        RECT 103.500 209.010 103.640 210.730 ;
        RECT 95.620 208.690 95.880 209.010 ;
        RECT 97.460 208.690 97.720 209.010 ;
        RECT 103.440 208.690 103.700 209.010 ;
        RECT 93.320 208.350 93.580 208.670 ;
        RECT 93.380 207.650 93.520 208.350 ;
        RECT 93.320 207.330 93.580 207.650 ;
        RECT 91.940 204.950 92.200 205.270 ;
        RECT 92.000 203.910 92.140 204.950 ;
        RECT 91.940 203.590 92.200 203.910 ;
        RECT 89.640 202.910 89.900 203.230 ;
        RECT 90.560 202.910 90.820 203.230 ;
        RECT 91.020 202.910 91.280 203.230 ;
        RECT 92.400 202.910 92.660 203.230 ;
        RECT 89.180 201.890 89.440 202.210 ;
        RECT 89.240 200.170 89.380 201.890 ;
        RECT 89.180 199.850 89.440 200.170 ;
        RECT 89.240 197.790 89.380 199.850 ;
        RECT 89.700 198.130 89.840 202.910 ;
        RECT 90.620 202.210 90.760 202.910 ;
        RECT 90.560 201.890 90.820 202.210 ;
        RECT 90.620 200.170 90.760 201.890 ;
        RECT 91.080 201.190 91.220 202.910 ;
        RECT 91.020 200.870 91.280 201.190 ;
        RECT 92.460 200.850 92.600 202.910 ;
        RECT 95.680 202.890 95.820 208.690 ;
        RECT 96.540 208.350 96.800 208.670 ;
        RECT 96.600 207.990 96.740 208.350 ;
        RECT 96.540 207.900 96.800 207.990 ;
        RECT 96.540 207.760 97.200 207.900 ;
        RECT 96.540 207.670 96.800 207.760 ;
        RECT 96.540 205.290 96.800 205.610 ;
        RECT 96.600 203.570 96.740 205.290 ;
        RECT 97.060 204.930 97.200 207.760 ;
        RECT 97.520 206.630 97.660 208.690 ;
        RECT 98.840 208.010 99.100 208.330 ;
        RECT 97.460 206.310 97.720 206.630 ;
        RECT 97.000 204.610 97.260 204.930 ;
        RECT 96.540 203.250 96.800 203.570 ;
        RECT 95.620 202.570 95.880 202.890 ;
        RECT 93.320 202.460 93.580 202.550 ;
        RECT 92.920 202.320 93.580 202.460 ;
        RECT 92.400 200.530 92.660 200.850 ;
        RECT 92.920 200.170 93.060 202.320 ;
        RECT 93.320 202.230 93.580 202.320 ;
        RECT 90.560 199.850 90.820 200.170 ;
        RECT 92.860 199.850 93.120 200.170 ;
        RECT 95.620 199.170 95.880 199.490 ;
        RECT 89.640 197.810 89.900 198.130 ;
        RECT 89.180 197.470 89.440 197.790 ;
        RECT 89.700 192.690 89.840 197.810 ;
        RECT 94.240 197.470 94.500 197.790 ;
        RECT 91.480 196.450 91.740 196.770 ;
        RECT 91.540 194.730 91.680 196.450 ;
        RECT 91.480 194.410 91.740 194.730 ;
        RECT 89.640 192.370 89.900 192.690 ;
        RECT 89.180 189.200 89.440 189.290 ;
        RECT 89.700 189.200 89.840 192.370 ;
        RECT 91.540 190.310 91.680 194.410 ;
        RECT 94.300 194.050 94.440 197.470 ;
        RECT 94.700 196.450 94.960 196.770 ;
        RECT 94.240 193.730 94.500 194.050 ;
        RECT 94.300 193.030 94.440 193.730 ;
        RECT 94.240 192.710 94.500 193.030 ;
        RECT 94.760 192.350 94.900 196.450 ;
        RECT 95.680 195.750 95.820 199.170 ;
        RECT 96.080 197.470 96.340 197.790 ;
        RECT 96.140 195.750 96.280 197.470 ;
        RECT 95.620 195.430 95.880 195.750 ;
        RECT 96.080 195.430 96.340 195.750 ;
        RECT 95.680 193.030 95.820 195.430 ;
        RECT 96.600 195.070 96.740 203.250 ;
        RECT 97.060 202.210 97.200 204.610 ;
        RECT 98.900 203.230 99.040 208.010 ;
        RECT 103.500 206.630 103.640 208.690 ;
        RECT 106.660 207.670 106.920 207.990 ;
        RECT 104.360 207.330 104.620 207.650 ;
        RECT 103.440 206.310 103.700 206.630 ;
        RECT 100.680 204.950 100.940 205.270 ;
        RECT 103.440 204.950 103.700 205.270 ;
        RECT 97.460 202.910 97.720 203.230 ;
        RECT 98.840 202.910 99.100 203.230 ;
        RECT 97.000 201.890 97.260 202.210 ;
        RECT 96.540 194.750 96.800 195.070 ;
        RECT 95.620 192.710 95.880 193.030 ;
        RECT 95.680 192.430 95.820 192.710 ;
        RECT 92.400 192.030 92.660 192.350 ;
        RECT 94.700 192.030 94.960 192.350 ;
        RECT 95.680 192.290 96.280 192.430 ;
        RECT 92.460 190.310 92.600 192.030 ;
        RECT 94.760 191.750 94.900 192.030 ;
        RECT 94.300 191.610 94.900 191.750 ;
        RECT 91.480 189.990 91.740 190.310 ;
        RECT 92.400 189.990 92.660 190.310 ;
        RECT 90.550 189.455 90.830 189.825 ;
        RECT 90.620 189.290 90.760 189.455 ;
        RECT 94.300 189.290 94.440 191.610 ;
        RECT 94.700 191.010 94.960 191.330 ;
        RECT 94.760 189.970 94.900 191.010 ;
        RECT 94.700 189.650 94.960 189.970 ;
        RECT 96.140 189.630 96.280 192.290 ;
        RECT 96.080 189.310 96.340 189.630 ;
        RECT 89.180 189.060 89.840 189.200 ;
        RECT 89.180 188.970 89.440 189.060 ;
        RECT 90.560 188.970 90.820 189.290 ;
        RECT 94.240 188.970 94.500 189.290 ;
        RECT 95.620 188.970 95.880 189.290 ;
        RECT 90.620 187.590 90.760 188.970 ;
        RECT 94.300 188.610 94.440 188.970 ;
        RECT 94.240 188.290 94.500 188.610 ;
        RECT 94.700 188.290 94.960 188.610 ;
        RECT 90.560 187.270 90.820 187.590 ;
        RECT 94.240 183.530 94.500 183.850 ;
        RECT 91.020 182.850 91.280 183.170 ;
        RECT 91.080 182.150 91.220 182.850 ;
        RECT 91.020 181.830 91.280 182.150 ;
        RECT 94.300 181.550 94.440 183.530 ;
        RECT 94.760 182.150 94.900 188.290 ;
        RECT 95.680 183.850 95.820 188.970 ;
        RECT 96.070 188.775 96.350 189.145 ;
        RECT 96.140 188.610 96.280 188.775 ;
        RECT 96.080 188.290 96.340 188.610 ;
        RECT 96.600 184.870 96.740 194.750 ;
        RECT 97.000 192.545 97.260 192.690 ;
        RECT 96.990 192.175 97.270 192.545 ;
        RECT 96.540 184.550 96.800 184.870 ;
        RECT 95.620 183.530 95.880 183.850 ;
        RECT 94.700 181.830 94.960 182.150 ;
        RECT 94.300 181.410 94.900 181.550 ;
        RECT 94.760 179.090 94.900 181.410 ;
        RECT 96.540 181.150 96.800 181.470 ;
        RECT 97.000 181.150 97.260 181.470 ;
        RECT 94.700 178.770 94.960 179.090 ;
        RECT 94.700 175.710 94.960 176.030 ;
        RECT 94.760 171.270 94.900 175.710 ;
        RECT 95.160 175.370 95.420 175.690 ;
        RECT 94.700 170.950 94.960 171.270 ;
        RECT 95.220 168.550 95.360 175.370 ;
        RECT 96.080 174.690 96.340 175.010 ;
        RECT 96.140 173.310 96.280 174.690 ;
        RECT 96.080 172.990 96.340 173.310 ;
        RECT 95.620 171.970 95.880 172.290 ;
        RECT 96.080 171.970 96.340 172.290 ;
        RECT 95.160 168.230 95.420 168.550 ;
        RECT 91.020 165.170 91.280 165.490 ;
        RECT 88.260 164.830 88.520 165.150 ;
        RECT 87.800 162.510 88.060 162.770 ;
        RECT 87.400 162.450 88.060 162.510 ;
        RECT 87.400 162.370 88.000 162.450 ;
        RECT 87.400 162.090 87.540 162.370 ;
        RECT 88.320 162.090 88.460 164.830 ;
        RECT 88.720 164.150 88.980 164.470 ;
        RECT 88.780 163.110 88.920 164.150 ;
        RECT 88.720 162.790 88.980 163.110 ;
        RECT 89.640 162.450 89.900 162.770 ;
        RECT 89.700 162.090 89.840 162.450 ;
        RECT 87.340 161.770 87.600 162.090 ;
        RECT 88.260 162.000 88.520 162.090 ;
        RECT 87.860 161.860 88.520 162.000 ;
        RECT 86.880 161.430 87.140 161.750 ;
        RECT 84.120 159.390 84.380 159.710 ;
        RECT 67.100 159.050 67.360 159.370 ;
        RECT 79.520 159.050 79.780 159.370 ;
        RECT 63.420 156.330 63.680 156.650 ;
        RECT 64.800 156.330 65.060 156.650 ;
        RECT 63.480 152.230 63.620 156.330 ;
        RECT 64.860 155.970 65.000 156.330 ;
        RECT 67.160 156.310 67.300 159.050 ;
        RECT 79.580 157.670 79.720 159.050 ;
        RECT 82.740 158.370 83.000 158.690 ;
        RECT 82.800 157.670 82.940 158.370 ;
        RECT 79.520 157.350 79.780 157.670 ;
        RECT 82.740 157.580 83.000 157.670 ;
        RECT 82.340 157.440 83.000 157.580 ;
        RECT 71.700 156.670 71.960 156.990 ;
        RECT 67.560 156.330 67.820 156.650 ;
        RECT 67.100 155.990 67.360 156.310 ;
        RECT 64.800 155.650 65.060 155.970 ;
        RECT 63.420 151.910 63.680 152.230 ;
        RECT 64.860 151.210 65.000 155.650 ;
        RECT 67.160 153.250 67.300 155.990 ;
        RECT 67.620 153.590 67.760 156.330 ;
        RECT 69.400 155.990 69.660 156.310 ;
        RECT 68.940 153.610 69.200 153.930 ;
        RECT 67.560 153.270 67.820 153.590 ;
        RECT 67.100 152.930 67.360 153.250 ;
        RECT 65.260 151.910 65.520 152.230 ;
        RECT 64.340 150.890 64.600 151.210 ;
        RECT 64.800 150.890 65.060 151.210 ;
        RECT 64.400 149.170 64.540 150.890 ;
        RECT 64.340 148.850 64.600 149.170 ;
        RECT 60.660 148.510 60.920 148.830 ;
        RECT 61.120 148.510 61.380 148.830 ;
        RECT 62.960 148.510 63.220 148.830 ;
        RECT 60.720 148.150 60.860 148.510 ;
        RECT 64.860 148.490 65.000 150.890 ;
        RECT 65.320 149.170 65.460 151.910 ;
        RECT 66.640 150.550 66.900 150.870 ;
        RECT 66.700 149.170 66.840 150.550 ;
        RECT 65.260 148.850 65.520 149.170 ;
        RECT 66.640 148.850 66.900 149.170 ;
        RECT 64.800 148.170 65.060 148.490 ;
        RECT 60.660 147.830 60.920 148.150 ;
        RECT 66.700 146.450 66.840 148.850 ;
        RECT 67.620 148.150 67.760 153.270 ;
        RECT 68.020 152.930 68.280 153.250 ;
        RECT 68.080 151.210 68.220 152.930 ;
        RECT 68.020 150.890 68.280 151.210 ;
        RECT 68.480 150.890 68.740 151.210 ;
        RECT 67.560 147.830 67.820 148.150 ;
        RECT 66.640 146.130 66.900 146.450 ;
        RECT 60.660 145.790 60.920 146.110 ;
        RECT 60.720 143.730 60.860 145.790 ;
        RECT 64.800 145.110 65.060 145.430 ;
        RECT 62.500 144.770 62.760 145.090 ;
        RECT 61.120 143.750 61.380 144.070 ;
        RECT 60.660 143.410 60.920 143.730 ;
        RECT 60.200 143.070 60.460 143.390 ;
        RECT 58.360 142.050 58.620 142.370 ;
        RECT 58.420 141.350 58.560 142.050 ;
        RECT 58.360 141.030 58.620 141.350 ;
        RECT 60.260 140.670 60.400 143.070 ;
        RECT 60.200 140.350 60.460 140.670 ;
        RECT 61.180 138.290 61.320 143.750 ;
        RECT 62.560 143.730 62.700 144.770 ;
        RECT 62.500 143.410 62.760 143.730 ;
        RECT 64.860 141.350 65.000 145.110 ;
        RECT 68.540 145.090 68.680 150.890 ;
        RECT 68.480 144.770 68.740 145.090 ;
        RECT 68.540 144.070 68.680 144.770 ;
        RECT 68.480 143.750 68.740 144.070 ;
        RECT 64.800 141.030 65.060 141.350 ;
        RECT 66.180 140.690 66.440 141.010 ;
        RECT 62.500 140.350 62.760 140.670 ;
        RECT 57.440 137.970 57.700 138.290 ;
        RECT 61.120 137.970 61.380 138.290 ;
        RECT 62.560 137.950 62.700 140.350 ;
        RECT 62.960 140.010 63.220 140.330 ;
        RECT 63.020 138.290 63.160 140.010 ;
        RECT 64.800 139.330 65.060 139.650 ;
        RECT 64.860 138.290 65.000 139.330 ;
        RECT 66.240 138.630 66.380 140.690 ;
        RECT 69.000 140.670 69.140 153.610 ;
        RECT 69.460 147.810 69.600 155.990 ;
        RECT 70.780 153.950 71.040 154.270 ;
        RECT 70.840 152.230 70.980 153.950 ;
        RECT 71.760 153.930 71.900 156.670 ;
        RECT 73.080 155.990 73.340 156.310 ;
        RECT 74.000 155.990 74.260 156.310 ;
        RECT 74.920 155.990 75.180 156.310 ;
        RECT 80.440 155.990 80.700 156.310 ;
        RECT 73.140 154.950 73.280 155.990 ;
        RECT 73.080 154.630 73.340 154.950 ;
        RECT 71.700 153.610 71.960 153.930 ;
        RECT 73.540 153.610 73.800 153.930 ;
        RECT 71.700 152.930 71.960 153.250 ;
        RECT 70.780 151.910 71.040 152.230 ;
        RECT 70.320 151.230 70.580 151.550 ;
        RECT 70.380 148.830 70.520 151.230 ;
        RECT 71.760 149.170 71.900 152.930 ;
        RECT 73.600 151.550 73.740 153.610 ;
        RECT 73.540 151.230 73.800 151.550 ;
        RECT 74.060 151.210 74.200 155.990 ;
        RECT 74.980 153.590 75.120 155.990 ;
        RECT 79.060 155.650 79.320 155.970 ;
        RECT 79.120 154.610 79.260 155.650 ;
        RECT 79.060 154.290 79.320 154.610 ;
        RECT 74.920 153.270 75.180 153.590 ;
        RECT 74.000 150.890 74.260 151.210 ;
        RECT 74.060 149.590 74.200 150.890 ;
        RECT 74.060 149.510 74.660 149.590 ;
        RECT 74.060 149.450 74.720 149.510 ;
        RECT 74.460 149.190 74.720 149.450 ;
        RECT 71.700 148.850 71.960 149.170 ;
        RECT 70.320 148.510 70.580 148.830 ;
        RECT 69.400 147.490 69.660 147.810 ;
        RECT 68.940 140.350 69.200 140.670 ;
        RECT 66.640 139.670 66.900 139.990 ;
        RECT 66.180 138.310 66.440 138.630 ;
        RECT 62.960 138.030 63.220 138.290 ;
        RECT 62.960 137.970 63.620 138.030 ;
        RECT 64.800 137.970 65.060 138.290 ;
        RECT 55.600 137.630 55.860 137.950 ;
        RECT 62.500 137.630 62.760 137.950 ;
        RECT 63.020 137.890 63.620 137.970 ;
        RECT 54.680 135.590 54.940 135.910 ;
        RECT 62.560 134.890 62.700 137.630 ;
        RECT 62.960 136.610 63.220 136.930 ;
        RECT 63.020 135.910 63.160 136.610 ;
        RECT 63.480 135.910 63.620 137.890 ;
        RECT 62.960 135.590 63.220 135.910 ;
        RECT 63.420 135.590 63.680 135.910 ;
        RECT 62.500 134.570 62.760 134.890 ;
        RECT 54.220 132.530 54.480 132.850 ;
        RECT 66.700 132.510 66.840 139.670 ;
        RECT 69.000 137.950 69.140 140.350 ;
        RECT 70.380 140.330 70.520 148.510 ;
        RECT 74.000 145.450 74.260 145.770 ;
        RECT 74.060 143.390 74.200 145.450 ;
        RECT 74.980 145.090 75.120 153.270 ;
        RECT 75.840 152.930 76.100 153.250 ;
        RECT 75.900 151.210 76.040 152.930 ;
        RECT 75.840 150.890 76.100 151.210 ;
        RECT 79.120 150.870 79.260 154.290 ;
        RECT 80.500 153.840 80.640 155.990 ;
        RECT 80.900 153.840 81.160 153.930 ;
        RECT 80.500 153.700 81.160 153.840 ;
        RECT 80.900 153.610 81.160 153.700 ;
        RECT 82.340 151.210 82.480 157.440 ;
        RECT 82.740 157.350 83.000 157.440 ;
        RECT 82.740 155.990 83.000 156.310 ;
        RECT 82.800 154.950 82.940 155.990 ;
        RECT 82.740 154.630 83.000 154.950 ;
        RECT 85.500 153.950 85.760 154.270 ;
        RECT 83.200 152.930 83.460 153.250 ;
        RECT 83.260 151.210 83.400 152.930 ;
        RECT 85.560 152.230 85.700 153.950 ;
        RECT 86.420 153.610 86.680 153.930 ;
        RECT 85.500 151.910 85.760 152.230 ;
        RECT 86.480 151.210 86.620 153.610 ;
        RECT 82.280 150.890 82.540 151.210 ;
        RECT 83.200 150.890 83.460 151.210 ;
        RECT 86.420 150.890 86.680 151.210 ;
        RECT 79.060 150.550 79.320 150.870 ;
        RECT 78.600 150.210 78.860 150.530 ;
        RECT 74.920 144.770 75.180 145.090 ;
        RECT 76.300 144.770 76.560 145.090 ;
        RECT 74.000 143.070 74.260 143.390 ;
        RECT 75.380 142.730 75.640 143.050 ;
        RECT 73.540 142.050 73.800 142.370 ;
        RECT 70.320 140.010 70.580 140.330 ;
        RECT 68.940 137.630 69.200 137.950 ;
        RECT 44.560 132.190 44.820 132.510 ;
        RECT 66.640 132.190 66.900 132.510 ;
        RECT 41.800 131.850 42.060 132.170 ;
        RECT 31.220 131.170 31.480 131.490 ;
        RECT 22.940 130.150 23.200 130.470 ;
        RECT 28.000 130.150 28.260 130.470 ;
        RECT 31.280 129.790 31.420 131.170 ;
        RECT 32.870 130.635 34.410 131.005 ;
        RECT 31.680 130.150 31.940 130.470 ;
        RECT 31.740 129.870 31.880 130.150 ;
        RECT 31.220 129.470 31.480 129.790 ;
        RECT 31.740 129.730 32.340 129.870 ;
        RECT 32.600 129.810 32.860 130.130 ;
        RECT 20.640 129.130 20.900 129.450 ;
        RECT 24.780 129.130 25.040 129.450 ;
        RECT 30.300 129.130 30.560 129.450 ;
        RECT 24.320 128.790 24.580 129.110 ;
        RECT 21.100 126.410 21.360 126.730 ;
        RECT 19.320 124.290 19.920 124.430 ;
        RECT 19.780 124.010 19.920 124.290 ;
        RECT 19.720 123.750 19.980 124.010 ;
        RECT 21.160 123.750 21.300 126.410 ;
        RECT 19.720 123.690 21.300 123.750 ;
        RECT 19.780 123.610 21.300 123.690 ;
        RECT 16.030 120.775 16.310 121.145 ;
        RECT 16.040 120.630 16.300 120.775 ;
        RECT 16.040 119.105 16.300 119.250 ;
        RECT 16.030 118.735 16.310 119.105 ;
        RECT 20.240 116.190 20.380 123.610 ;
        RECT 22.020 123.350 22.280 123.670 ;
        RECT 22.080 122.310 22.220 123.350 ;
        RECT 22.020 121.990 22.280 122.310 ;
        RECT 24.380 121.630 24.520 128.790 ;
        RECT 24.840 126.730 24.980 129.130 ;
        RECT 30.360 127.750 30.500 129.130 ;
        RECT 31.220 128.790 31.480 129.110 ;
        RECT 30.300 127.430 30.560 127.750 ;
        RECT 26.160 126.750 26.420 127.070 ;
        RECT 24.780 126.410 25.040 126.730 ;
        RECT 26.220 125.030 26.360 126.750 ;
        RECT 26.160 124.710 26.420 125.030 ;
        RECT 30.360 123.330 30.500 127.430 ;
        RECT 31.280 124.690 31.420 128.790 ;
        RECT 32.200 127.070 32.340 129.730 ;
        RECT 32.660 127.750 32.800 129.810 ;
        RECT 66.700 129.110 66.840 132.190 ;
        RECT 66.640 128.790 66.900 129.110 ;
        RECT 36.170 127.915 37.710 128.285 ;
        RECT 32.600 127.430 32.860 127.750 ;
        RECT 32.140 126.750 32.400 127.070 ;
        RECT 65.260 126.750 65.520 127.070 ;
        RECT 31.680 125.730 31.940 126.050 ;
        RECT 31.220 124.370 31.480 124.690 ;
        RECT 26.160 123.010 26.420 123.330 ;
        RECT 30.300 123.010 30.560 123.330 ;
        RECT 26.220 121.970 26.360 123.010 ;
        RECT 26.160 121.650 26.420 121.970 ;
        RECT 24.320 121.310 24.580 121.630 ;
        RECT 22.020 118.250 22.280 118.570 ;
        RECT 21.100 117.570 21.360 117.890 ;
        RECT 20.180 115.870 20.440 116.190 ;
        RECT 19.260 114.850 19.520 115.170 ;
        RECT 19.320 113.470 19.460 114.850 ;
        RECT 19.260 113.150 19.520 113.470 ;
        RECT 20.240 111.430 20.380 115.870 ;
        RECT 21.160 115.025 21.300 117.570 ;
        RECT 21.090 114.655 21.370 115.025 ;
        RECT 21.560 112.470 21.820 112.790 ;
        RECT 21.620 111.430 21.760 112.470 ;
        RECT 22.080 112.450 22.220 118.250 ;
        RECT 22.020 112.130 22.280 112.450 ;
        RECT 22.080 111.430 22.220 112.130 ;
        RECT 24.380 111.430 24.520 121.310 ;
        RECT 25.700 118.250 25.960 118.570 ;
        RECT 25.760 116.870 25.900 118.250 ;
        RECT 26.620 117.910 26.880 118.230 ;
        RECT 25.700 116.550 25.960 116.870 ;
        RECT 26.160 115.870 26.420 116.190 ;
        RECT 26.220 115.170 26.360 115.870 ;
        RECT 26.160 114.850 26.420 115.170 ;
        RECT 26.220 113.130 26.360 114.850 ;
        RECT 26.160 112.810 26.420 113.130 ;
        RECT 20.180 111.110 20.440 111.430 ;
        RECT 21.560 111.110 21.820 111.430 ;
        RECT 22.020 111.110 22.280 111.430 ;
        RECT 24.320 111.110 24.580 111.430 ;
        RECT 16.030 110.575 16.310 110.945 ;
        RECT 16.040 110.430 16.300 110.575 ;
        RECT 20.180 110.430 20.440 110.750 ;
        RECT 20.240 108.225 20.380 110.430 ;
        RECT 24.380 108.270 24.520 111.110 ;
        RECT 26.220 110.410 26.360 112.810 ;
        RECT 26.680 110.750 26.820 117.910 ;
        RECT 31.280 115.850 31.420 124.370 ;
        RECT 31.740 124.010 31.880 125.730 ;
        RECT 31.680 123.690 31.940 124.010 ;
        RECT 31.680 117.570 31.940 117.890 ;
        RECT 31.740 116.190 31.880 117.570 ;
        RECT 31.680 115.870 31.940 116.190 ;
        RECT 31.220 115.530 31.480 115.850 ;
        RECT 29.840 114.850 30.100 115.170 ;
        RECT 28.920 113.830 29.180 114.150 ;
        RECT 27.540 112.130 27.800 112.450 ;
        RECT 26.620 110.430 26.880 110.750 ;
        RECT 26.160 110.090 26.420 110.410 ;
        RECT 20.170 107.855 20.450 108.225 ;
        RECT 24.380 108.130 24.980 108.270 ;
        RECT 24.320 104.990 24.580 105.310 ;
        RECT 23.860 104.650 24.120 104.970 ;
        RECT 16.040 104.145 16.300 104.290 ;
        RECT 16.030 103.775 16.310 104.145 ;
        RECT 20.180 102.950 20.440 103.270 ;
        RECT 18.330 101.055 18.610 101.425 ;
        RECT 18.400 100.550 18.540 101.055 ;
        RECT 18.340 100.230 18.600 100.550 ;
        RECT 20.240 99.870 20.380 102.950 ;
        RECT 20.180 99.550 20.440 99.870 ;
        RECT 22.020 99.550 22.280 99.870 ;
        RECT 18.330 97.655 18.610 98.025 ;
        RECT 16.950 94.255 17.230 94.625 ;
        RECT 17.020 93.750 17.160 94.255 ;
        RECT 16.960 93.430 17.220 93.750 ;
        RECT 18.400 93.410 18.540 97.655 ;
        RECT 19.260 95.810 19.520 96.130 ;
        RECT 19.320 94.430 19.460 95.810 ;
        RECT 22.080 94.430 22.220 99.550 ;
        RECT 23.920 94.430 24.060 104.650 ;
        RECT 24.380 103.270 24.520 104.990 ;
        RECT 24.320 102.950 24.580 103.270 ;
        RECT 24.840 97.830 24.980 108.130 ;
        RECT 26.220 104.880 26.360 110.090 ;
        RECT 27.600 105.650 27.740 112.130 ;
        RECT 28.000 109.410 28.260 109.730 ;
        RECT 27.540 105.330 27.800 105.650 ;
        RECT 27.080 104.880 27.340 104.970 ;
        RECT 26.220 104.740 27.340 104.880 ;
        RECT 27.080 104.650 27.340 104.740 ;
        RECT 25.700 103.970 25.960 104.290 ;
        RECT 25.760 102.250 25.900 103.970 ;
        RECT 27.140 102.250 27.280 104.650 ;
        RECT 27.600 102.590 27.740 105.330 ;
        RECT 27.540 102.270 27.800 102.590 ;
        RECT 25.700 101.930 25.960 102.250 ;
        RECT 27.080 101.930 27.340 102.250 ;
        RECT 27.140 98.850 27.280 101.930 ;
        RECT 27.080 98.530 27.340 98.850 ;
        RECT 24.780 97.510 25.040 97.830 ;
        RECT 27.140 96.810 27.280 98.530 ;
        RECT 28.060 96.810 28.200 109.410 ;
        RECT 28.980 107.690 29.120 113.830 ;
        RECT 29.900 112.790 30.040 114.850 ;
        RECT 29.840 112.470 30.100 112.790 ;
        RECT 29.380 110.430 29.640 110.750 ;
        RECT 28.920 107.370 29.180 107.690 ;
        RECT 28.920 106.920 29.180 107.010 ;
        RECT 29.440 106.920 29.580 110.430 ;
        RECT 29.900 109.730 30.040 112.470 ;
        RECT 30.300 110.430 30.560 110.750 ;
        RECT 29.840 109.410 30.100 109.730 ;
        RECT 29.900 107.690 30.040 109.410 ;
        RECT 29.840 107.370 30.100 107.690 ;
        RECT 28.920 106.780 29.580 106.920 ;
        RECT 28.920 106.690 29.180 106.780 ;
        RECT 28.980 99.530 29.120 106.690 ;
        RECT 30.360 106.070 30.500 110.430 ;
        RECT 29.440 105.930 30.500 106.070 ;
        RECT 28.920 99.270 29.180 99.530 ;
        RECT 28.520 99.210 29.180 99.270 ;
        RECT 28.520 99.130 29.120 99.210 ;
        RECT 27.080 96.490 27.340 96.810 ;
        RECT 28.000 96.490 28.260 96.810 ;
        RECT 25.700 96.150 25.960 96.470 ;
        RECT 25.760 95.110 25.900 96.150 ;
        RECT 25.700 94.790 25.960 95.110 ;
        RECT 19.260 94.110 19.520 94.430 ;
        RECT 22.020 94.110 22.280 94.430 ;
        RECT 23.860 94.110 24.120 94.430 ;
        RECT 25.700 94.110 25.960 94.430 ;
        RECT 18.340 93.090 18.600 93.410 ;
        RECT 25.760 89.670 25.900 94.110 ;
        RECT 26.160 93.090 26.420 93.410 ;
        RECT 25.700 89.350 25.960 89.670 ;
        RECT 15.120 85.950 15.380 86.270 ;
        RECT 11.900 85.270 12.160 85.590 ;
        RECT 11.960 77.700 12.100 85.270 ;
        RECT 15.180 77.700 15.320 85.950 ;
        RECT 18.340 85.610 18.600 85.930 ;
        RECT 24.780 85.610 25.040 85.930 ;
        RECT 18.400 77.700 18.540 85.610 ;
        RECT 21.560 84.930 21.820 85.250 ;
        RECT 21.620 77.700 21.760 84.930 ;
        RECT 24.840 77.700 24.980 85.610 ;
        RECT 25.760 85.590 25.900 89.350 ;
        RECT 26.220 89.330 26.360 93.090 ;
        RECT 27.140 91.370 27.280 96.490 ;
        RECT 28.520 93.750 28.660 99.130 ;
        RECT 28.920 94.450 29.180 94.770 ;
        RECT 28.460 93.430 28.720 93.750 ;
        RECT 27.540 93.090 27.800 93.410 ;
        RECT 27.600 91.370 27.740 93.090 ;
        RECT 27.080 91.050 27.340 91.370 ;
        RECT 27.540 91.050 27.800 91.370 ;
        RECT 26.620 90.710 26.880 91.030 ;
        RECT 26.680 89.670 26.820 90.710 ;
        RECT 26.620 89.350 26.880 89.670 ;
        RECT 26.160 89.010 26.420 89.330 ;
        RECT 27.140 88.650 27.280 91.050 ;
        RECT 27.600 89.330 27.740 91.050 ;
        RECT 28.460 90.370 28.720 90.690 ;
        RECT 28.520 89.670 28.660 90.370 ;
        RECT 28.460 89.350 28.720 89.670 ;
        RECT 27.540 89.010 27.800 89.330 ;
        RECT 27.080 88.330 27.340 88.650 ;
        RECT 27.600 85.590 27.740 89.010 ;
        RECT 28.520 85.930 28.660 89.350 ;
        RECT 28.980 86.950 29.120 94.450 ;
        RECT 29.440 94.090 29.580 105.930 ;
        RECT 30.760 104.990 31.020 105.310 ;
        RECT 30.820 103.270 30.960 104.990 ;
        RECT 30.760 102.950 31.020 103.270 ;
        RECT 30.760 101.250 31.020 101.570 ;
        RECT 30.820 100.550 30.960 101.250 ;
        RECT 30.760 100.230 31.020 100.550 ;
        RECT 29.840 96.490 30.100 96.810 ;
        RECT 29.380 93.770 29.640 94.090 ;
        RECT 29.440 88.650 29.580 93.770 ;
        RECT 29.380 88.330 29.640 88.650 ;
        RECT 29.900 86.950 30.040 96.490 ;
        RECT 30.820 89.670 30.960 100.230 ;
        RECT 31.280 97.830 31.420 115.530 ;
        RECT 32.200 112.790 32.340 126.750 ;
        RECT 32.870 125.195 34.410 125.565 ;
        RECT 65.320 125.030 65.460 126.750 ;
        RECT 66.180 125.730 66.440 126.050 ;
        RECT 65.260 124.710 65.520 125.030 ;
        RECT 62.040 123.690 62.300 124.010 ;
        RECT 32.600 123.350 32.860 123.670 ;
        RECT 35.820 123.350 36.080 123.670 ;
        RECT 32.660 121.290 32.800 123.350 ;
        RECT 34.900 123.010 35.160 123.330 ;
        RECT 32.600 120.970 32.860 121.290 ;
        RECT 32.870 119.755 34.410 120.125 ;
        RECT 34.960 115.850 35.100 123.010 ;
        RECT 35.360 115.870 35.620 116.190 ;
        RECT 34.900 115.530 35.160 115.850 ;
        RECT 32.870 114.315 34.410 114.685 ;
        RECT 34.960 112.870 35.100 115.530 ;
        RECT 35.420 114.150 35.560 115.870 ;
        RECT 35.360 113.830 35.620 114.150 ;
        RECT 32.140 112.470 32.400 112.790 ;
        RECT 34.500 112.730 35.100 112.870 ;
        RECT 34.500 110.410 34.640 112.730 ;
        RECT 34.900 112.130 35.160 112.450 ;
        RECT 34.440 110.090 34.700 110.410 ;
        RECT 34.960 110.070 35.100 112.130 ;
        RECT 35.420 111.090 35.560 113.830 ;
        RECT 35.880 111.430 36.020 123.350 ;
        RECT 36.170 122.475 37.710 122.845 ;
        RECT 62.100 121.630 62.240 123.690 ;
        RECT 64.800 123.350 65.060 123.670 ;
        RECT 62.040 121.310 62.300 121.630 ;
        RECT 64.860 119.590 65.000 123.350 ;
        RECT 64.800 119.270 65.060 119.590 ;
        RECT 66.240 118.910 66.380 125.730 ;
        RECT 66.700 121.970 66.840 128.790 ;
        RECT 67.100 126.750 67.360 127.070 ;
        RECT 68.480 126.750 68.740 127.070 ;
        RECT 67.160 126.050 67.300 126.750 ;
        RECT 67.100 125.730 67.360 126.050 ;
        RECT 67.160 124.010 67.300 125.730 ;
        RECT 68.540 125.030 68.680 126.750 ;
        RECT 68.480 124.710 68.740 125.030 ;
        RECT 67.100 123.690 67.360 124.010 ;
        RECT 68.480 123.010 68.740 123.330 ;
        RECT 66.640 121.650 66.900 121.970 ;
        RECT 66.640 120.970 66.900 121.290 ;
        RECT 66.180 118.590 66.440 118.910 ;
        RECT 36.170 117.035 37.710 117.405 ;
        RECT 36.170 111.595 37.710 111.965 ;
        RECT 35.820 111.110 36.080 111.430 ;
        RECT 35.360 110.770 35.620 111.090 ;
        RECT 35.360 110.090 35.620 110.410 ;
        RECT 34.900 109.750 35.160 110.070 ;
        RECT 32.870 108.875 34.410 109.245 ;
        RECT 32.140 105.670 32.400 105.990 ;
        RECT 32.200 102.250 32.340 105.670 ;
        RECT 32.870 103.435 34.410 103.805 ;
        RECT 32.140 101.930 32.400 102.250 ;
        RECT 32.870 97.995 34.410 98.365 ;
        RECT 31.220 97.510 31.480 97.830 ;
        RECT 35.420 97.490 35.560 110.090 ;
        RECT 36.170 106.155 37.710 106.525 ;
        RECT 66.700 105.310 66.840 120.970 ;
        RECT 68.540 117.890 68.680 123.010 ;
        RECT 69.000 118.570 69.140 137.630 ;
        RECT 70.380 137.610 70.520 140.010 ;
        RECT 73.600 138.290 73.740 142.050 ;
        RECT 73.540 137.970 73.800 138.290 ;
        RECT 70.320 137.290 70.580 137.610 ;
        RECT 70.380 135.870 70.520 137.290 ;
        RECT 75.440 135.910 75.580 142.730 ;
        RECT 76.360 139.650 76.500 144.770 ;
        RECT 78.660 144.070 78.800 150.210 ;
        RECT 86.940 147.810 87.080 161.430 ;
        RECT 87.860 161.410 88.000 161.860 ;
        RECT 88.260 161.770 88.520 161.860 ;
        RECT 89.640 161.770 89.900 162.090 ;
        RECT 87.800 161.090 88.060 161.410 ;
        RECT 88.260 161.090 88.520 161.410 ;
        RECT 87.860 158.690 88.000 161.090 ;
        RECT 88.320 159.905 88.460 161.090 ;
        RECT 88.720 160.070 88.980 160.390 ;
        RECT 88.250 159.535 88.530 159.905 ;
        RECT 88.260 159.050 88.520 159.370 ;
        RECT 87.800 158.370 88.060 158.690 ;
        RECT 88.320 153.250 88.460 159.050 ;
        RECT 88.780 154.270 88.920 160.070 ;
        RECT 89.180 159.730 89.440 160.050 ;
        RECT 88.720 153.950 88.980 154.270 ;
        RECT 88.260 152.930 88.520 153.250 ;
        RECT 88.320 152.230 88.460 152.930 ;
        RECT 88.260 151.910 88.520 152.230 ;
        RECT 89.240 151.210 89.380 159.730 ;
        RECT 89.700 159.710 89.840 161.770 ;
        RECT 89.640 159.390 89.900 159.710 ;
        RECT 91.080 151.210 91.220 165.170 ;
        RECT 92.400 162.790 92.660 163.110 ;
        RECT 92.460 159.710 92.600 162.790 ;
        RECT 92.400 159.390 92.660 159.710 ;
        RECT 93.320 153.610 93.580 153.930 ;
        RECT 89.180 150.890 89.440 151.210 ;
        RECT 91.020 150.890 91.280 151.210 ;
        RECT 92.860 150.550 93.120 150.870 ;
        RECT 88.260 150.210 88.520 150.530 ;
        RECT 87.340 148.170 87.600 148.490 ;
        RECT 86.880 147.490 87.140 147.810 ;
        RECT 79.060 145.450 79.320 145.770 ;
        RECT 79.980 145.450 80.240 145.770 ;
        RECT 78.600 143.750 78.860 144.070 ;
        RECT 78.140 142.730 78.400 143.050 ;
        RECT 76.760 142.050 77.020 142.370 ;
        RECT 76.820 141.350 76.960 142.050 ;
        RECT 76.760 141.030 77.020 141.350 ;
        RECT 78.200 141.010 78.340 142.730 ;
        RECT 78.140 140.690 78.400 141.010 ;
        RECT 77.220 140.350 77.480 140.670 ;
        RECT 76.300 139.330 76.560 139.650 ;
        RECT 69.920 135.730 70.520 135.870 ;
        RECT 69.920 132.170 70.060 135.730 ;
        RECT 75.380 135.590 75.640 135.910 ;
        RECT 72.160 134.570 72.420 134.890 ;
        RECT 69.860 131.850 70.120 132.170 ;
        RECT 69.920 127.070 70.060 131.850 ;
        RECT 70.320 129.470 70.580 129.790 ;
        RECT 70.380 128.770 70.520 129.470 ;
        RECT 70.320 128.450 70.580 128.770 ;
        RECT 69.860 126.750 70.120 127.070 ;
        RECT 72.220 124.350 72.360 134.570 ;
        RECT 77.280 132.850 77.420 140.350 ;
        RECT 78.200 133.190 78.340 140.690 ;
        RECT 79.120 139.990 79.260 145.450 ;
        RECT 79.520 144.770 79.780 145.090 ;
        RECT 79.580 143.050 79.720 144.770 ;
        RECT 79.520 142.730 79.780 143.050 ;
        RECT 79.580 140.330 79.720 142.730 ;
        RECT 79.520 140.010 79.780 140.330 ;
        RECT 78.600 139.670 78.860 139.990 ;
        RECT 79.060 139.670 79.320 139.990 ;
        RECT 78.660 138.290 78.800 139.670 ;
        RECT 79.120 138.630 79.260 139.670 ;
        RECT 79.520 139.390 79.780 139.650 ;
        RECT 80.040 139.390 80.180 145.450 ;
        RECT 83.660 144.770 83.920 145.090 ;
        RECT 80.440 143.750 80.700 144.070 ;
        RECT 80.500 140.330 80.640 143.750 ;
        RECT 83.720 142.370 83.860 144.770 ;
        RECT 86.420 143.410 86.680 143.730 ;
        RECT 85.960 143.070 86.220 143.390 ;
        RECT 83.660 142.050 83.920 142.370 ;
        RECT 83.720 140.670 83.860 142.050 ;
        RECT 86.020 141.350 86.160 143.070 ;
        RECT 86.480 141.350 86.620 143.410 ;
        RECT 85.960 141.030 86.220 141.350 ;
        RECT 86.420 141.030 86.680 141.350 ;
        RECT 83.660 140.350 83.920 140.670 ;
        RECT 80.440 140.010 80.700 140.330 ;
        RECT 81.820 139.670 82.080 139.990 ;
        RECT 79.520 139.330 80.180 139.390 ;
        RECT 79.580 139.250 80.180 139.330 ;
        RECT 79.060 138.310 79.320 138.630 ;
        RECT 78.600 137.970 78.860 138.290 ;
        RECT 78.660 135.570 78.800 137.970 ;
        RECT 79.120 137.610 79.260 138.310 ;
        RECT 79.060 137.290 79.320 137.610 ;
        RECT 79.580 137.270 79.720 139.250 ;
        RECT 79.980 137.630 80.240 137.950 ;
        RECT 79.520 136.950 79.780 137.270 ;
        RECT 78.600 135.250 78.860 135.570 ;
        RECT 79.580 134.890 79.720 136.950 ;
        RECT 80.040 135.910 80.180 137.630 ;
        RECT 81.880 137.610 82.020 139.670 ;
        RECT 81.820 137.290 82.080 137.610 ;
        RECT 82.280 137.290 82.540 137.610 ;
        RECT 79.980 135.590 80.240 135.910 ;
        RECT 79.520 134.570 79.780 134.890 ;
        RECT 78.140 132.870 78.400 133.190 ;
        RECT 77.220 132.760 77.480 132.850 ;
        RECT 77.220 132.620 77.880 132.760 ;
        RECT 77.220 132.530 77.480 132.620 ;
        RECT 76.300 131.850 76.560 132.170 ;
        RECT 76.360 130.470 76.500 131.850 ;
        RECT 72.620 130.150 72.880 130.470 ;
        RECT 76.300 130.150 76.560 130.470 ;
        RECT 72.160 124.030 72.420 124.350 ;
        RECT 72.220 122.310 72.360 124.030 ;
        RECT 72.160 121.990 72.420 122.310 ;
        RECT 70.780 121.310 71.040 121.630 ;
        RECT 70.840 119.590 70.980 121.310 ;
        RECT 70.780 119.270 71.040 119.590 ;
        RECT 72.680 118.910 72.820 130.150 ;
        RECT 73.540 129.810 73.800 130.130 ;
        RECT 73.600 127.750 73.740 129.810 ;
        RECT 74.000 129.470 74.260 129.790 ;
        RECT 73.540 127.430 73.800 127.750 ;
        RECT 74.060 124.010 74.200 129.470 ;
        RECT 76.360 126.050 76.500 130.150 ;
        RECT 77.220 129.130 77.480 129.450 ;
        RECT 77.280 127.070 77.420 129.130 ;
        RECT 77.740 128.770 77.880 132.620 ;
        RECT 81.880 132.170 82.020 137.290 ;
        RECT 82.340 135.910 82.480 137.290 ;
        RECT 82.280 135.590 82.540 135.910 ;
        RECT 83.720 135.870 83.860 140.350 ;
        RECT 86.420 139.330 86.680 139.650 ;
        RECT 86.480 136.930 86.620 139.330 ;
        RECT 85.500 136.610 85.760 136.930 ;
        RECT 86.420 136.610 86.680 136.930 ;
        RECT 83.260 135.730 83.860 135.870 ;
        RECT 82.740 132.190 83.000 132.510 ;
        RECT 81.820 131.850 82.080 132.170 ;
        RECT 82.800 129.450 82.940 132.190 ;
        RECT 82.740 129.130 83.000 129.450 ;
        RECT 77.680 128.450 77.940 128.770 ;
        RECT 77.740 127.070 77.880 128.450 ;
        RECT 82.800 127.150 82.940 129.130 ;
        RECT 82.340 127.070 82.940 127.150 ;
        RECT 77.220 126.750 77.480 127.070 ;
        RECT 77.680 126.750 77.940 127.070 ;
        RECT 82.280 127.010 82.940 127.070 ;
        RECT 82.280 126.750 82.540 127.010 ;
        RECT 76.300 125.730 76.560 126.050 ;
        RECT 76.360 125.030 76.500 125.730 ;
        RECT 77.280 125.030 77.420 126.750 ;
        RECT 80.440 126.470 80.700 126.730 ;
        RECT 80.440 126.410 82.020 126.470 ;
        RECT 80.500 126.390 82.020 126.410 ;
        RECT 80.500 126.330 82.080 126.390 ;
        RECT 81.820 126.070 82.080 126.330 ;
        RECT 79.980 125.730 80.240 126.050 ;
        RECT 82.280 125.730 82.540 126.050 ;
        RECT 80.040 125.030 80.180 125.730 ;
        RECT 76.300 124.710 76.560 125.030 ;
        RECT 77.220 124.710 77.480 125.030 ;
        RECT 79.980 124.710 80.240 125.030 ;
        RECT 74.000 123.690 74.260 124.010 ;
        RECT 73.080 120.290 73.340 120.610 ;
        RECT 77.220 120.290 77.480 120.610 ;
        RECT 72.620 118.590 72.880 118.910 ;
        RECT 68.940 118.250 69.200 118.570 ;
        RECT 73.140 118.230 73.280 120.290 ;
        RECT 77.280 118.230 77.420 120.290 ;
        RECT 82.340 118.910 82.480 125.730 ;
        RECT 82.740 121.310 83.000 121.630 ;
        RECT 82.800 119.590 82.940 121.310 ;
        RECT 82.740 119.270 83.000 119.590 ;
        RECT 82.280 118.590 82.540 118.910 ;
        RECT 73.080 117.910 73.340 118.230 ;
        RECT 77.220 117.910 77.480 118.230 ;
        RECT 68.480 117.570 68.740 117.890 ;
        RECT 71.700 117.570 71.960 117.890 ;
        RECT 66.640 104.990 66.900 105.310 ;
        RECT 66.700 102.250 66.840 104.990 ;
        RECT 68.480 102.610 68.740 102.930 ;
        RECT 61.580 101.930 61.840 102.250 ;
        RECT 66.640 101.930 66.900 102.250 ;
        RECT 36.170 100.715 37.710 101.085 ;
        RECT 35.360 97.230 35.620 97.490 ;
        RECT 34.500 97.170 35.620 97.230 ;
        RECT 34.500 97.090 35.560 97.170 ;
        RECT 34.500 96.810 34.640 97.090 ;
        RECT 61.120 96.830 61.380 97.150 ;
        RECT 32.600 96.490 32.860 96.810 ;
        RECT 34.440 96.490 34.700 96.810 ;
        RECT 35.360 96.490 35.620 96.810 ;
        RECT 31.220 96.150 31.480 96.470 ;
        RECT 31.280 94.430 31.420 96.150 ;
        RECT 31.220 94.110 31.480 94.430 ;
        RECT 32.140 94.340 32.400 94.430 ;
        RECT 31.740 94.200 32.400 94.340 ;
        RECT 31.740 91.790 31.880 94.200 ;
        RECT 32.140 94.110 32.400 94.200 ;
        RECT 32.660 93.320 32.800 96.490 ;
        RECT 33.980 95.810 34.240 96.130 ;
        RECT 33.520 94.110 33.780 94.430 ;
        RECT 33.580 93.410 33.720 94.110 ;
        RECT 34.040 93.410 34.180 95.810 ;
        RECT 35.420 94.770 35.560 96.490 ;
        RECT 35.820 95.810 36.080 96.130 ;
        RECT 35.360 94.450 35.620 94.770 ;
        RECT 35.360 93.770 35.620 94.090 ;
        RECT 32.200 93.180 32.800 93.320 ;
        RECT 32.200 92.390 32.340 93.180 ;
        RECT 33.520 93.090 33.780 93.410 ;
        RECT 33.980 93.090 34.240 93.410 ;
        RECT 34.900 93.090 35.160 93.410 ;
        RECT 32.870 92.555 34.410 92.925 ;
        RECT 32.140 92.070 32.400 92.390 ;
        RECT 31.740 91.650 32.800 91.790 ;
        RECT 32.660 91.370 32.800 91.650 ;
        RECT 32.140 91.050 32.400 91.370 ;
        RECT 32.600 91.050 32.860 91.370 ;
        RECT 33.980 91.050 34.240 91.370 ;
        RECT 31.220 90.370 31.480 90.690 ;
        RECT 30.760 89.350 31.020 89.670 ;
        RECT 31.280 88.990 31.420 90.370 ;
        RECT 31.220 88.670 31.480 88.990 ;
        RECT 28.920 86.630 29.180 86.950 ;
        RECT 29.840 86.630 30.100 86.950 ;
        RECT 32.200 86.860 32.340 91.050 ;
        RECT 32.660 87.970 32.800 91.050 ;
        RECT 33.520 90.710 33.780 91.030 ;
        RECT 33.580 88.990 33.720 90.710 ;
        RECT 34.040 89.670 34.180 91.050 ;
        RECT 33.980 89.350 34.240 89.670 ;
        RECT 33.520 88.670 33.780 88.990 ;
        RECT 32.600 87.650 32.860 87.970 ;
        RECT 32.870 87.115 34.410 87.485 ;
        RECT 32.200 86.720 33.720 86.860 ;
        RECT 33.580 85.930 33.720 86.720 ;
        RECT 34.960 86.610 35.100 93.090 ;
        RECT 35.420 91.710 35.560 93.770 ;
        RECT 35.360 91.390 35.620 91.710 ;
        RECT 35.360 90.370 35.620 90.690 ;
        RECT 35.420 89.330 35.560 90.370 ;
        RECT 35.360 89.010 35.620 89.330 ;
        RECT 35.360 88.560 35.620 88.650 ;
        RECT 35.880 88.560 36.020 95.810 ;
        RECT 36.170 95.275 37.710 95.645 ;
        RECT 61.180 94.770 61.320 96.830 ;
        RECT 36.740 94.450 37.000 94.770 ;
        RECT 61.120 94.450 61.380 94.770 ;
        RECT 36.800 91.030 36.940 94.450 ;
        RECT 61.640 94.430 61.780 101.930 ;
        RECT 64.800 101.590 65.060 101.910 ;
        RECT 64.860 100.550 65.000 101.590 ;
        RECT 64.800 100.230 65.060 100.550 ;
        RECT 68.540 100.210 68.680 102.610 ;
        RECT 71.240 102.270 71.500 102.590 ;
        RECT 70.320 101.250 70.580 101.570 ;
        RECT 70.780 101.250 71.040 101.570 ;
        RECT 67.100 99.890 67.360 100.210 ;
        RECT 68.480 99.890 68.740 100.210 ;
        RECT 67.160 97.150 67.300 99.890 ;
        RECT 69.400 97.170 69.660 97.490 ;
        RECT 67.100 96.830 67.360 97.150 ;
        RECT 68.480 96.490 68.740 96.810 ;
        RECT 64.340 95.810 64.600 96.130 ;
        RECT 67.100 95.810 67.360 96.130 ;
        RECT 64.400 94.770 64.540 95.810 ;
        RECT 64.340 94.450 64.600 94.770 ;
        RECT 38.580 94.110 38.840 94.430 ;
        RECT 39.960 94.110 40.220 94.430 ;
        RECT 41.340 94.110 41.600 94.430 ;
        RECT 41.800 94.110 42.060 94.430 ;
        RECT 61.580 94.110 61.840 94.430 ;
        RECT 64.800 94.110 65.060 94.430 ;
        RECT 38.120 93.090 38.380 93.410 ;
        RECT 36.740 90.710 37.000 91.030 ;
        RECT 36.170 89.835 37.710 90.205 ;
        RECT 37.660 88.670 37.920 88.990 ;
        RECT 35.360 88.420 36.020 88.560 ;
        RECT 35.360 88.330 35.620 88.420 ;
        RECT 36.280 88.330 36.540 88.650 ;
        RECT 36.340 86.950 36.480 88.330 ;
        RECT 36.740 87.650 37.000 87.970 ;
        RECT 36.800 86.950 36.940 87.650 ;
        RECT 36.280 86.630 36.540 86.950 ;
        RECT 36.740 86.630 37.000 86.950 ;
        RECT 37.720 86.610 37.860 88.670 ;
        RECT 38.180 86.610 38.320 93.090 ;
        RECT 38.640 88.990 38.780 94.110 ;
        RECT 39.500 91.390 39.760 91.710 ;
        RECT 39.560 91.110 39.700 91.390 ;
        RECT 39.100 90.970 39.700 91.110 ;
        RECT 38.580 88.670 38.840 88.990 ;
        RECT 39.100 87.970 39.240 90.970 ;
        RECT 40.020 90.690 40.160 94.110 ;
        RECT 40.880 93.770 41.140 94.090 ;
        RECT 40.420 91.050 40.680 91.370 ;
        RECT 39.960 90.430 40.220 90.690 ;
        RECT 39.560 90.370 40.220 90.430 ;
        RECT 39.560 90.290 40.160 90.370 ;
        RECT 39.560 88.990 39.700 90.290 ;
        RECT 39.500 88.670 39.760 88.990 ;
        RECT 39.040 87.650 39.300 87.970 ;
        RECT 34.900 86.290 35.160 86.610 ;
        RECT 37.660 86.290 37.920 86.610 ;
        RECT 38.120 86.290 38.380 86.610 ;
        RECT 28.460 85.610 28.720 85.930 ;
        RECT 31.220 85.610 31.480 85.930 ;
        RECT 33.520 85.610 33.780 85.930 ;
        RECT 34.900 85.840 35.160 85.930 ;
        RECT 34.500 85.700 35.160 85.840 ;
        RECT 25.700 85.270 25.960 85.590 ;
        RECT 27.540 85.270 27.800 85.590 ;
        RECT 28.000 84.930 28.260 85.250 ;
        RECT 28.060 77.700 28.200 84.930 ;
        RECT 31.280 77.700 31.420 85.610 ;
        RECT 33.580 84.230 33.720 85.610 ;
        RECT 33.520 83.910 33.780 84.230 ;
        RECT 34.500 77.700 34.640 85.700 ;
        RECT 34.900 85.610 35.160 85.700 ;
        RECT 38.120 85.610 38.380 85.930 ;
        RECT 36.170 84.395 37.710 84.765 ;
        RECT 38.180 80.230 38.320 85.610 ;
        RECT 39.100 85.250 39.240 87.650 ;
        RECT 39.560 86.950 39.700 88.670 ;
        RECT 40.480 88.650 40.620 91.050 ;
        RECT 40.940 91.030 41.080 93.770 ;
        RECT 41.400 92.050 41.540 94.110 ;
        RECT 41.340 91.730 41.600 92.050 ;
        RECT 40.880 90.710 41.140 91.030 ;
        RECT 40.940 88.990 41.080 90.710 ;
        RECT 41.860 89.670 42.000 94.110 ;
        RECT 43.640 93.430 43.900 93.750 ;
        RECT 42.260 92.070 42.520 92.390 ;
        RECT 41.800 89.350 42.060 89.670 ;
        RECT 42.320 88.990 42.460 92.070 ;
        RECT 43.700 89.670 43.840 93.430 ;
        RECT 44.560 93.090 44.820 93.410 ;
        RECT 58.820 93.090 59.080 93.410 ;
        RECT 43.640 89.350 43.900 89.670 ;
        RECT 44.620 88.990 44.760 93.090 ;
        RECT 48.240 91.730 48.500 92.050 ;
        RECT 46.860 91.050 47.120 91.370 ;
        RECT 45.940 90.370 46.200 90.690 ;
        RECT 46.000 88.990 46.140 90.370 ;
        RECT 40.880 88.670 41.140 88.990 ;
        RECT 42.260 88.670 42.520 88.990 ;
        RECT 44.560 88.670 44.820 88.990 ;
        RECT 45.940 88.670 46.200 88.990 ;
        RECT 40.420 88.330 40.680 88.650 ;
        RECT 40.940 86.950 41.080 88.670 ;
        RECT 39.500 86.630 39.760 86.950 ;
        RECT 40.880 86.630 41.140 86.950 ;
        RECT 42.320 86.610 42.460 88.670 ;
        RECT 42.260 86.290 42.520 86.610 ;
        RECT 40.880 85.610 41.140 85.930 ;
        RECT 44.100 85.610 44.360 85.930 ;
        RECT 39.040 84.930 39.300 85.250 ;
        RECT 37.720 80.090 38.320 80.230 ;
        RECT 37.720 77.700 37.860 80.090 ;
        RECT 40.940 77.700 41.080 85.610 ;
        RECT 44.160 77.700 44.300 85.610 ;
        RECT 46.000 85.590 46.140 88.670 ;
        RECT 46.920 87.970 47.060 91.050 ;
        RECT 48.300 89.670 48.440 91.730 ;
        RECT 58.880 91.030 59.020 93.090 ;
        RECT 61.640 92.390 61.780 94.110 ;
        RECT 61.580 92.070 61.840 92.390 ;
        RECT 61.640 91.370 61.780 92.070 ;
        RECT 61.580 91.050 61.840 91.370 ;
        RECT 58.820 90.710 59.080 91.030 ;
        RECT 48.240 89.350 48.500 89.670 ;
        RECT 61.640 89.330 61.780 91.050 ;
        RECT 61.580 89.010 61.840 89.330 ;
        RECT 56.980 88.670 57.240 88.990 ;
        RECT 62.040 88.670 62.300 88.990 ;
        RECT 46.860 87.650 47.120 87.970 ;
        RECT 48.700 87.650 48.960 87.970 ;
        RECT 48.760 86.950 48.900 87.650 ;
        RECT 48.700 86.630 48.960 86.950 ;
        RECT 47.320 85.610 47.580 85.930 ;
        RECT 50.540 85.610 50.800 85.930 ;
        RECT 53.760 85.610 54.020 85.930 ;
        RECT 45.940 85.270 46.200 85.590 ;
        RECT 47.380 77.700 47.520 85.610 ;
        RECT 47.780 84.930 48.040 85.250 ;
        RECT 47.840 84.230 47.980 84.930 ;
        RECT 47.780 83.910 48.040 84.230 ;
        RECT 50.600 77.700 50.740 85.610 ;
        RECT 53.820 77.700 53.960 85.610 ;
        RECT 57.040 77.700 57.180 88.670 ;
        RECT 62.100 86.950 62.240 88.670 ;
        RECT 62.040 86.630 62.300 86.950 ;
        RECT 60.200 86.290 60.460 86.610 ;
        RECT 57.900 85.610 58.160 85.930 ;
        RECT 57.960 84.230 58.100 85.610 ;
        RECT 57.900 83.910 58.160 84.230 ;
        RECT 60.260 77.700 60.400 86.290 ;
        RECT 64.860 85.590 65.000 94.110 ;
        RECT 66.180 93.090 66.440 93.410 ;
        RECT 66.240 85.590 66.380 93.090 ;
        RECT 67.160 86.610 67.300 95.810 ;
        RECT 68.540 92.390 68.680 96.490 ;
        RECT 68.940 95.810 69.200 96.130 ;
        RECT 68.480 92.070 68.740 92.390 ;
        RECT 68.480 91.050 68.740 91.370 ;
        RECT 68.020 90.710 68.280 91.030 ;
        RECT 67.560 89.350 67.820 89.670 ;
        RECT 67.100 86.290 67.360 86.610 ;
        RECT 67.620 85.930 67.760 89.350 ;
        RECT 68.080 86.950 68.220 90.710 ;
        RECT 68.540 87.570 68.680 91.050 ;
        RECT 69.000 89.670 69.140 95.810 ;
        RECT 69.460 95.110 69.600 97.170 ;
        RECT 69.400 94.790 69.660 95.110 ;
        RECT 70.380 91.370 70.520 101.250 ;
        RECT 70.840 99.190 70.980 101.250 ;
        RECT 70.780 98.870 71.040 99.190 ;
        RECT 71.300 97.150 71.440 102.270 ;
        RECT 71.760 99.530 71.900 117.570 ;
        RECT 73.140 108.790 73.280 117.910 ;
        RECT 80.440 111.110 80.700 111.430 ;
        RECT 79.060 110.430 79.320 110.750 ;
        RECT 74.000 110.090 74.260 110.410 ;
        RECT 72.680 108.650 73.280 108.790 ;
        RECT 72.680 102.250 72.820 108.650 ;
        RECT 73.080 107.710 73.340 108.030 ;
        RECT 73.140 105.990 73.280 107.710 ;
        RECT 74.060 107.010 74.200 110.090 ;
        RECT 76.300 109.410 76.560 109.730 ;
        RECT 76.360 107.350 76.500 109.410 ;
        RECT 76.300 107.030 76.560 107.350 ;
        RECT 73.540 106.690 73.800 107.010 ;
        RECT 74.000 106.690 74.260 107.010 ;
        RECT 73.080 105.670 73.340 105.990 ;
        RECT 73.600 105.650 73.740 106.690 ;
        RECT 73.540 105.330 73.800 105.650 ;
        RECT 74.060 102.930 74.200 106.690 ;
        RECT 79.120 104.290 79.260 110.430 ;
        RECT 79.980 109.750 80.240 110.070 ;
        RECT 80.040 107.010 80.180 109.750 ;
        RECT 79.980 106.690 80.240 107.010 ;
        RECT 80.040 105.990 80.180 106.690 ;
        RECT 79.980 105.670 80.240 105.990 ;
        RECT 77.680 103.970 77.940 104.290 ;
        RECT 79.060 103.970 79.320 104.290 ;
        RECT 74.000 102.610 74.260 102.930 ;
        RECT 72.620 101.930 72.880 102.250 ;
        RECT 74.060 101.990 74.200 102.610 ;
        RECT 73.600 101.850 74.200 101.990 ;
        RECT 71.700 99.210 71.960 99.530 ;
        RECT 71.240 96.830 71.500 97.150 ;
        RECT 70.780 94.790 71.040 95.110 ;
        RECT 70.840 94.625 70.980 94.790 ;
        RECT 70.770 94.255 71.050 94.625 ;
        RECT 71.300 93.830 71.440 96.830 ;
        RECT 71.760 94.625 71.900 99.210 ;
        RECT 72.160 96.150 72.420 96.470 ;
        RECT 73.080 96.150 73.340 96.470 ;
        RECT 72.220 94.770 72.360 96.150 ;
        RECT 73.140 95.110 73.280 96.150 ;
        RECT 73.080 94.790 73.340 95.110 ;
        RECT 71.690 94.255 71.970 94.625 ;
        RECT 72.160 94.450 72.420 94.770 ;
        RECT 71.700 93.830 71.960 94.090 ;
        RECT 71.300 93.770 71.960 93.830 ;
        RECT 71.300 93.690 71.900 93.770 ;
        RECT 71.240 92.070 71.500 92.390 ;
        RECT 70.320 91.050 70.580 91.370 ;
        RECT 69.860 90.710 70.120 91.030 ;
        RECT 68.940 89.350 69.200 89.670 ;
        RECT 69.000 88.310 69.140 89.350 ;
        RECT 68.940 87.990 69.200 88.310 ;
        RECT 69.400 87.650 69.660 87.970 ;
        RECT 68.540 87.430 69.140 87.570 ;
        RECT 68.020 86.630 68.280 86.950 ;
        RECT 67.560 85.610 67.820 85.930 ;
        RECT 63.420 85.270 63.680 85.590 ;
        RECT 64.800 85.270 65.060 85.590 ;
        RECT 66.180 85.270 66.440 85.590 ;
        RECT 63.480 77.700 63.620 85.270 ;
        RECT 66.640 84.930 66.900 85.250 ;
        RECT 66.700 77.700 66.840 84.930 ;
        RECT 69.000 84.230 69.140 87.430 ;
        RECT 69.460 86.610 69.600 87.650 ;
        RECT 69.400 86.290 69.660 86.610 ;
        RECT 68.940 83.910 69.200 84.230 ;
        RECT 69.920 77.700 70.060 90.710 ;
        RECT 71.300 87.570 71.440 92.070 ;
        RECT 72.220 91.110 72.360 94.450 ;
        RECT 73.140 91.370 73.280 94.790 ;
        RECT 73.600 94.430 73.740 101.850 ;
        RECT 74.460 96.830 74.720 97.150 ;
        RECT 74.000 94.790 74.260 95.110 ;
        RECT 73.540 94.110 73.800 94.430 ;
        RECT 71.760 90.970 72.360 91.110 ;
        RECT 73.080 91.050 73.340 91.370 ;
        RECT 71.760 88.990 71.900 90.970 ;
        RECT 72.160 90.370 72.420 90.690 ;
        RECT 72.220 89.670 72.360 90.370 ;
        RECT 72.160 89.350 72.420 89.670 ;
        RECT 71.700 88.670 71.960 88.990 ;
        RECT 73.540 88.670 73.800 88.990 ;
        RECT 72.620 88.330 72.880 88.650 ;
        RECT 71.300 87.430 71.900 87.570 ;
        RECT 71.230 86.095 71.510 86.465 ;
        RECT 71.760 86.270 71.900 87.430 ;
        RECT 72.680 86.270 72.820 88.330 ;
        RECT 71.300 85.930 71.440 86.095 ;
        RECT 71.700 85.950 71.960 86.270 ;
        RECT 72.620 85.950 72.880 86.270 ;
        RECT 73.600 85.930 73.740 88.670 ;
        RECT 74.060 88.650 74.200 94.790 ;
        RECT 74.520 89.330 74.660 96.830 ;
        RECT 75.380 96.150 75.640 96.470 ;
        RECT 74.460 89.010 74.720 89.330 ;
        RECT 75.440 88.990 75.580 96.150 ;
        RECT 75.840 93.090 76.100 93.410 ;
        RECT 75.900 91.030 76.040 93.090 ;
        RECT 75.840 90.710 76.100 91.030 ;
        RECT 75.380 88.670 75.640 88.990 ;
        RECT 74.000 88.330 74.260 88.650 ;
        RECT 77.740 85.930 77.880 103.970 ;
        RECT 79.120 102.590 79.260 103.970 ;
        RECT 79.060 102.270 79.320 102.590 ;
        RECT 78.140 101.930 78.400 102.250 ;
        RECT 78.200 99.190 78.340 101.930 ;
        RECT 78.140 98.870 78.400 99.190 ;
        RECT 78.200 94.430 78.340 98.870 ;
        RECT 79.520 98.530 79.780 98.850 ;
        RECT 79.580 94.770 79.720 98.530 ;
        RECT 79.520 94.450 79.780 94.770 ;
        RECT 78.140 94.110 78.400 94.430 ;
        RECT 78.140 93.430 78.400 93.750 ;
        RECT 78.200 90.690 78.340 93.430 ;
        RECT 78.140 90.370 78.400 90.690 ;
        RECT 78.200 85.930 78.340 90.370 ;
        RECT 80.040 85.930 80.180 105.670 ;
        RECT 80.500 105.650 80.640 111.110 ;
        RECT 80.900 107.370 81.160 107.690 ;
        RECT 80.440 105.330 80.700 105.650 ;
        RECT 80.960 94.430 81.100 107.370 ;
        RECT 83.260 98.850 83.400 135.730 ;
        RECT 85.560 134.890 85.700 136.610 ;
        RECT 85.500 134.570 85.760 134.890 ;
        RECT 85.960 132.530 86.220 132.850 ;
        RECT 85.500 132.190 85.760 132.510 ;
        RECT 85.560 130.470 85.700 132.190 ;
        RECT 85.500 130.150 85.760 130.470 ;
        RECT 86.020 129.450 86.160 132.530 ;
        RECT 86.420 131.850 86.680 132.170 ;
        RECT 85.960 129.130 86.220 129.450 ;
        RECT 86.020 127.070 86.160 129.130 ;
        RECT 85.960 126.750 86.220 127.070 ;
        RECT 84.580 125.730 84.840 126.050 ;
        RECT 84.640 124.350 84.780 125.730 ;
        RECT 84.580 124.030 84.840 124.350 ;
        RECT 86.480 124.010 86.620 131.850 ;
        RECT 86.940 129.110 87.080 147.490 ;
        RECT 87.400 146.790 87.540 148.170 ;
        RECT 87.340 146.470 87.600 146.790 ;
        RECT 87.800 140.010 88.060 140.330 ;
        RECT 87.860 138.630 88.000 140.010 ;
        RECT 88.320 139.990 88.460 150.210 ;
        RECT 92.920 149.510 93.060 150.550 ;
        RECT 92.860 149.190 93.120 149.510 ;
        RECT 90.560 143.410 90.820 143.730 ;
        RECT 90.620 140.670 90.760 143.410 ;
        RECT 90.560 140.350 90.820 140.670 ;
        RECT 88.260 139.670 88.520 139.990 ;
        RECT 87.800 138.310 88.060 138.630 ;
        RECT 87.800 137.290 88.060 137.610 ;
        RECT 87.340 136.610 87.600 136.930 ;
        RECT 87.400 134.890 87.540 136.610 ;
        RECT 87.860 135.230 88.000 137.290 ;
        RECT 87.800 134.910 88.060 135.230 ;
        RECT 87.340 134.570 87.600 134.890 ;
        RECT 87.400 132.510 87.540 134.570 ;
        RECT 87.340 132.190 87.600 132.510 ;
        RECT 87.340 131.170 87.600 131.490 ;
        RECT 87.400 129.790 87.540 131.170 ;
        RECT 87.340 129.470 87.600 129.790 ;
        RECT 86.880 128.790 87.140 129.110 ;
        RECT 87.860 127.150 88.000 134.910 ;
        RECT 89.640 134.230 89.900 134.550 ;
        RECT 89.700 133.190 89.840 134.230 ;
        RECT 89.640 132.870 89.900 133.190 ;
        RECT 90.100 131.850 90.360 132.170 ;
        RECT 90.160 129.450 90.300 131.850 ;
        RECT 93.380 129.450 93.520 153.610 ;
        RECT 94.240 151.910 94.500 152.230 ;
        RECT 94.300 146.110 94.440 151.910 ;
        RECT 95.680 149.510 95.820 171.970 ;
        RECT 96.140 167.530 96.280 171.970 ;
        RECT 96.080 167.210 96.340 167.530 ;
        RECT 96.080 150.210 96.340 150.530 ;
        RECT 95.620 149.190 95.880 149.510 ;
        RECT 94.240 145.790 94.500 146.110 ;
        RECT 93.780 145.110 94.040 145.430 ;
        RECT 93.840 144.070 93.980 145.110 ;
        RECT 93.780 143.750 94.040 144.070 ;
        RECT 93.840 143.050 93.980 143.750 ;
        RECT 94.300 143.730 94.440 145.790 ;
        RECT 94.700 145.110 94.960 145.430 ;
        RECT 94.240 143.410 94.500 143.730 ;
        RECT 93.780 142.730 94.040 143.050 ;
        RECT 94.760 142.710 94.900 145.110 ;
        RECT 94.700 142.390 94.960 142.710 ;
        RECT 94.240 142.050 94.500 142.370 ;
        RECT 94.300 140.330 94.440 142.050 ;
        RECT 94.240 140.010 94.500 140.330 ;
        RECT 95.160 133.890 95.420 134.210 ;
        RECT 95.220 133.190 95.360 133.890 ;
        RECT 95.160 132.870 95.420 133.190 ;
        RECT 90.100 129.130 90.360 129.450 ;
        RECT 93.320 129.130 93.580 129.450 ;
        RECT 89.640 128.790 89.900 129.110 ;
        RECT 88.260 128.450 88.520 128.770 ;
        RECT 88.320 127.410 88.460 128.450 ;
        RECT 87.400 127.070 88.000 127.150 ;
        RECT 88.260 127.090 88.520 127.410 ;
        RECT 87.340 127.010 88.000 127.070 ;
        RECT 87.340 126.750 87.600 127.010 ;
        RECT 87.860 124.350 88.000 127.010 ;
        RECT 87.800 124.030 88.060 124.350 ;
        RECT 86.420 123.690 86.680 124.010 ;
        RECT 86.480 118.570 86.620 123.690 ;
        RECT 86.880 123.010 87.140 123.330 ;
        RECT 86.940 121.630 87.080 123.010 ;
        RECT 87.860 121.970 88.000 124.030 ;
        RECT 87.800 121.650 88.060 121.970 ;
        RECT 86.880 121.310 87.140 121.630 ;
        RECT 86.420 118.250 86.680 118.570 ;
        RECT 86.420 117.570 86.680 117.890 ;
        RECT 85.960 112.470 86.220 112.790 ;
        RECT 83.660 110.770 83.920 111.090 ;
        RECT 83.720 105.650 83.860 110.770 ;
        RECT 85.500 110.090 85.760 110.410 ;
        RECT 84.120 109.410 84.380 109.730 ;
        RECT 83.660 105.330 83.920 105.650 ;
        RECT 83.200 98.530 83.460 98.850 ;
        RECT 83.720 97.150 83.860 105.330 ;
        RECT 84.180 102.930 84.320 109.410 ;
        RECT 84.580 107.030 84.840 107.350 ;
        RECT 84.640 103.270 84.780 107.030 ;
        RECT 85.040 106.690 85.300 107.010 ;
        RECT 85.100 105.310 85.240 106.690 ;
        RECT 85.040 104.990 85.300 105.310 ;
        RECT 84.580 102.950 84.840 103.270 ;
        RECT 84.120 102.610 84.380 102.930 ;
        RECT 83.660 96.830 83.920 97.150 ;
        RECT 85.100 96.470 85.240 104.990 ;
        RECT 85.040 96.150 85.300 96.470 ;
        RECT 81.820 95.810 82.080 96.130 ;
        RECT 81.880 94.430 82.020 95.810 ;
        RECT 80.900 94.110 81.160 94.430 ;
        RECT 81.820 94.110 82.080 94.430 ;
        RECT 80.960 91.370 81.100 94.110 ;
        RECT 85.100 91.710 85.240 96.150 ;
        RECT 85.560 93.410 85.700 110.090 ;
        RECT 86.020 96.810 86.160 112.470 ;
        RECT 86.480 111.430 86.620 117.570 ;
        RECT 86.880 115.870 87.140 116.190 ;
        RECT 86.420 111.110 86.680 111.430 ;
        RECT 86.420 107.600 86.680 107.690 ;
        RECT 86.940 107.600 87.080 115.870 ;
        RECT 87.860 115.850 88.000 121.650 ;
        RECT 89.700 118.570 89.840 128.790 ;
        RECT 90.560 128.450 90.820 128.770 ;
        RECT 91.020 128.450 91.280 128.770 ;
        RECT 90.620 126.050 90.760 128.450 ;
        RECT 90.560 125.730 90.820 126.050 ;
        RECT 91.080 124.010 91.220 128.450 ;
        RECT 91.020 123.690 91.280 124.010 ;
        RECT 89.640 118.250 89.900 118.570 ;
        RECT 88.720 117.910 88.980 118.230 ;
        RECT 88.780 116.190 88.920 117.910 ;
        RECT 89.700 116.190 89.840 118.250 ;
        RECT 93.380 116.950 93.520 129.130 ;
        RECT 94.700 128.450 94.960 128.770 ;
        RECT 93.780 125.730 94.040 126.050 ;
        RECT 93.840 124.350 93.980 125.730 ;
        RECT 93.780 124.030 94.040 124.350 ;
        RECT 94.760 123.330 94.900 128.450 ;
        RECT 94.700 123.010 94.960 123.330 ;
        RECT 93.380 116.810 93.980 116.950 ;
        RECT 88.720 115.870 88.980 116.190 ;
        RECT 89.640 115.870 89.900 116.190 ;
        RECT 87.800 115.530 88.060 115.850 ;
        RECT 93.320 115.530 93.580 115.850 ;
        RECT 91.940 113.830 92.200 114.150 ;
        RECT 88.720 113.490 88.980 113.810 ;
        RECT 88.260 112.130 88.520 112.450 ;
        RECT 87.800 109.750 88.060 110.070 ;
        RECT 86.420 107.460 87.080 107.600 ;
        RECT 86.420 107.370 86.680 107.460 ;
        RECT 86.940 105.310 87.080 107.460 ;
        RECT 86.880 104.990 87.140 105.310 ;
        RECT 86.420 104.650 86.680 104.970 ;
        RECT 87.860 104.710 88.000 109.750 ;
        RECT 88.320 105.310 88.460 112.130 ;
        RECT 88.780 108.710 88.920 113.490 ;
        RECT 90.100 111.110 90.360 111.430 ;
        RECT 89.180 110.430 89.440 110.750 ;
        RECT 88.720 108.390 88.980 108.710 ;
        RECT 89.240 107.010 89.380 110.430 ;
        RECT 89.640 107.370 89.900 107.690 ;
        RECT 89.180 106.690 89.440 107.010 ;
        RECT 88.260 104.990 88.520 105.310 ;
        RECT 86.480 103.270 86.620 104.650 ;
        RECT 86.940 104.630 88.000 104.710 ;
        RECT 86.880 104.570 88.000 104.630 ;
        RECT 86.880 104.310 87.140 104.570 ;
        RECT 86.420 102.950 86.680 103.270 ;
        RECT 86.420 98.870 86.680 99.190 ;
        RECT 86.480 96.810 86.620 98.870 ;
        RECT 87.860 97.150 88.000 104.570 ;
        RECT 89.240 101.910 89.380 106.690 ;
        RECT 89.700 102.250 89.840 107.370 ;
        RECT 90.160 107.010 90.300 111.110 ;
        RECT 92.000 110.750 92.140 113.830 ;
        RECT 93.380 113.470 93.520 115.530 ;
        RECT 93.320 113.150 93.580 113.470 ;
        RECT 93.840 110.750 93.980 116.810 ;
        RECT 91.940 110.660 92.200 110.750 ;
        RECT 91.940 110.520 93.060 110.660 ;
        RECT 91.940 110.430 92.200 110.520 ;
        RECT 90.100 106.690 90.360 107.010 ;
        RECT 89.640 101.930 89.900 102.250 ;
        RECT 89.180 101.590 89.440 101.910 ;
        RECT 89.700 99.270 89.840 101.930 ;
        RECT 90.560 101.590 90.820 101.910 ;
        RECT 89.240 99.130 89.840 99.270 ;
        RECT 87.800 96.830 88.060 97.150 ;
        RECT 85.960 96.490 86.220 96.810 ;
        RECT 86.420 96.490 86.680 96.810 ;
        RECT 86.020 94.770 86.160 96.490 ;
        RECT 87.340 95.810 87.600 96.130 ;
        RECT 85.960 94.450 86.220 94.770 ;
        RECT 85.500 93.090 85.760 93.410 ;
        RECT 85.040 91.390 85.300 91.710 ;
        RECT 80.900 91.050 81.160 91.370 ;
        RECT 86.020 91.110 86.160 94.450 ;
        RECT 87.400 93.410 87.540 95.810 ;
        RECT 87.860 95.110 88.000 96.830 ;
        RECT 87.800 94.790 88.060 95.110 ;
        RECT 87.340 93.090 87.600 93.410 ;
        RECT 87.800 93.090 88.060 93.410 ;
        RECT 82.740 90.710 83.000 91.030 ;
        RECT 86.020 90.970 87.080 91.110 ;
        RECT 82.800 88.990 82.940 90.710 ;
        RECT 85.960 89.010 86.220 89.330 ;
        RECT 82.740 88.670 83.000 88.990 ;
        RECT 86.020 86.950 86.160 89.010 ;
        RECT 85.960 86.630 86.220 86.950 ;
        RECT 86.940 86.270 87.080 90.970 ;
        RECT 87.400 86.270 87.540 93.090 ;
        RECT 87.860 86.610 88.000 93.090 ;
        RECT 89.240 90.690 89.380 99.130 ;
        RECT 89.640 98.530 89.900 98.850 ;
        RECT 89.700 95.110 89.840 98.530 ;
        RECT 90.620 97.230 90.760 101.590 ;
        RECT 91.940 101.250 92.200 101.570 ;
        RECT 90.160 97.090 91.680 97.230 ;
        RECT 90.160 96.470 90.300 97.090 ;
        RECT 90.560 96.490 90.820 96.810 ;
        RECT 90.100 96.150 90.360 96.470 ;
        RECT 89.640 94.790 89.900 95.110 ;
        RECT 90.100 94.790 90.360 95.110 ;
        RECT 89.640 90.710 89.900 91.030 ;
        RECT 89.180 90.370 89.440 90.690 ;
        RECT 89.700 86.950 89.840 90.710 ;
        RECT 90.160 89.185 90.300 94.790 ;
        RECT 90.620 92.390 90.760 96.490 ;
        RECT 90.560 92.070 90.820 92.390 ;
        RECT 91.540 89.670 91.680 97.090 ;
        RECT 91.480 89.350 91.740 89.670 ;
        RECT 90.090 88.815 90.370 89.185 ;
        RECT 90.160 88.310 90.300 88.815 ;
        RECT 90.100 87.990 90.360 88.310 ;
        RECT 89.640 86.630 89.900 86.950 ;
        RECT 87.800 86.290 88.060 86.610 ;
        RECT 86.880 85.950 87.140 86.270 ;
        RECT 87.340 85.950 87.600 86.270 ;
        RECT 92.000 85.930 92.140 101.250 ;
        RECT 92.920 96.810 93.060 110.520 ;
        RECT 93.780 110.430 94.040 110.750 ;
        RECT 93.840 108.370 93.980 110.430 ;
        RECT 95.160 110.090 95.420 110.410 ;
        RECT 95.220 108.710 95.360 110.090 ;
        RECT 95.160 108.390 95.420 108.710 ;
        RECT 93.780 108.050 94.040 108.370 ;
        RECT 95.620 108.050 95.880 108.370 ;
        RECT 95.160 107.710 95.420 108.030 ;
        RECT 93.780 106.690 94.040 107.010 ;
        RECT 93.840 104.290 93.980 106.690 ;
        RECT 94.700 105.330 94.960 105.650 ;
        RECT 93.780 103.970 94.040 104.290 ;
        RECT 93.840 102.250 93.980 103.970 ;
        RECT 93.780 101.930 94.040 102.250 ;
        RECT 93.840 100.550 93.980 101.930 ;
        RECT 94.760 100.630 94.900 105.330 ;
        RECT 95.220 104.290 95.360 107.710 ;
        RECT 95.680 105.310 95.820 108.050 ;
        RECT 95.620 104.990 95.880 105.310 ;
        RECT 95.160 103.970 95.420 104.290 ;
        RECT 93.780 100.230 94.040 100.550 ;
        RECT 94.760 100.490 95.360 100.630 ;
        RECT 94.700 98.530 94.960 98.850 ;
        RECT 94.240 97.510 94.500 97.830 ;
        RECT 92.860 96.490 93.120 96.810 ;
        RECT 92.860 94.790 93.120 95.110 ;
        RECT 92.920 94.090 93.060 94.790 ;
        RECT 93.780 94.110 94.040 94.430 ;
        RECT 92.860 93.770 93.120 94.090 ;
        RECT 92.400 92.070 92.660 92.390 ;
        RECT 92.460 88.650 92.600 92.070 ;
        RECT 93.840 92.050 93.980 94.110 ;
        RECT 93.780 91.730 94.040 92.050 ;
        RECT 93.320 90.710 93.580 91.030 ;
        RECT 92.850 88.815 93.130 89.185 ;
        RECT 93.380 88.990 93.520 90.710 ;
        RECT 94.300 90.690 94.440 97.510 ;
        RECT 94.240 90.370 94.500 90.690 ;
        RECT 92.860 88.670 93.120 88.815 ;
        RECT 93.320 88.670 93.580 88.990 ;
        RECT 94.230 88.815 94.510 89.185 ;
        RECT 94.760 88.990 94.900 98.530 ;
        RECT 95.220 94.090 95.360 100.490 ;
        RECT 96.140 96.810 96.280 150.210 ;
        RECT 96.600 148.150 96.740 181.150 ;
        RECT 97.060 175.350 97.200 181.150 ;
        RECT 97.520 175.430 97.660 202.910 ;
        RECT 98.380 201.890 98.640 202.210 ;
        RECT 98.440 200.170 98.580 201.890 ;
        RECT 98.900 200.850 99.040 202.910 ;
        RECT 99.760 202.230 100.020 202.550 ;
        RECT 98.840 200.530 99.100 200.850 ;
        RECT 99.820 200.170 99.960 202.230 ;
        RECT 100.740 201.190 100.880 204.950 ;
        RECT 102.980 202.570 103.240 202.890 ;
        RECT 100.680 200.870 100.940 201.190 ;
        RECT 98.380 199.850 98.640 200.170 ;
        RECT 99.760 199.850 100.020 200.170 ;
        RECT 97.920 195.430 98.180 195.750 ;
        RECT 97.980 188.950 98.120 195.430 ;
        RECT 99.300 194.070 99.560 194.390 ;
        RECT 99.360 193.030 99.500 194.070 ;
        RECT 101.600 193.730 101.860 194.050 ;
        RECT 99.300 192.710 99.560 193.030 ;
        RECT 99.300 192.030 99.560 192.350 ;
        RECT 98.380 191.010 98.640 191.330 ;
        RECT 98.440 189.290 98.580 191.010 ;
        RECT 98.380 188.970 98.640 189.290 ;
        RECT 98.840 188.970 99.100 189.290 ;
        RECT 99.360 189.030 99.500 192.030 ;
        RECT 99.760 191.690 100.020 192.010 ;
        RECT 99.820 189.970 99.960 191.690 ;
        RECT 99.760 189.650 100.020 189.970 ;
        RECT 100.220 189.310 100.480 189.630 ;
        RECT 101.130 189.455 101.410 189.825 ;
        RECT 100.280 189.030 100.420 189.310 ;
        RECT 101.200 189.290 101.340 189.455 ;
        RECT 97.920 188.630 98.180 188.950 ;
        RECT 98.900 187.590 99.040 188.970 ;
        RECT 99.360 188.890 100.420 189.030 ;
        RECT 101.140 188.970 101.400 189.290 ;
        RECT 101.660 188.950 101.800 193.730 ;
        RECT 103.040 193.030 103.180 202.570 ;
        RECT 103.500 199.830 103.640 204.950 ;
        RECT 104.420 203.230 104.560 207.330 ;
        RECT 106.720 203.230 106.860 207.670 ;
        RECT 107.120 204.950 107.380 205.270 ;
        RECT 107.180 203.910 107.320 204.950 ;
        RECT 107.120 203.590 107.380 203.910 ;
        RECT 104.360 202.910 104.620 203.230 ;
        RECT 106.660 202.910 106.920 203.230 ;
        RECT 103.440 199.510 103.700 199.830 ;
        RECT 102.980 192.710 103.240 193.030 ;
        RECT 102.510 192.175 102.790 192.545 ;
        RECT 102.520 192.030 102.780 192.175 ;
        RECT 102.980 188.970 103.240 189.290 ;
        RECT 98.840 187.270 99.100 187.590 ;
        RECT 98.380 186.590 98.640 186.910 ;
        RECT 98.840 186.820 99.100 186.910 ;
        RECT 99.360 186.820 99.500 188.890 ;
        RECT 100.680 188.630 100.940 188.950 ;
        RECT 101.600 188.630 101.860 188.950 ;
        RECT 100.220 188.290 100.480 188.610 ;
        RECT 98.840 186.680 99.500 186.820 ;
        RECT 98.840 186.590 99.100 186.680 ;
        RECT 97.920 180.810 98.180 181.130 ;
        RECT 97.980 179.430 98.120 180.810 ;
        RECT 97.920 179.110 98.180 179.430 ;
        RECT 98.440 176.030 98.580 186.590 ;
        RECT 99.760 184.550 100.020 184.870 ;
        RECT 99.820 178.750 99.960 184.550 ;
        RECT 100.280 181.130 100.420 188.290 ;
        RECT 100.740 187.500 100.880 188.630 ;
        RECT 102.060 188.290 102.320 188.610 ;
        RECT 102.520 188.290 102.780 188.610 ;
        RECT 101.140 187.500 101.400 187.590 ;
        RECT 100.740 187.360 101.400 187.500 ;
        RECT 100.740 186.570 100.880 187.360 ;
        RECT 101.140 187.270 101.400 187.360 ;
        RECT 102.120 186.910 102.260 188.290 ;
        RECT 102.580 187.250 102.720 188.290 ;
        RECT 102.520 186.930 102.780 187.250 ;
        RECT 101.600 186.590 101.860 186.910 ;
        RECT 102.060 186.590 102.320 186.910 ;
        RECT 100.680 186.250 100.940 186.570 ;
        RECT 101.660 184.870 101.800 186.590 ;
        RECT 103.040 184.870 103.180 188.970 ;
        RECT 101.600 184.550 101.860 184.870 ;
        RECT 102.980 184.550 103.240 184.870 ;
        RECT 101.660 184.170 101.800 184.550 ;
        RECT 103.500 184.190 103.640 199.510 ;
        RECT 106.200 194.070 106.460 194.390 ;
        RECT 103.900 193.730 104.160 194.050 ;
        RECT 103.960 192.690 104.100 193.730 ;
        RECT 103.900 192.370 104.160 192.690 ;
        RECT 106.260 192.350 106.400 194.070 ;
        RECT 106.200 192.030 106.460 192.350 ;
        RECT 107.180 192.010 107.320 203.590 ;
        RECT 108.040 200.190 108.300 200.510 ;
        RECT 108.100 197.790 108.240 200.190 ;
        RECT 108.040 197.470 108.300 197.790 ;
        RECT 108.100 195.150 108.240 197.470 ;
        RECT 108.500 197.130 108.760 197.450 ;
        RECT 107.640 195.010 108.240 195.150 ;
        RECT 107.640 193.030 107.780 195.010 ;
        RECT 108.040 194.410 108.300 194.730 ;
        RECT 107.580 192.710 107.840 193.030 ;
        RECT 103.900 191.690 104.160 192.010 ;
        RECT 104.820 191.690 105.080 192.010 ;
        RECT 105.280 191.690 105.540 192.010 ;
        RECT 107.120 191.690 107.380 192.010 ;
        RECT 103.960 187.590 104.100 191.690 ;
        RECT 104.880 190.310 105.020 191.690 ;
        RECT 104.820 189.990 105.080 190.310 ;
        RECT 105.340 189.145 105.480 191.690 ;
        RECT 106.660 191.010 106.920 191.330 ;
        RECT 105.730 189.455 106.010 189.825 ;
        RECT 105.800 189.290 105.940 189.455 ;
        RECT 106.720 189.290 106.860 191.010 ;
        RECT 107.580 189.310 107.840 189.630 ;
        RECT 105.270 188.775 105.550 189.145 ;
        RECT 105.740 188.970 106.000 189.290 ;
        RECT 106.660 188.970 106.920 189.290 ;
        RECT 105.280 188.290 105.540 188.610 ;
        RECT 105.340 187.590 105.480 188.290 ;
        RECT 103.900 187.270 104.160 187.590 ;
        RECT 105.280 187.270 105.540 187.590 ;
        RECT 106.720 186.570 106.860 188.970 ;
        RECT 106.660 186.250 106.920 186.570 ;
        RECT 107.640 184.190 107.780 189.310 ;
        RECT 108.100 186.910 108.240 194.410 ;
        RECT 108.560 194.050 108.700 197.130 ;
        RECT 114.940 194.070 115.200 194.390 ;
        RECT 108.500 193.730 108.760 194.050 ;
        RECT 108.560 189.970 108.700 193.730 ;
        RECT 115.000 193.030 115.140 194.070 ;
        RECT 114.940 192.710 115.200 193.030 ;
        RECT 120.920 192.030 121.180 192.350 ;
        RECT 108.500 189.650 108.760 189.970 ;
        RECT 117.240 188.970 117.500 189.290 ;
        RECT 110.340 188.290 110.600 188.610 ;
        RECT 110.400 187.250 110.540 188.290 ;
        RECT 110.340 186.930 110.600 187.250 ;
        RECT 108.040 186.590 108.300 186.910 ;
        RECT 108.100 184.190 108.240 186.590 ;
        RECT 117.300 185.890 117.440 188.970 ;
        RECT 118.160 188.630 118.420 188.950 ;
        RECT 117.240 185.570 117.500 185.890 ;
        RECT 118.220 184.870 118.360 188.630 ;
        RECT 120.980 187.590 121.120 192.030 ;
        RECT 124.600 188.970 124.860 189.290 ;
        RECT 125.060 188.970 125.320 189.290 ;
        RECT 122.300 188.290 122.560 188.610 ;
        RECT 120.920 187.270 121.180 187.590 ;
        RECT 120.920 186.250 121.180 186.570 ;
        RECT 114.940 184.550 115.200 184.870 ;
        RECT 118.160 184.550 118.420 184.870 ;
        RECT 101.660 184.030 102.260 184.170 ;
        RECT 102.120 181.470 102.260 184.030 ;
        RECT 103.440 183.870 103.700 184.190 ;
        RECT 107.580 183.870 107.840 184.190 ;
        RECT 108.040 183.870 108.300 184.190 ;
        RECT 102.060 181.150 102.320 181.470 ;
        RECT 100.220 180.810 100.480 181.130 ;
        RECT 103.500 180.790 103.640 183.870 ;
        RECT 106.660 182.850 106.920 183.170 ;
        RECT 106.720 182.150 106.860 182.850 ;
        RECT 106.660 181.830 106.920 182.150 ;
        RECT 107.640 181.130 107.780 183.870 ;
        RECT 108.100 181.810 108.240 183.870 ;
        RECT 108.500 183.190 108.760 183.510 ;
        RECT 108.560 182.150 108.700 183.190 ;
        RECT 108.500 181.830 108.760 182.150 ;
        RECT 111.720 181.830 111.980 182.150 ;
        RECT 108.040 181.490 108.300 181.810 ;
        RECT 107.580 180.810 107.840 181.130 ;
        RECT 103.440 180.470 103.700 180.790 ;
        RECT 102.520 180.130 102.780 180.450 ;
        RECT 102.580 178.750 102.720 180.130 ;
        RECT 103.500 178.750 103.640 180.470 ;
        RECT 99.760 178.430 100.020 178.750 ;
        RECT 102.520 178.430 102.780 178.750 ;
        RECT 103.440 178.430 103.700 178.750 ;
        RECT 99.820 176.030 99.960 178.430 ;
        RECT 101.140 178.090 101.400 178.410 ;
        RECT 110.340 178.090 110.600 178.410 ;
        RECT 110.800 178.090 111.060 178.410 ;
        RECT 98.380 175.710 98.640 176.030 ;
        RECT 99.760 175.710 100.020 176.030 ;
        RECT 97.000 175.030 97.260 175.350 ;
        RECT 97.520 175.290 98.120 175.430 ;
        RECT 97.460 174.690 97.720 175.010 ;
        RECT 97.520 171.270 97.660 174.690 ;
        RECT 97.460 170.950 97.720 171.270 ;
        RECT 97.000 170.270 97.260 170.590 ;
        RECT 97.060 168.550 97.200 170.270 ;
        RECT 97.000 168.230 97.260 168.550 ;
        RECT 97.000 161.090 97.260 161.410 ;
        RECT 97.060 160.050 97.200 161.090 ;
        RECT 97.000 159.730 97.260 160.050 ;
        RECT 97.060 156.990 97.200 159.730 ;
        RECT 97.980 157.670 98.120 175.290 ;
        RECT 98.440 173.990 98.580 175.710 ;
        RECT 98.380 173.670 98.640 173.990 ;
        RECT 101.200 173.310 101.340 178.090 ;
        RECT 107.580 177.410 107.840 177.730 ;
        RECT 108.500 177.410 108.760 177.730 ;
        RECT 105.280 175.370 105.540 175.690 ;
        RECT 102.980 174.690 103.240 175.010 ;
        RECT 103.040 173.310 103.180 174.690 ;
        RECT 98.380 172.990 98.640 173.310 ;
        RECT 101.140 172.990 101.400 173.310 ;
        RECT 102.980 172.990 103.240 173.310 ;
        RECT 98.440 170.250 98.580 172.990 ;
        RECT 100.680 170.270 100.940 170.590 ;
        RECT 105.340 170.370 105.480 175.370 ;
        RECT 105.740 174.690 106.000 175.010 ;
        RECT 105.800 172.970 105.940 174.690 ;
        RECT 105.740 172.650 106.000 172.970 ;
        RECT 106.660 172.650 106.920 172.970 ;
        RECT 98.380 169.930 98.640 170.250 ;
        RECT 99.760 167.210 100.020 167.530 ;
        RECT 99.820 165.150 99.960 167.210 ;
        RECT 100.220 165.510 100.480 165.830 ;
        RECT 98.840 164.830 99.100 165.150 ;
        RECT 99.760 164.830 100.020 165.150 ;
        RECT 98.900 163.110 99.040 164.830 ;
        RECT 98.840 162.790 99.100 163.110 ;
        RECT 98.900 159.710 99.040 162.790 ;
        RECT 99.820 159.905 99.960 164.830 ;
        RECT 98.840 159.390 99.100 159.710 ;
        RECT 99.300 159.390 99.560 159.710 ;
        RECT 99.750 159.535 100.030 159.905 ;
        RECT 100.280 159.710 100.420 165.510 ;
        RECT 100.740 162.090 100.880 170.270 ;
        RECT 104.420 170.230 105.480 170.370 ;
        RECT 103.900 167.550 104.160 167.870 ;
        RECT 103.440 166.870 103.700 167.190 ;
        RECT 101.140 162.110 101.400 162.430 ;
        RECT 100.680 161.770 100.940 162.090 ;
        RECT 100.680 160.070 100.940 160.390 ;
        RECT 99.760 159.390 100.020 159.535 ;
        RECT 100.220 159.390 100.480 159.710 ;
        RECT 99.360 158.690 99.500 159.390 ;
        RECT 100.740 159.030 100.880 160.070 ;
        RECT 100.680 158.710 100.940 159.030 ;
        RECT 99.300 158.370 99.560 158.690 ;
        RECT 97.920 157.350 98.180 157.670 ;
        RECT 97.000 156.670 97.260 156.990 ;
        RECT 97.460 156.330 97.720 156.650 ;
        RECT 97.520 151.890 97.660 156.330 ;
        RECT 101.200 154.270 101.340 162.110 ;
        RECT 102.980 161.770 103.240 162.090 ;
        RECT 103.040 160.390 103.180 161.770 ;
        RECT 102.980 160.070 103.240 160.390 ;
        RECT 101.140 153.950 101.400 154.270 ;
        RECT 101.200 152.230 101.340 153.950 ;
        RECT 101.140 151.910 101.400 152.230 ;
        RECT 97.460 151.570 97.720 151.890 ;
        RECT 97.920 150.890 98.180 151.210 ;
        RECT 97.460 150.210 97.720 150.530 ;
        RECT 97.520 148.490 97.660 150.210 ;
        RECT 97.980 148.490 98.120 150.890 ;
        RECT 98.380 148.510 98.640 148.830 ;
        RECT 101.140 148.510 101.400 148.830 ;
        RECT 102.980 148.510 103.240 148.830 ;
        RECT 97.460 148.170 97.720 148.490 ;
        RECT 97.920 148.170 98.180 148.490 ;
        RECT 96.540 147.830 96.800 148.150 ;
        RECT 97.520 145.770 97.660 148.170 ;
        RECT 97.460 145.450 97.720 145.770 ;
        RECT 98.440 145.090 98.580 148.510 ;
        RECT 98.380 144.770 98.640 145.090 ;
        RECT 98.440 143.390 98.580 144.770 ;
        RECT 101.200 143.390 101.340 148.510 ;
        RECT 97.000 143.070 97.260 143.390 ;
        RECT 98.380 143.070 98.640 143.390 ;
        RECT 101.140 143.070 101.400 143.390 ;
        RECT 97.060 135.910 97.200 143.070 ;
        RECT 101.200 141.350 101.340 143.070 ;
        RECT 101.140 141.030 101.400 141.350 ;
        RECT 102.520 140.690 102.780 141.010 ;
        RECT 98.840 140.010 99.100 140.330 ;
        RECT 98.900 137.950 99.040 140.010 ;
        RECT 101.600 139.330 101.860 139.650 ;
        RECT 101.660 138.290 101.800 139.330 ;
        RECT 101.600 137.970 101.860 138.290 ;
        RECT 97.460 137.630 97.720 137.950 ;
        RECT 98.840 137.630 99.100 137.950 ;
        RECT 99.760 137.630 100.020 137.950 ;
        RECT 97.000 135.590 97.260 135.910 ;
        RECT 96.540 117.570 96.800 117.890 ;
        RECT 96.600 116.530 96.740 117.570 ;
        RECT 96.540 116.210 96.800 116.530 ;
        RECT 96.540 109.410 96.800 109.730 ;
        RECT 96.600 105.220 96.740 109.410 ;
        RECT 97.520 105.990 97.660 137.630 ;
        RECT 98.900 134.890 99.040 137.630 ;
        RECT 99.820 135.570 99.960 137.630 ;
        RECT 102.580 135.910 102.720 140.690 ;
        RECT 103.040 140.330 103.180 148.510 ;
        RECT 102.980 140.010 103.240 140.330 ;
        RECT 102.520 135.590 102.780 135.910 ;
        RECT 99.760 135.310 100.020 135.570 ;
        RECT 99.760 135.250 100.420 135.310 ;
        RECT 99.820 135.170 100.420 135.250 ;
        RECT 98.840 134.570 99.100 134.890 ;
        RECT 99.760 134.570 100.020 134.890 ;
        RECT 98.900 130.130 99.040 134.570 ;
        RECT 98.840 129.810 99.100 130.130 ;
        RECT 98.840 123.690 99.100 124.010 ;
        RECT 98.380 123.010 98.640 123.330 ;
        RECT 98.440 118.230 98.580 123.010 ;
        RECT 98.900 121.290 99.040 123.690 ;
        RECT 98.840 120.970 99.100 121.290 ;
        RECT 98.380 117.910 98.640 118.230 ;
        RECT 99.300 117.570 99.560 117.890 ;
        RECT 99.360 113.130 99.500 117.570 ;
        RECT 99.300 112.810 99.560 113.130 ;
        RECT 97.460 105.670 97.720 105.990 ;
        RECT 97.460 105.220 97.720 105.310 ;
        RECT 96.600 105.080 97.720 105.220 ;
        RECT 97.460 104.990 97.720 105.080 ;
        RECT 96.540 102.270 96.800 102.590 ;
        RECT 96.080 96.490 96.340 96.810 ;
        RECT 95.160 93.770 95.420 94.090 ;
        RECT 95.220 91.710 95.360 93.770 ;
        RECT 95.160 91.390 95.420 91.710 ;
        RECT 95.620 91.280 95.880 91.370 ;
        RECT 96.140 91.280 96.280 96.490 ;
        RECT 96.600 96.130 96.740 102.270 ;
        RECT 97.520 101.910 97.660 104.990 ;
        RECT 98.380 103.970 98.640 104.290 ;
        RECT 98.440 102.590 98.580 103.970 ;
        RECT 98.380 102.270 98.640 102.590 ;
        RECT 97.460 101.590 97.720 101.910 ;
        RECT 99.820 96.470 99.960 134.570 ;
        RECT 100.280 129.790 100.420 135.170 ;
        RECT 101.600 134.570 101.860 134.890 ;
        RECT 100.220 129.470 100.480 129.790 ;
        RECT 101.660 119.250 101.800 134.570 ;
        RECT 102.520 132.080 102.780 132.170 ;
        RECT 103.500 132.080 103.640 166.870 ;
        RECT 103.960 165.490 104.100 167.550 ;
        RECT 104.420 166.850 104.560 170.230 ;
        RECT 105.280 167.210 105.540 167.530 ;
        RECT 105.800 167.270 105.940 172.650 ;
        RECT 106.720 168.550 106.860 172.650 ;
        RECT 107.120 169.250 107.380 169.570 ;
        RECT 107.640 169.425 107.780 177.410 ;
        RECT 108.040 175.710 108.300 176.030 ;
        RECT 108.100 173.310 108.240 175.710 ;
        RECT 108.040 172.990 108.300 173.310 ;
        RECT 108.100 170.590 108.240 172.990 ;
        RECT 108.560 171.270 108.700 177.410 ;
        RECT 110.400 176.710 110.540 178.090 ;
        RECT 110.340 176.390 110.600 176.710 ;
        RECT 110.340 175.710 110.600 176.030 ;
        RECT 108.500 170.950 108.760 171.270 ;
        RECT 108.040 170.270 108.300 170.590 ;
        RECT 106.660 168.230 106.920 168.550 ;
        RECT 107.180 168.460 107.320 169.250 ;
        RECT 107.570 169.055 107.850 169.425 ;
        RECT 108.100 168.745 108.240 170.270 ;
        RECT 107.580 168.460 107.840 168.550 ;
        RECT 107.180 168.320 107.840 168.460 ;
        RECT 108.030 168.375 108.310 168.745 ;
        RECT 107.580 168.230 107.840 168.320 ;
        RECT 108.040 167.950 108.300 168.210 ;
        RECT 107.640 167.890 108.300 167.950 ;
        RECT 107.640 167.810 108.240 167.890 ;
        RECT 104.360 166.530 104.620 166.850 ;
        RECT 105.340 166.705 105.480 167.210 ;
        RECT 105.800 167.130 105.985 167.270 ;
        RECT 105.845 167.100 105.985 167.130 ;
        RECT 105.845 166.960 106.400 167.100 ;
        RECT 105.270 166.335 105.550 166.705 ;
        RECT 105.280 165.510 105.540 165.830 ;
        RECT 103.900 165.170 104.160 165.490 ;
        RECT 105.340 160.390 105.480 165.510 ;
        RECT 106.260 164.550 106.400 166.960 ;
        RECT 107.640 166.850 107.780 167.810 ;
        RECT 108.500 167.550 108.760 167.870 ;
        RECT 108.030 167.015 108.310 167.385 ;
        RECT 107.580 166.530 107.840 166.850 ;
        RECT 108.100 165.150 108.240 167.015 ;
        RECT 108.560 165.490 108.700 167.550 ;
        RECT 110.400 166.705 110.540 175.710 ;
        RECT 110.860 171.270 111.000 178.090 ;
        RECT 111.260 175.710 111.520 176.030 ;
        RECT 110.800 170.950 111.060 171.270 ;
        RECT 111.320 168.550 111.460 175.710 ;
        RECT 111.260 168.230 111.520 168.550 ;
        RECT 110.800 166.870 111.060 167.190 ;
        RECT 110.330 166.335 110.610 166.705 ;
        RECT 108.500 165.170 108.760 165.490 ;
        RECT 108.040 164.830 108.300 165.150 ;
        RECT 110.400 164.810 110.540 166.335 ;
        RECT 106.260 164.410 106.860 164.550 ;
        RECT 110.340 164.490 110.600 164.810 ;
        RECT 106.200 163.810 106.460 164.130 ;
        RECT 105.280 160.070 105.540 160.390 ;
        RECT 106.260 160.050 106.400 163.810 ;
        RECT 106.720 160.390 106.860 164.410 ;
        RECT 108.500 163.810 108.760 164.130 ;
        RECT 107.120 162.450 107.380 162.770 ;
        RECT 106.660 160.070 106.920 160.390 ;
        RECT 106.200 159.730 106.460 160.050 ;
        RECT 106.720 159.710 106.860 160.070 ;
        RECT 107.180 159.710 107.320 162.450 ;
        RECT 108.560 159.710 108.700 163.810 ;
        RECT 110.400 163.470 110.540 164.490 ;
        RECT 109.940 163.330 110.540 163.470 ;
        RECT 109.940 161.410 110.080 163.330 ;
        RECT 110.340 162.790 110.600 163.110 ;
        RECT 109.880 161.090 110.140 161.410 ;
        RECT 110.400 159.710 110.540 162.790 ;
        RECT 106.660 159.390 106.920 159.710 ;
        RECT 107.120 159.390 107.380 159.710 ;
        RECT 108.500 159.390 108.760 159.710 ;
        RECT 110.340 159.390 110.600 159.710 ;
        RECT 109.880 156.330 110.140 156.650 ;
        RECT 109.940 154.950 110.080 156.330 ;
        RECT 109.880 154.630 110.140 154.950 ;
        RECT 108.030 152.055 108.310 152.425 ;
        RECT 108.040 151.910 108.300 152.055 ;
        RECT 109.940 151.890 110.080 154.630 ;
        RECT 109.880 151.570 110.140 151.890 ;
        RECT 110.860 151.550 111.000 166.870 ;
        RECT 111.320 165.490 111.460 168.230 ;
        RECT 111.260 165.170 111.520 165.490 ;
        RECT 110.800 151.230 111.060 151.550 ;
        RECT 104.360 150.550 104.620 150.870 ;
        RECT 108.500 150.550 108.760 150.870 ;
        RECT 104.420 149.510 104.560 150.550 ;
        RECT 104.360 149.190 104.620 149.510 ;
        RECT 108.040 148.850 108.300 149.170 ;
        RECT 106.200 148.510 106.460 148.830 ;
        RECT 103.900 147.490 104.160 147.810 ;
        RECT 103.960 143.730 104.100 147.490 ;
        RECT 106.260 146.790 106.400 148.510 ;
        RECT 108.100 146.790 108.240 148.850 ;
        RECT 108.560 148.490 108.700 150.550 ;
        RECT 108.500 148.170 108.760 148.490 ;
        RECT 111.780 146.790 111.920 181.830 ;
        RECT 115.000 181.470 115.140 184.550 ;
        RECT 120.980 184.190 121.120 186.250 ;
        RECT 120.920 183.870 121.180 184.190 ;
        RECT 118.620 183.530 118.880 183.850 ;
        RECT 116.320 182.850 116.580 183.170 ;
        RECT 116.380 182.150 116.520 182.850 ;
        RECT 118.680 182.150 118.820 183.530 ;
        RECT 120.000 182.850 120.260 183.170 ;
        RECT 116.320 181.830 116.580 182.150 ;
        RECT 118.620 181.830 118.880 182.150 ;
        RECT 114.940 181.150 115.200 181.470 ;
        RECT 117.240 181.150 117.500 181.470 ;
        RECT 116.320 180.470 116.580 180.790 ;
        RECT 115.860 177.750 116.120 178.070 ;
        RECT 112.180 177.410 112.440 177.730 ;
        RECT 112.240 167.870 112.380 177.410 ;
        RECT 114.020 176.390 114.280 176.710 ;
        RECT 114.080 172.290 114.220 176.390 ;
        RECT 115.400 175.030 115.660 175.350 ;
        RECT 115.460 173.990 115.600 175.030 ;
        RECT 115.400 173.670 115.660 173.990 ;
        RECT 114.480 172.650 114.740 172.970 ;
        RECT 114.020 171.970 114.280 172.290 ;
        RECT 114.080 168.210 114.220 171.970 ;
        RECT 114.020 167.890 114.280 168.210 ;
        RECT 112.180 167.550 112.440 167.870 ;
        RECT 114.540 166.850 114.680 172.650 ;
        RECT 114.940 170.950 115.200 171.270 ;
        RECT 115.000 167.530 115.140 170.950 ;
        RECT 115.460 170.590 115.600 173.670 ;
        RECT 115.400 170.270 115.660 170.590 ;
        RECT 114.940 167.210 115.200 167.530 ;
        RECT 114.480 166.530 114.740 166.850 ;
        RECT 113.100 164.830 113.360 165.150 ;
        RECT 112.640 164.490 112.900 164.810 ;
        RECT 112.700 163.110 112.840 164.490 ;
        RECT 113.160 163.110 113.300 164.830 ;
        RECT 115.000 164.810 115.140 167.210 ;
        RECT 115.400 165.170 115.660 165.490 ;
        RECT 114.940 164.490 115.200 164.810 ;
        RECT 112.640 162.790 112.900 163.110 ;
        RECT 113.100 162.790 113.360 163.110 ;
        RECT 112.700 162.430 112.840 162.790 ;
        RECT 112.640 162.110 112.900 162.430 ;
        RECT 113.160 159.710 113.300 162.790 ;
        RECT 115.000 162.770 115.140 164.490 ;
        RECT 114.940 162.450 115.200 162.770 ;
        RECT 115.460 162.090 115.600 165.170 ;
        RECT 115.400 161.770 115.660 162.090 ;
        RECT 113.100 159.390 113.360 159.710 ;
        RECT 115.460 159.370 115.600 161.770 ;
        RECT 115.920 160.390 116.060 177.750 ;
        RECT 116.380 167.190 116.520 180.470 ;
        RECT 116.320 166.870 116.580 167.190 ;
        RECT 115.860 160.070 116.120 160.390 ;
        RECT 115.400 159.050 115.660 159.370 ;
        RECT 113.560 158.710 113.820 159.030 ;
        RECT 113.620 157.670 113.760 158.710 ;
        RECT 115.860 158.370 116.120 158.690 ;
        RECT 113.560 157.350 113.820 157.670 ;
        RECT 112.630 156.815 112.910 157.185 ;
        RECT 112.700 154.610 112.840 156.815 ;
        RECT 115.920 156.650 116.060 158.370 ;
        RECT 115.860 156.330 116.120 156.650 ;
        RECT 116.320 155.990 116.580 156.310 ;
        RECT 114.020 155.650 114.280 155.970 ;
        RECT 116.380 155.825 116.520 155.990 ;
        RECT 112.640 154.290 112.900 154.610 ;
        RECT 114.080 154.270 114.220 155.650 ;
        RECT 116.310 155.455 116.590 155.825 ;
        RECT 117.300 154.350 117.440 181.150 ;
        RECT 118.680 179.430 118.820 181.830 ;
        RECT 118.620 179.110 118.880 179.430 ;
        RECT 117.700 170.270 117.960 170.590 ;
        RECT 118.610 170.415 118.890 170.785 ;
        RECT 118.620 170.270 118.880 170.415 ;
        RECT 117.760 167.870 117.900 170.270 ;
        RECT 118.160 169.590 118.420 169.910 ;
        RECT 117.700 167.550 117.960 167.870 ;
        RECT 117.760 165.490 117.900 167.550 ;
        RECT 118.220 167.270 118.360 169.590 ;
        RECT 118.680 168.210 118.820 170.270 ;
        RECT 119.530 169.735 119.810 170.105 ;
        RECT 119.600 168.550 119.740 169.735 ;
        RECT 119.540 168.230 119.800 168.550 ;
        RECT 118.620 167.890 118.880 168.210 ;
        RECT 118.620 167.270 118.880 167.530 ;
        RECT 118.220 167.210 118.880 167.270 ;
        RECT 119.080 167.210 119.340 167.530 ;
        RECT 118.220 167.130 118.820 167.210 ;
        RECT 117.700 165.170 117.960 165.490 ;
        RECT 117.700 164.490 117.960 164.810 ;
        RECT 117.760 157.330 117.900 164.490 ;
        RECT 118.160 163.810 118.420 164.130 ;
        RECT 118.220 162.090 118.360 163.810 ;
        RECT 118.680 162.510 118.820 167.130 ;
        RECT 119.140 163.110 119.280 167.210 ;
        RECT 119.080 162.790 119.340 163.110 ;
        RECT 119.540 162.790 119.800 163.110 ;
        RECT 119.600 162.510 119.740 162.790 ;
        RECT 118.680 162.370 119.740 162.510 ;
        RECT 118.160 161.770 118.420 162.090 ;
        RECT 118.220 160.390 118.360 161.770 ;
        RECT 118.680 161.410 118.820 162.370 ;
        RECT 118.620 161.090 118.880 161.410 ;
        RECT 118.160 160.070 118.420 160.390 ;
        RECT 118.680 159.710 118.820 161.090 ;
        RECT 118.620 159.390 118.880 159.710 ;
        RECT 119.080 159.390 119.340 159.710 ;
        RECT 118.160 158.370 118.420 158.690 ;
        RECT 117.700 157.010 117.960 157.330 ;
        RECT 117.700 156.330 117.960 156.650 ;
        RECT 117.760 154.950 117.900 156.330 ;
        RECT 117.700 154.630 117.960 154.950 ;
        RECT 114.020 153.950 114.280 154.270 ;
        RECT 116.320 153.950 116.580 154.270 ;
        RECT 117.300 154.210 117.900 154.350 ;
        RECT 115.860 153.610 116.120 153.930 ;
        RECT 116.380 153.785 116.520 153.950 ;
        RECT 112.180 153.270 112.440 153.590 ;
        RECT 112.240 151.210 112.380 153.270 ;
        RECT 115.400 152.930 115.660 153.250 ;
        RECT 112.640 151.230 112.900 151.550 ;
        RECT 112.180 150.890 112.440 151.210 ;
        RECT 106.200 146.470 106.460 146.790 ;
        RECT 108.040 146.470 108.300 146.790 ;
        RECT 111.720 146.470 111.980 146.790 ;
        RECT 112.180 145.450 112.440 145.770 ;
        RECT 112.240 143.730 112.380 145.450 ;
        RECT 103.900 143.410 104.160 143.730 ;
        RECT 112.180 143.410 112.440 143.730 ;
        RECT 102.520 131.940 103.640 132.080 ;
        RECT 102.520 131.850 102.780 131.940 ;
        RECT 102.580 127.750 102.720 131.850 ;
        RECT 103.960 131.830 104.100 143.410 ;
        RECT 104.820 143.070 105.080 143.390 ;
        RECT 104.880 138.630 105.020 143.070 ;
        RECT 112.240 143.050 112.380 143.410 ;
        RECT 109.420 142.730 109.680 143.050 ;
        RECT 112.180 142.730 112.440 143.050 ;
        RECT 106.200 140.690 106.460 141.010 ;
        RECT 104.820 138.310 105.080 138.630 ;
        RECT 105.740 138.310 106.000 138.630 ;
        RECT 105.800 137.950 105.940 138.310 ;
        RECT 105.740 137.630 106.000 137.950 ;
        RECT 105.800 135.230 105.940 137.630 ;
        RECT 106.260 135.910 106.400 140.690 ;
        RECT 106.660 139.330 106.920 139.650 ;
        RECT 106.720 138.290 106.860 139.330 ;
        RECT 106.660 137.970 106.920 138.290 ;
        RECT 109.480 137.950 109.620 142.730 ;
        RECT 109.420 137.630 109.680 137.950 ;
        RECT 106.200 135.590 106.460 135.910 ;
        RECT 105.740 134.910 106.000 135.230 ;
        RECT 105.280 132.870 105.540 133.190 ;
        RECT 104.360 132.530 104.620 132.850 ;
        RECT 103.900 131.510 104.160 131.830 ;
        RECT 103.960 130.470 104.100 131.510 ;
        RECT 103.900 130.150 104.160 130.470 ;
        RECT 103.440 129.810 103.700 130.130 ;
        RECT 102.520 127.430 102.780 127.750 ;
        RECT 103.500 124.350 103.640 129.810 ;
        RECT 104.420 129.450 104.560 132.530 ;
        RECT 104.360 129.130 104.620 129.450 ;
        RECT 104.420 124.350 104.560 129.130 ;
        RECT 104.820 128.450 105.080 128.770 ;
        RECT 104.880 127.410 105.020 128.450 ;
        RECT 104.820 127.090 105.080 127.410 ;
        RECT 103.440 124.030 103.700 124.350 ;
        RECT 104.360 124.030 104.620 124.350 ;
        RECT 103.500 122.310 103.640 124.030 ;
        RECT 103.440 121.990 103.700 122.310 ;
        RECT 102.520 120.290 102.780 120.610 ;
        RECT 101.600 118.930 101.860 119.250 ;
        RECT 102.580 118.230 102.720 120.290 ;
        RECT 103.500 118.910 103.640 121.990 ;
        RECT 104.420 121.970 104.560 124.030 ;
        RECT 104.360 121.650 104.620 121.970 ;
        RECT 103.440 118.590 103.700 118.910 ;
        RECT 102.060 117.910 102.320 118.230 ;
        RECT 102.520 117.910 102.780 118.230 ;
        RECT 102.120 116.870 102.260 117.910 ;
        RECT 103.900 117.570 104.160 117.890 ;
        RECT 102.060 116.550 102.320 116.870 ;
        RECT 101.600 114.850 101.860 115.170 ;
        RECT 101.660 111.430 101.800 114.850 ;
        RECT 102.120 113.130 102.260 116.550 ;
        RECT 103.960 116.190 104.100 117.570 ;
        RECT 104.420 116.530 104.560 121.650 ;
        RECT 104.360 116.210 104.620 116.530 ;
        RECT 103.900 115.870 104.160 116.190 ;
        RECT 103.960 113.130 104.100 115.870 ;
        RECT 104.420 113.130 104.560 116.210 ;
        RECT 102.060 112.810 102.320 113.130 ;
        RECT 103.900 112.810 104.160 113.130 ;
        RECT 104.360 112.810 104.620 113.130 ;
        RECT 101.600 111.110 101.860 111.430 ;
        RECT 102.120 110.830 102.260 112.810 ;
        RECT 102.120 110.750 102.720 110.830 ;
        RECT 103.960 110.750 104.100 112.810 ;
        RECT 104.420 111.090 104.560 112.810 ;
        RECT 105.340 111.430 105.480 132.870 ;
        RECT 109.420 132.190 109.680 132.510 ;
        RECT 107.120 131.170 107.380 131.490 ;
        RECT 108.500 131.170 108.760 131.490 ;
        RECT 107.180 129.790 107.320 131.170 ;
        RECT 107.120 129.470 107.380 129.790 ;
        RECT 105.740 129.130 106.000 129.450 ;
        RECT 105.800 114.150 105.940 129.130 ;
        RECT 108.560 127.410 108.700 131.170 ;
        RECT 108.500 127.090 108.760 127.410 ;
        RECT 107.120 121.990 107.380 122.310 ;
        RECT 107.180 121.630 107.320 121.990 ;
        RECT 109.480 121.970 109.620 132.190 ;
        RECT 110.340 131.850 110.600 132.170 ;
        RECT 110.400 130.470 110.540 131.850 ;
        RECT 110.340 130.150 110.600 130.470 ;
        RECT 112.700 129.790 112.840 151.230 ;
        RECT 115.460 151.210 115.600 152.930 ;
        RECT 115.920 152.230 116.060 153.610 ;
        RECT 116.310 153.415 116.590 153.785 ;
        RECT 115.860 151.910 116.120 152.230 ;
        RECT 116.780 151.570 117.040 151.890 ;
        RECT 115.400 150.890 115.660 151.210 ;
        RECT 114.940 149.190 115.200 149.510 ;
        RECT 115.000 148.490 115.140 149.190 ;
        RECT 115.460 148.830 115.600 150.890 ;
        RECT 115.400 148.510 115.660 148.830 ;
        RECT 114.940 148.170 115.200 148.490 ;
        RECT 115.460 148.230 115.600 148.510 ;
        RECT 115.460 148.090 116.060 148.230 ;
        RECT 115.920 147.810 116.060 148.090 ;
        RECT 114.940 147.490 115.200 147.810 ;
        RECT 115.400 147.490 115.660 147.810 ;
        RECT 115.860 147.490 116.120 147.810 ;
        RECT 115.000 146.450 115.140 147.490 ;
        RECT 114.940 146.130 115.200 146.450 ;
        RECT 115.460 145.770 115.600 147.490 ;
        RECT 116.840 146.110 116.980 151.570 ;
        RECT 117.240 150.210 117.500 150.530 ;
        RECT 117.300 148.830 117.440 150.210 ;
        RECT 117.240 148.510 117.500 148.830 ;
        RECT 117.240 147.830 117.500 148.150 ;
        RECT 116.780 145.790 117.040 146.110 ;
        RECT 115.400 145.450 115.660 145.770 ;
        RECT 115.860 144.770 116.120 145.090 ;
        RECT 115.920 142.905 116.060 144.770 ;
        RECT 117.300 143.390 117.440 147.830 ;
        RECT 117.240 143.070 117.500 143.390 ;
        RECT 115.850 142.535 116.130 142.905 ;
        RECT 114.940 134.910 115.200 135.230 ;
        RECT 114.020 133.890 114.280 134.210 ;
        RECT 113.560 132.190 113.820 132.510 ;
        RECT 112.640 129.470 112.900 129.790 ;
        RECT 111.720 129.130 111.980 129.450 ;
        RECT 111.780 127.410 111.920 129.130 ;
        RECT 112.700 127.750 112.840 129.470 ;
        RECT 112.640 127.430 112.900 127.750 ;
        RECT 111.720 127.090 111.980 127.410 ;
        RECT 111.780 124.010 111.920 127.090 ;
        RECT 113.620 125.030 113.760 132.190 ;
        RECT 113.560 124.710 113.820 125.030 ;
        RECT 111.720 123.690 111.980 124.010 ;
        RECT 109.420 121.650 109.680 121.970 ;
        RECT 106.660 121.310 106.920 121.630 ;
        RECT 107.120 121.310 107.380 121.630 ;
        RECT 108.040 121.310 108.300 121.630 ;
        RECT 111.250 121.455 111.530 121.825 ;
        RECT 111.780 121.630 111.920 123.690 ;
        RECT 105.740 113.830 106.000 114.150 ;
        RECT 105.280 111.110 105.540 111.430 ;
        RECT 104.360 110.770 104.620 111.090 ;
        RECT 105.340 110.830 105.480 111.110 ;
        RECT 101.600 110.430 101.860 110.750 ;
        RECT 102.120 110.690 102.780 110.750 ;
        RECT 102.520 110.430 102.780 110.690 ;
        RECT 103.900 110.430 104.160 110.750 ;
        RECT 100.680 107.370 100.940 107.690 ;
        RECT 101.140 107.370 101.400 107.690 ;
        RECT 100.740 104.630 100.880 107.370 ;
        RECT 101.200 105.990 101.340 107.370 ;
        RECT 101.660 105.990 101.800 110.430 ;
        RECT 104.420 110.070 104.560 110.770 ;
        RECT 104.880 110.690 105.480 110.830 ;
        RECT 104.360 109.750 104.620 110.070 ;
        RECT 104.880 107.690 105.020 110.690 ;
        RECT 105.280 110.090 105.540 110.410 ;
        RECT 106.200 110.090 106.460 110.410 ;
        RECT 104.820 107.370 105.080 107.690 ;
        RECT 103.440 106.690 103.700 107.010 ;
        RECT 101.140 105.670 101.400 105.990 ;
        RECT 101.600 105.670 101.860 105.990 ;
        RECT 101.660 105.310 101.800 105.670 ;
        RECT 101.600 104.990 101.860 105.310 ;
        RECT 102.980 104.990 103.240 105.310 ;
        RECT 100.680 104.310 100.940 104.630 ;
        RECT 103.040 103.270 103.180 104.990 ;
        RECT 102.980 102.950 103.240 103.270 ;
        RECT 103.500 102.930 103.640 106.690 ;
        RECT 105.340 105.310 105.480 110.090 ;
        RECT 106.260 108.710 106.400 110.090 ;
        RECT 106.200 108.390 106.460 108.710 ;
        RECT 105.280 104.990 105.540 105.310 ;
        RECT 103.440 102.610 103.700 102.930 ;
        RECT 101.140 102.270 101.400 102.590 ;
        RECT 99.760 96.150 100.020 96.470 ;
        RECT 96.540 95.810 96.800 96.130 ;
        RECT 99.300 95.810 99.560 96.130 ;
        RECT 95.620 91.140 96.280 91.280 ;
        RECT 95.620 91.050 95.880 91.140 ;
        RECT 99.360 88.990 99.500 95.810 ;
        RECT 101.200 94.430 101.340 102.270 ;
        RECT 103.900 99.210 104.160 99.530 ;
        RECT 103.440 96.830 103.700 97.150 ;
        RECT 102.060 95.810 102.320 96.130 ;
        RECT 101.140 94.110 101.400 94.430 ;
        RECT 92.400 88.390 92.660 88.650 ;
        RECT 93.780 88.390 94.040 88.650 ;
        RECT 92.400 88.330 94.040 88.390 ;
        RECT 92.460 88.250 93.980 88.330 ;
        RECT 94.300 85.930 94.440 88.815 ;
        RECT 94.700 88.670 94.960 88.990 ;
        RECT 99.300 88.670 99.560 88.990 ;
        RECT 97.460 88.330 97.720 88.650 ;
        RECT 100.680 88.560 100.940 88.650 ;
        RECT 101.200 88.560 101.340 94.110 ;
        RECT 101.600 90.710 101.860 91.030 ;
        RECT 101.660 89.670 101.800 90.710 ;
        RECT 101.600 89.350 101.860 89.670 ;
        RECT 100.680 88.420 101.340 88.560 ;
        RECT 100.680 88.330 100.940 88.420 ;
        RECT 95.160 87.650 95.420 87.970 ;
        RECT 95.220 86.610 95.360 87.650 ;
        RECT 95.160 86.290 95.420 86.610 ;
        RECT 95.620 86.290 95.880 86.610 ;
        RECT 71.240 85.610 71.500 85.930 ;
        RECT 73.540 85.610 73.800 85.930 ;
        RECT 77.680 85.610 77.940 85.930 ;
        RECT 78.140 85.610 78.400 85.930 ;
        RECT 79.980 85.610 80.240 85.930 ;
        RECT 91.940 85.610 92.200 85.930 ;
        RECT 94.240 85.610 94.500 85.930 ;
        RECT 89.180 85.270 89.440 85.590 ;
        RECT 92.400 85.270 92.660 85.590 ;
        RECT 73.080 84.930 73.340 85.250 ;
        RECT 76.300 84.930 76.560 85.250 ;
        RECT 79.520 84.930 79.780 85.250 ;
        RECT 82.740 84.930 83.000 85.250 ;
        RECT 85.960 84.930 86.220 85.250 ;
        RECT 73.140 77.700 73.280 84.930 ;
        RECT 76.360 77.700 76.500 84.930 ;
        RECT 79.580 77.700 79.720 84.930 ;
        RECT 82.800 77.700 82.940 84.930 ;
        RECT 86.020 77.700 86.160 84.930 ;
        RECT 89.240 77.700 89.380 85.270 ;
        RECT 92.460 77.700 92.600 85.270 ;
        RECT 95.680 77.700 95.820 86.290 ;
        RECT 97.520 85.930 97.660 88.330 ;
        RECT 102.120 88.310 102.260 95.810 ;
        RECT 103.500 95.110 103.640 96.830 ;
        RECT 103.960 96.470 104.100 99.210 ;
        RECT 103.900 96.150 104.160 96.470 ;
        RECT 103.960 95.110 104.100 96.150 ;
        RECT 104.360 95.810 104.620 96.130 ;
        RECT 103.440 94.790 103.700 95.110 ;
        RECT 103.900 94.790 104.160 95.110 ;
        RECT 102.980 93.090 103.240 93.410 ;
        RECT 103.040 91.710 103.180 93.090 ;
        RECT 104.420 92.390 104.560 95.810 ;
        RECT 104.360 92.070 104.620 92.390 ;
        RECT 102.980 91.390 103.240 91.710 ;
        RECT 102.060 87.990 102.320 88.310 ;
        RECT 103.040 85.930 103.180 91.390 ;
        RECT 104.420 91.370 104.560 92.070 ;
        RECT 105.340 92.050 105.480 104.990 ;
        RECT 105.740 96.830 106.000 97.150 ;
        RECT 105.800 94.430 105.940 96.830 ;
        RECT 105.740 94.110 106.000 94.430 ;
        RECT 106.720 92.390 106.860 121.310 ;
        RECT 107.180 115.590 107.320 121.310 ;
        RECT 108.100 120.610 108.240 121.310 ;
        RECT 111.320 121.290 111.460 121.455 ;
        RECT 111.720 121.310 111.980 121.630 ;
        RECT 112.180 121.310 112.440 121.630 ;
        RECT 111.260 120.970 111.520 121.290 ;
        RECT 108.040 120.290 108.300 120.610 ;
        RECT 108.100 118.910 108.240 120.290 ;
        RECT 112.240 119.590 112.380 121.310 ;
        RECT 112.180 119.270 112.440 119.590 ;
        RECT 108.040 118.590 108.300 118.910 ;
        RECT 108.960 117.910 109.220 118.230 ;
        RECT 113.550 118.055 113.830 118.425 ;
        RECT 113.560 117.910 113.820 118.055 ;
        RECT 108.490 115.590 108.770 115.705 ;
        RECT 107.180 115.450 108.770 115.590 ;
        RECT 108.490 115.335 108.770 115.450 ;
        RECT 108.560 113.470 108.700 115.335 ;
        RECT 108.500 113.150 108.760 113.470 ;
        RECT 109.020 111.090 109.160 117.910 ;
        RECT 113.620 113.550 113.760 117.910 ;
        RECT 114.080 115.590 114.220 133.890 ;
        RECT 114.480 129.020 114.740 129.110 ;
        RECT 115.000 129.020 115.140 134.910 ;
        RECT 114.480 128.880 115.140 129.020 ;
        RECT 114.480 128.790 114.740 128.880 ;
        RECT 115.000 118.910 115.140 128.880 ;
        RECT 115.400 126.070 115.660 126.390 ;
        RECT 115.460 125.030 115.600 126.070 ;
        RECT 115.400 124.710 115.660 125.030 ;
        RECT 115.460 118.910 115.600 124.710 ;
        RECT 114.940 118.590 115.200 118.910 ;
        RECT 115.400 118.590 115.660 118.910 ;
        RECT 115.000 116.190 115.140 118.590 ;
        RECT 115.920 116.870 116.060 142.535 ;
        RECT 117.760 137.950 117.900 154.210 ;
        RECT 118.220 148.830 118.360 158.370 ;
        RECT 118.680 157.330 118.820 159.390 ;
        RECT 118.620 157.010 118.880 157.330 ;
        RECT 119.140 157.185 119.280 159.390 ;
        RECT 119.070 156.815 119.350 157.185 ;
        RECT 118.620 156.330 118.880 156.650 ;
        RECT 118.680 154.270 118.820 156.330 ;
        RECT 119.080 155.650 119.340 155.970 ;
        RECT 118.620 153.950 118.880 154.270 ;
        RECT 118.680 152.230 118.820 153.950 ;
        RECT 118.620 151.910 118.880 152.230 ;
        RECT 119.140 151.745 119.280 155.650 ;
        RECT 119.540 154.290 119.800 154.610 ;
        RECT 119.070 151.375 119.350 151.745 ;
        RECT 119.600 151.210 119.740 154.290 ;
        RECT 119.540 150.890 119.800 151.210 ;
        RECT 118.160 148.510 118.420 148.830 ;
        RECT 118.620 148.510 118.880 148.830 ;
        RECT 118.220 147.810 118.360 148.510 ;
        RECT 118.160 147.490 118.420 147.810 ;
        RECT 118.220 145.430 118.360 147.490 ;
        RECT 118.160 145.110 118.420 145.430 ;
        RECT 118.680 141.010 118.820 148.510 ;
        RECT 119.540 148.170 119.800 148.490 ;
        RECT 119.600 146.790 119.740 148.170 ;
        RECT 119.540 146.470 119.800 146.790 ;
        RECT 119.080 145.450 119.340 145.770 ;
        RECT 119.140 144.070 119.280 145.450 ;
        RECT 119.080 143.750 119.340 144.070 ;
        RECT 118.620 140.690 118.880 141.010 ;
        RECT 119.540 140.010 119.800 140.330 ;
        RECT 117.700 137.630 117.960 137.950 ;
        RECT 116.320 136.610 116.580 136.930 ;
        RECT 117.700 136.610 117.960 136.930 ;
        RECT 116.380 134.550 116.520 136.610 ;
        RECT 116.320 134.230 116.580 134.550 ;
        RECT 117.760 132.510 117.900 136.610 ;
        RECT 117.700 132.190 117.960 132.510 ;
        RECT 118.620 131.510 118.880 131.830 ;
        RECT 116.780 128.790 117.040 129.110 ;
        RECT 116.840 127.750 116.980 128.790 ;
        RECT 116.780 127.430 117.040 127.750 ;
        RECT 118.680 127.070 118.820 131.510 ;
        RECT 117.700 126.750 117.960 127.070 ;
        RECT 118.620 126.750 118.880 127.070 ;
        RECT 117.760 119.590 117.900 126.750 ;
        RECT 118.680 124.350 118.820 126.750 ;
        RECT 119.600 126.050 119.740 140.010 ;
        RECT 120.060 130.470 120.200 182.850 ;
        RECT 120.980 180.790 121.120 183.870 ;
        RECT 120.920 180.470 121.180 180.790 ;
        RECT 122.360 178.410 122.500 188.290 ;
        RECT 123.680 186.930 123.940 187.250 ;
        RECT 123.740 181.810 123.880 186.930 ;
        RECT 123.680 181.490 123.940 181.810 ;
        RECT 123.740 178.750 123.880 181.490 ;
        RECT 124.140 181.150 124.400 181.470 ;
        RECT 124.200 179.430 124.340 181.150 ;
        RECT 124.140 179.110 124.400 179.430 ;
        RECT 123.680 178.430 123.940 178.750 ;
        RECT 122.300 178.090 122.560 178.410 ;
        RECT 123.680 175.370 123.940 175.690 ;
        RECT 123.740 173.990 123.880 175.370 ;
        RECT 123.680 173.670 123.940 173.990 ;
        RECT 123.680 172.650 123.940 172.970 ;
        RECT 123.740 168.065 123.880 172.650 ;
        RECT 124.140 171.970 124.400 172.290 ;
        RECT 120.450 167.695 120.730 168.065 ;
        RECT 123.670 167.695 123.950 168.065 ;
        RECT 124.200 167.870 124.340 171.970 ;
        RECT 120.520 162.770 120.660 167.695 ;
        RECT 124.140 167.550 124.400 167.870 ;
        RECT 121.840 166.870 122.100 167.190 ;
        RECT 121.900 165.490 122.040 166.870 ;
        RECT 122.760 166.530 123.020 166.850 ;
        RECT 121.840 165.170 122.100 165.490 ;
        RECT 120.460 162.680 120.720 162.770 ;
        RECT 120.460 162.540 121.580 162.680 ;
        RECT 120.460 162.450 120.720 162.540 ;
        RECT 120.460 161.770 120.720 162.090 ;
        RECT 121.440 161.830 121.580 162.540 ;
        RECT 121.900 162.510 122.040 165.170 ;
        RECT 121.900 162.370 122.500 162.510 ;
        RECT 122.360 162.090 122.500 162.370 ;
        RECT 120.520 159.710 120.660 161.770 ;
        RECT 121.440 161.690 122.040 161.830 ;
        RECT 122.300 161.770 122.560 162.090 ;
        RECT 121.380 161.090 121.640 161.410 ;
        RECT 120.460 159.390 120.720 159.710 ;
        RECT 120.520 156.650 120.660 159.390 ;
        RECT 121.440 159.110 121.580 161.090 ;
        RECT 120.980 158.970 121.580 159.110 ;
        RECT 120.460 156.330 120.720 156.650 ;
        RECT 120.450 153.415 120.730 153.785 ;
        RECT 120.520 148.830 120.660 153.415 ;
        RECT 120.460 148.510 120.720 148.830 ;
        RECT 120.980 146.450 121.120 158.970 ;
        RECT 121.380 158.545 121.640 158.690 ;
        RECT 121.370 158.175 121.650 158.545 ;
        RECT 121.440 154.270 121.580 158.175 ;
        RECT 121.380 153.950 121.640 154.270 ;
        RECT 121.440 153.590 121.580 153.950 ;
        RECT 121.380 153.270 121.640 153.590 ;
        RECT 121.440 149.025 121.580 153.270 ;
        RECT 121.900 151.210 122.040 161.690 ;
        RECT 122.300 153.950 122.560 154.270 ;
        RECT 121.840 150.890 122.100 151.210 ;
        RECT 122.360 150.385 122.500 153.950 ;
        RECT 122.820 152.990 122.960 166.530 ;
        RECT 123.680 165.510 123.940 165.830 ;
        RECT 123.220 164.830 123.480 165.150 ;
        RECT 123.280 161.410 123.420 164.830 ;
        RECT 123.740 162.770 123.880 165.510 ;
        RECT 124.200 164.130 124.340 167.550 ;
        RECT 124.660 166.850 124.800 188.970 ;
        RECT 125.120 184.870 125.260 188.970 ;
        RECT 126.900 188.630 127.160 188.950 ;
        RECT 125.520 186.590 125.780 186.910 ;
        RECT 125.060 184.550 125.320 184.870 ;
        RECT 125.580 184.170 125.720 186.590 ;
        RECT 125.120 184.030 125.720 184.170 ;
        RECT 124.600 166.530 124.860 166.850 ;
        RECT 124.140 163.810 124.400 164.130 ;
        RECT 123.680 162.450 123.940 162.770 ;
        RECT 123.220 161.090 123.480 161.410 ;
        RECT 123.280 160.050 123.420 161.090 ;
        RECT 123.220 159.730 123.480 160.050 ;
        RECT 123.740 158.690 123.880 162.450 ;
        RECT 124.130 162.255 124.410 162.625 ;
        RECT 124.660 162.430 124.800 166.530 ;
        RECT 124.200 162.090 124.340 162.255 ;
        RECT 124.600 162.110 124.860 162.430 ;
        RECT 124.140 161.770 124.400 162.090 ;
        RECT 124.660 159.370 124.800 162.110 ;
        RECT 124.600 159.050 124.860 159.370 ;
        RECT 123.680 158.370 123.940 158.690 ;
        RECT 124.140 157.350 124.400 157.670 ;
        RECT 123.680 156.330 123.940 156.650 ;
        RECT 123.740 154.270 123.880 156.330 ;
        RECT 123.680 153.950 123.940 154.270 ;
        RECT 123.740 153.250 123.880 153.950 ;
        RECT 122.820 152.850 123.420 152.990 ;
        RECT 123.680 152.930 123.940 153.250 ;
        RECT 122.290 150.015 122.570 150.385 ;
        RECT 122.760 150.210 123.020 150.530 ;
        RECT 121.370 148.655 121.650 149.025 ;
        RECT 122.820 148.910 122.960 150.210 ;
        RECT 123.280 149.510 123.420 152.850 ;
        RECT 124.200 151.550 124.340 157.350 ;
        RECT 124.660 156.310 124.800 159.050 ;
        RECT 124.600 155.990 124.860 156.310 ;
        RECT 124.600 152.930 124.860 153.250 ;
        RECT 124.140 151.230 124.400 151.550 ;
        RECT 124.200 150.530 124.340 151.230 ;
        RECT 124.140 150.210 124.400 150.530 ;
        RECT 123.220 149.190 123.480 149.510 ;
        RECT 122.360 148.770 122.960 148.910 ;
        RECT 123.280 148.910 123.420 149.190 ;
        RECT 123.280 148.830 124.340 148.910 ;
        RECT 123.280 148.770 124.400 148.830 ;
        RECT 120.920 146.130 121.180 146.450 ;
        RECT 120.980 145.510 121.120 146.130 ;
        RECT 120.520 145.370 121.120 145.510 ;
        RECT 120.520 143.050 120.660 145.370 ;
        RECT 120.920 144.770 121.180 145.090 ;
        RECT 120.460 142.730 120.720 143.050 ;
        RECT 120.460 137.630 120.720 137.950 ;
        RECT 120.520 133.190 120.660 137.630 ;
        RECT 120.460 132.870 120.720 133.190 ;
        RECT 120.000 130.150 120.260 130.470 ;
        RECT 120.980 130.130 121.120 144.770 ;
        RECT 121.440 143.390 121.580 148.655 ;
        RECT 122.360 147.810 122.500 148.770 ;
        RECT 124.140 148.510 124.400 148.770 ;
        RECT 122.760 147.830 123.020 148.150 ;
        RECT 122.300 147.490 122.560 147.810 ;
        RECT 121.380 143.070 121.640 143.390 ;
        RECT 122.300 143.070 122.560 143.390 ;
        RECT 121.440 140.330 121.580 143.070 ;
        RECT 121.380 140.010 121.640 140.330 ;
        RECT 121.840 140.010 122.100 140.330 ;
        RECT 121.900 134.890 122.040 140.010 ;
        RECT 121.840 134.570 122.100 134.890 ;
        RECT 122.360 134.210 122.500 143.070 ;
        RECT 122.820 140.670 122.960 147.830 ;
        RECT 124.140 147.490 124.400 147.810 ;
        RECT 124.200 146.450 124.340 147.490 ;
        RECT 124.140 146.130 124.400 146.450 ;
        RECT 123.680 143.300 123.940 143.390 ;
        RECT 124.660 143.300 124.800 152.930 ;
        RECT 123.680 143.160 124.800 143.300 ;
        RECT 123.680 143.070 123.940 143.160 ;
        RECT 122.760 140.350 123.020 140.670 ;
        RECT 123.220 140.240 123.480 140.330 ;
        RECT 123.740 140.240 123.880 143.070 ;
        RECT 124.140 140.240 124.400 140.330 ;
        RECT 123.220 140.100 124.400 140.240 ;
        RECT 123.220 140.010 123.480 140.100 ;
        RECT 124.140 140.010 124.400 140.100 ;
        RECT 124.600 135.870 124.860 135.910 ;
        RECT 125.120 135.870 125.260 184.030 ;
        RECT 126.960 179.430 127.100 188.630 ;
        RECT 131.960 188.290 132.220 188.610 ;
        RECT 127.360 187.270 127.620 187.590 ;
        RECT 127.420 184.190 127.560 187.270 ;
        RECT 132.020 184.870 132.160 188.290 ;
        RECT 132.420 186.590 132.680 186.910 ;
        RECT 134.260 186.590 134.520 186.910 ;
        RECT 132.480 184.870 132.620 186.590 ;
        RECT 132.880 185.910 133.140 186.230 ;
        RECT 131.960 184.550 132.220 184.870 ;
        RECT 132.420 184.550 132.680 184.870 ;
        RECT 127.360 183.870 127.620 184.190 ;
        RECT 132.420 183.870 132.680 184.190 ;
        RECT 131.040 183.530 131.300 183.850 ;
        RECT 127.820 182.850 128.080 183.170 ;
        RECT 130.120 182.850 130.380 183.170 ;
        RECT 127.880 182.150 128.020 182.850 ;
        RECT 127.820 181.830 128.080 182.150 ;
        RECT 128.740 181.490 129.000 181.810 ;
        RECT 128.280 180.130 128.540 180.450 ;
        RECT 126.900 179.110 127.160 179.430 ;
        RECT 126.440 178.770 126.700 179.090 ;
        RECT 125.520 177.750 125.780 178.070 ;
        RECT 125.980 177.750 126.240 178.070 ;
        RECT 125.580 172.630 125.720 177.750 ;
        RECT 126.040 176.710 126.180 177.750 ;
        RECT 125.980 176.390 126.240 176.710 ;
        RECT 126.500 176.370 126.640 178.770 ;
        RECT 127.360 178.430 127.620 178.750 ;
        RECT 126.440 176.050 126.700 176.370 ;
        RECT 125.520 172.310 125.780 172.630 ;
        RECT 126.500 172.290 126.640 176.050 ;
        RECT 126.900 174.690 127.160 175.010 ;
        RECT 126.440 171.970 126.700 172.290 ;
        RECT 126.500 171.270 126.640 171.970 ;
        RECT 126.440 170.950 126.700 171.270 ;
        RECT 126.440 170.270 126.700 170.590 ;
        RECT 125.970 168.375 126.250 168.745 ;
        RECT 125.980 168.230 126.240 168.375 ;
        RECT 125.520 167.890 125.780 168.210 ;
        RECT 125.580 167.530 125.720 167.890 ;
        RECT 125.520 167.210 125.780 167.530 ;
        RECT 125.580 165.490 125.720 167.210 ;
        RECT 126.500 165.830 126.640 170.270 ;
        RECT 126.960 167.190 127.100 174.690 ;
        RECT 126.900 166.870 127.160 167.190 ;
        RECT 126.440 165.510 126.700 165.830 ;
        RECT 127.420 165.490 127.560 178.430 ;
        RECT 128.340 178.410 128.480 180.130 ;
        RECT 128.800 178.830 128.940 181.490 ;
        RECT 128.800 178.690 129.400 178.830 ;
        RECT 129.660 178.770 129.920 179.090 ;
        RECT 128.280 178.090 128.540 178.410 ;
        RECT 127.820 177.750 128.080 178.070 ;
        RECT 127.880 175.010 128.020 177.750 ;
        RECT 128.800 176.110 128.940 178.690 ;
        RECT 129.260 178.410 129.400 178.690 ;
        RECT 129.720 178.410 129.860 178.770 ;
        RECT 129.200 178.090 129.460 178.410 ;
        RECT 129.660 178.090 129.920 178.410 ;
        RECT 129.200 177.410 129.460 177.730 ;
        RECT 129.260 176.370 129.400 177.410 ;
        RECT 129.660 176.390 129.920 176.710 ;
        RECT 128.340 175.970 128.940 176.110 ;
        RECT 129.200 176.050 129.460 176.370 ;
        RECT 128.340 175.690 128.480 175.970 ;
        RECT 128.280 175.370 128.540 175.690 ;
        RECT 127.820 174.690 128.080 175.010 ;
        RECT 127.880 168.630 128.020 174.690 ;
        RECT 129.260 173.990 129.400 176.050 ;
        RECT 129.200 173.670 129.460 173.990 ;
        RECT 128.280 172.650 128.540 172.970 ;
        RECT 128.340 172.290 128.480 172.650 ;
        RECT 128.730 172.455 129.010 172.825 ;
        RECT 128.800 172.290 128.940 172.455 ;
        RECT 128.280 171.970 128.540 172.290 ;
        RECT 128.740 171.970 129.000 172.290 ;
        RECT 128.340 170.590 128.480 171.970 ;
        RECT 128.800 170.670 128.940 171.970 ;
        RECT 129.260 171.270 129.400 173.670 ;
        RECT 129.720 171.270 129.860 176.390 ;
        RECT 130.180 175.350 130.320 182.850 ;
        RECT 130.580 177.750 130.840 178.070 ;
        RECT 130.640 175.690 130.780 177.750 ;
        RECT 130.580 175.370 130.840 175.690 ;
        RECT 130.120 175.030 130.380 175.350 ;
        RECT 129.200 170.950 129.460 171.270 ;
        RECT 129.660 170.950 129.920 171.270 ;
        RECT 128.280 170.270 128.540 170.590 ;
        RECT 128.800 170.530 129.400 170.670 ;
        RECT 127.880 168.490 128.480 168.630 ;
        RECT 127.820 167.890 128.080 168.210 ;
        RECT 127.880 167.530 128.020 167.890 ;
        RECT 127.820 167.210 128.080 167.530 ;
        RECT 128.340 167.270 128.480 168.490 ;
        RECT 125.520 165.170 125.780 165.490 ;
        RECT 127.360 165.170 127.620 165.490 ;
        RECT 125.980 164.490 126.240 164.810 ;
        RECT 126.040 160.390 126.180 164.490 ;
        RECT 127.420 161.830 127.560 165.170 ;
        RECT 127.880 162.625 128.020 167.210 ;
        RECT 128.340 167.130 128.940 167.270 ;
        RECT 128.800 166.850 128.940 167.130 ;
        RECT 128.280 166.530 128.540 166.850 ;
        RECT 128.740 166.530 129.000 166.850 ;
        RECT 127.810 162.255 128.090 162.625 ;
        RECT 128.340 162.430 128.480 166.530 ;
        RECT 129.260 165.910 129.400 170.530 ;
        RECT 130.180 170.370 130.320 175.030 ;
        RECT 130.640 172.145 130.780 175.370 ;
        RECT 130.570 171.775 130.850 172.145 ;
        RECT 130.640 170.930 130.780 171.775 ;
        RECT 130.580 170.610 130.840 170.930 ;
        RECT 130.180 170.230 130.780 170.370 ;
        RECT 129.660 169.590 129.920 169.910 ;
        RECT 130.120 169.590 130.380 169.910 ;
        RECT 129.720 169.425 129.860 169.590 ;
        RECT 129.650 169.055 129.930 169.425 ;
        RECT 130.180 168.550 130.320 169.590 ;
        RECT 130.120 168.230 130.380 168.550 ;
        RECT 130.120 166.870 130.380 167.190 ;
        RECT 129.260 165.770 129.860 165.910 ;
        RECT 129.200 164.830 129.460 165.150 ;
        RECT 128.740 163.810 129.000 164.130 ;
        RECT 128.800 162.770 128.940 163.810 ;
        RECT 128.740 162.450 129.000 162.770 ;
        RECT 127.820 162.110 128.080 162.255 ;
        RECT 128.280 162.110 128.540 162.430 ;
        RECT 126.960 161.750 127.560 161.830 ;
        RECT 126.900 161.690 127.560 161.750 ;
        RECT 126.900 161.430 127.160 161.690 ;
        RECT 127.820 161.430 128.080 161.750 ;
        RECT 125.980 160.070 126.240 160.390 ;
        RECT 127.880 157.670 128.020 161.430 ;
        RECT 129.260 161.410 129.400 164.830 ;
        RECT 129.200 161.090 129.460 161.410 ;
        RECT 128.740 159.620 129.000 159.710 ;
        RECT 129.260 159.620 129.400 161.090 ;
        RECT 128.740 159.480 129.400 159.620 ;
        RECT 128.740 159.390 129.000 159.480 ;
        RECT 129.200 158.710 129.460 159.030 ;
        RECT 127.820 157.350 128.080 157.670 ;
        RECT 125.970 156.815 126.250 157.185 ;
        RECT 126.040 151.550 126.180 156.815 ;
        RECT 127.820 156.670 128.080 156.990 ;
        RECT 127.880 154.610 128.020 156.670 ;
        RECT 128.740 156.560 129.000 156.650 ;
        RECT 129.260 156.560 129.400 158.710 ;
        RECT 129.720 156.990 129.860 165.770 ;
        RECT 130.180 164.470 130.320 166.870 ;
        RECT 130.640 165.490 130.780 170.230 ;
        RECT 131.100 170.105 131.240 183.530 ;
        RECT 131.960 181.150 132.220 181.470 ;
        RECT 131.500 178.770 131.760 179.090 ;
        RECT 131.560 176.030 131.700 178.770 ;
        RECT 132.020 178.410 132.160 181.150 ;
        RECT 131.960 178.090 132.220 178.410 ;
        RECT 132.020 176.710 132.160 178.090 ;
        RECT 132.480 178.070 132.620 183.870 ;
        RECT 132.940 179.430 133.080 185.910 ;
        RECT 133.800 183.530 134.060 183.850 ;
        RECT 133.860 182.150 134.000 183.530 ;
        RECT 134.320 182.150 134.460 186.590 ;
        RECT 133.800 181.830 134.060 182.150 ;
        RECT 134.260 181.830 134.520 182.150 ;
        RECT 132.880 179.110 133.140 179.430 ;
        RECT 132.420 177.750 132.680 178.070 ;
        RECT 131.960 176.390 132.220 176.710 ;
        RECT 132.020 176.225 132.160 176.390 ;
        RECT 131.500 175.710 131.760 176.030 ;
        RECT 131.950 175.855 132.230 176.225 ;
        RECT 131.560 170.250 131.700 175.710 ;
        RECT 132.480 175.350 132.620 177.750 ;
        RECT 132.940 176.710 133.080 179.110 ;
        RECT 132.880 176.390 133.140 176.710 ;
        RECT 132.940 176.030 134.000 176.110 ;
        RECT 132.940 175.970 134.060 176.030 ;
        RECT 132.420 175.030 132.680 175.350 ;
        RECT 131.960 174.690 132.220 175.010 ;
        RECT 132.020 172.970 132.160 174.690 ;
        RECT 131.960 172.650 132.220 172.970 ;
        RECT 132.480 172.030 132.620 175.030 ;
        RECT 132.940 172.290 133.080 175.970 ;
        RECT 133.800 175.710 134.060 175.970 ;
        RECT 133.340 175.370 133.600 175.690 ;
        RECT 134.320 175.430 134.460 181.830 ;
        RECT 140.700 181.150 140.960 181.470 ;
        RECT 137.480 180.130 137.740 180.450 ;
        RECT 137.540 178.410 137.680 180.130 ;
        RECT 140.760 179.430 140.900 181.150 ;
        RECT 140.700 179.110 140.960 179.430 ;
        RECT 137.480 178.090 137.740 178.410 ;
        RECT 142.080 178.090 142.340 178.410 ;
        RECT 143.920 178.090 144.180 178.410 ;
        RECT 135.640 177.750 135.900 178.070 ;
        RECT 135.700 176.710 135.840 177.750 ;
        RECT 135.640 176.390 135.900 176.710 ;
        RECT 134.710 175.855 134.990 176.225 ;
        RECT 137.540 176.030 137.680 178.090 ;
        RECT 140.700 177.410 140.960 177.730 ;
        RECT 134.720 175.710 134.980 175.855 ;
        RECT 136.560 175.710 136.820 176.030 ;
        RECT 137.480 175.710 137.740 176.030 ;
        RECT 137.940 175.710 138.200 176.030 ;
        RECT 138.860 175.710 139.120 176.030 ;
        RECT 133.400 173.650 133.540 175.370 ;
        RECT 134.320 175.290 134.920 175.430 ;
        RECT 133.340 173.330 133.600 173.650 ;
        RECT 133.340 172.650 133.600 172.970 ;
        RECT 133.800 172.650 134.060 172.970 ;
        RECT 134.260 172.650 134.520 172.970 ;
        RECT 132.020 171.890 132.620 172.030 ;
        RECT 132.880 171.970 133.140 172.290 ;
        RECT 131.030 169.735 131.310 170.105 ;
        RECT 131.500 169.930 131.760 170.250 ;
        RECT 131.040 169.250 131.300 169.570 ;
        RECT 131.100 168.210 131.240 169.250 ;
        RECT 131.040 167.890 131.300 168.210 ;
        RECT 131.500 167.210 131.760 167.530 ;
        RECT 130.580 165.170 130.840 165.490 ;
        RECT 131.030 164.975 131.310 165.345 ;
        RECT 131.040 164.830 131.300 164.975 ;
        RECT 130.120 164.150 130.380 164.470 ;
        RECT 130.180 162.090 130.320 164.150 ;
        RECT 131.040 162.450 131.300 162.770 ;
        RECT 130.120 161.770 130.380 162.090 ;
        RECT 130.180 159.710 130.320 161.770 ;
        RECT 131.100 161.410 131.240 162.450 ;
        RECT 130.580 161.090 130.840 161.410 ;
        RECT 131.040 161.090 131.300 161.410 ;
        RECT 130.120 159.390 130.380 159.710 ;
        RECT 130.180 158.690 130.320 159.390 ;
        RECT 130.120 158.370 130.380 158.690 ;
        RECT 129.660 156.670 129.920 156.990 ;
        RECT 130.640 156.650 130.780 161.090 ;
        RECT 128.740 156.420 129.400 156.560 ;
        RECT 128.740 156.330 129.000 156.420 ;
        RECT 130.580 156.330 130.840 156.650 ;
        RECT 131.040 156.330 131.300 156.650 ;
        RECT 128.280 155.990 128.540 156.310 ;
        RECT 129.660 155.990 129.920 156.310 ;
        RECT 127.820 154.290 128.080 154.610 ;
        RECT 127.820 153.610 128.080 153.930 ;
        RECT 127.880 152.230 128.020 153.610 ;
        RECT 127.820 151.910 128.080 152.230 ;
        RECT 126.440 151.630 126.700 151.890 ;
        RECT 128.340 151.630 128.480 155.990 ;
        RECT 128.740 155.710 129.000 155.970 ;
        RECT 128.740 155.650 129.400 155.710 ;
        RECT 128.800 155.570 129.400 155.650 ;
        RECT 126.440 151.570 128.480 151.630 ;
        RECT 125.980 151.230 126.240 151.550 ;
        RECT 126.500 151.490 128.480 151.570 ;
        RECT 125.520 150.550 125.780 150.870 ;
        RECT 125.580 148.830 125.720 150.550 ;
        RECT 125.520 148.510 125.780 148.830 ;
        RECT 125.580 145.510 125.720 148.510 ;
        RECT 126.040 148.490 126.180 151.230 ;
        RECT 126.440 150.890 126.700 151.210 ;
        RECT 127.820 150.890 128.080 151.210 ;
        RECT 125.980 148.170 126.240 148.490 ;
        RECT 126.500 146.110 126.640 150.890 ;
        RECT 127.880 150.530 128.020 150.890 ;
        RECT 127.820 150.210 128.080 150.530 ;
        RECT 128.340 148.830 128.480 151.490 ;
        RECT 128.280 148.510 128.540 148.830 ;
        RECT 127.360 148.170 127.620 148.490 ;
        RECT 126.440 145.790 126.700 146.110 ;
        RECT 125.580 145.370 126.180 145.510 ;
        RECT 125.520 144.770 125.780 145.090 ;
        RECT 125.580 143.390 125.720 144.770 ;
        RECT 125.520 143.070 125.780 143.390 ;
        RECT 126.040 140.330 126.180 145.370 ;
        RECT 126.900 144.770 127.160 145.090 ;
        RECT 126.960 141.350 127.100 144.770 ;
        RECT 127.420 144.070 127.560 148.170 ;
        RECT 127.360 143.750 127.620 144.070 ;
        RECT 126.900 141.030 127.160 141.350 ;
        RECT 128.740 140.350 129.000 140.670 ;
        RECT 125.980 140.010 126.240 140.330 ;
        RECT 128.800 138.290 128.940 140.350 ;
        RECT 128.740 137.970 129.000 138.290 ;
        RECT 129.260 137.950 129.400 155.570 ;
        RECT 129.720 154.950 129.860 155.990 ;
        RECT 129.660 154.630 129.920 154.950 ;
        RECT 130.570 154.095 130.850 154.465 ;
        RECT 130.640 153.590 130.780 154.095 ;
        RECT 131.100 153.785 131.240 156.330 ;
        RECT 130.580 153.270 130.840 153.590 ;
        RECT 131.030 153.415 131.310 153.785 ;
        RECT 131.100 151.550 131.240 153.415 ;
        RECT 131.040 151.230 131.300 151.550 ;
        RECT 131.560 151.210 131.700 167.210 ;
        RECT 132.020 164.665 132.160 171.890 ;
        RECT 132.940 170.590 133.080 171.970 ;
        RECT 133.400 171.270 133.540 172.650 ;
        RECT 133.340 170.950 133.600 171.270 ;
        RECT 133.400 170.785 133.540 170.950 ;
        RECT 132.880 170.270 133.140 170.590 ;
        RECT 133.330 170.415 133.610 170.785 ;
        RECT 133.860 170.590 134.000 172.650 ;
        RECT 134.320 170.590 134.460 172.650 ;
        RECT 134.780 170.590 134.920 175.290 ;
        RECT 135.640 175.030 135.900 175.350 ;
        RECT 135.700 172.970 135.840 175.030 ;
        RECT 136.620 175.010 136.760 175.710 ;
        RECT 136.100 174.690 136.360 175.010 ;
        RECT 136.560 174.690 136.820 175.010 ;
        RECT 136.160 173.650 136.300 174.690 ;
        RECT 136.100 173.330 136.360 173.650 ;
        RECT 135.640 172.650 135.900 172.970 ;
        RECT 132.420 169.590 132.680 169.910 ;
        RECT 132.880 169.590 133.140 169.910 ;
        RECT 132.480 169.425 132.620 169.590 ;
        RECT 132.410 169.055 132.690 169.425 ;
        RECT 131.950 164.295 132.230 164.665 ;
        RECT 131.960 163.810 132.220 164.130 ;
        RECT 132.020 159.710 132.160 163.810 ;
        RECT 132.480 163.110 132.620 169.055 ;
        RECT 132.940 168.065 133.080 169.590 ;
        RECT 132.870 167.695 133.150 168.065 ;
        RECT 132.940 167.190 133.080 167.695 ;
        RECT 132.880 166.870 133.140 167.190 ;
        RECT 133.400 165.345 133.540 170.415 ;
        RECT 133.800 170.270 134.060 170.590 ;
        RECT 134.260 170.270 134.520 170.590 ;
        RECT 134.720 170.270 134.980 170.590 ;
        RECT 134.260 168.230 134.520 168.550 ;
        RECT 134.320 167.270 134.460 168.230 ;
        RECT 134.780 168.210 134.920 170.270 ;
        RECT 135.180 169.930 135.440 170.250 ;
        RECT 135.240 169.570 135.380 169.930 ;
        RECT 135.180 169.250 135.440 169.570 ;
        RECT 135.640 169.250 135.900 169.570 ;
        RECT 134.720 167.890 134.980 168.210 ;
        RECT 135.700 167.870 135.840 169.250 ;
        RECT 136.620 168.745 136.760 174.690 ;
        RECT 137.020 169.590 137.280 169.910 ;
        RECT 136.100 168.230 136.360 168.550 ;
        RECT 136.550 168.375 136.830 168.745 ;
        RECT 135.640 167.550 135.900 167.870 ;
        RECT 136.160 167.270 136.300 168.230 ;
        RECT 137.080 167.530 137.220 169.590 ;
        RECT 134.320 167.130 134.920 167.270 ;
        RECT 133.800 166.530 134.060 166.850 ;
        RECT 134.260 166.530 134.520 166.850 ;
        RECT 133.330 164.975 133.610 165.345 ;
        RECT 132.420 162.790 132.680 163.110 ;
        RECT 133.860 162.090 134.000 166.530 ;
        RECT 133.800 161.770 134.060 162.090 ;
        RECT 132.420 161.430 132.680 161.750 ;
        RECT 133.340 161.430 133.600 161.750 ;
        RECT 132.480 160.390 132.620 161.430 ;
        RECT 132.420 160.300 132.680 160.390 ;
        RECT 132.420 160.160 133.080 160.300 ;
        RECT 132.420 160.070 132.680 160.160 ;
        RECT 131.960 159.390 132.220 159.710 ;
        RECT 132.420 159.390 132.680 159.710 ;
        RECT 132.480 158.545 132.620 159.390 ;
        RECT 132.940 159.110 133.080 160.160 ;
        RECT 133.400 159.710 133.540 161.430 ;
        RECT 133.800 160.070 134.060 160.390 ;
        RECT 133.860 159.710 134.000 160.070 ;
        RECT 133.340 159.390 133.600 159.710 ;
        RECT 133.800 159.390 134.060 159.710 ;
        RECT 132.940 158.970 133.540 159.110 ;
        RECT 132.410 158.175 132.690 158.545 ;
        RECT 132.880 158.370 133.140 158.690 ;
        RECT 132.410 156.815 132.690 157.185 ;
        RECT 132.420 156.670 132.680 156.815 ;
        RECT 132.940 154.950 133.080 158.370 ;
        RECT 132.880 154.630 133.140 154.950 ;
        RECT 132.420 153.950 132.680 154.270 ;
        RECT 132.480 152.230 132.620 153.950 ;
        RECT 133.400 153.250 133.540 158.970 ;
        RECT 133.800 158.710 134.060 159.030 ;
        RECT 133.340 152.930 133.600 153.250 ;
        RECT 132.420 151.910 132.680 152.230 ;
        RECT 129.660 150.890 129.920 151.210 ;
        RECT 131.500 150.890 131.760 151.210 ;
        RECT 129.720 149.510 129.860 150.890 ;
        RECT 129.660 149.190 129.920 149.510 ;
        RECT 129.660 148.510 129.920 148.830 ;
        RECT 130.110 148.740 130.390 149.025 ;
        RECT 131.500 148.850 131.760 149.170 ;
        RECT 130.110 148.655 130.780 148.740 ;
        RECT 130.120 148.600 130.780 148.655 ;
        RECT 130.120 148.510 130.380 148.600 ;
        RECT 129.720 141.010 129.860 148.510 ;
        RECT 130.120 147.490 130.380 147.810 ;
        RECT 129.660 140.690 129.920 141.010 ;
        RECT 130.180 140.330 130.320 147.490 ;
        RECT 130.640 140.330 130.780 148.600 ;
        RECT 131.040 145.790 131.300 146.110 ;
        RECT 131.100 144.070 131.240 145.790 ;
        RECT 131.040 143.750 131.300 144.070 ;
        RECT 130.120 140.010 130.380 140.330 ;
        RECT 130.580 140.010 130.840 140.330 ;
        RECT 130.120 139.330 130.380 139.650 ;
        RECT 129.200 137.630 129.460 137.950 ;
        RECT 124.600 135.730 125.260 135.870 ;
        RECT 124.600 135.590 124.860 135.730 ;
        RECT 125.120 134.890 125.260 135.730 ;
        RECT 125.060 134.570 125.320 134.890 ;
        RECT 128.280 134.230 128.540 134.550 ;
        RECT 122.300 133.890 122.560 134.210 ;
        RECT 128.340 133.190 128.480 134.230 ;
        RECT 128.280 132.870 128.540 133.190 ;
        RECT 129.200 132.190 129.460 132.510 ;
        RECT 122.300 131.850 122.560 132.170 ;
        RECT 120.920 130.040 121.180 130.130 ;
        RECT 120.920 129.900 121.580 130.040 ;
        RECT 120.920 129.810 121.180 129.900 ;
        RECT 120.920 129.130 121.180 129.450 ;
        RECT 119.540 125.730 119.800 126.050 ;
        RECT 118.620 124.030 118.880 124.350 ;
        RECT 119.600 122.070 119.740 125.730 ;
        RECT 119.600 121.930 120.200 122.070 ;
        RECT 117.700 119.270 117.960 119.590 ;
        RECT 120.060 118.570 120.200 121.930 ;
        RECT 120.980 118.570 121.120 129.130 ;
        RECT 121.440 127.410 121.580 129.900 ;
        RECT 122.360 127.750 122.500 131.850 ;
        RECT 129.260 130.470 129.400 132.190 ;
        RECT 127.360 130.150 127.620 130.470 ;
        RECT 129.200 130.150 129.460 130.470 ;
        RECT 122.760 128.790 123.020 129.110 ;
        RECT 122.300 127.430 122.560 127.750 ;
        RECT 121.380 127.090 121.640 127.410 ;
        RECT 122.820 125.030 122.960 128.790 ;
        RECT 127.420 127.070 127.560 130.150 ;
        RECT 130.180 129.790 130.320 139.330 ;
        RECT 130.640 138.290 130.780 140.010 ;
        RECT 130.580 137.970 130.840 138.290 ;
        RECT 131.560 135.870 131.700 148.850 ;
        RECT 133.400 148.830 133.540 152.930 ;
        RECT 133.860 151.550 134.000 158.710 ;
        RECT 134.320 156.650 134.460 166.530 ;
        RECT 134.780 162.090 134.920 167.130 ;
        RECT 135.700 167.130 136.300 167.270 ;
        RECT 137.020 167.210 137.280 167.530 ;
        RECT 135.180 164.830 135.440 165.150 ;
        RECT 134.720 161.770 134.980 162.090 ;
        RECT 134.720 161.090 134.980 161.410 ;
        RECT 134.260 156.330 134.520 156.650 ;
        RECT 134.260 153.950 134.520 154.270 ;
        RECT 133.800 151.230 134.060 151.550 ;
        RECT 133.860 148.830 134.000 151.230 ;
        RECT 133.340 148.510 133.600 148.830 ;
        RECT 133.800 148.510 134.060 148.830 ;
        RECT 133.860 146.110 134.000 148.510 ;
        RECT 133.800 145.790 134.060 146.110 ;
        RECT 133.860 143.730 134.000 145.790 ;
        RECT 133.800 143.410 134.060 143.730 ;
        RECT 131.960 139.330 132.220 139.650 ;
        RECT 131.100 135.730 131.700 135.870 ;
        RECT 130.580 133.890 130.840 134.210 ;
        RECT 130.640 132.510 130.780 133.890 ;
        RECT 130.580 132.190 130.840 132.510 ;
        RECT 130.120 129.470 130.380 129.790 ;
        RECT 127.360 126.750 127.620 127.070 ;
        RECT 123.220 125.730 123.480 126.050 ;
        RECT 122.760 124.710 123.020 125.030 ;
        RECT 123.280 124.350 123.420 125.730 ;
        RECT 128.280 124.370 128.540 124.690 ;
        RECT 123.220 124.030 123.480 124.350 ;
        RECT 126.440 120.970 126.700 121.290 ;
        RECT 121.380 120.290 121.640 120.610 ;
        RECT 118.160 118.250 118.420 118.570 ;
        RECT 120.000 118.250 120.260 118.570 ;
        RECT 120.920 118.250 121.180 118.570 ;
        RECT 115.860 116.550 116.120 116.870 ;
        RECT 118.220 116.530 118.360 118.250 ;
        RECT 119.540 117.910 119.800 118.230 ;
        RECT 118.160 116.210 118.420 116.530 ;
        RECT 114.940 115.870 115.200 116.190 ;
        RECT 114.080 115.450 114.680 115.590 ;
        RECT 116.320 115.530 116.580 115.850 ;
        RECT 114.020 114.850 114.280 115.170 ;
        RECT 113.160 113.410 113.760 113.550 ;
        RECT 110.800 112.810 111.060 113.130 ;
        RECT 108.960 111.000 109.220 111.090 ;
        RECT 108.960 110.860 109.620 111.000 ;
        RECT 108.960 110.770 109.220 110.860 ;
        RECT 108.960 110.090 109.220 110.410 ;
        RECT 108.500 107.710 108.760 108.030 ;
        RECT 108.040 107.370 108.300 107.690 ;
        RECT 108.100 105.650 108.240 107.370 ;
        RECT 108.040 105.330 108.300 105.650 ;
        RECT 108.100 104.290 108.240 105.330 ;
        RECT 108.560 104.630 108.700 107.710 ;
        RECT 109.020 107.010 109.160 110.090 ;
        RECT 108.960 106.690 109.220 107.010 ;
        RECT 108.500 104.310 108.760 104.630 ;
        RECT 108.040 103.970 108.300 104.290 ;
        RECT 107.120 93.770 107.380 94.090 ;
        RECT 106.660 92.070 106.920 92.390 ;
        RECT 105.280 91.730 105.540 92.050 ;
        RECT 107.180 91.370 107.320 93.770 ;
        RECT 104.360 91.050 104.620 91.370 ;
        RECT 107.120 91.050 107.380 91.370 ;
        RECT 104.420 85.930 104.560 91.050 ;
        RECT 104.820 90.710 105.080 91.030 ;
        RECT 107.580 90.710 107.840 91.030 ;
        RECT 104.880 87.970 105.020 90.710 ;
        RECT 107.640 89.670 107.780 90.710 ;
        RECT 107.580 89.350 107.840 89.670 ;
        RECT 104.820 87.650 105.080 87.970 ;
        RECT 97.460 85.610 97.720 85.930 ;
        RECT 102.980 85.610 103.240 85.930 ;
        RECT 104.360 85.610 104.620 85.930 ;
        RECT 98.840 84.930 99.100 85.250 ;
        RECT 102.060 84.930 102.320 85.250 ;
        RECT 98.900 77.700 99.040 84.930 ;
        RECT 102.120 77.700 102.260 84.930 ;
        RECT 104.880 83.890 105.020 87.650 ;
        RECT 108.100 85.930 108.240 103.970 ;
        RECT 108.560 97.150 108.700 104.310 ;
        RECT 109.480 102.250 109.620 110.860 ;
        RECT 109.880 109.410 110.140 109.730 ;
        RECT 109.940 102.930 110.080 109.410 ;
        RECT 110.340 107.030 110.600 107.350 ;
        RECT 110.400 103.270 110.540 107.030 ;
        RECT 110.340 102.950 110.600 103.270 ;
        RECT 109.880 102.610 110.140 102.930 ;
        RECT 109.420 101.930 109.680 102.250 ;
        RECT 109.480 100.210 109.620 101.930 ;
        RECT 109.420 99.890 109.680 100.210 ;
        RECT 108.960 98.870 109.220 99.190 ;
        RECT 108.500 96.830 108.760 97.150 ;
        RECT 108.500 95.810 108.760 96.130 ;
        RECT 108.560 88.310 108.700 95.810 ;
        RECT 109.020 95.110 109.160 98.870 ;
        RECT 109.420 98.530 109.680 98.850 ;
        RECT 108.960 94.790 109.220 95.110 ;
        RECT 109.480 94.770 109.620 98.530 ;
        RECT 110.340 95.810 110.600 96.130 ;
        RECT 110.400 94.770 110.540 95.810 ;
        RECT 109.420 94.450 109.680 94.770 ;
        RECT 110.340 94.450 110.600 94.770 ;
        RECT 110.860 89.330 111.000 112.810 ;
        RECT 111.260 106.690 111.520 107.010 ;
        RECT 111.320 105.310 111.460 106.690 ;
        RECT 111.260 104.990 111.520 105.310 ;
        RECT 110.800 89.010 111.060 89.330 ;
        RECT 108.500 87.990 108.760 88.310 ;
        RECT 111.320 85.930 111.460 104.990 ;
        RECT 112.640 99.890 112.900 100.210 ;
        RECT 111.720 98.530 111.980 98.850 ;
        RECT 111.780 97.490 111.920 98.530 ;
        RECT 111.720 97.170 111.980 97.490 ;
        RECT 112.700 89.330 112.840 99.890 ;
        RECT 113.160 96.470 113.300 113.410 ;
        RECT 113.560 112.810 113.820 113.130 ;
        RECT 113.620 108.710 113.760 112.810 ;
        RECT 114.080 110.070 114.220 114.850 ;
        RECT 114.020 109.750 114.280 110.070 ;
        RECT 113.560 108.390 113.820 108.710 ;
        RECT 114.540 102.250 114.680 115.450 ;
        RECT 115.400 113.830 115.660 114.150 ;
        RECT 114.940 112.470 115.200 112.790 ;
        RECT 115.000 111.430 115.140 112.470 ;
        RECT 115.460 112.450 115.600 113.830 ;
        RECT 116.380 113.130 116.520 115.530 ;
        RECT 116.320 112.810 116.580 113.130 ;
        RECT 115.400 112.130 115.660 112.450 ;
        RECT 114.940 111.110 115.200 111.430 ;
        RECT 119.080 109.410 119.340 109.730 ;
        RECT 114.940 105.330 115.200 105.650 ;
        RECT 114.480 102.160 114.740 102.250 ;
        RECT 114.080 102.020 114.740 102.160 ;
        RECT 114.080 99.530 114.220 102.020 ;
        RECT 114.480 101.930 114.740 102.020 ;
        RECT 114.480 101.250 114.740 101.570 ;
        RECT 114.020 99.210 114.280 99.530 ;
        RECT 114.540 97.830 114.680 101.250 ;
        RECT 114.480 97.510 114.740 97.830 ;
        RECT 115.000 97.490 115.140 105.330 ;
        RECT 116.780 104.650 117.040 104.970 ;
        RECT 116.840 99.870 116.980 104.650 ;
        RECT 118.620 101.590 118.880 101.910 ;
        RECT 117.700 101.250 117.960 101.570 ;
        RECT 116.780 99.550 117.040 99.870 ;
        RECT 114.940 97.170 115.200 97.490 ;
        RECT 116.840 96.810 116.980 99.550 ;
        RECT 117.760 99.190 117.900 101.250 ;
        RECT 118.680 100.550 118.820 101.590 ;
        RECT 118.160 100.230 118.420 100.550 ;
        RECT 118.620 100.230 118.880 100.550 ;
        RECT 117.700 98.870 117.960 99.190 ;
        RECT 117.240 97.170 117.500 97.490 ;
        RECT 114.940 96.490 115.200 96.810 ;
        RECT 116.780 96.490 117.040 96.810 ;
        RECT 113.100 96.150 113.360 96.470 ;
        RECT 115.000 90.690 115.140 96.490 ;
        RECT 115.400 95.810 115.660 96.130 ;
        RECT 116.780 95.810 117.040 96.130 ;
        RECT 113.100 90.370 113.360 90.690 ;
        RECT 114.940 90.370 115.200 90.690 ;
        RECT 112.640 89.010 112.900 89.330 ;
        RECT 113.160 85.930 113.300 90.370 ;
        RECT 113.560 88.330 113.820 88.650 ;
        RECT 113.620 86.610 113.760 88.330 ;
        RECT 115.460 86.950 115.600 95.810 ;
        RECT 116.840 94.430 116.980 95.810 ;
        RECT 117.300 94.770 117.440 97.170 ;
        RECT 118.220 97.150 118.360 100.230 ;
        RECT 118.160 96.830 118.420 97.150 ;
        RECT 117.700 94.790 117.960 95.110 ;
        RECT 117.240 94.450 117.500 94.770 ;
        RECT 116.780 94.110 117.040 94.430 ;
        RECT 116.840 93.750 116.980 94.110 ;
        RECT 116.780 93.430 117.040 93.750 ;
        RECT 116.320 93.090 116.580 93.410 ;
        RECT 115.860 90.710 116.120 91.030 ;
        RECT 115.920 89.670 116.060 90.710 ;
        RECT 115.860 89.350 116.120 89.670 ;
        RECT 115.400 86.630 115.660 86.950 ;
        RECT 116.380 86.610 116.520 93.090 ;
        RECT 117.760 89.670 117.900 94.790 ;
        RECT 118.160 90.370 118.420 90.690 ;
        RECT 118.220 89.670 118.360 90.370 ;
        RECT 117.700 89.350 117.960 89.670 ;
        RECT 118.160 89.350 118.420 89.670 ;
        RECT 118.220 87.570 118.360 89.350 ;
        RECT 119.140 88.650 119.280 109.410 ;
        RECT 119.600 97.830 119.740 117.910 ;
        RECT 120.460 116.210 120.720 116.530 ;
        RECT 120.000 113.490 120.260 113.810 ;
        RECT 119.540 97.510 119.800 97.830 ;
        RECT 119.080 88.330 119.340 88.650 ;
        RECT 120.060 87.570 120.200 113.490 ;
        RECT 120.520 113.130 120.660 116.210 ;
        RECT 120.460 112.810 120.720 113.130 ;
        RECT 120.980 110.750 121.120 118.250 ;
        RECT 121.440 118.230 121.580 120.290 ;
        RECT 125.060 118.250 125.320 118.570 ;
        RECT 121.380 117.910 121.640 118.230 ;
        RECT 125.120 116.530 125.260 118.250 ;
        RECT 125.060 116.210 125.320 116.530 ;
        RECT 124.600 112.470 124.860 112.790 ;
        RECT 123.680 110.770 123.940 111.090 ;
        RECT 120.920 110.430 121.180 110.750 ;
        RECT 123.740 108.710 123.880 110.770 ;
        RECT 123.680 108.390 123.940 108.710 ;
        RECT 124.660 108.030 124.800 112.470 ;
        RECT 125.060 108.050 125.320 108.370 ;
        RECT 122.300 107.710 122.560 108.030 ;
        RECT 124.600 107.710 124.860 108.030 ;
        RECT 122.360 104.970 122.500 107.710 ;
        RECT 124.140 106.690 124.400 107.010 ;
        RECT 124.200 105.650 124.340 106.690 ;
        RECT 125.120 105.990 125.260 108.050 ;
        RECT 126.500 108.030 126.640 120.970 ;
        RECT 126.900 120.630 127.160 120.950 ;
        RECT 126.960 116.870 127.100 120.630 ;
        RECT 128.340 116.870 128.480 124.370 ;
        RECT 128.740 123.690 129.000 124.010 ;
        RECT 128.800 119.590 128.940 123.690 ;
        RECT 129.200 121.990 129.460 122.310 ;
        RECT 129.260 121.825 129.400 121.990 ;
        RECT 129.190 121.455 129.470 121.825 ;
        RECT 130.180 121.630 130.320 129.470 ;
        RECT 131.100 124.690 131.240 135.730 ;
        RECT 131.500 126.750 131.760 127.070 ;
        RECT 131.040 124.370 131.300 124.690 ;
        RECT 130.580 123.350 130.840 123.670 ;
        RECT 130.120 121.310 130.380 121.630 ;
        RECT 130.640 121.290 130.780 123.350 ;
        RECT 130.580 120.970 130.840 121.290 ;
        RECT 128.740 119.270 129.000 119.590 ;
        RECT 130.640 118.910 130.780 120.970 ;
        RECT 130.580 118.590 130.840 118.910 ;
        RECT 129.200 117.570 129.460 117.890 ;
        RECT 126.900 116.550 127.160 116.870 ;
        RECT 128.280 116.550 128.540 116.870 ;
        RECT 126.440 107.710 126.700 108.030 ;
        RECT 125.060 105.670 125.320 105.990 ;
        RECT 124.140 105.330 124.400 105.650 ;
        RECT 122.300 104.650 122.560 104.970 ;
        RECT 122.360 102.250 122.500 104.650 ;
        RECT 124.600 102.950 124.860 103.270 ;
        RECT 122.300 101.930 122.560 102.250 ;
        RECT 120.920 94.110 121.180 94.430 ;
        RECT 118.220 87.430 118.820 87.570 ;
        RECT 113.560 86.290 113.820 86.610 ;
        RECT 116.320 86.290 116.580 86.610 ;
        RECT 118.160 86.290 118.420 86.610 ;
        RECT 108.040 85.610 108.300 85.930 ;
        RECT 111.260 85.610 111.520 85.930 ;
        RECT 113.100 85.610 113.360 85.930 ;
        RECT 114.940 85.270 115.200 85.590 ;
        RECT 105.280 84.930 105.540 85.250 ;
        RECT 108.500 84.930 108.760 85.250 ;
        RECT 111.720 84.930 111.980 85.250 ;
        RECT 104.820 83.570 105.080 83.890 ;
        RECT 105.340 77.700 105.480 84.930 ;
        RECT 108.560 77.700 108.700 84.930 ;
        RECT 111.780 77.700 111.920 84.930 ;
        RECT 115.000 77.700 115.140 85.270 ;
        RECT 116.320 84.930 116.580 85.250 ;
        RECT 116.380 84.230 116.520 84.930 ;
        RECT 116.320 83.910 116.580 84.230 ;
        RECT 118.220 77.700 118.360 86.290 ;
        RECT 118.680 86.270 118.820 87.430 ;
        RECT 119.600 87.430 120.200 87.570 ;
        RECT 118.620 85.950 118.880 86.270 ;
        RECT 118.680 85.590 118.820 85.950 ;
        RECT 119.600 85.930 119.740 87.430 ;
        RECT 120.000 86.630 120.260 86.950 ;
        RECT 120.060 85.930 120.200 86.630 ;
        RECT 120.980 85.930 121.120 94.110 ;
        RECT 124.660 94.090 124.800 102.950 ;
        RECT 126.500 102.590 126.640 107.710 ;
        RECT 126.440 102.270 126.700 102.590 ;
        RECT 126.500 97.150 126.640 102.270 ;
        RECT 126.440 96.830 126.700 97.150 ;
        RECT 128.340 95.190 128.480 116.550 ;
        RECT 129.260 116.190 129.400 117.570 ;
        RECT 129.200 115.870 129.460 116.190 ;
        RECT 131.040 114.850 131.300 115.170 ;
        RECT 129.200 112.810 129.460 113.130 ;
        RECT 130.580 112.810 130.840 113.130 ;
        RECT 128.740 109.410 129.000 109.730 ;
        RECT 128.800 108.710 128.940 109.410 ;
        RECT 128.740 108.390 129.000 108.710 ;
        RECT 129.260 105.650 129.400 112.810 ;
        RECT 129.660 112.130 129.920 112.450 ;
        RECT 129.200 105.330 129.460 105.650 ;
        RECT 129.720 104.710 129.860 112.130 ;
        RECT 130.640 111.430 130.780 112.810 ;
        RECT 131.100 112.790 131.240 114.850 ;
        RECT 131.560 114.150 131.700 126.750 ;
        RECT 132.020 122.310 132.160 139.330 ;
        RECT 132.880 137.970 133.140 138.290 ;
        RECT 132.420 136.610 132.680 136.930 ;
        RECT 132.480 132.170 132.620 136.610 ;
        RECT 132.940 135.870 133.080 137.970 ;
        RECT 133.860 137.950 134.000 143.410 ;
        RECT 134.320 141.350 134.460 153.950 ;
        RECT 134.780 148.910 134.920 161.090 ;
        RECT 135.240 156.650 135.380 164.830 ;
        RECT 135.180 156.330 135.440 156.650 ;
        RECT 135.240 155.970 135.380 156.330 ;
        RECT 135.180 155.650 135.440 155.970 ;
        RECT 135.700 154.465 135.840 167.130 ;
        RECT 137.540 165.490 137.680 175.710 ;
        RECT 138.000 173.650 138.140 175.710 ;
        RECT 138.920 173.990 139.060 175.710 ;
        RECT 138.860 173.670 139.120 173.990 ;
        RECT 137.940 173.330 138.200 173.650 ;
        RECT 140.760 172.970 140.900 177.410 ;
        RECT 137.940 172.650 138.200 172.970 ;
        RECT 140.700 172.650 140.960 172.970 ;
        RECT 142.140 172.825 142.280 178.090 ;
        RECT 143.980 176.370 144.120 178.090 ;
        RECT 143.920 176.050 144.180 176.370 ;
        RECT 138.000 172.145 138.140 172.650 ;
        RECT 138.400 172.310 138.660 172.630 ;
        RECT 137.930 171.775 138.210 172.145 ;
        RECT 138.460 170.590 138.600 172.310 ;
        RECT 140.760 170.590 140.900 172.650 ;
        RECT 142.070 172.455 142.350 172.825 ;
        RECT 143.980 170.930 144.120 176.050 ;
        RECT 143.920 170.610 144.180 170.930 ;
        RECT 138.400 170.270 138.660 170.590 ;
        RECT 140.700 170.270 140.960 170.590 ;
        RECT 145.300 167.210 145.560 167.530 ;
        RECT 145.360 166.025 145.500 167.210 ;
        RECT 145.290 165.655 145.570 166.025 ;
        RECT 137.480 165.170 137.740 165.490 ;
        RECT 137.940 164.830 138.200 165.150 ;
        RECT 143.920 164.830 144.180 165.150 ;
        RECT 136.560 164.150 136.820 164.470 ;
        RECT 136.620 162.430 136.760 164.150 ;
        RECT 138.000 163.110 138.140 164.830 ;
        RECT 143.460 163.810 143.720 164.130 ;
        RECT 137.940 162.790 138.200 163.110 ;
        RECT 136.560 162.110 136.820 162.430 ;
        RECT 143.520 162.090 143.660 163.810 ;
        RECT 143.460 161.770 143.720 162.090 ;
        RECT 138.860 161.430 139.120 161.750 ;
        RECT 136.100 161.090 136.360 161.410 ;
        RECT 135.630 154.095 135.910 154.465 ;
        RECT 135.180 152.930 135.440 153.250 ;
        RECT 135.240 151.210 135.380 152.930 ;
        RECT 135.180 150.890 135.440 151.210 ;
        RECT 134.780 148.770 135.380 148.910 ;
        RECT 134.260 141.030 134.520 141.350 ;
        RECT 134.720 139.330 134.980 139.650 ;
        RECT 134.780 138.290 134.920 139.330 ;
        RECT 134.720 137.970 134.980 138.290 ;
        RECT 133.800 137.630 134.060 137.950 ;
        RECT 132.940 135.730 133.540 135.870 ;
        RECT 132.420 131.850 132.680 132.170 ;
        RECT 132.420 131.170 132.680 131.490 ;
        RECT 132.480 130.130 132.620 131.170 ;
        RECT 132.420 129.810 132.680 130.130 ;
        RECT 133.400 126.980 133.540 135.730 ;
        RECT 134.260 134.230 134.520 134.550 ;
        RECT 134.320 133.190 134.460 134.230 ;
        RECT 134.260 132.870 134.520 133.190 ;
        RECT 135.240 131.830 135.380 148.770 ;
        RECT 136.160 140.670 136.300 161.090 ;
        RECT 137.020 159.390 137.280 159.710 ;
        RECT 137.080 157.670 137.220 159.390 ;
        RECT 137.020 157.350 137.280 157.670 ;
        RECT 137.940 155.650 138.200 155.970 ;
        RECT 136.560 153.950 136.820 154.270 ;
        RECT 136.620 149.510 136.760 153.950 ;
        RECT 138.000 153.250 138.140 155.650 ;
        RECT 137.940 152.930 138.200 153.250 ;
        RECT 138.920 152.990 139.060 161.430 ;
        RECT 139.780 161.090 140.040 161.410 ;
        RECT 139.840 160.390 139.980 161.090 ;
        RECT 139.780 160.070 140.040 160.390 ;
        RECT 142.540 158.370 142.800 158.690 ;
        RECT 142.600 156.990 142.740 158.370 ;
        RECT 142.540 156.670 142.800 156.990 ;
        RECT 140.700 154.290 140.960 154.610 ;
        RECT 138.920 152.850 139.520 152.990 ;
        RECT 138.860 151.910 139.120 152.230 ;
        RECT 136.560 149.190 136.820 149.510 ;
        RECT 137.480 147.490 137.740 147.810 ;
        RECT 137.540 145.430 137.680 147.490 ;
        RECT 137.480 145.110 137.740 145.430 ;
        RECT 137.540 143.390 137.680 145.110 ;
        RECT 138.920 144.070 139.060 151.910 ;
        RECT 138.860 143.750 139.120 144.070 ;
        RECT 137.480 143.070 137.740 143.390 ;
        RECT 136.100 140.350 136.360 140.670 ;
        RECT 136.100 134.230 136.360 134.550 ;
        RECT 136.160 132.850 136.300 134.230 ;
        RECT 139.380 132.850 139.520 152.850 ;
        RECT 140.760 152.230 140.900 154.290 ;
        RECT 143.520 154.270 143.660 161.770 ;
        RECT 143.980 154.950 144.120 164.830 ;
        RECT 144.840 163.810 145.100 164.130 ;
        RECT 144.900 162.625 145.040 163.810 ;
        RECT 144.830 162.255 145.110 162.625 ;
        RECT 144.380 159.730 144.640 160.050 ;
        RECT 143.920 154.630 144.180 154.950 ;
        RECT 144.440 154.350 144.580 159.730 ;
        RECT 144.830 158.855 145.110 159.225 ;
        RECT 144.840 158.710 145.100 158.855 ;
        RECT 144.830 155.455 145.110 155.825 ;
        RECT 144.900 154.950 145.040 155.455 ;
        RECT 144.840 154.630 145.100 154.950 ;
        RECT 143.460 153.950 143.720 154.270 ;
        RECT 143.980 154.210 144.580 154.350 ;
        RECT 143.000 153.270 143.260 153.590 ;
        RECT 143.060 152.425 143.200 153.270 ;
        RECT 140.700 151.910 140.960 152.230 ;
        RECT 142.990 152.055 143.270 152.425 ;
        RECT 143.450 151.375 143.730 151.745 ;
        RECT 143.980 151.550 144.120 154.210 ;
        RECT 144.830 154.095 145.110 154.465 ;
        RECT 145.300 154.290 145.560 154.610 ;
        RECT 143.460 151.230 143.720 151.375 ;
        RECT 143.920 151.230 144.180 151.550 ;
        RECT 141.160 150.210 141.420 150.530 ;
        RECT 143.000 150.210 143.260 150.530 ;
        RECT 141.220 149.170 141.360 150.210 ;
        RECT 141.160 148.850 141.420 149.170 ;
        RECT 141.620 147.490 141.880 147.810 ;
        RECT 141.680 145.770 141.820 147.490 ;
        RECT 143.060 146.790 143.200 150.210 ;
        RECT 144.900 148.490 145.040 154.095 ;
        RECT 145.360 149.025 145.500 154.290 ;
        RECT 145.290 148.655 145.570 149.025 ;
        RECT 143.920 148.170 144.180 148.490 ;
        RECT 144.840 148.170 145.100 148.490 ;
        RECT 143.000 146.470 143.260 146.790 ;
        RECT 143.460 146.130 143.720 146.450 ;
        RECT 141.620 145.450 141.880 145.770 ;
        RECT 142.080 144.770 142.340 145.090 ;
        RECT 142.140 143.390 142.280 144.770 ;
        RECT 143.000 143.750 143.260 144.070 ;
        RECT 140.240 143.300 140.500 143.390 ;
        RECT 139.840 143.160 140.500 143.300 ;
        RECT 139.840 138.630 139.980 143.160 ;
        RECT 140.240 143.070 140.500 143.160 ;
        RECT 142.080 143.070 142.340 143.390 ;
        RECT 143.060 142.225 143.200 143.750 ;
        RECT 142.990 141.855 143.270 142.225 ;
        RECT 143.520 140.330 143.660 146.130 ;
        RECT 143.980 144.070 144.120 148.170 ;
        RECT 144.830 145.255 145.110 145.625 ;
        RECT 143.920 143.750 144.180 144.070 ;
        RECT 143.920 142.730 144.180 143.050 ;
        RECT 143.980 140.330 144.120 142.730 ;
        RECT 144.900 141.350 145.040 145.255 ;
        RECT 144.840 141.030 145.100 141.350 ;
        RECT 140.240 140.010 140.500 140.330 ;
        RECT 143.460 140.010 143.720 140.330 ;
        RECT 143.920 140.010 144.180 140.330 ;
        RECT 140.300 138.630 140.440 140.010 ;
        RECT 139.780 138.310 140.040 138.630 ;
        RECT 140.240 138.310 140.500 138.630 ;
        RECT 144.830 138.455 145.110 138.825 ;
        RECT 144.840 138.310 145.100 138.455 ;
        RECT 143.000 136.610 143.260 136.930 ;
        RECT 143.060 135.425 143.200 136.610 ;
        RECT 142.080 134.910 142.340 135.230 ;
        RECT 142.990 135.055 143.270 135.425 ;
        RECT 141.160 133.890 141.420 134.210 ;
        RECT 141.220 133.190 141.360 133.890 ;
        RECT 141.160 132.870 141.420 133.190 ;
        RECT 136.100 132.530 136.360 132.850 ;
        RECT 139.320 132.530 139.580 132.850 ;
        RECT 135.640 132.190 135.900 132.510 ;
        RECT 135.180 131.510 135.440 131.830 ;
        RECT 135.700 129.450 135.840 132.190 ;
        RECT 134.720 129.130 134.980 129.450 ;
        RECT 135.640 129.130 135.900 129.450 ;
        RECT 134.780 127.750 134.920 129.130 ;
        RECT 136.160 128.770 136.300 132.530 ;
        RECT 136.560 129.810 136.820 130.130 ;
        RECT 136.100 128.450 136.360 128.770 ;
        RECT 136.620 128.510 136.760 129.810 ;
        RECT 137.020 129.360 137.280 129.450 ;
        RECT 137.020 129.220 139.060 129.360 ;
        RECT 137.020 129.130 137.280 129.220 ;
        RECT 134.720 127.430 134.980 127.750 ;
        RECT 133.800 126.980 134.060 127.070 ;
        RECT 133.400 126.840 134.060 126.980 ;
        RECT 131.960 121.990 132.220 122.310 ;
        RECT 131.960 120.290 132.220 120.610 ;
        RECT 132.420 120.290 132.680 120.610 ;
        RECT 132.020 116.870 132.160 120.290 ;
        RECT 132.480 119.250 132.620 120.290 ;
        RECT 132.420 118.930 132.680 119.250 ;
        RECT 131.960 116.550 132.220 116.870 ;
        RECT 131.500 113.830 131.760 114.150 ;
        RECT 133.400 113.470 133.540 126.840 ;
        RECT 133.800 126.750 134.060 126.840 ;
        RECT 134.260 121.310 134.520 121.630 ;
        RECT 133.800 120.630 134.060 120.950 ;
        RECT 133.860 114.150 134.000 120.630 ;
        RECT 133.800 113.830 134.060 114.150 ;
        RECT 133.340 113.150 133.600 113.470 ;
        RECT 131.040 112.470 131.300 112.790 ;
        RECT 130.580 111.110 130.840 111.430 ;
        RECT 133.400 110.750 133.540 113.150 ;
        RECT 134.320 111.090 134.460 121.310 ;
        RECT 134.780 118.570 134.920 127.430 ;
        RECT 136.160 126.730 136.300 128.450 ;
        RECT 136.620 128.370 137.220 128.510 ;
        RECT 136.560 126.750 136.820 127.070 ;
        RECT 136.100 126.410 136.360 126.730 ;
        RECT 135.640 125.730 135.900 126.050 ;
        RECT 135.700 124.690 135.840 125.730 ;
        RECT 135.640 124.370 135.900 124.690 ;
        RECT 135.180 120.630 135.440 120.950 ;
        RECT 135.240 118.570 135.380 120.630 ;
        RECT 136.160 119.250 136.300 126.410 ;
        RECT 136.620 125.030 136.760 126.750 ;
        RECT 136.560 124.710 136.820 125.030 ;
        RECT 136.560 123.010 136.820 123.330 ;
        RECT 136.100 118.930 136.360 119.250 ;
        RECT 134.720 118.250 134.980 118.570 ;
        RECT 135.180 118.250 135.440 118.570 ;
        RECT 135.240 117.890 135.380 118.250 ;
        RECT 135.180 117.570 135.440 117.890 ;
        RECT 136.100 113.150 136.360 113.470 ;
        RECT 136.160 111.430 136.300 113.150 ;
        RECT 136.100 111.110 136.360 111.430 ;
        RECT 134.260 110.770 134.520 111.090 ;
        RECT 133.340 110.430 133.600 110.750 ;
        RECT 132.880 110.090 133.140 110.410 ;
        RECT 131.500 107.370 131.760 107.690 ;
        RECT 129.260 104.570 129.860 104.710 ;
        RECT 128.740 95.810 129.000 96.130 ;
        RECT 126.960 95.110 128.480 95.190 ;
        RECT 126.900 95.050 128.480 95.110 ;
        RECT 126.900 94.790 127.160 95.050 ;
        RECT 128.800 94.770 128.940 95.810 ;
        RECT 128.740 94.450 129.000 94.770 ;
        RECT 123.680 93.770 123.940 94.090 ;
        RECT 124.600 93.770 124.860 94.090 ;
        RECT 123.740 92.390 123.880 93.770 ;
        RECT 123.680 92.070 123.940 92.390 ;
        RECT 122.760 91.050 123.020 91.370 ;
        RECT 122.820 89.330 122.960 91.050 ;
        RECT 124.140 90.710 124.400 91.030 ;
        RECT 122.760 89.010 123.020 89.330 ;
        RECT 119.540 85.610 119.800 85.930 ;
        RECT 120.000 85.610 120.260 85.930 ;
        RECT 120.920 85.610 121.180 85.930 ;
        RECT 118.620 85.270 118.880 85.590 ;
        RECT 119.080 85.270 119.340 85.590 ;
        RECT 121.380 85.270 121.640 85.590 ;
        RECT 119.140 83.890 119.280 85.270 ;
        RECT 119.080 83.570 119.340 83.890 ;
        RECT 121.440 77.700 121.580 85.270 ;
        RECT 124.200 84.230 124.340 90.710 ;
        RECT 124.660 86.270 124.800 93.770 ;
        RECT 125.980 92.070 126.240 92.390 ;
        RECT 126.040 86.950 126.180 92.070 ;
        RECT 129.260 88.310 129.400 104.570 ;
        RECT 131.040 98.870 131.300 99.190 ;
        RECT 129.660 98.530 129.920 98.850 ;
        RECT 129.720 96.470 129.860 98.530 ;
        RECT 131.100 97.490 131.240 98.870 ;
        RECT 130.580 97.170 130.840 97.490 ;
        RECT 131.040 97.170 131.300 97.490 ;
        RECT 129.660 96.150 129.920 96.470 ;
        RECT 129.200 87.990 129.460 88.310 ;
        RECT 129.720 87.970 129.860 96.150 ;
        RECT 130.120 90.370 130.380 90.690 ;
        RECT 130.180 88.990 130.320 90.370 ;
        RECT 130.640 89.670 130.780 97.170 ;
        RECT 131.100 94.770 131.240 97.170 ;
        RECT 131.560 96.810 131.700 107.370 ;
        RECT 132.940 104.970 133.080 110.090 ;
        RECT 134.320 107.690 134.460 110.770 ;
        RECT 136.620 110.660 136.760 123.010 ;
        RECT 137.080 118.910 137.220 128.370 ;
        RECT 137.480 121.990 137.740 122.310 ;
        RECT 137.020 118.590 137.280 118.910 ;
        RECT 137.080 115.705 137.220 118.590 ;
        RECT 137.010 115.335 137.290 115.705 ;
        RECT 136.620 110.520 137.220 110.660 ;
        RECT 136.100 110.090 136.360 110.410 ;
        RECT 136.160 108.370 136.300 110.090 ;
        RECT 136.560 109.750 136.820 110.070 ;
        RECT 136.620 108.710 136.760 109.750 ;
        RECT 136.560 108.390 136.820 108.710 ;
        RECT 136.100 108.050 136.360 108.370 ;
        RECT 134.260 107.370 134.520 107.690 ;
        RECT 132.880 104.650 133.140 104.970 ;
        RECT 132.940 103.270 133.080 104.650 ;
        RECT 133.340 103.970 133.600 104.290 ;
        RECT 132.880 102.950 133.140 103.270 ;
        RECT 133.400 102.930 133.540 103.970 ;
        RECT 133.340 102.610 133.600 102.930 ;
        RECT 136.160 102.590 136.300 108.050 ;
        RECT 136.560 103.970 136.820 104.290 ;
        RECT 136.100 102.270 136.360 102.590 ;
        RECT 136.160 99.870 136.300 102.270 ;
        RECT 132.420 99.550 132.680 99.870 ;
        RECT 135.640 99.550 135.900 99.870 ;
        RECT 136.100 99.550 136.360 99.870 ;
        RECT 131.500 96.490 131.760 96.810 ;
        RECT 131.040 94.450 131.300 94.770 ;
        RECT 131.040 91.730 131.300 92.050 ;
        RECT 130.580 89.350 130.840 89.670 ;
        RECT 130.120 88.670 130.380 88.990 ;
        RECT 130.120 87.990 130.380 88.310 ;
        RECT 129.660 87.650 129.920 87.970 ;
        RECT 130.180 87.570 130.320 87.990 ;
        RECT 130.180 87.430 130.780 87.570 ;
        RECT 125.980 86.630 126.240 86.950 ;
        RECT 125.060 86.290 125.320 86.610 ;
        RECT 124.600 85.950 124.860 86.270 ;
        RECT 124.140 83.910 124.400 84.230 ;
        RECT 125.120 79.550 125.260 86.290 ;
        RECT 126.040 85.930 126.180 86.630 ;
        RECT 130.640 85.930 130.780 87.430 ;
        RECT 131.100 86.950 131.240 91.730 ;
        RECT 131.500 87.990 131.760 88.310 ;
        RECT 131.560 87.825 131.700 87.990 ;
        RECT 131.490 87.455 131.770 87.825 ;
        RECT 131.040 86.630 131.300 86.950 ;
        RECT 131.040 86.180 131.300 86.270 ;
        RECT 131.560 86.180 131.700 87.455 ;
        RECT 131.040 86.040 131.700 86.180 ;
        RECT 131.040 85.950 131.300 86.040 ;
        RECT 132.480 85.930 132.620 99.550 ;
        RECT 133.800 99.210 134.060 99.530 ;
        RECT 133.860 97.150 134.000 99.210 ;
        RECT 133.800 96.830 134.060 97.150 ;
        RECT 133.860 94.090 134.000 96.830 ;
        RECT 135.700 96.810 135.840 99.550 ;
        RECT 135.640 96.490 135.900 96.810 ;
        RECT 133.800 93.770 134.060 94.090 ;
        RECT 133.340 93.090 133.600 93.410 ;
        RECT 132.880 90.370 133.140 90.690 ;
        RECT 132.940 89.670 133.080 90.370 ;
        RECT 133.400 89.670 133.540 93.090 ;
        RECT 133.860 91.710 134.000 93.770 ;
        RECT 136.160 93.750 136.300 99.550 ;
        RECT 136.620 99.190 136.760 103.970 ;
        RECT 136.560 98.870 136.820 99.190 ;
        RECT 137.080 97.910 137.220 110.520 ;
        RECT 137.540 107.690 137.680 121.990 ;
        RECT 138.400 120.970 138.660 121.290 ;
        RECT 138.460 115.510 138.600 120.970 ;
        RECT 138.400 115.190 138.660 115.510 ;
        RECT 137.480 107.370 137.740 107.690 ;
        RECT 137.540 105.990 137.680 107.370 ;
        RECT 137.480 105.670 137.740 105.990 ;
        RECT 137.540 105.310 137.680 105.670 ;
        RECT 137.480 104.990 137.740 105.310 ;
        RECT 137.940 104.650 138.200 104.970 ;
        RECT 138.000 101.570 138.140 104.650 ;
        RECT 137.940 101.250 138.200 101.570 ;
        RECT 137.080 97.770 137.680 97.910 ;
        RECT 136.560 97.170 136.820 97.490 ;
        RECT 136.620 95.110 136.760 97.170 ;
        RECT 137.020 96.830 137.280 97.150 ;
        RECT 136.560 94.790 136.820 95.110 ;
        RECT 136.100 93.430 136.360 93.750 ;
        RECT 136.160 92.390 136.300 93.430 ;
        RECT 136.100 92.070 136.360 92.390 ;
        RECT 136.160 91.790 136.300 92.070 ;
        RECT 133.800 91.390 134.060 91.710 ;
        RECT 136.160 91.650 136.760 91.790 ;
        RECT 132.880 89.350 133.140 89.670 ;
        RECT 133.340 89.350 133.600 89.670 ;
        RECT 125.980 85.610 126.240 85.930 ;
        RECT 130.580 85.610 130.840 85.930 ;
        RECT 132.420 85.610 132.680 85.930 ;
        RECT 131.040 85.270 131.300 85.590 ;
        RECT 127.820 80.170 128.080 80.490 ;
        RECT 124.660 79.410 125.260 79.550 ;
        RECT 124.660 77.700 124.800 79.410 ;
        RECT 127.880 77.700 128.020 80.170 ;
        RECT 131.100 77.700 131.240 85.270 ;
        RECT 132.940 85.250 133.080 89.350 ;
        RECT 133.860 88.310 134.000 91.390 ;
        RECT 135.180 89.350 135.440 89.670 ;
        RECT 133.800 87.990 134.060 88.310 ;
        RECT 135.240 85.930 135.380 89.350 ;
        RECT 136.620 88.990 136.760 91.650 ;
        RECT 137.080 91.370 137.220 96.830 ;
        RECT 137.540 95.110 137.680 97.770 ;
        RECT 138.000 96.810 138.140 101.250 ;
        RECT 137.940 96.490 138.200 96.810 ;
        RECT 138.400 96.150 138.660 96.470 ;
        RECT 138.460 95.110 138.600 96.150 ;
        RECT 137.480 94.790 137.740 95.110 ;
        RECT 138.400 94.790 138.660 95.110 ;
        RECT 137.540 93.830 137.680 94.790 ;
        RECT 137.540 93.690 138.140 93.830 ;
        RECT 137.480 93.090 137.740 93.410 ;
        RECT 137.020 91.050 137.280 91.370 ;
        RECT 136.100 88.670 136.360 88.990 ;
        RECT 136.560 88.670 136.820 88.990 ;
        RECT 135.180 85.785 135.440 85.930 ;
        RECT 135.170 85.415 135.450 85.785 ;
        RECT 135.640 85.610 135.900 85.930 ;
        RECT 132.880 84.930 133.140 85.250 ;
        RECT 135.700 83.890 135.840 85.610 ;
        RECT 135.640 83.570 135.900 83.890 ;
        RECT 136.160 80.490 136.300 88.670 ;
        RECT 136.560 88.220 136.820 88.310 ;
        RECT 136.560 88.080 137.220 88.220 ;
        RECT 136.560 87.990 136.820 88.080 ;
        RECT 136.550 87.455 136.830 87.825 ;
        RECT 136.620 85.930 136.760 87.455 ;
        RECT 136.560 85.610 136.820 85.930 ;
        RECT 137.080 85.840 137.220 88.080 ;
        RECT 137.540 86.610 137.680 93.090 ;
        RECT 138.000 90.690 138.140 93.690 ;
        RECT 137.940 90.370 138.200 90.690 ;
        RECT 138.920 86.950 139.060 129.220 ;
        RECT 139.380 123.330 139.520 132.530 ;
        RECT 142.140 132.510 142.280 134.910 ;
        RECT 142.080 132.190 142.340 132.510 ;
        RECT 140.700 131.850 140.960 132.170 ;
        RECT 140.760 126.050 140.900 131.850 ;
        RECT 144.380 131.510 144.640 131.830 ;
        RECT 144.830 131.655 145.110 132.025 ;
        RECT 144.840 131.510 145.100 131.655 ;
        RECT 144.440 130.470 144.580 131.510 ;
        RECT 144.380 130.150 144.640 130.470 ;
        RECT 144.440 127.070 144.580 130.150 ;
        RECT 144.830 128.255 145.110 128.625 ;
        RECT 144.900 127.750 145.040 128.255 ;
        RECT 144.840 127.430 145.100 127.750 ;
        RECT 144.380 126.750 144.640 127.070 ;
        RECT 143.920 126.070 144.180 126.390 ;
        RECT 140.700 125.730 140.960 126.050 ;
        RECT 139.320 123.010 139.580 123.330 ;
        RECT 140.760 121.290 140.900 125.730 ;
        RECT 143.980 124.010 144.120 126.070 ;
        RECT 144.830 124.855 145.110 125.225 ;
        RECT 144.840 124.710 145.100 124.855 ;
        RECT 142.080 123.690 142.340 124.010 ;
        RECT 143.920 123.690 144.180 124.010 ;
        RECT 142.140 121.970 142.280 123.690 ;
        RECT 143.000 123.010 143.260 123.330 ;
        RECT 142.080 121.650 142.340 121.970 ;
        RECT 143.060 121.825 143.200 123.010 ;
        RECT 142.990 121.455 143.270 121.825 ;
        RECT 140.700 120.970 140.960 121.290 ;
        RECT 140.700 118.250 140.960 118.570 ;
        RECT 139.320 115.190 139.580 115.510 ;
        RECT 139.380 112.790 139.520 115.190 ;
        RECT 139.780 113.150 140.040 113.470 ;
        RECT 139.320 112.470 139.580 112.790 ;
        RECT 139.320 109.470 139.580 109.730 ;
        RECT 139.840 109.470 139.980 113.150 ;
        RECT 139.320 109.410 139.980 109.470 ;
        RECT 139.380 109.330 139.980 109.410 ;
        RECT 139.840 108.030 139.980 109.330 ;
        RECT 139.780 107.710 140.040 108.030 ;
        RECT 139.840 105.990 139.980 107.710 ;
        RECT 140.760 107.010 140.900 118.250 ;
        RECT 144.830 118.055 145.110 118.425 ;
        RECT 143.920 117.570 144.180 117.890 ;
        RECT 143.000 115.190 143.260 115.510 ;
        RECT 143.060 115.025 143.200 115.190 ;
        RECT 142.990 114.655 143.270 115.025 ;
        RECT 141.620 113.490 141.880 113.810 ;
        RECT 141.680 107.690 141.820 113.490 ;
        RECT 143.980 113.130 144.120 117.570 ;
        RECT 144.900 116.870 145.040 118.055 ;
        RECT 144.840 116.550 145.100 116.870 ;
        RECT 143.920 112.810 144.180 113.130 ;
        RECT 142.540 112.130 142.800 112.450 ;
        RECT 143.000 112.130 143.260 112.450 ;
        RECT 144.840 112.130 145.100 112.450 ;
        RECT 142.600 107.690 142.740 112.130 ;
        RECT 143.060 108.225 143.200 112.130 ;
        RECT 144.900 111.625 145.040 112.130 ;
        RECT 144.830 111.255 145.110 111.625 ;
        RECT 144.380 109.410 144.640 109.730 ;
        RECT 142.990 107.855 143.270 108.225 ;
        RECT 144.440 108.030 144.580 109.410 ;
        RECT 144.380 107.710 144.640 108.030 ;
        RECT 141.620 107.370 141.880 107.690 ;
        RECT 142.540 107.370 142.800 107.690 ;
        RECT 143.460 107.370 143.720 107.690 ;
        RECT 140.700 106.690 140.960 107.010 ;
        RECT 141.160 106.690 141.420 107.010 ;
        RECT 139.780 105.670 140.040 105.990 ;
        RECT 139.780 104.650 140.040 104.970 ;
        RECT 139.320 104.310 139.580 104.630 ;
        RECT 139.380 94.090 139.520 104.310 ;
        RECT 139.320 93.770 139.580 94.090 ;
        RECT 139.840 93.750 139.980 104.650 ;
        RECT 141.220 96.130 141.360 106.690 ;
        RECT 141.160 95.810 141.420 96.130 ;
        RECT 141.680 94.340 141.820 107.370 ;
        RECT 143.520 105.650 143.660 107.370 ;
        RECT 143.460 105.330 143.720 105.650 ;
        RECT 142.080 104.650 142.340 104.970 ;
        RECT 142.140 100.550 142.280 104.650 ;
        RECT 142.540 101.990 142.800 102.250 ;
        RECT 142.540 101.930 143.200 101.990 ;
        RECT 142.600 101.850 143.200 101.930 ;
        RECT 142.080 100.230 142.340 100.550 ;
        RECT 142.140 96.810 142.280 100.230 ;
        RECT 142.080 96.490 142.340 96.810 ;
        RECT 142.080 94.340 142.340 94.430 ;
        RECT 141.680 94.200 142.340 94.340 ;
        RECT 142.080 94.110 142.340 94.200 ;
        RECT 139.780 93.430 140.040 93.750 ;
        RECT 141.160 93.430 141.420 93.750 ;
        RECT 139.840 89.670 139.980 93.430 ;
        RECT 141.220 92.390 141.360 93.430 ;
        RECT 141.160 92.070 141.420 92.390 ;
        RECT 139.780 89.350 140.040 89.670 ;
        RECT 141.220 89.330 141.360 92.070 ;
        RECT 141.620 90.370 141.880 90.690 ;
        RECT 141.160 89.010 141.420 89.330 ;
        RECT 139.780 88.670 140.040 88.990 ;
        RECT 139.840 86.950 139.980 88.670 ;
        RECT 140.230 87.455 140.510 87.825 ;
        RECT 138.860 86.630 139.120 86.950 ;
        RECT 139.780 86.630 140.040 86.950 ;
        RECT 137.480 86.290 137.740 86.610 ;
        RECT 138.400 85.950 138.660 86.270 ;
        RECT 137.480 85.840 137.740 85.930 ;
        RECT 137.080 85.700 137.740 85.840 ;
        RECT 137.480 85.610 137.740 85.700 ;
        RECT 136.100 80.170 136.360 80.490 ;
        RECT 138.460 79.550 138.600 85.950 ;
        RECT 140.300 85.930 140.440 87.455 ;
        RECT 141.680 86.610 141.820 90.370 ;
        RECT 141.620 86.290 141.880 86.610 ;
        RECT 143.060 85.930 143.200 101.850 ;
        RECT 143.520 99.870 143.660 105.330 ;
        RECT 144.440 105.310 144.580 107.710 ;
        RECT 145.300 105.670 145.560 105.990 ;
        RECT 144.380 104.990 144.640 105.310 ;
        RECT 144.830 104.455 145.110 104.825 ;
        RECT 144.840 104.310 145.100 104.455 ;
        RECT 144.840 101.425 145.100 101.570 ;
        RECT 144.830 101.055 145.110 101.425 ;
        RECT 143.460 99.550 143.720 99.870 ;
        RECT 144.840 98.530 145.100 98.850 ;
        RECT 144.900 98.025 145.040 98.530 ;
        RECT 144.830 97.655 145.110 98.025 ;
        RECT 143.920 94.110 144.180 94.430 ;
        RECT 143.980 90.690 144.120 94.110 ;
        RECT 144.380 93.090 144.640 93.410 ;
        RECT 143.920 90.370 144.180 90.690 ;
        RECT 143.980 89.670 144.120 90.370 ;
        RECT 143.920 89.350 144.180 89.670 ;
        RECT 144.440 87.570 144.580 93.090 ;
        RECT 145.360 91.710 145.500 105.670 ;
        RECT 147.140 96.150 147.400 96.470 ;
        RECT 145.300 91.390 145.560 91.710 ;
        RECT 144.840 87.650 145.100 87.970 ;
        RECT 143.980 87.430 144.580 87.570 ;
        RECT 140.240 85.610 140.500 85.930 ;
        RECT 142.080 85.785 142.340 85.930 ;
        RECT 142.070 85.415 142.350 85.785 ;
        RECT 143.000 85.610 143.260 85.930 ;
        RECT 143.000 84.930 143.260 85.250 ;
        RECT 140.700 79.830 140.960 80.150 ;
        RECT 134.260 79.150 134.520 79.470 ;
        RECT 137.540 79.410 138.600 79.550 ;
        RECT 134.320 77.700 134.460 79.150 ;
        RECT 137.540 77.700 137.680 79.410 ;
        RECT 140.760 77.700 140.900 79.830 ;
        RECT 143.060 79.470 143.200 84.930 ;
        RECT 143.000 79.150 143.260 79.470 ;
        RECT 143.980 77.700 144.120 87.430 ;
        RECT 144.900 80.150 145.040 87.650 ;
        RECT 144.840 79.830 145.100 80.150 ;
        RECT 147.200 77.700 147.340 96.150 ;
        RECT 150.360 95.810 150.620 96.130 ;
        RECT 150.420 77.700 150.560 95.810 ;
        RECT 11.890 73.700 12.170 77.700 ;
        RECT 15.110 73.700 15.390 77.700 ;
        RECT 18.330 73.700 18.610 77.700 ;
        RECT 21.550 73.700 21.830 77.700 ;
        RECT 24.770 73.700 25.050 77.700 ;
        RECT 27.990 73.700 28.270 77.700 ;
        RECT 31.210 73.700 31.490 77.700 ;
        RECT 34.430 73.700 34.710 77.700 ;
        RECT 37.650 73.700 37.930 77.700 ;
        RECT 40.870 73.700 41.150 77.700 ;
        RECT 44.090 73.700 44.370 77.700 ;
        RECT 47.310 73.700 47.590 77.700 ;
        RECT 50.530 73.700 50.810 77.700 ;
        RECT 53.750 73.700 54.030 77.700 ;
        RECT 56.970 73.700 57.250 77.700 ;
        RECT 60.190 73.700 60.470 77.700 ;
        RECT 63.410 73.700 63.690 77.700 ;
        RECT 66.630 73.700 66.910 77.700 ;
        RECT 69.850 73.700 70.130 77.700 ;
        RECT 73.070 73.700 73.350 77.700 ;
        RECT 76.290 73.700 76.570 77.700 ;
        RECT 79.510 73.700 79.790 77.700 ;
        RECT 82.730 73.700 83.010 77.700 ;
        RECT 85.950 73.700 86.230 77.700 ;
        RECT 89.170 73.700 89.450 77.700 ;
        RECT 92.390 73.700 92.670 77.700 ;
        RECT 95.610 73.700 95.890 77.700 ;
        RECT 98.830 73.700 99.110 77.700 ;
        RECT 102.050 73.700 102.330 77.700 ;
        RECT 105.270 73.700 105.550 77.700 ;
        RECT 108.490 73.700 108.770 77.700 ;
        RECT 111.710 73.700 111.990 77.700 ;
        RECT 114.930 73.700 115.210 77.700 ;
        RECT 118.150 73.700 118.430 77.700 ;
        RECT 121.370 73.700 121.650 77.700 ;
        RECT 124.590 73.700 124.870 77.700 ;
        RECT 127.810 73.700 128.090 77.700 ;
        RECT 131.030 73.700 131.310 77.700 ;
        RECT 134.250 73.700 134.530 77.700 ;
        RECT 137.470 73.700 137.750 77.700 ;
        RECT 140.690 73.700 140.970 77.700 ;
        RECT 143.910 73.700 144.190 77.700 ;
        RECT 147.130 73.700 147.410 77.700 ;
        RECT 150.350 73.700 150.630 77.700 ;
      LAYER met3 ;
        RECT 32.850 212.255 34.430 212.585 ;
        RECT 36.150 209.535 37.730 209.865 ;
        RECT 32.850 206.815 34.430 207.145 ;
        RECT 36.150 204.095 37.730 204.425 ;
        RECT 32.850 201.375 34.430 201.705 ;
        RECT 36.150 198.655 37.730 198.985 ;
        RECT 32.850 195.935 34.430 196.265 ;
        RECT 36.150 193.215 37.730 193.545 ;
        RECT 96.965 192.510 97.295 192.525 ;
        RECT 102.485 192.510 102.815 192.525 ;
        RECT 96.965 192.210 102.815 192.510 ;
        RECT 96.965 192.195 97.295 192.210 ;
        RECT 102.485 192.195 102.815 192.210 ;
        RECT 39.005 191.150 39.335 191.165 ;
        RECT 52.345 191.150 52.675 191.165 ;
        RECT 65.685 191.150 66.015 191.165 ;
        RECT 39.005 190.850 66.015 191.150 ;
        RECT 39.005 190.835 39.335 190.850 ;
        RECT 52.345 190.835 52.675 190.850 ;
        RECT 65.685 190.835 66.015 190.850 ;
        RECT 32.850 190.495 34.430 190.825 ;
        RECT 11.800 189.790 15.800 189.940 ;
        RECT 18.765 189.790 19.095 189.805 ;
        RECT 11.800 189.490 19.095 189.790 ;
        RECT 11.800 189.340 15.800 189.490 ;
        RECT 18.765 189.475 19.095 189.490 ;
        RECT 90.525 189.790 90.855 189.805 ;
        RECT 101.105 189.790 101.435 189.805 ;
        RECT 105.705 189.790 106.035 189.805 ;
        RECT 90.525 189.490 106.035 189.790 ;
        RECT 90.525 189.475 90.855 189.490 ;
        RECT 101.105 189.475 101.435 189.490 ;
        RECT 105.705 189.475 106.035 189.490 ;
        RECT 96.045 189.110 96.375 189.125 ;
        RECT 105.245 189.110 105.575 189.125 ;
        RECT 96.045 188.810 105.575 189.110 ;
        RECT 96.045 188.795 96.375 188.810 ;
        RECT 105.245 188.795 105.575 188.810 ;
        RECT 36.150 187.775 37.730 188.105 ;
        RECT 32.850 185.055 34.430 185.385 ;
        RECT 36.150 182.335 37.730 182.665 ;
        RECT 32.850 179.615 34.430 179.945 ;
        RECT 36.150 176.895 37.730 177.225 ;
        RECT 131.925 176.190 132.255 176.205 ;
        RECT 134.685 176.190 135.015 176.205 ;
        RECT 131.925 175.890 135.015 176.190 ;
        RECT 131.925 175.875 132.255 175.890 ;
        RECT 134.685 175.875 135.015 175.890 ;
        RECT 32.850 174.175 34.430 174.505 ;
        RECT 128.705 172.790 129.035 172.805 ;
        RECT 142.045 172.790 142.375 172.805 ;
        RECT 128.705 172.490 142.375 172.790 ;
        RECT 128.705 172.475 129.035 172.490 ;
        RECT 142.045 172.475 142.375 172.490 ;
        RECT 130.545 172.110 130.875 172.125 ;
        RECT 137.905 172.110 138.235 172.125 ;
        RECT 130.545 171.810 138.235 172.110 ;
        RECT 130.545 171.795 130.875 171.810 ;
        RECT 137.905 171.795 138.235 171.810 ;
        RECT 36.150 171.455 37.730 171.785 ;
        RECT 118.585 170.750 118.915 170.765 ;
        RECT 133.305 170.750 133.635 170.765 ;
        RECT 118.585 170.450 133.635 170.750 ;
        RECT 118.585 170.435 118.915 170.450 ;
        RECT 133.305 170.435 133.635 170.450 ;
        RECT 119.505 170.070 119.835 170.085 ;
        RECT 131.005 170.070 131.335 170.085 ;
        RECT 119.505 169.770 131.335 170.070 ;
        RECT 119.505 169.755 119.835 169.770 ;
        RECT 131.005 169.755 131.335 169.770 ;
        RECT 107.545 169.400 107.875 169.405 ;
        RECT 107.545 169.390 108.130 169.400 ;
        RECT 129.625 169.390 129.955 169.405 ;
        RECT 132.385 169.390 132.715 169.405 ;
        RECT 107.545 169.090 108.330 169.390 ;
        RECT 129.625 169.090 132.715 169.390 ;
        RECT 107.545 169.080 108.130 169.090 ;
        RECT 107.545 169.075 107.875 169.080 ;
        RECT 129.625 169.075 129.955 169.090 ;
        RECT 132.385 169.075 132.715 169.090 ;
        RECT 32.850 168.735 34.430 169.065 ;
        RECT 108.005 168.710 108.335 168.725 ;
        RECT 107.790 168.395 108.335 168.710 ;
        RECT 125.945 168.710 126.275 168.725 ;
        RECT 136.525 168.710 136.855 168.725 ;
        RECT 125.945 168.410 136.855 168.710 ;
        RECT 125.945 168.395 126.275 168.410 ;
        RECT 136.525 168.395 136.855 168.410 ;
        RECT 107.790 167.365 108.090 168.395 ;
        RECT 120.425 168.030 120.755 168.045 ;
        RECT 123.645 168.030 123.975 168.045 ;
        RECT 132.845 168.030 133.175 168.045 ;
        RECT 120.425 167.730 133.175 168.030 ;
        RECT 120.425 167.715 120.755 167.730 ;
        RECT 123.645 167.715 123.975 167.730 ;
        RECT 132.845 167.715 133.175 167.730 ;
        RECT 107.790 167.050 108.335 167.365 ;
        RECT 108.005 167.035 108.335 167.050 ;
        RECT 105.245 166.670 105.575 166.685 ;
        RECT 110.305 166.670 110.635 166.685 ;
        RECT 105.245 166.370 110.635 166.670 ;
        RECT 105.245 166.355 105.575 166.370 ;
        RECT 110.305 166.355 110.635 166.370 ;
        RECT 36.150 166.015 37.730 166.345 ;
        RECT 145.265 165.990 145.595 166.005 ;
        RECT 148.805 165.990 152.805 166.140 ;
        RECT 145.265 165.690 152.805 165.990 ;
        RECT 145.265 165.675 145.595 165.690 ;
        RECT 148.805 165.540 152.805 165.690 ;
        RECT 131.005 165.310 131.335 165.325 ;
        RECT 133.305 165.310 133.635 165.325 ;
        RECT 131.005 165.010 133.635 165.310 ;
        RECT 131.005 164.995 131.335 165.010 ;
        RECT 133.305 164.995 133.635 165.010 ;
        RECT 131.925 164.630 132.255 164.645 ;
        RECT 132.590 164.630 132.970 164.640 ;
        RECT 131.925 164.330 132.970 164.630 ;
        RECT 131.925 164.315 132.255 164.330 ;
        RECT 132.590 164.320 132.970 164.330 ;
        RECT 32.850 163.295 34.430 163.625 ;
        RECT 124.105 162.590 124.435 162.605 ;
        RECT 127.785 162.590 128.115 162.605 ;
        RECT 124.105 162.290 128.115 162.590 ;
        RECT 124.105 162.275 124.435 162.290 ;
        RECT 127.785 162.275 128.115 162.290 ;
        RECT 144.805 162.590 145.135 162.605 ;
        RECT 148.805 162.590 152.805 162.740 ;
        RECT 144.805 162.290 152.805 162.590 ;
        RECT 144.805 162.275 145.135 162.290 ;
        RECT 148.805 162.140 152.805 162.290 ;
        RECT 36.150 160.575 37.730 160.905 ;
        RECT 88.225 159.870 88.555 159.885 ;
        RECT 99.725 159.870 100.055 159.885 ;
        RECT 88.225 159.570 100.055 159.870 ;
        RECT 88.225 159.555 88.555 159.570 ;
        RECT 99.725 159.555 100.055 159.570 ;
        RECT 144.805 159.190 145.135 159.205 ;
        RECT 148.805 159.190 152.805 159.340 ;
        RECT 144.805 158.890 152.805 159.190 ;
        RECT 144.805 158.875 145.135 158.890 ;
        RECT 148.805 158.740 152.805 158.890 ;
        RECT 121.345 158.510 121.675 158.525 ;
        RECT 132.385 158.510 132.715 158.525 ;
        RECT 121.345 158.210 132.715 158.510 ;
        RECT 121.345 158.195 121.675 158.210 ;
        RECT 132.385 158.195 132.715 158.210 ;
        RECT 32.850 157.855 34.430 158.185 ;
        RECT 112.605 157.150 112.935 157.165 ;
        RECT 119.045 157.150 119.375 157.165 ;
        RECT 125.945 157.150 126.275 157.165 ;
        RECT 132.385 157.160 132.715 157.165 ;
        RECT 132.385 157.150 132.970 157.160 ;
        RECT 112.605 156.850 132.970 157.150 ;
        RECT 112.605 156.835 112.935 156.850 ;
        RECT 119.045 156.835 119.375 156.850 ;
        RECT 125.945 156.835 126.275 156.850 ;
        RECT 132.385 156.840 132.970 156.850 ;
        RECT 132.385 156.835 132.715 156.840 ;
        RECT 116.285 155.800 116.615 155.805 ;
        RECT 116.030 155.790 116.615 155.800 ;
        RECT 115.830 155.490 116.615 155.790 ;
        RECT 116.030 155.480 116.615 155.490 ;
        RECT 116.285 155.475 116.615 155.480 ;
        RECT 144.805 155.790 145.135 155.805 ;
        RECT 148.805 155.790 152.805 155.940 ;
        RECT 144.805 155.490 152.805 155.790 ;
        RECT 144.805 155.475 145.135 155.490 ;
        RECT 36.150 155.135 37.730 155.465 ;
        RECT 148.805 155.340 152.805 155.490 ;
        RECT 130.545 154.430 130.875 154.445 ;
        RECT 135.605 154.430 135.935 154.445 ;
        RECT 144.805 154.430 145.135 154.445 ;
        RECT 130.545 154.130 145.135 154.430 ;
        RECT 130.545 154.115 130.875 154.130 ;
        RECT 135.605 154.115 135.935 154.130 ;
        RECT 144.805 154.115 145.135 154.130 ;
        RECT 116.285 153.750 116.615 153.765 ;
        RECT 120.425 153.750 120.755 153.765 ;
        RECT 131.005 153.750 131.335 153.765 ;
        RECT 116.285 153.450 131.335 153.750 ;
        RECT 116.285 153.435 116.615 153.450 ;
        RECT 120.425 153.435 120.755 153.450 ;
        RECT 131.005 153.435 131.335 153.450 ;
        RECT 16.005 153.070 16.335 153.085 ;
        RECT 15.790 152.755 16.335 153.070 ;
        RECT 15.790 152.540 16.090 152.755 ;
        RECT 11.800 152.090 16.090 152.540 ;
        RECT 32.850 152.415 34.430 152.745 ;
        RECT 108.005 152.400 108.335 152.405 ;
        RECT 107.750 152.390 108.335 152.400 ;
        RECT 107.550 152.090 108.335 152.390 ;
        RECT 11.800 151.940 15.800 152.090 ;
        RECT 107.750 152.080 108.335 152.090 ;
        RECT 108.005 152.075 108.335 152.080 ;
        RECT 142.965 152.390 143.295 152.405 ;
        RECT 148.805 152.390 152.805 152.540 ;
        RECT 142.965 152.090 152.805 152.390 ;
        RECT 142.965 152.075 143.295 152.090 ;
        RECT 148.805 151.940 152.805 152.090 ;
        RECT 119.045 151.710 119.375 151.725 ;
        RECT 143.425 151.710 143.755 151.725 ;
        RECT 119.045 151.410 143.755 151.710 ;
        RECT 119.045 151.395 119.375 151.410 ;
        RECT 143.425 151.395 143.755 151.410 ;
        RECT 122.265 150.360 122.595 150.365 ;
        RECT 122.265 150.350 122.850 150.360 ;
        RECT 122.265 150.050 123.050 150.350 ;
        RECT 122.265 150.040 122.850 150.050 ;
        RECT 122.265 150.035 122.595 150.040 ;
        RECT 11.780 149.580 15.780 149.710 ;
        RECT 36.150 149.695 37.730 150.025 ;
        RECT 11.780 149.110 16.330 149.580 ;
        RECT 14.990 149.080 16.330 149.110 ;
        RECT 121.345 148.990 121.675 149.005 ;
        RECT 130.085 148.990 130.415 149.005 ;
        RECT 121.345 148.690 130.415 148.990 ;
        RECT 121.345 148.675 121.675 148.690 ;
        RECT 130.085 148.675 130.415 148.690 ;
        RECT 145.265 148.990 145.595 149.005 ;
        RECT 148.805 148.990 152.805 149.140 ;
        RECT 145.265 148.690 152.805 148.990 ;
        RECT 145.265 148.675 145.595 148.690 ;
        RECT 148.805 148.540 152.805 148.690 ;
        RECT 32.850 146.975 34.430 147.305 ;
        RECT 144.805 145.590 145.135 145.605 ;
        RECT 148.805 145.590 152.805 145.740 ;
        RECT 144.805 145.290 152.805 145.590 ;
        RECT 144.805 145.275 145.135 145.290 ;
        RECT 148.805 145.140 152.805 145.290 ;
        RECT 36.150 144.255 37.730 144.585 ;
        RECT 115.825 142.880 116.155 142.885 ;
        RECT 115.825 142.870 116.410 142.880 ;
        RECT 115.600 142.570 116.410 142.870 ;
        RECT 115.825 142.560 116.410 142.570 ;
        RECT 115.825 142.555 116.155 142.560 ;
        RECT 142.965 142.190 143.295 142.205 ;
        RECT 148.805 142.190 152.805 142.340 ;
        RECT 142.965 141.890 152.805 142.190 ;
        RECT 142.965 141.875 143.295 141.890 ;
        RECT 32.850 141.535 34.430 141.865 ;
        RECT 148.805 141.740 152.805 141.890 ;
        RECT 36.150 138.815 37.730 139.145 ;
        RECT 144.805 138.790 145.135 138.805 ;
        RECT 148.805 138.790 152.805 138.940 ;
        RECT 144.805 138.490 152.805 138.790 ;
        RECT 144.805 138.475 145.135 138.490 ;
        RECT 148.805 138.340 152.805 138.490 ;
        RECT 32.850 136.095 34.430 136.425 ;
        RECT 11.800 135.390 15.800 135.540 ;
        RECT 19.225 135.390 19.555 135.405 ;
        RECT 11.800 135.090 19.555 135.390 ;
        RECT 11.800 134.940 15.800 135.090 ;
        RECT 19.225 135.075 19.555 135.090 ;
        RECT 142.965 135.390 143.295 135.405 ;
        RECT 148.805 135.390 152.805 135.540 ;
        RECT 142.965 135.090 152.805 135.390 ;
        RECT 142.965 135.075 143.295 135.090 ;
        RECT 148.805 134.940 152.805 135.090 ;
        RECT 36.150 133.375 37.730 133.705 ;
        RECT 16.005 132.670 16.335 132.685 ;
        RECT 15.790 132.355 16.335 132.670 ;
        RECT 15.790 132.140 16.090 132.355 ;
        RECT 11.800 131.690 16.090 132.140 ;
        RECT 144.805 131.990 145.135 132.005 ;
        RECT 148.805 131.990 152.805 132.140 ;
        RECT 144.805 131.690 152.805 131.990 ;
        RECT 11.800 131.540 15.800 131.690 ;
        RECT 144.805 131.675 145.135 131.690 ;
        RECT 148.805 131.540 152.805 131.690 ;
        RECT 32.850 130.655 34.430 130.985 ;
        RECT 11.800 128.590 15.800 128.740 ;
        RECT 16.465 128.590 16.795 128.605 ;
        RECT 11.800 128.290 16.795 128.590 ;
        RECT 11.800 128.140 15.800 128.290 ;
        RECT 16.465 128.275 16.795 128.290 ;
        RECT 144.805 128.590 145.135 128.605 ;
        RECT 148.805 128.590 152.805 128.740 ;
        RECT 144.805 128.290 152.805 128.590 ;
        RECT 144.805 128.275 145.135 128.290 ;
        RECT 36.150 127.935 37.730 128.265 ;
        RECT 148.805 128.140 152.805 128.290 ;
        RECT 16.005 125.870 16.335 125.885 ;
        RECT 15.790 125.555 16.335 125.870 ;
        RECT 15.790 125.340 16.090 125.555 ;
        RECT 11.800 124.890 16.090 125.340 ;
        RECT 32.850 125.215 34.430 125.545 ;
        RECT 144.805 125.190 145.135 125.205 ;
        RECT 148.805 125.190 152.805 125.340 ;
        RECT 144.805 124.890 152.805 125.190 ;
        RECT 11.800 124.740 15.800 124.890 ;
        RECT 144.805 124.875 145.135 124.890 ;
        RECT 148.805 124.740 152.805 124.890 ;
        RECT 36.150 122.495 37.730 122.825 ;
        RECT 11.800 121.790 15.800 121.940 ;
        RECT 111.225 121.790 111.555 121.805 ;
        RECT 129.165 121.790 129.495 121.805 ;
        RECT 11.800 121.340 16.090 121.790 ;
        RECT 111.225 121.490 129.495 121.790 ;
        RECT 111.225 121.475 111.555 121.490 ;
        RECT 129.165 121.475 129.495 121.490 ;
        RECT 142.965 121.790 143.295 121.805 ;
        RECT 148.805 121.790 152.805 121.940 ;
        RECT 142.965 121.490 152.805 121.790 ;
        RECT 142.965 121.475 143.295 121.490 ;
        RECT 148.805 121.340 152.805 121.490 ;
        RECT 15.790 121.125 16.090 121.340 ;
        RECT 15.790 120.810 16.335 121.125 ;
        RECT 16.005 120.795 16.335 120.810 ;
        RECT 32.850 119.775 34.430 120.105 ;
        RECT 16.005 119.070 16.335 119.085 ;
        RECT 15.790 118.755 16.335 119.070 ;
        RECT 15.790 118.540 16.090 118.755 ;
        RECT 11.800 118.090 16.090 118.540 ;
        RECT 113.525 118.390 113.855 118.405 ;
        RECT 122.470 118.390 122.850 118.400 ;
        RECT 113.525 118.090 122.850 118.390 ;
        RECT 11.800 117.940 15.800 118.090 ;
        RECT 113.525 118.075 113.855 118.090 ;
        RECT 122.470 118.080 122.850 118.090 ;
        RECT 144.805 118.390 145.135 118.405 ;
        RECT 148.805 118.390 152.805 118.540 ;
        RECT 144.805 118.090 152.805 118.390 ;
        RECT 144.805 118.075 145.135 118.090 ;
        RECT 148.805 117.940 152.805 118.090 ;
        RECT 36.150 117.055 37.730 117.385 ;
        RECT 108.465 115.670 108.795 115.685 ;
        RECT 136.985 115.670 137.315 115.685 ;
        RECT 108.465 115.370 137.315 115.670 ;
        RECT 108.465 115.355 108.795 115.370 ;
        RECT 136.985 115.355 137.315 115.370 ;
        RECT 11.800 114.990 15.800 115.140 ;
        RECT 21.065 114.990 21.395 115.005 ;
        RECT 11.800 114.690 21.395 114.990 ;
        RECT 11.800 114.540 15.800 114.690 ;
        RECT 21.065 114.675 21.395 114.690 ;
        RECT 142.965 114.990 143.295 115.005 ;
        RECT 148.805 114.990 152.805 115.140 ;
        RECT 142.965 114.690 152.805 114.990 ;
        RECT 142.965 114.675 143.295 114.690 ;
        RECT 32.850 114.335 34.430 114.665 ;
        RECT 148.805 114.540 152.805 114.690 ;
        RECT 11.800 111.590 15.800 111.740 ;
        RECT 36.150 111.615 37.730 111.945 ;
        RECT 144.805 111.590 145.135 111.605 ;
        RECT 148.805 111.590 152.805 111.740 ;
        RECT 11.800 111.140 16.090 111.590 ;
        RECT 144.805 111.290 152.805 111.590 ;
        RECT 144.805 111.275 145.135 111.290 ;
        RECT 148.805 111.140 152.805 111.290 ;
        RECT 15.790 110.925 16.090 111.140 ;
        RECT 15.790 110.610 16.335 110.925 ;
        RECT 16.005 110.595 16.335 110.610 ;
        RECT 32.850 108.895 34.430 109.225 ;
        RECT 11.800 108.190 15.800 108.340 ;
        RECT 20.145 108.190 20.475 108.205 ;
        RECT 11.800 107.890 20.475 108.190 ;
        RECT 11.800 107.740 15.800 107.890 ;
        RECT 20.145 107.875 20.475 107.890 ;
        RECT 142.965 108.190 143.295 108.205 ;
        RECT 148.805 108.190 152.805 108.340 ;
        RECT 142.965 107.890 152.805 108.190 ;
        RECT 142.965 107.875 143.295 107.890 ;
        RECT 148.805 107.740 152.805 107.890 ;
        RECT 36.150 106.175 37.730 106.505 ;
        RECT 11.800 104.790 15.800 104.940 ;
        RECT 144.805 104.790 145.135 104.805 ;
        RECT 148.805 104.790 152.805 104.940 ;
        RECT 11.800 104.340 16.090 104.790 ;
        RECT 144.805 104.490 152.805 104.790 ;
        RECT 144.805 104.475 145.135 104.490 ;
        RECT 148.805 104.340 152.805 104.490 ;
        RECT 15.790 104.125 16.090 104.340 ;
        RECT 15.790 103.810 16.335 104.125 ;
        RECT 16.005 103.795 16.335 103.810 ;
        RECT 32.850 103.455 34.430 103.785 ;
        RECT 11.800 101.390 15.800 101.540 ;
        RECT 18.305 101.390 18.635 101.405 ;
        RECT 11.800 101.090 18.635 101.390 ;
        RECT 11.800 100.940 15.800 101.090 ;
        RECT 18.305 101.075 18.635 101.090 ;
        RECT 144.805 101.390 145.135 101.405 ;
        RECT 148.805 101.390 152.805 101.540 ;
        RECT 144.805 101.090 152.805 101.390 ;
        RECT 144.805 101.075 145.135 101.090 ;
        RECT 36.150 100.735 37.730 101.065 ;
        RECT 148.805 100.940 152.805 101.090 ;
        RECT 11.800 97.990 15.800 98.140 ;
        RECT 32.850 98.015 34.430 98.345 ;
        RECT 18.305 97.990 18.635 98.005 ;
        RECT 11.800 97.690 18.635 97.990 ;
        RECT 11.800 97.540 15.800 97.690 ;
        RECT 18.305 97.675 18.635 97.690 ;
        RECT 144.805 97.990 145.135 98.005 ;
        RECT 148.805 97.990 152.805 98.140 ;
        RECT 144.805 97.690 152.805 97.990 ;
        RECT 144.805 97.675 145.135 97.690 ;
        RECT 148.805 97.540 152.805 97.690 ;
        RECT 36.150 95.295 37.730 95.625 ;
        RECT 11.800 94.590 15.800 94.740 ;
        RECT 16.925 94.590 17.255 94.605 ;
        RECT 70.745 94.600 71.075 94.605 ;
        RECT 70.745 94.590 71.330 94.600 ;
        RECT 71.665 94.590 71.995 94.605 ;
        RECT 11.800 94.290 17.255 94.590 ;
        RECT 70.520 94.290 71.995 94.590 ;
        RECT 11.800 94.140 15.800 94.290 ;
        RECT 16.925 94.275 17.255 94.290 ;
        RECT 70.745 94.280 71.330 94.290 ;
        RECT 70.745 94.275 71.075 94.280 ;
        RECT 71.665 94.275 71.995 94.290 ;
        RECT 32.850 92.575 34.430 92.905 ;
        RECT 36.150 89.855 37.730 90.185 ;
        RECT 90.065 89.150 90.395 89.165 ;
        RECT 92.825 89.150 93.155 89.165 ;
        RECT 94.205 89.150 94.535 89.165 ;
        RECT 90.065 88.850 94.535 89.150 ;
        RECT 90.065 88.835 90.395 88.850 ;
        RECT 92.825 88.835 93.155 88.850 ;
        RECT 94.205 88.835 94.535 88.850 ;
        RECT 131.465 87.790 131.795 87.805 ;
        RECT 136.525 87.790 136.855 87.805 ;
        RECT 140.205 87.790 140.535 87.805 ;
        RECT 131.465 87.490 140.535 87.790 ;
        RECT 131.465 87.475 131.795 87.490 ;
        RECT 136.525 87.475 136.855 87.490 ;
        RECT 140.205 87.475 140.535 87.490 ;
        RECT 32.850 87.135 34.430 87.465 ;
        RECT 71.205 86.440 71.535 86.445 ;
        RECT 70.950 86.430 71.535 86.440 ;
        RECT 70.950 86.130 71.760 86.430 ;
        RECT 70.950 86.120 71.535 86.130 ;
        RECT 71.205 86.115 71.535 86.120 ;
        RECT 135.145 85.750 135.475 85.765 ;
        RECT 142.045 85.750 142.375 85.765 ;
        RECT 135.145 85.450 142.375 85.750 ;
        RECT 135.145 85.435 135.475 85.450 ;
        RECT 142.045 85.435 142.375 85.450 ;
        RECT 36.150 84.415 37.730 84.745 ;
      LAYER met4 ;
        RECT 32.840 84.340 34.440 212.660 ;
        RECT 36.140 84.340 37.740 212.660 ;
        RECT 107.775 169.075 108.105 169.405 ;
        RECT 107.790 152.405 108.090 169.075 ;
        RECT 132.615 164.315 132.945 164.645 ;
        RECT 132.630 157.165 132.930 164.315 ;
        RECT 132.615 156.835 132.945 157.165 ;
        RECT 116.055 155.475 116.385 155.805 ;
        RECT 107.775 152.075 108.105 152.405 ;
        RECT 116.070 142.885 116.370 155.475 ;
        RECT 122.495 150.035 122.825 150.365 ;
        RECT 116.055 142.555 116.385 142.885 ;
        RECT 122.510 118.405 122.810 150.035 ;
        RECT 122.495 118.075 122.825 118.405 ;
        RECT 70.975 94.275 71.305 94.605 ;
        RECT 70.990 86.445 71.290 94.275 ;
        RECT 70.975 86.115 71.305 86.445 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

