VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 240.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 29.854000 ;
    ANTENNADIFFAREA 365.205353 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 29.854000 ;
    ANTENNADIFFAREA 365.205353 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 29.854000 ;
    ANTENNADIFFAREA 365.205353 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 29.854000 ;
    ANTENNADIFFAREA 365.205353 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 108.065 217.595 108.875 217.735 ;
        RECT 107.875 217.425 108.875 217.595 ;
        RECT 108.065 216.365 108.875 217.425 ;
        RECT 108.065 216.215 108.875 216.355 ;
        RECT 107.875 216.045 108.875 216.215 ;
        RECT 108.065 210.845 108.875 216.045 ;
        RECT 108.065 210.695 108.875 210.835 ;
        RECT 107.875 210.525 108.875 210.695 ;
        RECT 108.065 207.165 108.875 210.525 ;
        RECT 107.905 206.900 108.015 207.020 ;
        RECT 108.065 206.555 108.745 206.695 ;
        RECT 107.875 206.385 108.745 206.555 ;
        RECT 108.065 206.210 108.745 206.385 ;
        RECT 108.065 204.865 108.975 206.210 ;
        RECT 108.150 204.415 108.935 204.845 ;
        RECT 107.905 204.140 108.015 204.260 ;
        RECT 108.065 202.590 108.975 203.935 ;
        RECT 108.065 202.415 108.745 202.590 ;
        RECT 107.875 202.245 108.745 202.415 ;
        RECT 108.065 202.105 108.745 202.245 ;
        RECT 108.065 201.955 108.745 202.095 ;
        RECT 107.875 201.785 108.745 201.955 ;
        RECT 108.065 198.580 108.745 201.785 ;
        RECT 108.065 197.670 108.965 198.580 ;
        RECT 108.065 196.135 108.745 197.670 ;
        RECT 108.065 194.785 108.975 196.135 ;
        RECT 108.065 193.390 108.975 194.735 ;
        RECT 108.065 193.215 108.745 193.390 ;
        RECT 107.875 193.045 108.745 193.215 ;
        RECT 108.065 192.905 108.745 193.045 ;
        RECT 107.910 192.585 108.020 192.745 ;
        RECT 108.150 191.535 108.935 191.965 ;
        RECT 107.910 191.205 108.020 191.365 ;
        RECT 108.065 190.455 108.745 190.595 ;
        RECT 107.875 190.285 108.745 190.455 ;
        RECT 108.065 190.110 108.745 190.285 ;
        RECT 108.065 188.765 108.975 190.110 ;
        RECT 108.065 187.705 108.845 188.755 ;
        RECT 107.875 187.535 108.845 187.705 ;
        RECT 108.065 187.385 108.845 187.535 ;
        RECT 107.910 187.065 108.020 187.225 ;
        RECT 108.065 186.315 108.745 186.455 ;
        RECT 107.875 186.145 108.745 186.315 ;
        RECT 108.065 184.635 108.745 186.145 ;
        RECT 108.065 183.705 108.975 184.635 ;
        RECT 107.905 183.440 108.015 183.560 ;
        RECT 108.065 182.175 108.875 183.235 ;
        RECT 107.875 182.005 108.875 182.175 ;
        RECT 108.065 181.865 108.875 182.005 ;
      LAYER nwell ;
        RECT 109.265 181.670 112.095 217.930 ;
      LAYER pwell ;
        RECT 112.485 217.595 113.295 217.735 ;
        RECT 113.505 217.595 114.315 217.735 ;
        RECT 112.485 217.425 114.315 217.595 ;
        RECT 112.485 216.365 113.295 217.425 ;
        RECT 113.505 216.365 114.315 217.425 ;
        RECT 112.385 215.010 113.295 216.355 ;
        RECT 112.615 214.835 113.295 215.010 ;
        RECT 113.505 214.965 114.415 216.315 ;
        RECT 112.615 214.665 113.485 214.835 ;
        RECT 112.615 214.525 113.295 214.665 ;
        RECT 113.340 214.205 113.450 214.365 ;
        RECT 112.385 213.180 113.295 213.595 ;
        RECT 113.505 213.430 114.185 214.965 ;
        RECT 112.385 213.010 113.485 213.180 ;
        RECT 112.385 212.665 113.295 213.010 ;
        RECT 112.615 209.695 113.295 212.665 ;
        RECT 113.505 212.520 114.405 213.430 ;
        RECT 112.485 209.315 113.295 209.455 ;
        RECT 113.505 209.315 114.185 212.520 ;
        RECT 112.485 209.145 114.185 209.315 ;
        RECT 112.485 205.785 113.295 209.145 ;
        RECT 113.505 209.005 114.185 209.145 ;
        RECT 113.505 208.855 114.315 208.995 ;
        RECT 113.315 208.685 114.315 208.855 ;
        RECT 112.485 205.635 113.295 205.775 ;
        RECT 112.485 205.465 113.485 205.635 ;
        RECT 112.485 204.405 113.295 205.465 ;
        RECT 113.505 205.325 114.315 208.685 ;
        RECT 113.345 205.060 113.455 205.180 ;
        RECT 113.590 204.415 114.375 204.845 ;
        RECT 112.385 203.005 113.295 204.355 ;
        RECT 113.505 204.255 114.185 204.395 ;
        RECT 113.315 204.085 114.185 204.255 ;
        RECT 112.615 201.470 113.295 203.005 ;
        RECT 112.395 200.560 113.295 201.470 ;
        RECT 112.615 197.355 113.295 200.560 ;
        RECT 112.615 197.185 113.485 197.355 ;
        RECT 112.615 197.045 113.295 197.185 ;
        RECT 112.385 196.620 113.295 197.035 ;
        RECT 112.385 196.450 113.485 196.620 ;
        RECT 112.385 196.105 113.295 196.450 ;
        RECT 112.615 193.135 113.295 196.105 ;
        RECT 113.505 195.290 114.185 204.085 ;
        RECT 113.505 195.055 114.315 195.195 ;
        RECT 113.315 194.885 114.315 195.055 ;
        RECT 113.505 193.825 114.315 194.885 ;
        RECT 113.505 193.675 114.285 193.815 ;
        RECT 113.315 193.505 114.285 193.675 ;
        RECT 113.340 192.585 113.450 192.745 ;
        RECT 113.505 192.445 114.285 193.505 ;
        RECT 113.505 192.295 114.285 192.435 ;
        RECT 113.315 192.125 114.285 192.295 ;
        RECT 112.425 191.535 113.210 191.965 ;
        RECT 112.385 190.500 113.295 191.420 ;
        RECT 113.505 191.065 114.285 192.125 ;
        RECT 113.505 190.915 114.285 191.055 ;
        RECT 113.315 190.745 114.285 190.915 ;
        RECT 112.615 188.155 113.295 190.500 ;
        RECT 113.505 189.685 114.285 190.745 ;
        RECT 113.505 189.535 114.285 189.675 ;
        RECT 113.315 189.365 114.285 189.535 ;
        RECT 113.505 188.305 114.285 189.365 ;
        RECT 112.615 187.985 113.485 188.155 ;
        RECT 112.615 187.955 113.295 187.985 ;
        RECT 113.340 187.525 113.450 187.685 ;
        RECT 113.505 187.240 114.415 188.275 ;
        RECT 113.315 187.070 114.415 187.240 ;
        RECT 113.505 186.925 114.415 187.070 ;
        RECT 112.385 184.475 113.295 186.915 ;
        RECT 113.505 186.775 114.415 186.835 ;
        RECT 113.315 186.605 114.415 186.775 ;
        RECT 112.385 184.305 113.485 184.475 ;
        RECT 112.385 184.165 113.295 184.305 ;
        RECT 113.340 183.845 113.450 184.005 ;
        RECT 113.505 183.385 114.415 186.605 ;
        RECT 112.485 182.175 113.295 183.235 ;
        RECT 113.505 182.175 114.315 183.235 ;
        RECT 112.485 182.005 114.315 182.175 ;
        RECT 112.485 181.865 113.295 182.005 ;
        RECT 113.505 181.865 114.315 182.005 ;
      LAYER nwell ;
        RECT 114.705 181.670 117.535 217.930 ;
      LAYER pwell ;
        RECT 117.925 217.595 118.735 217.735 ;
        RECT 118.945 217.595 119.755 217.735 ;
        RECT 117.925 217.425 119.755 217.595 ;
        RECT 117.925 216.365 118.735 217.425 ;
        RECT 118.945 216.365 119.755 217.425 ;
        RECT 117.825 215.010 118.735 216.355 ;
        RECT 118.945 216.215 119.625 216.355 ;
        RECT 118.755 216.045 119.625 216.215 ;
        RECT 118.055 214.835 118.735 215.010 ;
        RECT 118.055 214.665 118.925 214.835 ;
        RECT 118.055 214.525 118.735 214.665 ;
        RECT 118.780 214.205 118.890 214.365 ;
        RECT 118.055 213.455 118.735 213.485 ;
        RECT 118.055 213.285 118.925 213.455 ;
        RECT 118.055 210.940 118.735 213.285 ;
        RECT 117.825 210.020 118.735 210.940 ;
        RECT 118.945 212.840 119.625 216.045 ;
        RECT 118.945 211.930 119.845 212.840 ;
        RECT 118.945 210.395 119.625 211.930 ;
        RECT 118.780 209.605 118.890 209.765 ;
        RECT 118.945 209.045 119.855 210.395 ;
        RECT 118.055 208.855 118.735 208.885 ;
        RECT 118.945 208.855 119.755 208.995 ;
        RECT 118.055 208.685 119.755 208.855 ;
        RECT 118.055 206.340 118.735 208.685 ;
        RECT 117.825 205.420 118.735 206.340 ;
        RECT 118.945 205.325 119.755 208.685 ;
        RECT 118.055 202.115 118.735 205.085 ;
        RECT 118.785 205.060 118.895 205.180 ;
        RECT 119.030 204.415 119.815 204.845 ;
        RECT 118.945 204.255 119.625 204.395 ;
        RECT 118.755 204.085 119.625 204.255 ;
        RECT 117.825 201.770 118.735 202.115 ;
        RECT 117.825 201.600 118.925 201.770 ;
        RECT 117.825 201.185 118.735 201.600 ;
        RECT 117.925 201.035 118.735 201.175 ;
        RECT 117.925 200.865 118.925 201.035 ;
        RECT 118.945 200.880 119.625 204.085 ;
        RECT 117.925 199.345 118.735 200.865 ;
        RECT 118.945 199.970 119.845 200.880 ;
        RECT 118.055 199.195 118.735 199.335 ;
        RECT 118.055 199.025 118.925 199.195 ;
        RECT 118.055 195.820 118.735 199.025 ;
        RECT 118.945 198.435 119.625 199.970 ;
        RECT 118.945 197.085 119.855 198.435 ;
        RECT 118.945 196.890 119.625 197.035 ;
        RECT 118.755 196.720 119.625 196.890 ;
        RECT 117.835 194.910 118.735 195.820 ;
        RECT 118.055 193.375 118.735 194.910 ;
        RECT 118.945 195.190 119.625 196.720 ;
        RECT 118.945 193.825 119.855 195.190 ;
        RECT 118.945 193.675 119.755 193.815 ;
        RECT 118.755 193.505 119.755 193.675 ;
        RECT 117.825 192.025 118.735 193.375 ;
        RECT 117.865 191.535 118.650 191.965 ;
        RECT 117.825 191.100 118.735 191.515 ;
        RECT 117.825 190.930 118.925 191.100 ;
        RECT 118.945 191.065 119.755 193.505 ;
        RECT 117.825 190.585 118.735 190.930 ;
        RECT 118.785 190.800 118.895 190.920 ;
        RECT 118.055 187.615 118.735 190.585 ;
        RECT 118.945 190.455 119.625 190.485 ;
        RECT 118.755 190.285 119.625 190.455 ;
        RECT 118.945 187.940 119.625 190.285 ;
        RECT 117.955 187.235 118.735 187.375 ;
        RECT 117.955 187.065 118.925 187.235 ;
        RECT 117.955 186.005 118.735 187.065 ;
        RECT 118.945 187.020 119.855 187.940 ;
        RECT 118.945 186.775 119.855 186.835 ;
        RECT 118.755 186.605 119.855 186.775 ;
        RECT 117.825 185.050 118.735 185.995 ;
        RECT 118.025 183.560 118.705 185.050 ;
        RECT 118.945 183.835 119.855 186.605 ;
        RECT 118.025 183.390 118.925 183.560 ;
        RECT 118.025 183.245 118.705 183.390 ;
        RECT 117.925 182.175 118.735 183.235 ;
        RECT 118.945 182.175 119.755 183.235 ;
        RECT 117.925 182.005 119.755 182.175 ;
        RECT 117.925 181.865 118.735 182.005 ;
        RECT 118.945 181.865 119.755 182.005 ;
      LAYER nwell ;
        RECT 120.145 181.670 122.975 217.930 ;
      LAYER pwell ;
        RECT 123.365 217.595 124.175 217.735 ;
        RECT 124.385 217.595 125.195 217.735 ;
        RECT 123.365 217.425 125.195 217.595 ;
        RECT 123.365 216.365 124.175 217.425 ;
        RECT 124.385 216.365 125.195 217.425 ;
        RECT 123.265 215.010 124.175 216.355 ;
        RECT 124.385 216.215 125.195 216.355 ;
        RECT 124.195 216.045 125.195 216.215 ;
        RECT 123.495 214.835 124.175 215.010 ;
        RECT 124.385 214.985 125.195 216.045 ;
        RECT 124.385 214.835 125.065 214.865 ;
        RECT 123.495 214.665 125.065 214.835 ;
        RECT 123.495 214.525 124.175 214.665 ;
        RECT 124.225 214.260 124.335 214.380 ;
        RECT 123.265 213.640 124.175 214.055 ;
        RECT 123.265 213.470 124.365 213.640 ;
        RECT 123.265 213.125 124.175 213.470 ;
        RECT 123.495 210.155 124.175 213.125 ;
        RECT 124.385 212.320 125.065 214.665 ;
        RECT 124.385 211.400 125.295 212.320 ;
        RECT 124.385 210.280 125.295 211.200 ;
        RECT 123.495 209.775 124.175 209.915 ;
        RECT 123.495 209.605 124.365 209.775 ;
        RECT 123.495 206.400 124.175 209.605 ;
        RECT 124.385 207.935 125.065 210.280 ;
        RECT 124.195 207.765 125.065 207.935 ;
        RECT 124.385 207.735 125.065 207.765 ;
        RECT 124.385 207.475 125.195 207.615 ;
        RECT 124.195 207.305 125.195 207.475 ;
        RECT 123.275 205.490 124.175 206.400 ;
        RECT 123.495 203.955 124.175 205.490 ;
        RECT 124.385 204.865 125.195 207.305 ;
        RECT 124.470 204.415 125.255 204.845 ;
        RECT 123.265 202.605 124.175 203.955 ;
        RECT 124.385 203.340 125.295 204.375 ;
        RECT 124.195 203.170 125.295 203.340 ;
        RECT 124.385 203.025 125.295 203.170 ;
        RECT 123.265 202.140 124.175 202.555 ;
        RECT 123.265 201.970 124.365 202.140 ;
        RECT 123.265 201.625 124.175 201.970 ;
        RECT 123.495 198.655 124.175 201.625 ;
        RECT 124.385 199.195 125.295 202.945 ;
        RECT 124.195 199.025 125.295 199.195 ;
        RECT 124.385 198.885 125.295 199.025 ;
        RECT 123.265 197.400 124.175 198.320 ;
        RECT 123.495 195.055 124.175 197.400 ;
        RECT 124.385 197.860 125.295 198.780 ;
        RECT 124.385 195.515 125.065 197.860 ;
        RECT 124.195 195.345 125.065 195.515 ;
        RECT 124.385 195.315 125.065 195.345 ;
        RECT 124.385 195.055 125.195 195.195 ;
        RECT 123.495 194.885 125.195 195.055 ;
        RECT 123.495 194.855 124.175 194.885 ;
        RECT 123.365 194.595 124.175 194.735 ;
        RECT 123.365 194.425 124.365 194.595 ;
        RECT 123.365 191.985 124.175 194.425 ;
        RECT 124.385 193.825 125.195 194.885 ;
        RECT 124.385 192.865 125.295 193.815 ;
        RECT 123.305 191.535 124.090 191.965 ;
        RECT 123.265 188.620 124.175 191.225 ;
        RECT 124.415 190.460 125.095 192.865 ;
        RECT 124.195 190.290 125.095 190.460 ;
        RECT 124.415 190.145 125.095 190.290 ;
        RECT 124.385 189.990 125.295 190.135 ;
        RECT 124.195 189.820 125.295 189.990 ;
        RECT 124.385 188.785 125.295 189.820 ;
        RECT 123.265 188.605 124.365 188.620 ;
        RECT 124.385 188.605 125.165 188.755 ;
        RECT 123.265 188.450 125.165 188.605 ;
        RECT 123.265 188.305 124.175 188.450 ;
        RECT 124.195 188.435 125.165 188.450 ;
        RECT 124.220 187.985 124.330 188.145 ;
        RECT 124.385 187.385 125.165 188.435 ;
        RECT 123.265 184.015 124.175 187.235 ;
        RECT 124.385 184.015 125.295 187.235 ;
        RECT 123.265 183.845 125.295 184.015 ;
        RECT 123.265 183.785 124.175 183.845 ;
        RECT 124.385 183.785 125.295 183.845 ;
        RECT 124.225 183.440 124.335 183.560 ;
        RECT 123.365 182.175 124.175 183.235 ;
        RECT 124.385 182.175 125.195 183.235 ;
        RECT 123.365 182.005 125.195 182.175 ;
        RECT 123.365 181.865 124.175 182.005 ;
        RECT 124.385 181.865 125.195 182.005 ;
      LAYER nwell ;
        RECT 125.585 181.670 128.415 217.930 ;
      LAYER pwell ;
        RECT 128.805 217.595 129.615 217.735 ;
        RECT 129.825 217.595 130.635 217.735 ;
        RECT 128.805 217.425 130.635 217.595 ;
        RECT 128.805 216.365 129.615 217.425 ;
        RECT 129.825 216.365 130.635 217.425 ;
        RECT 128.705 214.965 129.615 216.315 ;
        RECT 129.825 215.940 130.735 216.355 ;
        RECT 129.635 215.770 130.735 215.940 ;
        RECT 128.935 213.430 129.615 214.965 ;
        RECT 128.715 212.520 129.615 213.430 ;
        RECT 128.935 209.315 129.615 212.520 ;
        RECT 129.825 215.425 130.735 215.770 ;
        RECT 129.825 212.455 130.505 215.425 ;
        RECT 129.825 212.075 130.505 212.215 ;
        RECT 129.635 211.905 130.505 212.075 ;
        RECT 128.935 209.145 129.805 209.315 ;
        RECT 128.935 209.005 129.615 209.145 ;
        RECT 128.805 208.855 129.615 208.995 ;
        RECT 128.805 208.685 129.805 208.855 ;
        RECT 129.825 208.700 130.505 211.905 ;
        RECT 128.805 206.245 129.615 208.685 ;
        RECT 129.825 207.790 130.725 208.700 ;
        RECT 129.825 206.255 130.505 207.790 ;
        RECT 129.665 205.980 129.775 206.100 ;
        RECT 128.935 205.635 129.615 205.775 ;
        RECT 128.935 205.465 129.805 205.635 ;
        RECT 128.935 196.670 129.615 205.465 ;
        RECT 129.825 204.905 130.735 206.255 ;
        RECT 129.910 204.415 130.695 204.845 ;
        RECT 129.825 204.255 130.505 204.395 ;
        RECT 129.635 204.085 130.505 204.255 ;
        RECT 129.825 200.880 130.505 204.085 ;
        RECT 129.825 199.970 130.725 200.880 ;
        RECT 129.825 198.435 130.505 199.970 ;
        RECT 129.825 197.085 130.735 198.435 ;
        RECT 129.665 196.780 129.775 196.900 ;
        RECT 128.705 195.560 129.615 196.480 ;
        RECT 128.935 193.215 129.615 195.560 ;
        RECT 129.825 195.210 130.735 196.575 ;
        RECT 129.825 193.680 130.505 195.210 ;
        RECT 129.635 193.510 130.505 193.680 ;
        RECT 129.825 193.365 130.505 193.510 ;
        RECT 128.935 193.045 129.805 193.215 ;
        RECT 128.935 193.015 129.615 193.045 ;
        RECT 129.660 192.585 129.770 192.745 ;
        RECT 129.825 192.295 130.735 192.355 ;
        RECT 129.635 192.125 130.735 192.295 ;
        RECT 128.745 191.535 129.530 191.965 ;
        RECT 128.905 191.380 129.585 191.505 ;
        RECT 128.905 191.210 129.805 191.380 ;
        RECT 128.905 190.180 129.585 191.210 ;
        RECT 128.705 189.225 129.615 190.180 ;
        RECT 129.825 189.355 130.735 192.125 ;
        RECT 128.805 189.075 129.615 189.215 ;
        RECT 128.805 189.070 129.805 189.075 ;
        RECT 129.825 189.070 130.735 189.215 ;
        RECT 128.805 188.905 130.735 189.070 ;
        RECT 128.805 186.465 129.615 188.905 ;
        RECT 129.635 188.900 130.735 188.905 ;
        RECT 129.825 187.865 130.735 188.900 ;
        RECT 129.665 187.580 129.775 187.700 ;
        RECT 129.825 187.235 130.735 187.295 ;
        RECT 129.635 187.065 130.735 187.235 ;
        RECT 129.665 186.200 129.775 186.320 ;
        RECT 128.705 184.940 129.615 185.975 ;
        RECT 128.705 184.770 129.805 184.940 ;
        RECT 128.705 184.625 129.615 184.770 ;
        RECT 128.835 183.555 129.615 184.615 ;
        RECT 129.825 183.845 130.735 187.065 ;
        RECT 129.665 183.555 129.775 183.560 ;
        RECT 128.835 183.385 129.805 183.555 ;
        RECT 128.835 183.245 129.615 183.385 ;
        RECT 128.805 182.175 129.615 183.235 ;
        RECT 129.825 182.175 130.635 183.235 ;
        RECT 128.805 182.005 130.635 182.175 ;
        RECT 128.805 181.865 129.615 182.005 ;
        RECT 129.825 181.865 130.635 182.005 ;
      LAYER nwell ;
        RECT 131.025 181.670 133.855 217.930 ;
      LAYER pwell ;
        RECT 134.245 217.595 135.055 217.735 ;
        RECT 135.265 217.595 136.075 217.735 ;
        RECT 134.245 217.425 136.075 217.595 ;
        RECT 134.245 216.365 135.055 217.425 ;
        RECT 135.265 216.365 136.075 217.425 ;
        RECT 134.145 215.010 135.055 216.355 ;
        RECT 135.265 216.215 135.945 216.355 ;
        RECT 135.075 216.045 135.945 216.215 ;
        RECT 134.375 214.835 135.055 215.010 ;
        RECT 134.375 214.665 135.245 214.835 ;
        RECT 134.375 214.525 135.055 214.665 ;
        RECT 134.145 214.100 135.055 214.515 ;
        RECT 134.145 213.930 135.245 214.100 ;
        RECT 134.145 213.585 135.055 213.930 ;
        RECT 134.375 210.615 135.055 213.585 ;
        RECT 135.265 212.840 135.945 216.045 ;
        RECT 135.265 211.930 136.165 212.840 ;
        RECT 135.265 210.395 135.945 211.930 ;
        RECT 134.245 210.235 135.055 210.375 ;
        RECT 134.245 210.065 135.245 210.235 ;
        RECT 134.245 209.005 135.055 210.065 ;
        RECT 135.265 209.045 136.175 210.395 ;
        RECT 134.375 200.115 135.055 208.910 ;
        RECT 135.265 207.980 136.175 208.900 ;
        RECT 135.265 205.635 135.945 207.980 ;
        RECT 135.075 205.465 135.945 205.635 ;
        RECT 135.265 205.435 135.945 205.465 ;
        RECT 135.105 205.060 135.215 205.180 ;
        RECT 135.350 204.415 136.135 204.845 ;
        RECT 135.265 203.980 136.175 204.395 ;
        RECT 135.075 203.810 136.175 203.980 ;
        RECT 135.265 203.465 136.175 203.810 ;
        RECT 135.265 200.495 135.945 203.465 ;
        RECT 135.105 200.115 135.215 200.120 ;
        RECT 134.375 199.945 135.245 200.115 ;
        RECT 134.375 199.805 135.055 199.945 ;
        RECT 134.145 198.780 135.055 199.700 ;
        RECT 135.075 199.650 135.245 199.655 ;
        RECT 135.075 199.485 135.945 199.650 ;
        RECT 134.375 196.435 135.055 198.780 ;
        RECT 135.265 198.745 135.945 199.485 ;
        RECT 135.265 197.815 136.175 198.745 ;
        RECT 135.265 196.435 136.175 197.485 ;
        RECT 134.375 196.265 136.175 196.435 ;
        RECT 134.375 196.235 135.055 196.265 ;
        RECT 135.265 196.135 136.175 196.265 ;
        RECT 134.245 195.975 135.055 196.115 ;
        RECT 135.265 195.975 135.945 196.115 ;
        RECT 134.245 195.805 135.945 195.975 ;
        RECT 134.245 194.745 135.055 195.805 ;
        RECT 134.345 194.590 135.025 194.735 ;
        RECT 134.345 194.420 135.245 194.590 ;
        RECT 134.345 192.930 135.025 194.420 ;
        RECT 134.145 191.985 135.055 192.930 ;
        RECT 135.265 192.600 135.945 195.805 ;
        RECT 134.185 191.535 134.970 191.965 ;
        RECT 135.265 191.690 136.165 192.600 ;
        RECT 134.145 191.375 135.055 191.435 ;
        RECT 134.145 191.205 135.245 191.375 ;
        RECT 134.145 187.985 135.055 191.205 ;
        RECT 135.265 190.155 135.945 191.690 ;
        RECT 135.265 188.805 136.175 190.155 ;
        RECT 135.105 188.500 135.215 188.620 ;
        RECT 135.075 188.150 135.245 188.155 ;
        RECT 135.075 187.985 135.945 188.150 ;
        RECT 134.145 187.695 135.055 187.755 ;
        RECT 134.145 187.525 135.245 187.695 ;
        RECT 134.145 184.305 135.055 187.525 ;
        RECT 135.265 187.245 135.945 187.985 ;
        RECT 135.265 186.315 136.175 187.245 ;
        RECT 135.265 185.855 136.045 185.995 ;
        RECT 135.075 185.685 136.045 185.855 ;
        RECT 135.265 184.625 136.045 185.685 ;
        RECT 135.100 183.845 135.210 184.005 ;
        RECT 135.265 183.565 136.045 184.615 ;
        RECT 135.075 183.395 136.045 183.565 ;
        RECT 135.265 183.245 136.045 183.395 ;
        RECT 134.245 182.175 135.055 183.235 ;
        RECT 135.265 182.175 136.075 183.235 ;
        RECT 134.245 182.005 136.075 182.175 ;
        RECT 134.245 181.865 135.055 182.005 ;
        RECT 135.265 181.865 136.075 182.005 ;
      LAYER nwell ;
        RECT 136.465 181.670 139.295 217.930 ;
      LAYER pwell ;
        RECT 139.685 217.595 140.495 217.735 ;
        RECT 140.705 217.595 141.515 217.735 ;
        RECT 139.685 217.425 141.515 217.595 ;
        RECT 139.685 216.365 140.495 217.425 ;
        RECT 140.705 216.365 141.515 217.425 ;
        RECT 139.685 216.215 140.495 216.355 ;
        RECT 140.705 216.215 141.515 216.355 ;
        RECT 139.685 216.045 141.515 216.215 ;
        RECT 139.685 212.685 140.495 216.045 ;
        RECT 140.545 212.420 140.655 212.540 ;
        RECT 139.585 210.825 140.495 212.175 ;
        RECT 140.705 210.845 141.515 216.045 ;
        RECT 139.815 209.290 140.495 210.825 ;
        RECT 140.550 210.525 140.660 210.685 ;
        RECT 140.705 209.775 141.385 209.915 ;
        RECT 140.515 209.605 141.385 209.775 ;
        RECT 139.595 208.380 140.495 209.290 ;
        RECT 139.815 205.175 140.495 208.380 ;
        RECT 140.705 209.430 141.385 209.605 ;
        RECT 140.705 208.085 141.615 209.430 ;
        RECT 140.705 205.175 141.615 207.945 ;
        RECT 139.815 205.005 141.615 205.175 ;
        RECT 139.815 204.865 140.495 205.005 ;
        RECT 140.705 204.945 141.615 205.005 ;
        RECT 139.815 204.715 140.495 204.855 ;
        RECT 139.815 204.545 140.685 204.715 ;
        RECT 139.815 201.340 140.495 204.545 ;
        RECT 140.790 204.415 141.575 204.845 ;
        RECT 140.550 204.085 140.660 204.245 ;
        RECT 140.705 203.335 141.385 203.365 ;
        RECT 140.515 203.165 141.385 203.335 ;
        RECT 139.595 200.430 140.495 201.340 ;
        RECT 139.815 198.895 140.495 200.430 ;
        RECT 140.705 200.820 141.385 203.165 ;
        RECT 140.705 199.900 141.615 200.820 ;
        RECT 140.550 199.485 140.660 199.645 ;
        RECT 139.585 197.545 140.495 198.895 ;
        RECT 140.705 197.530 141.615 198.875 ;
        RECT 140.705 197.355 141.385 197.530 ;
        RECT 140.515 197.185 141.385 197.355 ;
        RECT 139.585 196.255 140.495 197.185 ;
        RECT 140.705 197.045 141.385 197.185 ;
        RECT 140.705 196.895 141.385 196.925 ;
        RECT 140.515 196.725 141.385 196.895 ;
        RECT 139.815 195.515 140.495 196.255 ;
        RECT 139.815 195.350 140.685 195.515 ;
        RECT 140.515 195.345 140.685 195.350 ;
        RECT 139.815 195.055 140.495 195.195 ;
        RECT 139.815 194.885 140.685 195.055 ;
        RECT 139.815 194.710 140.495 194.885 ;
        RECT 139.585 193.365 140.495 194.710 ;
        RECT 140.705 194.380 141.385 196.725 ;
        RECT 140.705 193.460 141.615 194.380 ;
        RECT 139.585 193.215 140.495 193.345 ;
        RECT 139.585 193.205 140.685 193.215 ;
        RECT 140.705 193.205 141.485 193.355 ;
        RECT 139.585 193.045 141.485 193.205 ;
        RECT 139.585 191.995 140.495 193.045 ;
        RECT 140.515 193.035 141.485 193.045 ;
        RECT 140.705 191.985 141.485 193.035 ;
        RECT 139.625 191.535 140.410 191.965 ;
        RECT 140.790 191.535 141.575 191.965 ;
        RECT 139.585 191.375 140.495 191.435 ;
        RECT 139.585 191.205 140.685 191.375 ;
        RECT 139.585 188.435 140.495 191.205 ;
        RECT 140.705 189.250 141.615 190.595 ;
        RECT 140.705 189.075 141.385 189.250 ;
        RECT 140.515 188.905 141.385 189.075 ;
        RECT 140.705 188.765 141.385 188.905 ;
        RECT 140.705 188.615 141.515 188.755 ;
        RECT 140.515 188.445 141.515 188.615 ;
        RECT 139.815 188.155 140.495 188.185 ;
        RECT 139.815 187.985 140.685 188.155 ;
        RECT 139.815 185.640 140.495 187.985 ;
        RECT 140.705 187.385 141.515 188.445 ;
        RECT 140.705 186.315 141.485 187.375 ;
        RECT 140.515 186.145 141.485 186.315 ;
        RECT 140.705 186.005 141.485 186.145 ;
        RECT 139.585 184.720 140.495 185.640 ;
        RECT 140.705 184.935 141.485 185.995 ;
        RECT 140.515 184.765 141.485 184.935 ;
        RECT 140.705 184.625 141.485 184.765 ;
        RECT 139.715 183.565 140.495 184.615 ;
        RECT 140.705 183.565 141.485 184.615 ;
        RECT 139.715 183.395 141.485 183.565 ;
        RECT 139.715 183.245 140.495 183.395 ;
        RECT 140.705 183.245 141.485 183.395 ;
        RECT 139.685 182.175 140.495 183.235 ;
        RECT 140.705 182.175 141.515 183.235 ;
        RECT 139.685 182.005 141.515 182.175 ;
        RECT 139.685 181.865 140.495 182.005 ;
        RECT 140.705 181.865 141.515 182.005 ;
      LAYER nwell ;
        RECT 141.905 181.670 143.510 217.930 ;
      LAYER pwell ;
        RECT 98.250 163.430 104.350 173.220 ;
        RECT 98.250 163.400 104.360 163.430 ;
        RECT 98.450 163.000 99.610 163.400 ;
        RECT 101.570 161.320 104.360 163.400 ;
      LAYER nwell ;
        RECT 99.460 159.210 104.300 161.320 ;
        RECT 105.580 160.980 115.770 173.230 ;
      LAYER pwell ;
        RECT 117.290 163.460 123.390 173.250 ;
        RECT 117.290 163.430 123.400 163.460 ;
        RECT 117.490 163.030 118.650 163.430 ;
        RECT 120.610 161.350 123.400 163.430 ;
      LAYER nwell ;
        RECT 118.500 159.240 123.340 161.350 ;
        RECT 124.620 161.010 134.810 173.260 ;
      LAYER pwell ;
        RECT 136.240 163.500 142.340 173.290 ;
        RECT 136.240 163.470 142.350 163.500 ;
        RECT 136.440 163.070 137.600 163.470 ;
        RECT 139.560 161.390 142.350 163.470 ;
      LAYER nwell ;
        RECT 137.450 159.280 142.290 161.390 ;
        RECT 143.570 161.050 153.760 173.300 ;
      LAYER pwell ;
        RECT 98.250 148.440 104.350 158.230 ;
        RECT 98.250 148.410 104.360 148.440 ;
        RECT 98.450 148.010 99.610 148.410 ;
        RECT 101.570 146.330 104.360 148.410 ;
      LAYER nwell ;
        RECT 99.460 144.220 104.300 146.330 ;
        RECT 105.580 145.990 115.770 158.240 ;
      LAYER pwell ;
        RECT 117.290 148.440 123.390 158.230 ;
        RECT 117.290 148.410 123.400 148.440 ;
        RECT 117.490 148.010 118.650 148.410 ;
        RECT 120.610 146.330 123.400 148.410 ;
      LAYER nwell ;
        RECT 118.500 144.220 123.340 146.330 ;
        RECT 124.620 145.990 134.810 158.240 ;
      LAYER pwell ;
        RECT 136.290 148.440 142.390 158.230 ;
        RECT 136.290 148.410 142.400 148.440 ;
        RECT 136.490 148.010 137.650 148.410 ;
        RECT 139.610 146.330 142.400 148.410 ;
      LAYER nwell ;
        RECT 137.500 144.220 142.340 146.330 ;
        RECT 143.620 145.990 153.810 158.240 ;
      LAYER pwell ;
        RECT 98.250 133.460 104.350 143.250 ;
        RECT 98.250 133.430 104.360 133.460 ;
        RECT 98.450 133.030 99.610 133.430 ;
        RECT 101.570 131.350 104.360 133.430 ;
      LAYER nwell ;
        RECT 99.460 129.240 104.300 131.350 ;
        RECT 105.580 131.010 115.770 143.260 ;
      LAYER pwell ;
        RECT 117.240 133.420 123.340 143.210 ;
        RECT 117.240 133.390 123.350 133.420 ;
        RECT 117.440 132.990 118.600 133.390 ;
        RECT 120.560 131.310 123.350 133.390 ;
      LAYER nwell ;
        RECT 118.450 129.200 123.290 131.310 ;
        RECT 124.570 130.970 134.760 143.220 ;
      LAYER pwell ;
        RECT 136.240 133.420 142.340 143.210 ;
        RECT 136.240 133.390 142.350 133.420 ;
        RECT 136.440 132.990 137.600 133.390 ;
        RECT 139.560 131.310 142.350 133.390 ;
      LAYER nwell ;
        RECT 137.450 129.200 142.290 131.310 ;
        RECT 143.570 130.970 153.760 143.220 ;
      LAYER pwell ;
        RECT 98.250 118.430 104.350 128.220 ;
        RECT 98.250 118.400 104.360 118.430 ;
        RECT 98.450 118.000 99.610 118.400 ;
        RECT 101.570 116.320 104.360 118.400 ;
      LAYER nwell ;
        RECT 99.460 114.210 104.300 116.320 ;
        RECT 105.580 115.980 115.770 128.230 ;
      LAYER pwell ;
        RECT 117.240 118.400 123.340 128.190 ;
        RECT 117.240 118.370 123.350 118.400 ;
        RECT 117.440 117.970 118.600 118.370 ;
        RECT 120.560 116.290 123.350 118.370 ;
      LAYER nwell ;
        RECT 118.450 114.180 123.290 116.290 ;
        RECT 124.570 115.950 134.760 128.200 ;
      LAYER pwell ;
        RECT 136.240 118.400 142.340 128.190 ;
        RECT 136.240 118.370 142.350 118.400 ;
        RECT 136.440 117.970 137.600 118.370 ;
        RECT 139.560 116.290 142.350 118.370 ;
      LAYER nwell ;
        RECT 137.450 114.180 142.290 116.290 ;
        RECT 143.570 115.950 153.760 128.200 ;
      LAYER pwell ;
        RECT 98.250 103.440 104.350 113.230 ;
        RECT 98.250 103.410 104.360 103.440 ;
        RECT 98.450 103.010 99.610 103.410 ;
        RECT 101.570 101.330 104.360 103.410 ;
      LAYER nwell ;
        RECT 99.460 99.220 104.300 101.330 ;
        RECT 105.580 100.990 115.770 113.240 ;
      LAYER pwell ;
        RECT 117.240 103.420 123.340 113.210 ;
        RECT 117.240 103.390 123.350 103.420 ;
        RECT 117.440 102.990 118.600 103.390 ;
        RECT 120.560 101.310 123.350 103.390 ;
      LAYER nwell ;
        RECT 118.450 99.200 123.290 101.310 ;
        RECT 124.570 100.970 134.760 113.220 ;
      LAYER pwell ;
        RECT 136.290 103.420 142.390 113.210 ;
        RECT 136.290 103.390 142.400 103.420 ;
        RECT 136.490 102.990 137.650 103.390 ;
        RECT 139.610 101.310 142.400 103.390 ;
      LAYER nwell ;
        RECT 137.500 99.200 142.340 101.310 ;
        RECT 143.620 100.970 153.810 113.220 ;
      LAYER pwell ;
        RECT 99.970 96.680 154.410 98.690 ;
        RECT 99.970 95.200 142.430 96.680 ;
      LAYER li1 ;
        RECT 107.875 217.655 108.045 217.740 ;
        RECT 110.595 217.655 110.765 217.740 ;
        RECT 113.315 217.655 113.485 217.740 ;
        RECT 116.035 217.655 116.205 217.740 ;
        RECT 118.755 217.655 118.925 217.740 ;
        RECT 121.475 217.655 121.645 217.740 ;
        RECT 124.195 217.655 124.365 217.740 ;
        RECT 126.915 217.655 127.085 217.740 ;
        RECT 129.635 217.655 129.805 217.740 ;
        RECT 132.355 217.655 132.525 217.740 ;
        RECT 135.075 217.655 135.245 217.740 ;
        RECT 137.795 217.655 137.965 217.740 ;
        RECT 140.515 217.655 140.685 217.740 ;
        RECT 143.235 217.655 143.405 217.740 ;
        RECT 107.875 217.135 109.335 217.655 ;
        RECT 107.875 216.445 108.795 217.135 ;
        RECT 109.505 216.965 111.855 217.655 ;
        RECT 112.025 217.135 114.775 217.655 ;
        RECT 108.965 216.445 112.395 216.965 ;
        RECT 112.565 216.445 114.235 217.135 ;
        RECT 114.945 216.965 117.295 217.655 ;
        RECT 117.465 217.135 120.215 217.655 ;
        RECT 114.405 216.445 117.835 216.965 ;
        RECT 118.005 216.445 119.675 217.135 ;
        RECT 120.385 216.965 122.735 217.655 ;
        RECT 122.905 217.135 125.655 217.655 ;
        RECT 119.845 216.445 123.275 216.965 ;
        RECT 123.445 216.445 125.115 217.135 ;
        RECT 125.825 216.965 128.175 217.655 ;
        RECT 128.345 217.135 131.095 217.655 ;
        RECT 125.285 216.445 128.715 216.965 ;
        RECT 128.885 216.445 130.555 217.135 ;
        RECT 131.265 216.965 133.615 217.655 ;
        RECT 133.785 217.135 136.535 217.655 ;
        RECT 130.725 216.445 134.155 216.965 ;
        RECT 134.325 216.445 135.995 217.135 ;
        RECT 136.705 216.965 139.055 217.655 ;
        RECT 139.225 217.135 141.975 217.655 ;
        RECT 136.165 216.445 139.595 216.965 ;
        RECT 139.765 216.445 141.435 217.135 ;
        RECT 142.145 216.965 143.405 217.655 ;
        RECT 141.605 216.445 143.405 216.965 ;
        RECT 107.875 216.275 108.045 216.445 ;
        RECT 110.595 216.275 110.765 216.445 ;
        RECT 107.875 214.690 108.590 216.275 ;
        RECT 110.160 216.270 110.765 216.275 ;
        RECT 113.315 216.270 113.485 216.445 ;
        RECT 110.160 216.010 111.915 216.270 ;
        RECT 112.475 216.010 113.485 216.270 ;
        RECT 114.140 216.225 114.975 216.275 ;
        RECT 110.160 215.410 110.765 216.010 ;
        RECT 110.935 215.665 113.145 215.835 ;
        RECT 110.935 215.580 111.840 215.665 ;
        RECT 112.570 215.580 113.145 215.665 ;
        RECT 113.315 215.725 113.485 216.010 ;
        RECT 113.705 216.215 114.975 216.225 ;
        RECT 116.035 216.270 116.205 216.445 ;
        RECT 118.755 216.270 118.925 216.445 ;
        RECT 121.475 216.270 121.645 216.445 ;
        RECT 124.195 216.275 124.365 216.445 ;
        RECT 126.915 216.275 127.085 216.445 ;
        RECT 124.195 216.270 125.655 216.275 ;
        RECT 113.705 216.105 115.820 216.215 ;
        RECT 113.705 216.050 114.265 216.105 ;
        RECT 114.845 216.060 115.820 216.105 ;
        RECT 113.705 215.895 114.225 216.050 ;
        RECT 113.315 215.555 114.095 215.725 ;
        RECT 112.075 215.410 112.405 215.495 ;
        RECT 113.315 215.410 113.485 215.555 ;
        RECT 110.160 215.080 111.525 215.410 ;
        RECT 111.695 215.240 112.765 215.410 ;
        RECT 107.875 214.350 109.420 214.690 ;
        RECT 107.875 210.930 108.590 214.350 ;
        RECT 110.160 213.005 110.765 215.080 ;
        RECT 111.695 214.865 111.865 215.240 ;
        RECT 110.935 214.695 111.865 214.865 ;
        RECT 112.045 214.605 112.415 214.960 ;
        RECT 112.595 214.865 112.765 215.240 ;
        RECT 112.935 215.080 113.485 215.410 ;
        RECT 114.395 215.385 114.725 215.935 ;
        RECT 114.895 215.885 115.820 216.060 ;
        RECT 116.035 216.010 117.355 216.270 ;
        RECT 117.915 216.010 118.925 216.270 ;
        RECT 119.185 216.015 119.645 216.185 ;
        RECT 116.035 215.715 116.205 216.010 ;
        RECT 118.755 215.845 118.925 216.010 ;
        RECT 115.025 215.545 116.205 215.715 ;
        RECT 116.375 215.665 118.585 215.835 ;
        RECT 116.375 215.580 117.280 215.665 ;
        RECT 118.010 215.580 118.585 215.665 ;
        RECT 112.595 214.695 113.145 214.865 ;
        RECT 113.315 214.795 113.485 215.080 ;
        RECT 113.700 215.375 114.725 215.385 ;
        RECT 116.035 215.410 116.205 215.545 ;
        RECT 118.755 215.515 119.305 215.845 ;
        RECT 119.475 215.750 119.645 216.015 ;
        RECT 119.815 215.920 120.465 216.270 ;
        RECT 120.635 216.015 121.305 216.185 ;
        RECT 120.635 215.750 120.805 216.015 ;
        RECT 121.475 216.010 122.795 216.270 ;
        RECT 123.355 216.010 125.655 216.270 ;
        RECT 121.475 215.845 121.645 216.010 ;
        RECT 119.475 215.520 120.805 215.750 ;
        RECT 120.975 215.515 121.645 215.845 ;
        RECT 121.815 215.665 124.025 215.835 ;
        RECT 121.815 215.580 122.720 215.665 ;
        RECT 123.450 215.580 124.025 215.665 ;
        RECT 124.195 215.755 125.655 216.010 ;
        RECT 117.515 215.410 117.845 215.495 ;
        RECT 118.755 215.410 118.925 215.515 ;
        RECT 113.700 215.185 115.865 215.375 ;
        RECT 113.700 215.055 114.225 215.185 ;
        RECT 114.930 215.035 115.865 215.185 ;
        RECT 116.035 215.080 116.965 215.410 ;
        RECT 117.135 215.240 118.205 215.410 ;
        RECT 113.315 214.585 114.015 214.795 ;
        RECT 110.935 213.340 113.145 213.510 ;
        RECT 110.935 213.175 111.905 213.340 ;
        RECT 112.575 213.255 113.145 213.340 ;
        RECT 112.075 213.085 112.405 213.170 ;
        RECT 113.315 213.085 113.485 214.585 ;
        RECT 114.395 214.310 114.725 215.015 ;
        RECT 114.930 214.480 115.305 215.035 ;
        RECT 116.035 214.805 116.205 215.080 ;
        RECT 117.135 214.865 117.305 215.240 ;
        RECT 115.535 214.490 116.205 214.805 ;
        RECT 116.375 214.695 117.305 214.865 ;
        RECT 117.485 214.605 117.855 214.960 ;
        RECT 118.035 214.865 118.205 215.240 ;
        RECT 118.375 215.080 118.925 215.410 ;
        RECT 121.475 215.410 121.645 215.515 ;
        RECT 122.955 215.410 123.285 215.495 ;
        RECT 124.195 215.410 125.115 215.755 ;
        RECT 125.825 215.715 127.085 216.275 ;
        RECT 128.145 216.225 128.980 216.275 ;
        RECT 128.145 216.215 129.415 216.225 ;
        RECT 127.300 216.105 129.415 216.215 ;
        RECT 127.300 216.060 128.275 216.105 ;
        RECT 127.300 215.885 128.225 216.060 ;
        RECT 128.855 216.050 129.415 216.105 ;
        RECT 125.825 215.585 128.095 215.715 ;
        RECT 119.185 215.160 121.305 215.345 ;
        RECT 118.755 214.905 118.925 215.080 ;
        RECT 121.475 215.080 122.405 215.410 ;
        RECT 122.575 215.240 123.645 215.410 ;
        RECT 118.035 214.695 118.585 214.865 ;
        RECT 118.755 214.655 119.385 214.905 ;
        RECT 119.555 214.710 120.505 214.990 ;
        RECT 121.475 214.920 121.645 215.080 ;
        RECT 121.015 214.655 121.645 214.920 ;
        RECT 122.575 214.865 122.745 215.240 ;
        RECT 121.815 214.695 122.745 214.865 ;
        RECT 113.765 214.140 115.735 214.310 ;
        RECT 113.765 213.525 113.935 214.140 ;
        RECT 114.105 213.650 115.395 213.970 ;
        RECT 114.105 213.505 114.435 213.650 ;
        RECT 110.160 212.870 111.905 213.005 ;
        RECT 112.075 212.915 112.745 213.085 ;
        RECT 108.910 212.835 111.905 212.870 ;
        RECT 108.910 212.520 110.765 212.835 ;
        RECT 112.075 212.665 112.405 212.690 ;
        RECT 110.160 210.930 110.765 212.520 ;
        RECT 107.875 210.755 108.045 210.930 ;
        RECT 110.595 210.755 110.765 210.930 ;
        RECT 107.875 209.105 109.335 210.755 ;
        RECT 109.505 210.465 110.765 210.755 ;
        RECT 110.935 212.495 112.405 212.665 ;
        RECT 110.935 210.805 111.105 212.495 ;
        RECT 112.575 212.330 112.745 212.915 ;
        RECT 112.915 212.770 113.485 213.085 ;
        RECT 113.765 213.120 113.935 213.355 ;
        RECT 114.645 213.290 115.365 213.480 ;
        RECT 115.565 213.425 115.735 214.140 ;
        RECT 115.535 213.120 115.865 213.200 ;
        RECT 113.765 212.950 115.865 213.120 ;
        RECT 112.915 212.755 113.985 212.770 ;
        RECT 113.315 212.400 113.985 212.755 ;
        RECT 114.165 212.490 114.465 212.950 ;
        RECT 116.035 212.945 116.205 214.490 ;
        RECT 116.375 213.115 117.055 213.400 ;
        RECT 116.035 212.780 116.665 212.945 ;
        RECT 114.645 212.610 114.975 212.780 ;
        RECT 115.235 212.675 116.665 212.780 ;
        RECT 115.235 212.610 116.205 212.675 ;
        RECT 112.575 212.325 113.145 212.330 ;
        RECT 111.275 212.155 113.145 212.325 ;
        RECT 111.275 211.200 111.445 212.155 ;
        RECT 111.615 211.815 112.585 211.985 ;
        RECT 111.615 211.165 111.785 211.815 ;
        RECT 112.780 211.800 113.145 212.155 ;
        RECT 112.805 211.610 112.975 211.615 ;
        RECT 111.985 211.335 113.145 211.610 ;
        RECT 111.615 210.975 113.145 211.165 ;
        RECT 110.935 210.635 111.960 210.805 ;
        RECT 113.315 210.795 113.485 212.400 ;
        RECT 114.165 212.290 114.495 212.490 ;
        RECT 114.715 212.440 114.975 212.610 ;
        RECT 114.715 212.270 115.760 212.440 ;
        RECT 114.715 212.080 114.885 212.270 ;
        RECT 113.765 211.910 114.885 212.080 ;
        RECT 113.765 211.405 113.935 211.910 ;
        RECT 115.055 211.740 115.420 212.100 ;
        RECT 114.135 211.570 115.420 211.740 ;
        RECT 114.135 211.215 114.355 211.570 ;
        RECT 113.765 211.045 113.935 211.210 ;
        RECT 114.525 211.160 115.120 211.400 ;
        RECT 115.590 211.335 115.760 212.270 ;
        RECT 113.765 210.990 114.205 211.045 ;
        RECT 115.310 210.990 115.865 211.125 ;
        RECT 113.765 210.875 115.865 210.990 ;
        RECT 116.035 210.885 116.205 212.610 ;
        RECT 116.835 212.655 117.055 213.115 ;
        RECT 117.225 212.825 117.785 213.515 ;
        RECT 117.955 213.115 118.585 213.400 ;
        RECT 117.955 212.655 118.125 213.115 ;
        RECT 118.755 212.960 118.925 214.655 ;
        RECT 119.515 214.485 120.880 214.540 ;
        RECT 119.205 214.370 121.305 214.485 ;
        RECT 119.205 214.315 119.645 214.370 ;
        RECT 119.205 214.150 119.375 214.315 ;
        RECT 120.750 214.235 121.305 214.370 ;
        RECT 119.205 213.450 119.375 213.955 ;
        RECT 119.575 213.790 119.795 214.145 ;
        RECT 119.965 213.960 120.560 214.200 ;
        RECT 119.575 213.620 120.860 213.790 ;
        RECT 119.205 213.280 120.325 213.450 ;
        RECT 120.155 213.090 120.325 213.280 ;
        RECT 120.495 213.260 120.860 213.620 ;
        RECT 121.030 213.090 121.200 214.025 ;
        RECT 118.755 212.945 119.425 212.960 ;
        RECT 118.295 212.675 119.425 212.945 ;
        RECT 116.835 212.445 118.125 212.655 ;
        RECT 118.755 212.590 119.425 212.675 ;
        RECT 119.605 212.870 119.935 213.070 ;
        RECT 120.155 212.920 121.200 213.090 ;
        RECT 121.475 213.465 121.645 214.655 ;
        RECT 122.925 214.605 123.295 214.960 ;
        RECT 123.475 214.865 123.645 215.240 ;
        RECT 123.815 215.080 125.115 215.410 ;
        RECT 124.195 215.065 125.115 215.080 ;
        RECT 125.285 215.545 128.095 215.585 ;
        RECT 125.285 215.065 127.085 215.545 ;
        RECT 128.395 215.385 128.725 215.935 ;
        RECT 128.895 215.895 129.415 216.050 ;
        RECT 129.635 215.845 129.805 216.445 ;
        RECT 132.355 216.270 132.525 216.445 ;
        RECT 135.075 216.270 135.245 216.445 ;
        RECT 137.795 216.275 137.965 216.445 ;
        RECT 140.515 216.275 140.685 216.445 ;
        RECT 143.235 216.275 143.405 216.445 ;
        RECT 129.975 216.100 132.185 216.270 ;
        RECT 129.975 216.015 130.545 216.100 ;
        RECT 131.215 215.935 132.185 216.100 ;
        RECT 132.355 216.010 133.675 216.270 ;
        RECT 134.235 216.010 135.245 216.270 ;
        RECT 135.505 216.015 135.965 216.185 ;
        RECT 130.715 215.845 131.045 215.930 ;
        RECT 129.635 215.725 130.205 215.845 ;
        RECT 129.025 215.555 130.205 215.725 ;
        RECT 129.635 215.515 130.205 215.555 ;
        RECT 130.375 215.675 131.045 215.845 ;
        RECT 132.355 215.765 132.525 216.010 ;
        RECT 135.075 215.845 135.245 216.010 ;
        RECT 128.395 215.375 129.420 215.385 ;
        RECT 123.475 214.695 124.025 214.865 ;
        RECT 124.195 214.325 124.365 215.065 ;
        RECT 124.535 214.495 125.165 214.780 ;
        RECT 124.195 214.055 124.825 214.325 ;
        RECT 121.815 213.800 124.025 213.970 ;
        RECT 121.815 213.635 122.785 213.800 ;
        RECT 123.455 213.715 124.025 213.800 ;
        RECT 122.955 213.545 123.285 213.630 ;
        RECT 124.195 213.545 124.365 214.055 ;
        RECT 124.995 214.035 125.165 214.495 ;
        RECT 125.335 214.205 125.895 214.895 ;
        RECT 126.915 214.805 127.085 215.065 ;
        RECT 127.255 215.185 129.420 215.375 ;
        RECT 127.255 215.035 128.190 215.185 ;
        RECT 128.895 215.055 129.420 215.185 ;
        RECT 126.065 214.495 126.745 214.780 ;
        RECT 126.065 214.035 126.285 214.495 ;
        RECT 126.915 214.490 127.585 214.805 ;
        RECT 126.915 214.325 127.085 214.490 ;
        RECT 127.815 214.480 128.190 215.035 ;
        RECT 126.455 214.055 127.085 214.325 ;
        RECT 128.395 214.310 128.725 215.015 ;
        RECT 129.635 214.795 129.805 215.515 ;
        RECT 130.375 215.090 130.545 215.675 ;
        RECT 131.215 215.595 132.525 215.765 ;
        RECT 130.715 215.425 131.045 215.450 ;
        RECT 130.715 215.255 132.185 215.425 ;
        RECT 129.105 214.585 129.805 214.795 ;
        RECT 124.995 213.825 126.285 214.035 ;
        RECT 121.475 213.295 122.785 213.465 ;
        RECT 122.955 213.375 123.625 213.545 ;
        RECT 116.375 211.875 118.585 212.275 ;
        RECT 116.375 211.405 117.055 211.685 ;
        RECT 116.835 211.010 117.055 211.405 ;
        RECT 117.225 211.180 117.785 211.875 ;
        RECT 117.955 211.405 118.585 211.685 ;
        RECT 117.955 211.010 118.125 211.405 ;
        RECT 114.075 210.820 115.440 210.875 ;
        RECT 109.505 210.295 111.525 210.465 ;
        RECT 109.505 209.375 110.765 210.295 ;
        RECT 111.115 209.885 111.525 210.060 ;
        RECT 111.770 210.055 111.960 210.635 ;
        RECT 112.335 210.065 112.505 210.775 ;
        RECT 112.780 210.705 113.485 210.795 ;
        RECT 116.035 210.705 116.665 210.885 ;
        RECT 112.780 210.455 113.945 210.705 ;
        RECT 112.780 210.285 113.485 210.455 ;
        RECT 114.115 210.370 115.065 210.650 ;
        RECT 115.575 210.560 116.665 210.705 ;
        RECT 116.835 210.560 118.125 211.010 ;
        RECT 118.755 210.885 118.925 212.590 ;
        RECT 119.605 212.410 119.905 212.870 ;
        RECT 120.155 212.750 120.415 212.920 ;
        RECT 121.475 212.750 121.645 213.295 ;
        RECT 122.955 213.125 123.285 213.150 ;
        RECT 120.085 212.580 120.415 212.750 ;
        RECT 120.675 212.580 121.645 212.750 ;
        RECT 119.205 212.240 121.305 212.410 ;
        RECT 119.205 212.005 119.375 212.240 ;
        RECT 120.975 212.160 121.305 212.240 ;
        RECT 120.085 211.880 120.805 212.070 ;
        RECT 119.205 211.220 119.375 211.835 ;
        RECT 119.545 211.710 119.875 211.855 ;
        RECT 119.545 211.390 120.835 211.710 ;
        RECT 121.005 211.220 121.175 211.935 ;
        RECT 119.205 211.050 121.175 211.220 ;
        RECT 118.295 210.775 118.925 210.885 ;
        RECT 118.295 210.565 119.455 210.775 ;
        RECT 118.295 210.560 118.925 210.565 ;
        RECT 115.575 210.440 116.205 210.560 ;
        RECT 117.515 210.455 117.845 210.560 ;
        RECT 112.335 209.885 113.110 210.065 ;
        RECT 111.115 209.820 113.110 209.885 ;
        RECT 113.315 209.845 113.485 210.285 ;
        RECT 113.745 210.015 115.865 210.200 ;
        RECT 116.035 209.845 116.205 210.440 ;
        RECT 116.375 210.285 117.345 210.390 ;
        RECT 118.015 210.285 118.585 210.390 ;
        RECT 116.375 210.005 118.585 210.285 ;
        RECT 111.115 209.545 112.505 209.820 ;
        RECT 113.315 209.515 113.865 209.845 ;
        RECT 114.035 209.610 115.365 209.840 ;
        RECT 113.315 209.375 113.485 209.515 ;
        RECT 107.875 207.245 108.815 209.105 ;
        RECT 109.505 208.935 111.855 209.375 ;
        RECT 108.985 207.555 111.855 208.935 ;
        RECT 112.025 208.915 113.485 209.375 ;
        RECT 114.035 209.345 114.205 209.610 ;
        RECT 113.745 209.175 114.205 209.345 ;
        RECT 114.375 209.090 115.025 209.440 ;
        RECT 115.195 209.345 115.365 209.610 ;
        RECT 115.535 209.515 116.205 209.845 ;
        RECT 115.195 209.175 115.865 209.345 ;
        RECT 116.035 208.915 116.205 209.515 ;
        RECT 118.755 209.805 118.925 210.560 ;
        RECT 119.835 210.345 120.165 211.050 ;
        RECT 121.475 210.925 121.645 212.580 ;
        RECT 121.815 212.955 123.285 213.125 ;
        RECT 121.815 211.265 121.985 212.955 ;
        RECT 123.455 212.790 123.625 213.375 ;
        RECT 123.795 213.215 124.365 213.545 ;
        RECT 124.535 213.255 126.745 213.655 ;
        RECT 123.455 212.785 124.025 212.790 ;
        RECT 122.155 212.615 124.025 212.785 ;
        RECT 122.155 211.660 122.325 212.615 ;
        RECT 122.495 212.275 123.465 212.445 ;
        RECT 122.495 211.625 122.665 212.275 ;
        RECT 123.660 212.260 124.025 212.615 ;
        RECT 124.195 212.265 124.365 213.215 ;
        RECT 124.535 212.785 125.165 213.065 ;
        RECT 124.995 212.390 125.165 212.785 ;
        RECT 125.335 212.560 125.895 213.255 ;
        RECT 126.065 212.785 126.745 213.065 ;
        RECT 126.065 212.390 126.285 212.785 ;
        RECT 123.685 212.070 123.855 212.075 ;
        RECT 122.865 211.795 124.025 212.070 ;
        RECT 124.195 211.940 124.825 212.265 ;
        RECT 124.995 211.940 126.285 212.390 ;
        RECT 126.915 212.780 127.085 214.055 ;
        RECT 127.385 214.140 129.355 214.310 ;
        RECT 127.385 213.425 127.555 214.140 ;
        RECT 127.725 213.650 129.015 213.970 ;
        RECT 128.685 213.505 129.015 213.650 ;
        RECT 129.185 213.525 129.355 214.140 ;
        RECT 129.635 213.555 129.805 214.585 ;
        RECT 129.975 215.085 130.545 215.090 ;
        RECT 129.975 214.915 131.845 215.085 ;
        RECT 129.975 214.560 130.340 214.915 ;
        RECT 130.535 214.575 131.505 214.745 ;
        RECT 130.145 214.370 130.315 214.375 ;
        RECT 129.975 214.095 131.135 214.370 ;
        RECT 131.335 213.925 131.505 214.575 ;
        RECT 131.675 213.960 131.845 214.915 ;
        RECT 129.975 213.735 131.505 213.925 ;
        RECT 132.015 213.565 132.185 215.255 ;
        RECT 127.755 213.290 128.475 213.480 ;
        RECT 127.255 213.120 127.585 213.200 ;
        RECT 129.185 213.120 129.355 213.355 ;
        RECT 127.255 212.950 129.355 213.120 ;
        RECT 129.635 213.045 130.340 213.555 ;
        RECT 126.915 212.610 127.885 212.780 ;
        RECT 128.145 212.610 128.475 212.780 ;
        RECT 126.915 212.265 127.085 212.610 ;
        RECT 128.145 212.440 128.405 212.610 ;
        RECT 128.655 212.490 128.955 212.950 ;
        RECT 129.635 212.770 129.805 213.045 ;
        RECT 130.615 212.825 130.785 213.535 ;
        RECT 126.455 211.940 127.085 212.265 ;
        RECT 122.495 211.435 124.025 211.625 ;
        RECT 121.815 211.095 122.840 211.265 ;
        RECT 124.195 211.255 124.365 211.940 ;
        RECT 125.275 211.835 125.605 211.940 ;
        RECT 124.535 211.665 125.105 211.770 ;
        RECT 125.775 211.665 126.745 211.770 ;
        RECT 124.535 211.385 126.745 211.665 ;
        RECT 120.370 210.325 120.745 210.880 ;
        RECT 121.475 210.870 122.405 210.925 ;
        RECT 120.975 210.755 122.405 210.870 ;
        RECT 120.975 210.555 121.645 210.755 ;
        RECT 119.140 210.175 119.665 210.305 ;
        RECT 120.370 210.175 121.305 210.325 ;
        RECT 119.140 209.985 121.305 210.175 ;
        RECT 119.140 209.975 120.165 209.985 ;
        RECT 118.755 209.635 119.535 209.805 ;
        RECT 118.755 208.915 118.925 209.635 ;
        RECT 119.145 209.310 119.665 209.465 ;
        RECT 119.835 209.425 120.165 209.975 ;
        RECT 121.475 209.815 121.645 210.555 ;
        RECT 121.995 210.345 122.405 210.520 ;
        RECT 122.650 210.515 122.840 211.095 ;
        RECT 123.215 210.525 123.385 211.235 ;
        RECT 123.660 210.745 124.365 211.255 ;
        RECT 124.535 210.935 126.745 211.215 ;
        RECT 124.535 210.830 125.105 210.935 ;
        RECT 125.775 210.830 126.745 210.935 ;
        RECT 124.195 210.660 124.365 210.745 ;
        RECT 125.275 210.660 125.605 210.765 ;
        RECT 126.915 210.705 127.085 211.940 ;
        RECT 127.360 212.270 128.405 212.440 ;
        RECT 128.625 212.290 128.955 212.490 ;
        RECT 129.135 212.400 129.805 212.770 ;
        RECT 130.010 212.645 130.785 212.825 ;
        RECT 131.160 213.395 132.185 213.565 ;
        RECT 132.355 215.410 132.525 215.595 ;
        RECT 132.695 215.665 134.905 215.835 ;
        RECT 132.695 215.580 133.600 215.665 ;
        RECT 134.330 215.580 134.905 215.665 ;
        RECT 135.075 215.515 135.625 215.845 ;
        RECT 135.795 215.750 135.965 216.015 ;
        RECT 136.135 215.920 136.785 216.270 ;
        RECT 136.955 216.015 137.625 216.185 ;
        RECT 136.955 215.750 137.125 216.015 ;
        RECT 137.795 215.845 139.055 216.275 ;
        RECT 135.795 215.520 137.125 215.750 ;
        RECT 137.295 215.515 139.055 215.845 ;
        RECT 133.835 215.410 134.165 215.495 ;
        RECT 135.075 215.410 135.245 215.515 ;
        RECT 132.355 215.080 133.285 215.410 ;
        RECT 133.455 215.240 134.525 215.410 ;
        RECT 132.355 213.925 132.525 215.080 ;
        RECT 133.455 214.865 133.625 215.240 ;
        RECT 132.695 214.695 133.625 214.865 ;
        RECT 133.805 214.605 134.175 214.960 ;
        RECT 134.355 214.865 134.525 215.240 ;
        RECT 134.695 215.080 135.245 215.410 ;
        RECT 135.505 215.160 137.625 215.345 ;
        RECT 135.075 214.905 135.245 215.080 ;
        RECT 134.355 214.695 134.905 214.865 ;
        RECT 135.075 214.655 135.705 214.905 ;
        RECT 135.875 214.710 136.825 214.990 ;
        RECT 137.795 214.920 139.055 215.515 ;
        RECT 137.335 214.655 139.055 214.920 ;
        RECT 132.695 214.260 134.905 214.430 ;
        RECT 132.695 214.095 133.665 214.260 ;
        RECT 134.335 214.175 134.905 214.260 ;
        RECT 133.835 214.005 134.165 214.090 ;
        RECT 135.075 214.005 135.245 214.655 ;
        RECT 135.835 214.485 137.200 214.540 ;
        RECT 135.525 214.370 137.625 214.485 ;
        RECT 135.525 214.315 135.965 214.370 ;
        RECT 135.525 214.150 135.695 214.315 ;
        RECT 137.070 214.235 137.625 214.370 ;
        RECT 137.795 214.455 139.055 214.655 ;
        RECT 139.225 214.690 141.230 216.275 ;
        RECT 139.225 214.625 142.060 214.690 ;
        RECT 132.355 213.755 133.665 213.925 ;
        RECT 133.835 213.835 134.505 214.005 ;
        RECT 131.160 212.815 131.350 213.395 ;
        RECT 132.355 213.225 132.525 213.755 ;
        RECT 133.835 213.585 134.165 213.610 ;
        RECT 131.595 213.055 132.525 213.225 ;
        RECT 131.595 212.645 132.005 212.820 ;
        RECT 130.010 212.580 132.005 212.645 ;
        RECT 127.360 211.335 127.530 212.270 ;
        RECT 127.700 211.740 128.065 212.100 ;
        RECT 128.235 212.080 128.405 212.270 ;
        RECT 128.235 211.910 129.355 212.080 ;
        RECT 127.700 211.570 128.985 211.740 ;
        RECT 128.000 211.160 128.595 211.400 ;
        RECT 128.765 211.215 128.985 211.570 ;
        RECT 129.185 211.405 129.355 211.910 ;
        RECT 129.635 211.705 129.805 212.400 ;
        RECT 130.615 212.305 132.005 212.580 ;
        RECT 130.065 211.875 130.525 212.045 ;
        RECT 129.635 211.375 130.185 211.705 ;
        RECT 130.355 211.610 130.525 211.875 ;
        RECT 130.695 211.780 131.345 212.130 ;
        RECT 131.515 211.875 132.185 212.045 ;
        RECT 131.515 211.610 131.685 211.875 ;
        RECT 132.355 211.705 132.525 213.055 ;
        RECT 130.355 211.380 131.685 211.610 ;
        RECT 131.855 211.385 132.525 211.705 ;
        RECT 132.695 213.415 134.165 213.585 ;
        RECT 132.695 211.725 132.865 213.415 ;
        RECT 134.335 213.250 134.505 213.835 ;
        RECT 134.675 213.675 135.245 214.005 ;
        RECT 134.335 213.245 134.905 213.250 ;
        RECT 133.035 213.075 134.905 213.245 ;
        RECT 133.035 212.120 133.205 213.075 ;
        RECT 133.375 212.735 134.345 212.905 ;
        RECT 133.375 212.085 133.545 212.735 ;
        RECT 134.540 212.720 134.905 213.075 ;
        RECT 135.075 212.960 135.245 213.675 ;
        RECT 135.525 213.450 135.695 213.955 ;
        RECT 135.895 213.790 136.115 214.145 ;
        RECT 136.285 213.960 136.880 214.200 ;
        RECT 135.895 213.620 137.180 213.790 ;
        RECT 135.525 213.280 136.645 213.450 ;
        RECT 136.475 213.090 136.645 213.280 ;
        RECT 136.815 213.260 137.180 213.620 ;
        RECT 137.350 213.090 137.520 214.025 ;
        RECT 135.075 212.590 135.745 212.960 ;
        RECT 135.925 212.870 136.255 213.070 ;
        RECT 136.475 212.920 137.520 213.090 ;
        RECT 134.565 212.530 134.735 212.535 ;
        RECT 133.745 212.255 134.905 212.530 ;
        RECT 133.375 211.895 134.905 212.085 ;
        RECT 132.695 211.555 133.720 211.725 ;
        RECT 135.075 211.715 135.245 212.590 ;
        RECT 135.925 212.410 136.225 212.870 ;
        RECT 136.475 212.750 136.735 212.920 ;
        RECT 137.795 212.765 139.575 214.455 ;
        RECT 139.745 214.350 142.060 214.625 ;
        RECT 139.745 212.765 141.230 214.350 ;
        RECT 142.800 212.870 143.405 216.275 ;
        RECT 137.795 212.750 137.965 212.765 ;
        RECT 136.405 212.580 136.735 212.750 ;
        RECT 136.995 212.580 137.965 212.750 ;
        RECT 135.525 212.240 137.625 212.410 ;
        RECT 135.525 212.005 135.695 212.240 ;
        RECT 137.295 212.160 137.625 212.240 ;
        RECT 136.405 211.880 137.125 212.070 ;
        RECT 131.855 211.375 133.285 211.385 ;
        RECT 127.255 210.990 127.810 211.125 ;
        RECT 129.185 211.045 129.355 211.210 ;
        RECT 128.915 210.990 129.355 211.045 ;
        RECT 127.255 210.875 129.355 210.990 ;
        RECT 127.680 210.820 129.045 210.875 ;
        RECT 129.635 210.765 129.805 211.375 ;
        RECT 132.355 211.215 133.285 211.375 ;
        RECT 130.065 211.020 132.185 211.205 ;
        RECT 129.635 210.705 130.265 210.765 ;
        RECT 126.915 210.660 127.545 210.705 ;
        RECT 123.215 210.345 123.990 210.525 ;
        RECT 121.995 210.280 123.990 210.345 ;
        RECT 124.195 210.335 124.825 210.660 ;
        RECT 121.995 210.005 123.385 210.280 ;
        RECT 120.465 209.645 121.645 209.815 ;
        RECT 119.145 209.255 119.705 209.310 ;
        RECT 120.335 209.300 121.260 209.475 ;
        RECT 120.285 209.255 121.260 209.300 ;
        RECT 119.145 209.145 121.260 209.255 ;
        RECT 121.475 209.405 121.645 209.645 ;
        RECT 121.815 209.575 122.485 209.745 ;
        RECT 119.145 209.135 120.415 209.145 ;
        RECT 119.580 209.085 120.415 209.135 ;
        RECT 121.475 209.075 122.145 209.405 ;
        RECT 122.315 209.310 122.485 209.575 ;
        RECT 122.655 209.480 123.305 209.830 ;
        RECT 123.475 209.575 123.935 209.745 ;
        RECT 123.475 209.310 123.645 209.575 ;
        RECT 124.195 209.405 124.365 210.335 ;
        RECT 124.995 210.210 126.285 210.660 ;
        RECT 126.455 210.440 127.545 210.660 ;
        RECT 126.455 210.335 127.085 210.440 ;
        RECT 128.055 210.370 129.005 210.650 ;
        RECT 129.175 210.515 130.265 210.705 ;
        RECT 130.435 210.570 131.385 210.850 ;
        RECT 132.355 210.780 132.525 211.215 ;
        RECT 131.895 210.515 132.525 210.780 ;
        RECT 129.175 210.455 129.805 210.515 ;
        RECT 124.995 209.815 125.165 210.210 ;
        RECT 124.535 209.535 125.165 209.815 ;
        RECT 122.315 209.080 123.645 209.310 ;
        RECT 123.815 209.075 124.365 209.405 ;
        RECT 125.335 209.345 125.895 210.040 ;
        RECT 126.065 209.815 126.285 210.210 ;
        RECT 126.915 209.845 127.085 210.335 ;
        RECT 127.255 210.015 129.375 210.200 ;
        RECT 129.635 209.845 129.805 210.455 ;
        RECT 130.395 210.345 131.760 210.400 ;
        RECT 130.085 210.230 132.185 210.345 ;
        RECT 130.085 210.175 130.525 210.230 ;
        RECT 130.085 210.010 130.255 210.175 ;
        RECT 131.630 210.095 132.185 210.230 ;
        RECT 132.355 210.295 132.525 210.515 ;
        RECT 132.875 210.805 133.285 210.980 ;
        RECT 133.530 210.975 133.720 211.555 ;
        RECT 134.095 210.985 134.265 211.695 ;
        RECT 134.540 211.205 135.245 211.715 ;
        RECT 134.095 210.805 134.870 210.985 ;
        RECT 132.875 210.740 134.870 210.805 ;
        RECT 135.075 210.775 135.245 211.205 ;
        RECT 135.525 211.220 135.695 211.835 ;
        RECT 135.865 211.710 136.195 211.855 ;
        RECT 135.865 211.390 137.155 211.710 ;
        RECT 137.325 211.220 137.495 211.935 ;
        RECT 135.525 211.050 137.495 211.220 ;
        RECT 137.795 211.575 137.965 212.580 ;
        RECT 139.025 212.085 139.860 212.135 ;
        RECT 139.025 212.075 140.295 212.085 ;
        RECT 138.180 211.965 140.295 212.075 ;
        RECT 138.180 211.920 139.155 211.965 ;
        RECT 138.180 211.745 139.105 211.920 ;
        RECT 139.735 211.910 140.295 211.965 ;
        RECT 137.795 211.405 138.975 211.575 ;
        RECT 132.875 210.465 134.265 210.740 ;
        RECT 135.075 210.565 135.775 210.775 ;
        RECT 135.075 210.295 135.245 210.565 ;
        RECT 136.155 210.345 136.485 211.050 ;
        RECT 136.690 210.325 137.065 210.880 ;
        RECT 137.795 210.870 137.965 211.405 ;
        RECT 139.275 211.245 139.605 211.795 ;
        RECT 139.775 211.755 140.295 211.910 ;
        RECT 140.515 211.585 141.230 212.765 ;
        RECT 141.550 212.520 143.405 212.870 ;
        RECT 139.905 211.415 141.230 211.585 ;
        RECT 139.275 211.235 140.300 211.245 ;
        RECT 138.135 211.045 140.300 211.235 ;
        RECT 138.135 210.895 139.070 211.045 ;
        RECT 139.775 210.915 140.300 211.045 ;
        RECT 140.515 210.930 141.230 211.415 ;
        RECT 142.800 210.930 143.405 212.520 ;
        RECT 137.295 210.665 137.965 210.870 ;
        RECT 137.295 210.555 138.465 210.665 ;
        RECT 137.795 210.350 138.465 210.555 ;
        RECT 126.065 209.535 126.745 209.815 ;
        RECT 126.915 209.515 127.585 209.845 ;
        RECT 127.755 209.610 129.085 209.840 ;
        RECT 121.475 208.915 121.645 209.075 ;
        RECT 112.025 207.725 114.775 208.915 ;
        RECT 108.985 207.245 112.375 207.555 ;
        RECT 107.875 206.140 108.045 207.245 ;
        RECT 108.215 206.355 108.765 206.525 ;
        RECT 107.875 205.810 108.425 206.140 ;
        RECT 108.595 205.980 108.765 206.355 ;
        RECT 108.945 206.260 109.315 206.615 ;
        RECT 109.495 206.355 110.425 206.525 ;
        RECT 109.495 205.980 109.665 206.355 ;
        RECT 110.595 206.140 112.375 207.245 ;
        RECT 108.595 205.810 109.665 205.980 ;
        RECT 109.835 205.865 112.375 206.140 ;
        RECT 112.545 207.265 114.775 207.725 ;
        RECT 114.945 208.345 116.205 208.915 ;
        RECT 116.375 208.515 117.055 208.800 ;
        RECT 114.945 208.075 116.665 208.345 ;
        RECT 112.545 205.865 114.255 207.265 ;
        RECT 114.945 207.095 116.205 208.075 ;
        RECT 116.835 208.055 117.055 208.515 ;
        RECT 117.225 208.225 117.785 208.915 ;
        RECT 117.955 208.515 118.585 208.800 ;
        RECT 117.955 208.055 118.125 208.515 ;
        RECT 118.755 208.345 120.215 208.915 ;
        RECT 118.295 208.075 120.215 208.345 ;
        RECT 116.835 207.845 118.125 208.055 ;
        RECT 116.375 207.275 118.585 207.675 ;
        RECT 109.835 205.810 110.765 205.865 ;
        RECT 107.875 205.210 108.045 205.810 ;
        RECT 108.955 205.725 109.285 205.810 ;
        RECT 110.595 205.695 110.765 205.810 ;
        RECT 113.315 205.695 114.255 205.865 ;
        RECT 108.215 205.555 108.790 205.640 ;
        RECT 109.520 205.555 110.425 205.640 ;
        RECT 108.215 205.385 110.425 205.555 ;
        RECT 110.595 205.210 111.855 205.695 ;
        RECT 107.875 204.950 108.885 205.210 ;
        RECT 109.445 205.005 111.855 205.210 ;
        RECT 112.025 205.405 114.255 205.695 ;
        RECT 114.425 206.285 116.205 207.095 ;
        RECT 116.375 206.805 117.055 207.085 ;
        RECT 116.835 206.410 117.055 206.805 ;
        RECT 117.225 206.580 117.785 207.275 ;
        RECT 118.755 207.265 120.215 208.075 ;
        RECT 120.385 208.480 121.645 208.915 ;
        RECT 121.815 208.720 123.935 208.905 ;
        RECT 120.385 208.215 122.105 208.480 ;
        RECT 122.615 208.270 123.565 208.550 ;
        RECT 124.195 208.545 124.365 209.075 ;
        RECT 124.535 208.945 126.745 209.345 ;
        RECT 126.915 208.915 127.085 209.515 ;
        RECT 127.755 209.345 127.925 209.610 ;
        RECT 127.255 209.175 127.925 209.345 ;
        RECT 128.095 209.090 128.745 209.440 ;
        RECT 128.915 209.345 129.085 209.610 ;
        RECT 129.255 209.515 129.805 209.845 ;
        RECT 128.915 209.175 129.375 209.345 ;
        RECT 129.635 208.915 129.805 209.515 ;
        RECT 130.085 209.310 130.255 209.815 ;
        RECT 130.455 209.650 130.675 210.005 ;
        RECT 130.845 209.820 131.440 210.060 ;
        RECT 130.455 209.480 131.740 209.650 ;
        RECT 130.085 209.140 131.205 209.310 ;
        RECT 131.035 208.950 131.205 209.140 ;
        RECT 131.375 209.120 131.740 209.480 ;
        RECT 131.910 208.950 132.080 209.885 ;
        RECT 124.995 208.565 126.285 208.775 ;
        RECT 124.195 208.465 124.825 208.545 ;
        RECT 123.735 208.275 124.825 208.465 ;
        RECT 123.735 208.215 124.365 208.275 ;
        RECT 117.955 206.805 118.585 207.085 ;
        RECT 117.955 206.410 118.125 206.805 ;
        RECT 114.425 205.960 116.665 206.285 ;
        RECT 116.835 205.960 118.125 206.410 ;
        RECT 118.755 206.285 119.695 207.265 ;
        RECT 120.385 207.095 121.645 208.215 ;
        RECT 122.240 208.045 123.605 208.100 ;
        RECT 121.815 207.930 123.915 208.045 ;
        RECT 121.815 207.795 122.370 207.930 ;
        RECT 123.475 207.875 123.915 207.930 ;
        RECT 118.295 205.960 119.695 206.285 ;
        RECT 114.425 205.405 116.205 205.960 ;
        RECT 117.515 205.855 117.845 205.960 ;
        RECT 116.375 205.685 117.345 205.790 ;
        RECT 118.015 205.685 118.585 205.790 ;
        RECT 116.375 205.405 118.585 205.685 ;
        RECT 118.755 205.405 119.695 205.960 ;
        RECT 119.865 206.310 121.645 207.095 ;
        RECT 121.920 206.650 122.090 207.585 ;
        RECT 122.560 207.520 123.155 207.760 ;
        RECT 123.745 207.710 123.915 207.875 ;
        RECT 123.325 207.350 123.545 207.705 ;
        RECT 124.195 207.535 124.365 208.215 ;
        RECT 124.995 208.105 125.165 208.565 ;
        RECT 124.535 207.820 125.165 208.105 ;
        RECT 125.335 207.705 125.895 208.395 ;
        RECT 126.065 208.105 126.285 208.565 ;
        RECT 126.915 208.545 128.175 208.915 ;
        RECT 126.455 208.275 128.175 208.545 ;
        RECT 126.065 207.820 126.745 208.105 ;
        RECT 126.915 207.535 128.175 208.275 ;
        RECT 128.345 208.820 129.805 208.915 ;
        RECT 128.345 208.450 130.305 208.820 ;
        RECT 130.485 208.730 130.815 208.930 ;
        RECT 131.035 208.780 132.080 208.950 ;
        RECT 132.355 209.605 133.615 210.295 ;
        RECT 133.785 209.805 135.245 210.295 ;
        RECT 135.460 210.175 135.985 210.305 ;
        RECT 136.690 210.175 137.625 210.325 ;
        RECT 135.460 209.985 137.625 210.175 ;
        RECT 135.460 209.975 136.485 209.985 ;
        RECT 133.785 209.775 135.855 209.805 ;
        RECT 134.325 209.635 135.855 209.775 ;
        RECT 132.355 209.085 134.155 209.605 ;
        RECT 134.325 209.085 135.245 209.635 ;
        RECT 135.465 209.310 135.985 209.465 ;
        RECT 136.155 209.425 136.485 209.975 ;
        RECT 137.795 209.815 137.965 210.350 ;
        RECT 138.695 210.340 139.070 210.895 ;
        RECT 139.275 210.170 139.605 210.875 ;
        RECT 140.515 210.655 140.685 210.930 ;
        RECT 139.985 210.445 140.685 210.655 ;
        RECT 136.785 209.645 137.965 209.815 ;
        RECT 135.465 209.255 136.025 209.310 ;
        RECT 136.655 209.300 137.580 209.475 ;
        RECT 136.605 209.255 137.580 209.300 ;
        RECT 135.465 209.145 137.580 209.255 ;
        RECT 135.465 209.135 136.735 209.145 ;
        RECT 135.900 209.085 136.735 209.135 ;
        RECT 132.355 208.825 132.525 209.085 ;
        RECT 135.075 208.825 135.245 209.085 ;
        RECT 128.345 207.705 129.805 208.450 ;
        RECT 130.485 208.270 130.785 208.730 ;
        RECT 131.035 208.610 131.295 208.780 ;
        RECT 132.355 208.610 133.270 208.825 ;
        RECT 130.965 208.440 131.295 208.610 ;
        RECT 131.555 208.555 133.270 208.610 ;
        RECT 131.555 208.440 132.525 208.555 ;
        RECT 130.085 208.100 132.185 208.270 ;
        RECT 130.085 207.865 130.255 208.100 ;
        RECT 131.855 208.020 132.185 208.100 ;
        RECT 130.965 207.740 131.685 207.930 ;
        RECT 132.355 207.925 132.525 208.440 ;
        RECT 133.440 208.385 134.425 208.825 ;
        RECT 134.595 208.525 135.245 208.825 ;
        RECT 135.415 208.635 137.625 208.915 ;
        RECT 135.415 208.530 135.985 208.635 ;
        RECT 136.655 208.530 137.625 208.635 ;
        RECT 137.795 208.640 137.965 209.645 ;
        RECT 138.265 210.000 140.235 210.170 ;
        RECT 138.265 209.285 138.435 210.000 ;
        RECT 138.605 209.510 139.895 209.830 ;
        RECT 139.565 209.365 139.895 209.510 ;
        RECT 140.065 209.385 140.235 210.000 ;
        RECT 140.515 209.360 140.685 210.445 ;
        RECT 140.855 209.575 141.405 209.745 ;
        RECT 138.635 209.150 139.355 209.340 ;
        RECT 138.135 208.980 138.465 209.060 ;
        RECT 140.065 208.980 140.235 209.215 ;
        RECT 138.135 208.810 140.235 208.980 ;
        RECT 140.515 209.030 141.065 209.360 ;
        RECT 141.235 209.200 141.405 209.575 ;
        RECT 141.585 209.480 141.955 209.835 ;
        RECT 142.135 209.575 143.065 209.745 ;
        RECT 142.135 209.200 142.305 209.575 ;
        RECT 143.235 209.360 143.405 210.930 ;
        RECT 141.235 209.030 142.305 209.200 ;
        RECT 142.475 209.030 143.405 209.360 ;
        RECT 132.700 208.355 134.425 208.385 ;
        RECT 135.075 208.360 135.245 208.525 ;
        RECT 137.795 208.470 138.765 208.640 ;
        RECT 139.025 208.470 139.355 208.640 ;
        RECT 136.155 208.360 136.485 208.465 ;
        RECT 137.795 208.360 137.965 208.470 ;
        RECT 132.700 208.095 134.880 208.355 ;
        RECT 122.260 207.180 123.545 207.350 ;
        RECT 122.260 206.820 122.625 207.180 ;
        RECT 123.745 207.010 123.915 207.515 ;
        RECT 122.795 206.840 123.915 207.010 ;
        RECT 122.795 206.650 122.965 206.840 ;
        RECT 121.920 206.480 122.965 206.650 ;
        RECT 122.705 206.310 122.965 206.480 ;
        RECT 123.185 206.430 123.515 206.630 ;
        RECT 124.195 206.520 125.655 207.535 ;
        RECT 119.865 206.140 122.445 206.310 ;
        RECT 122.705 206.140 123.035 206.310 ;
        RECT 119.865 205.405 121.645 206.140 ;
        RECT 123.215 205.970 123.515 206.430 ;
        RECT 123.695 206.325 125.655 206.520 ;
        RECT 125.825 206.325 128.695 207.535 ;
        RECT 128.865 206.635 129.805 207.705 ;
        RECT 130.085 207.080 130.255 207.695 ;
        RECT 130.425 207.570 130.755 207.715 ;
        RECT 130.425 207.250 131.715 207.570 ;
        RECT 131.885 207.080 132.055 207.795 ;
        RECT 130.085 206.910 132.055 207.080 ;
        RECT 132.355 207.670 133.255 207.925 ;
        RECT 132.355 207.055 132.530 207.670 ;
        RECT 133.440 207.660 134.425 208.095 ;
        RECT 135.075 208.035 135.705 208.360 ;
        RECT 135.075 207.925 135.245 208.035 ;
        RECT 134.595 207.665 135.245 207.925 ;
        RECT 133.440 207.485 133.665 207.660 ;
        RECT 132.700 207.225 133.665 207.485 ;
        RECT 128.865 206.425 130.335 206.635 ;
        RECT 128.865 206.325 129.805 206.425 ;
        RECT 123.695 206.150 125.135 206.325 ;
        RECT 125.825 206.155 127.085 206.325 ;
        RECT 121.815 205.800 123.915 205.970 ;
        RECT 121.815 205.720 122.145 205.800 ;
        RECT 112.025 205.175 113.485 205.405 ;
        RECT 109.445 204.950 112.395 205.005 ;
        RECT 107.875 204.775 108.045 204.950 ;
        RECT 110.595 204.775 112.395 204.950 ;
        RECT 107.875 204.485 108.770 204.775 ;
        RECT 109.430 204.485 112.395 204.775 ;
        RECT 112.565 204.775 113.485 205.175 ;
        RECT 116.035 204.775 116.205 205.405 ;
        RECT 112.565 204.485 114.210 204.775 ;
        RECT 114.870 204.485 116.205 204.775 ;
        RECT 116.555 204.960 117.945 205.235 ;
        RECT 116.555 204.895 118.550 204.960 ;
        RECT 116.555 204.720 116.965 204.895 ;
        RECT 107.875 203.850 108.045 204.485 ;
        RECT 110.595 203.850 110.765 204.485 ;
        RECT 113.315 204.315 113.485 204.485 ;
        RECT 116.035 204.315 116.965 204.485 ;
        RECT 111.825 204.265 112.660 204.315 ;
        RECT 111.825 204.255 113.095 204.265 ;
        RECT 110.980 204.145 113.095 204.255 ;
        RECT 110.980 204.100 111.955 204.145 ;
        RECT 110.980 203.925 111.905 204.100 ;
        RECT 112.535 204.090 113.095 204.145 ;
        RECT 107.875 203.590 108.885 203.850 ;
        RECT 109.445 203.755 110.765 203.850 ;
        RECT 109.445 203.590 111.775 203.755 ;
        RECT 107.875 202.990 108.045 203.590 ;
        RECT 110.595 203.585 111.775 203.590 ;
        RECT 108.215 203.245 110.425 203.415 ;
        RECT 108.215 203.160 108.790 203.245 ;
        RECT 109.520 203.160 110.425 203.245 ;
        RECT 108.955 202.990 109.285 203.075 ;
        RECT 110.595 202.990 110.765 203.585 ;
        RECT 112.075 203.425 112.405 203.975 ;
        RECT 112.575 203.935 113.095 204.090 ;
        RECT 113.315 204.010 113.995 204.315 ;
        RECT 113.315 203.765 113.485 204.010 ;
        RECT 114.165 204.000 114.725 204.315 ;
        RECT 116.035 204.305 116.205 204.315 ;
        RECT 115.225 204.010 116.205 204.305 ;
        RECT 117.210 204.145 117.400 204.725 ;
        RECT 112.705 203.595 113.485 203.765 ;
        RECT 112.075 203.415 113.100 203.425 ;
        RECT 110.935 203.225 113.100 203.415 ;
        RECT 110.935 203.075 111.870 203.225 ;
        RECT 112.575 203.095 113.100 203.225 ;
        RECT 113.315 203.410 113.485 203.595 ;
        RECT 113.665 203.585 115.865 203.830 ;
        RECT 113.665 203.580 114.725 203.585 ;
        RECT 113.315 203.150 114.010 203.410 ;
        RECT 107.875 202.660 108.425 202.990 ;
        RECT 108.595 202.820 109.665 202.990 ;
        RECT 107.875 201.585 108.045 202.660 ;
        RECT 108.595 202.445 108.765 202.820 ;
        RECT 108.215 202.275 108.765 202.445 ;
        RECT 108.945 202.185 109.315 202.540 ;
        RECT 109.495 202.445 109.665 202.820 ;
        RECT 109.835 202.845 110.765 202.990 ;
        RECT 109.835 202.660 111.265 202.845 ;
        RECT 110.595 202.530 111.265 202.660 ;
        RECT 109.495 202.275 110.425 202.445 ;
        RECT 108.305 201.755 108.765 201.925 ;
        RECT 107.875 201.255 108.425 201.585 ;
        RECT 108.595 201.490 108.765 201.755 ;
        RECT 108.935 201.660 109.585 202.010 ;
        RECT 109.755 201.755 110.425 201.925 ;
        RECT 109.755 201.490 109.925 201.755 ;
        RECT 110.595 201.585 110.765 202.530 ;
        RECT 111.495 202.520 111.870 203.075 ;
        RECT 112.075 202.350 112.405 203.055 ;
        RECT 113.315 202.835 113.485 203.150 ;
        RECT 114.475 202.970 114.725 203.580 ;
        RECT 116.035 203.410 116.205 204.010 ;
        RECT 115.225 203.150 116.205 203.410 ;
        RECT 112.785 202.625 113.485 202.835 ;
        RECT 113.665 202.720 115.860 202.970 ;
        RECT 113.315 202.550 113.485 202.625 ;
        RECT 108.595 201.260 109.925 201.490 ;
        RECT 110.095 201.255 110.765 201.585 ;
        RECT 111.065 202.180 113.035 202.350 ;
        RECT 111.065 201.465 111.235 202.180 ;
        RECT 111.405 201.690 112.695 202.010 ;
        RECT 112.365 201.545 112.695 201.690 ;
        RECT 112.865 201.565 113.035 202.180 ;
        RECT 113.315 202.290 114.045 202.550 ;
        RECT 113.315 201.690 113.485 202.290 ;
        RECT 113.680 201.860 114.305 202.120 ;
        RECT 111.435 201.330 112.155 201.520 ;
        RECT 113.315 201.430 113.965 201.690 ;
        RECT 107.875 200.645 108.045 201.255 ;
        RECT 108.305 200.900 110.425 201.085 ;
        RECT 110.595 200.820 110.765 201.255 ;
        RECT 110.935 201.160 111.265 201.240 ;
        RECT 112.865 201.160 113.035 201.395 ;
        RECT 110.935 200.990 113.035 201.160 ;
        RECT 107.875 200.395 108.505 200.645 ;
        RECT 108.675 200.450 109.625 200.730 ;
        RECT 110.595 200.660 111.565 200.820 ;
        RECT 110.135 200.650 111.565 200.660 ;
        RECT 111.825 200.650 112.155 200.820 ;
        RECT 110.135 200.395 110.765 200.650 ;
        RECT 111.825 200.480 112.085 200.650 ;
        RECT 112.335 200.530 112.635 200.990 ;
        RECT 113.315 200.830 113.485 201.430 ;
        RECT 114.135 201.260 114.305 201.860 ;
        RECT 113.680 201.000 114.305 201.260 ;
        RECT 113.315 200.810 113.965 200.830 ;
        RECT 107.875 198.700 108.045 200.395 ;
        RECT 108.635 200.225 110.000 200.280 ;
        RECT 108.325 200.110 110.425 200.225 ;
        RECT 108.325 200.055 108.765 200.110 ;
        RECT 108.325 199.890 108.495 200.055 ;
        RECT 109.870 199.975 110.425 200.110 ;
        RECT 108.325 199.190 108.495 199.695 ;
        RECT 108.695 199.530 108.915 199.885 ;
        RECT 109.085 199.700 109.680 199.940 ;
        RECT 108.695 199.360 109.980 199.530 ;
        RECT 108.325 199.020 109.445 199.190 ;
        RECT 109.275 198.830 109.445 199.020 ;
        RECT 109.615 199.000 109.980 199.360 ;
        RECT 110.150 198.830 110.320 199.765 ;
        RECT 107.875 198.330 108.545 198.700 ;
        RECT 108.725 198.610 109.055 198.810 ;
        RECT 109.275 198.660 110.320 198.830 ;
        RECT 110.595 198.745 110.765 200.395 ;
        RECT 111.040 200.310 112.085 200.480 ;
        RECT 112.305 200.330 112.635 200.530 ;
        RECT 112.815 200.570 113.965 200.810 ;
        RECT 112.815 200.440 113.485 200.570 ;
        RECT 111.040 199.375 111.210 200.310 ;
        RECT 111.380 199.780 111.745 200.140 ;
        RECT 111.915 200.120 112.085 200.310 ;
        RECT 111.915 199.950 113.035 200.120 ;
        RECT 111.380 199.610 112.665 199.780 ;
        RECT 111.680 199.200 112.275 199.440 ;
        RECT 112.445 199.255 112.665 199.610 ;
        RECT 112.865 199.445 113.035 199.950 ;
        RECT 113.315 199.970 113.485 200.440 ;
        RECT 114.135 200.400 114.305 201.000 ;
        RECT 113.680 200.140 114.305 200.400 ;
        RECT 113.315 199.725 113.965 199.970 ;
        RECT 110.935 199.030 111.490 199.165 ;
        RECT 112.865 199.085 113.035 199.250 ;
        RECT 112.595 199.030 113.035 199.085 ;
        RECT 110.935 198.915 113.035 199.030 ;
        RECT 113.315 199.110 113.485 199.725 ;
        RECT 114.135 199.555 114.305 200.140 ;
        RECT 113.680 199.280 114.305 199.555 ;
        RECT 111.360 198.860 112.725 198.915 ;
        RECT 113.315 198.865 113.965 199.110 ;
        RECT 113.315 198.745 113.485 198.865 ;
        RECT 107.875 196.515 108.045 198.330 ;
        RECT 108.725 198.150 109.025 198.610 ;
        RECT 109.275 198.490 109.535 198.660 ;
        RECT 110.595 198.490 111.225 198.745 ;
        RECT 109.205 198.320 109.535 198.490 ;
        RECT 109.795 198.480 111.225 198.490 ;
        RECT 109.795 198.320 110.765 198.480 ;
        RECT 111.735 198.410 112.685 198.690 ;
        RECT 112.855 198.495 113.485 198.745 ;
        RECT 114.135 198.695 114.305 199.280 ;
        RECT 108.325 197.980 110.425 198.150 ;
        RECT 108.325 197.745 108.495 197.980 ;
        RECT 110.095 197.900 110.425 197.980 ;
        RECT 110.595 197.885 110.765 198.320 ;
        RECT 113.315 198.255 113.485 198.495 ;
        RECT 113.680 198.435 114.305 198.695 ;
        RECT 110.935 198.055 113.055 198.240 ;
        RECT 113.315 198.005 113.965 198.255 ;
        RECT 113.315 197.885 113.485 198.005 ;
        RECT 109.205 197.620 109.925 197.810 ;
        RECT 108.325 196.960 108.495 197.575 ;
        RECT 108.665 197.450 108.995 197.595 ;
        RECT 108.665 197.130 109.955 197.450 ;
        RECT 110.125 196.960 110.295 197.675 ;
        RECT 108.325 196.790 110.295 196.960 ;
        RECT 110.595 197.555 111.265 197.885 ;
        RECT 111.435 197.650 112.765 197.880 ;
        RECT 107.875 196.305 108.575 196.515 ;
        RECT 107.875 195.545 108.045 196.305 ;
        RECT 108.955 196.085 109.285 196.790 ;
        RECT 109.490 196.065 109.865 196.620 ;
        RECT 110.595 196.610 110.765 197.555 ;
        RECT 111.435 197.385 111.605 197.650 ;
        RECT 110.935 197.215 111.605 197.385 ;
        RECT 111.775 197.130 112.425 197.480 ;
        RECT 112.595 197.385 112.765 197.650 ;
        RECT 112.935 197.555 113.485 197.885 ;
        RECT 114.135 197.835 114.305 198.435 ;
        RECT 113.680 197.575 114.305 197.835 ;
        RECT 113.315 197.395 113.485 197.555 ;
        RECT 112.595 197.215 113.055 197.385 ;
        RECT 113.315 197.145 113.965 197.395 ;
        RECT 110.935 196.780 113.145 196.950 ;
        RECT 110.935 196.615 111.905 196.780 ;
        RECT 112.575 196.695 113.145 196.780 ;
        RECT 110.095 196.445 110.765 196.610 ;
        RECT 112.075 196.525 112.405 196.610 ;
        RECT 113.315 196.535 113.485 197.145 ;
        RECT 114.135 196.975 114.305 197.575 ;
        RECT 113.680 196.715 114.305 196.975 ;
        RECT 114.135 196.540 114.305 196.715 ;
        RECT 114.475 196.710 114.725 202.720 ;
        RECT 116.035 202.550 116.205 203.150 ;
        RECT 115.235 202.290 116.205 202.550 ;
        RECT 114.895 201.860 115.860 202.120 ;
        RECT 116.030 201.945 116.205 202.290 ;
        RECT 116.375 203.975 117.400 204.145 ;
        RECT 117.775 204.715 118.550 204.895 ;
        RECT 118.755 204.775 118.925 205.405 ;
        RECT 121.475 204.775 121.645 205.405 ;
        RECT 117.775 204.005 117.945 204.715 ;
        RECT 118.755 204.495 119.650 204.775 ;
        RECT 118.220 204.485 119.650 204.495 ;
        RECT 120.310 204.485 121.645 204.775 ;
        RECT 121.945 204.780 122.115 205.495 ;
        RECT 122.315 205.440 123.035 205.630 ;
        RECT 123.745 205.565 123.915 205.800 ;
        RECT 123.245 205.270 123.575 205.415 ;
        RECT 122.285 204.950 123.575 205.270 ;
        RECT 123.745 204.780 123.915 205.395 ;
        RECT 121.945 204.610 123.915 204.780 ;
        RECT 124.195 204.945 125.135 206.150 ;
        RECT 125.305 205.685 127.085 206.155 ;
        RECT 129.635 205.695 129.805 206.325 ;
        RECT 130.715 206.205 131.045 206.910 ;
        RECT 132.355 206.810 133.255 207.055 ;
        RECT 131.250 206.185 131.625 206.740 ;
        RECT 132.355 206.730 132.530 206.810 ;
        RECT 131.855 206.415 132.530 206.730 ;
        RECT 133.425 206.625 133.665 207.225 ;
        RECT 132.355 206.195 132.530 206.415 ;
        RECT 132.700 206.365 133.665 206.625 ;
        RECT 130.020 206.035 130.545 206.165 ;
        RECT 131.250 206.035 132.185 206.185 ;
        RECT 130.020 205.845 132.185 206.035 ;
        RECT 132.355 205.950 133.255 206.195 ;
        RECT 130.020 205.835 131.045 205.845 ;
        RECT 125.305 205.390 127.895 205.685 ;
        RECT 125.305 204.945 127.085 205.390 ;
        RECT 128.395 205.380 128.955 205.695 ;
        RECT 129.125 205.665 129.805 205.695 ;
        RECT 129.125 205.495 130.415 205.665 ;
        RECT 129.125 205.390 129.805 205.495 ;
        RECT 127.255 204.965 129.455 205.210 ;
        RECT 124.195 204.775 124.365 204.945 ;
        RECT 126.915 204.790 127.085 204.945 ;
        RECT 128.395 204.960 129.455 204.965 ;
        RECT 126.915 204.775 127.895 204.790 ;
        RECT 118.220 203.985 118.925 204.485 ;
        RECT 121.475 204.430 121.645 204.485 ;
        RECT 119.185 204.055 119.645 204.225 ;
        RECT 116.375 202.285 116.545 203.975 ;
        RECT 118.755 203.885 118.925 203.985 ;
        RECT 117.055 203.615 118.585 203.805 ;
        RECT 116.715 202.625 116.885 203.580 ;
        RECT 117.055 202.965 117.225 203.615 ;
        RECT 118.755 203.555 119.305 203.885 ;
        RECT 119.475 203.790 119.645 204.055 ;
        RECT 119.815 203.960 120.465 204.310 ;
        RECT 120.635 204.055 121.305 204.225 ;
        RECT 121.475 204.115 122.145 204.430 ;
        RECT 120.635 203.790 120.805 204.055 ;
        RECT 121.475 203.885 121.645 204.115 ;
        RECT 122.375 203.885 122.750 204.440 ;
        RECT 122.955 203.905 123.285 204.610 ;
        RECT 124.195 204.485 125.090 204.775 ;
        RECT 125.750 204.530 127.895 204.775 ;
        RECT 125.750 204.485 127.085 204.530 ;
        RECT 124.195 204.335 124.365 204.485 ;
        RECT 123.665 204.305 124.365 204.335 ;
        RECT 123.665 204.125 125.175 204.305 ;
        RECT 124.195 204.035 125.175 204.125 ;
        RECT 119.475 203.560 120.805 203.790 ;
        RECT 120.975 203.555 121.645 203.885 ;
        RECT 117.425 203.170 118.585 203.445 ;
        RECT 117.565 203.165 117.735 203.170 ;
        RECT 117.055 202.795 118.025 202.965 ;
        RECT 118.220 202.625 118.585 202.980 ;
        RECT 116.715 202.455 118.585 202.625 ;
        RECT 118.015 202.450 118.585 202.455 ;
        RECT 118.755 202.945 118.925 203.555 ;
        RECT 119.185 203.200 121.305 203.385 ;
        RECT 121.475 203.375 121.645 203.555 ;
        RECT 121.815 203.735 122.750 203.885 ;
        RECT 123.455 203.735 123.980 203.865 ;
        RECT 121.815 203.545 123.980 203.735 ;
        RECT 122.955 203.535 123.980 203.545 ;
        RECT 121.475 203.205 122.655 203.375 ;
        RECT 118.755 202.695 119.385 202.945 ;
        RECT 119.555 202.750 120.505 203.030 ;
        RECT 121.475 202.960 121.645 203.205 ;
        RECT 121.015 202.695 121.645 202.960 ;
        RECT 121.860 202.860 122.785 203.035 ;
        RECT 122.955 202.985 123.285 203.535 ;
        RECT 124.195 203.365 124.365 204.035 ;
        RECT 125.355 203.965 125.605 204.315 ;
        RECT 126.915 204.305 127.085 204.485 ;
        RECT 128.395 204.350 128.645 204.960 ;
        RECT 129.635 204.790 129.805 205.390 ;
        RECT 130.025 205.170 130.545 205.325 ;
        RECT 130.715 205.285 131.045 205.835 ;
        RECT 132.355 205.675 132.530 205.950 ;
        RECT 133.425 205.765 133.665 206.365 ;
        RECT 131.345 205.505 132.530 205.675 ;
        RECT 132.700 205.505 133.665 205.765 ;
        RECT 132.355 205.335 132.530 205.505 ;
        RECT 130.025 205.115 130.585 205.170 ;
        RECT 131.215 205.160 132.140 205.335 ;
        RECT 131.165 205.115 132.140 205.160 ;
        RECT 130.025 205.005 132.140 205.115 ;
        RECT 132.355 205.090 133.255 205.335 ;
        RECT 130.025 204.995 131.295 205.005 ;
        RECT 130.460 204.945 131.295 204.995 ;
        RECT 129.110 204.775 129.805 204.790 ;
        RECT 132.355 204.775 132.530 205.090 ;
        RECT 133.425 204.920 133.665 205.505 ;
        RECT 129.110 204.530 130.530 204.775 ;
        RECT 129.635 204.485 130.530 204.530 ;
        RECT 131.190 204.490 132.530 204.775 ;
        RECT 132.700 204.660 133.665 204.920 ;
        RECT 131.190 204.485 133.255 204.490 ;
        RECT 125.775 203.975 127.085 204.305 ;
        RECT 127.260 204.100 129.455 204.350 ;
        RECT 126.915 203.930 127.085 203.975 ;
        RECT 124.535 203.795 125.175 203.865 ;
        RECT 124.535 203.625 125.945 203.795 ;
        RECT 124.535 203.535 125.175 203.625 ;
        RECT 123.585 203.195 125.175 203.365 ;
        RECT 124.195 203.125 125.175 203.195 ;
        RECT 123.455 202.870 123.975 203.025 ;
        RECT 121.860 202.815 122.835 202.860 ;
        RECT 123.415 202.815 123.975 202.870 ;
        RECT 121.860 202.705 123.975 202.815 ;
        RECT 116.375 202.115 117.845 202.285 ;
        RECT 117.515 202.090 117.845 202.115 ;
        RECT 114.895 201.260 115.135 201.860 ;
        RECT 116.030 201.775 117.345 201.945 ;
        RECT 118.015 201.865 118.185 202.450 ;
        RECT 118.755 202.025 118.925 202.695 ;
        RECT 119.515 202.525 120.880 202.580 ;
        RECT 119.205 202.410 121.305 202.525 ;
        RECT 119.205 202.355 119.645 202.410 ;
        RECT 119.205 202.190 119.375 202.355 ;
        RECT 120.750 202.275 121.305 202.410 ;
        RECT 116.030 201.690 116.205 201.775 ;
        RECT 115.305 201.430 116.205 201.690 ;
        RECT 117.515 201.695 118.185 201.865 ;
        RECT 118.355 201.695 118.925 202.025 ;
        RECT 117.515 201.610 117.845 201.695 ;
        RECT 114.895 201.000 115.860 201.260 ;
        RECT 116.030 201.095 116.205 201.430 ;
        RECT 116.375 201.440 117.345 201.605 ;
        RECT 118.015 201.440 118.585 201.525 ;
        RECT 116.375 201.270 118.585 201.440 ;
        RECT 118.755 201.095 118.925 201.695 ;
        RECT 119.205 201.490 119.375 201.995 ;
        RECT 119.575 201.830 119.795 202.185 ;
        RECT 119.965 202.000 120.560 202.240 ;
        RECT 119.575 201.660 120.860 201.830 ;
        RECT 119.205 201.320 120.325 201.490 ;
        RECT 120.155 201.130 120.325 201.320 ;
        RECT 120.495 201.300 120.860 201.660 ;
        RECT 121.030 201.130 121.200 202.065 ;
        RECT 114.895 200.400 115.135 201.000 ;
        RECT 116.030 200.830 117.295 201.095 ;
        RECT 115.305 200.570 117.295 200.830 ;
        RECT 114.895 200.140 115.860 200.400 ;
        RECT 116.030 200.175 117.295 200.570 ;
        RECT 117.465 201.000 118.925 201.095 ;
        RECT 117.465 200.630 119.425 201.000 ;
        RECT 119.605 200.910 119.935 201.110 ;
        RECT 120.155 200.960 121.200 201.130 ;
        RECT 121.475 201.965 121.645 202.695 ;
        RECT 122.705 202.695 123.975 202.705 ;
        RECT 122.705 202.645 123.540 202.695 ;
        RECT 121.815 202.300 124.025 202.470 ;
        RECT 121.815 202.135 122.785 202.300 ;
        RECT 123.455 202.215 124.025 202.300 ;
        RECT 124.195 202.335 124.365 203.125 ;
        RECT 125.355 203.105 125.605 203.455 ;
        RECT 125.775 203.445 125.945 203.625 ;
        RECT 126.915 203.670 127.885 203.930 ;
        RECT 125.775 203.115 126.730 203.445 ;
        RECT 126.915 203.070 127.090 203.670 ;
        RECT 127.260 203.240 128.225 203.500 ;
        RECT 124.535 202.505 125.185 202.835 ;
        RECT 122.955 202.045 123.285 202.130 ;
        RECT 124.195 202.045 124.825 202.335 ;
        RECT 121.475 201.795 122.785 201.965 ;
        RECT 122.955 201.875 123.625 202.045 ;
        RECT 117.465 200.345 118.925 200.630 ;
        RECT 119.605 200.450 119.905 200.910 ;
        RECT 120.155 200.790 120.415 200.960 ;
        RECT 121.475 200.790 121.645 201.795 ;
        RECT 122.955 201.625 123.285 201.650 ;
        RECT 120.085 200.620 120.415 200.790 ;
        RECT 120.675 200.620 121.645 200.790 ;
        RECT 114.895 199.540 115.135 200.140 ;
        RECT 116.030 199.970 117.815 200.175 ;
        RECT 115.305 199.710 117.815 199.970 ;
        RECT 114.895 199.280 115.860 199.540 ;
        RECT 116.030 199.425 117.815 199.710 ;
        RECT 117.985 199.425 118.925 200.345 ;
        RECT 119.205 200.280 121.305 200.450 ;
        RECT 119.205 200.045 119.375 200.280 ;
        RECT 120.975 200.200 121.305 200.280 ;
        RECT 120.085 199.920 120.805 200.110 ;
        RECT 114.895 198.695 115.135 199.280 ;
        RECT 116.030 199.110 116.205 199.425 ;
        RECT 115.305 198.865 116.205 199.110 ;
        RECT 116.375 198.995 117.045 199.165 ;
        RECT 116.030 198.825 116.205 198.865 ;
        RECT 114.895 198.435 115.860 198.695 ;
        RECT 116.030 198.495 116.705 198.825 ;
        RECT 116.875 198.730 117.045 198.995 ;
        RECT 117.215 198.900 117.865 199.250 ;
        RECT 118.035 198.995 118.495 199.165 ;
        RECT 118.035 198.730 118.205 198.995 ;
        RECT 118.755 198.825 118.925 199.425 ;
        RECT 119.205 199.260 119.375 199.875 ;
        RECT 119.545 199.750 119.875 199.895 ;
        RECT 119.545 199.430 120.835 199.750 ;
        RECT 121.005 199.260 121.175 199.975 ;
        RECT 119.205 199.090 121.175 199.260 ;
        RECT 121.475 199.425 121.645 200.620 ;
        RECT 121.815 201.455 123.285 201.625 ;
        RECT 121.815 199.765 121.985 201.455 ;
        RECT 123.455 201.290 123.625 201.875 ;
        RECT 123.795 202.005 124.825 202.045 ;
        RECT 123.795 201.715 124.365 202.005 ;
        RECT 125.015 201.790 125.185 202.505 ;
        RECT 125.355 202.365 125.605 202.875 ;
        RECT 126.915 202.815 127.815 203.070 ;
        RECT 125.795 202.810 127.815 202.815 ;
        RECT 125.795 202.485 127.090 202.810 ;
        RECT 127.985 202.640 128.225 203.240 ;
        RECT 126.915 202.210 127.090 202.485 ;
        RECT 127.260 202.380 128.225 202.640 ;
        RECT 123.455 201.285 124.025 201.290 ;
        RECT 122.155 201.115 124.025 201.285 ;
        RECT 122.155 200.160 122.325 201.115 ;
        RECT 122.495 200.775 123.465 200.945 ;
        RECT 122.495 200.125 122.665 200.775 ;
        RECT 123.660 200.760 124.025 201.115 ;
        RECT 124.195 201.260 124.365 201.715 ;
        RECT 124.535 201.460 125.185 201.790 ;
        RECT 125.355 201.785 126.670 202.155 ;
        RECT 126.915 201.950 127.815 202.210 ;
        RECT 124.195 200.930 124.825 201.260 ;
        RECT 123.005 200.570 123.175 200.575 ;
        RECT 122.865 200.295 124.025 200.570 ;
        RECT 122.495 199.935 124.025 200.125 ;
        RECT 124.195 199.765 124.365 200.930 ;
        RECT 125.015 200.705 125.185 201.460 ;
        RECT 125.355 201.285 126.670 201.615 ;
        RECT 126.915 201.350 127.090 201.950 ;
        RECT 127.985 201.780 128.225 202.380 ;
        RECT 127.260 201.520 128.225 201.780 ;
        RECT 126.915 201.090 127.815 201.350 ;
        RECT 125.355 200.745 126.670 201.075 ;
        RECT 124.695 200.535 125.185 200.705 ;
        RECT 124.550 200.035 125.185 200.365 ;
        RECT 125.355 200.155 125.565 200.575 ;
        RECT 126.915 200.490 127.090 201.090 ;
        RECT 127.985 200.920 128.225 201.520 ;
        RECT 127.260 200.660 128.225 200.920 ;
        RECT 125.735 200.225 126.745 200.475 ;
        RECT 126.915 200.245 127.815 200.490 ;
        RECT 124.995 199.985 125.185 200.035 ;
        RECT 125.735 199.985 126.025 200.225 ;
        RECT 126.915 200.055 127.090 200.245 ;
        RECT 127.985 200.075 128.225 200.660 ;
        RECT 121.815 199.595 122.840 199.765 ;
        RECT 124.195 199.755 124.825 199.765 ;
        RECT 121.475 199.255 122.405 199.425 ;
        RECT 116.875 198.500 118.205 198.730 ;
        RECT 118.375 198.815 118.925 198.825 ;
        RECT 118.375 198.605 119.455 198.815 ;
        RECT 118.375 198.495 118.925 198.605 ;
        RECT 114.895 197.835 115.135 198.435 ;
        RECT 116.030 198.250 116.205 198.495 ;
        RECT 115.305 198.005 116.205 198.250 ;
        RECT 116.375 198.140 118.495 198.325 ;
        RECT 116.030 197.900 116.205 198.005 ;
        RECT 114.895 197.575 115.860 197.835 ;
        RECT 116.030 197.635 116.665 197.900 ;
        RECT 117.175 197.690 118.125 197.970 ;
        RECT 118.755 197.885 118.925 198.495 ;
        RECT 119.835 198.385 120.165 199.090 ;
        RECT 120.370 198.365 120.745 198.920 ;
        RECT 121.475 198.910 121.645 199.255 ;
        RECT 120.975 198.595 121.645 198.910 ;
        RECT 119.140 198.215 119.665 198.345 ;
        RECT 120.370 198.215 121.305 198.365 ;
        RECT 119.140 198.025 121.305 198.215 ;
        RECT 119.140 198.015 120.165 198.025 ;
        RECT 118.295 197.845 118.925 197.885 ;
        RECT 118.295 197.675 119.535 197.845 ;
        RECT 118.295 197.635 118.925 197.675 ;
        RECT 114.895 196.975 115.135 197.575 ;
        RECT 116.030 197.390 116.205 197.635 ;
        RECT 116.800 197.465 118.165 197.520 ;
        RECT 115.305 197.145 116.205 197.390 ;
        RECT 116.375 197.350 118.475 197.465 ;
        RECT 116.375 197.215 116.930 197.350 ;
        RECT 118.035 197.295 118.475 197.350 ;
        RECT 114.895 196.715 115.860 196.975 ;
        RECT 114.895 196.540 115.120 196.715 ;
        RECT 113.315 196.525 113.965 196.535 ;
        RECT 110.095 196.295 111.905 196.445 ;
        RECT 112.075 196.355 112.745 196.525 ;
        RECT 110.595 196.275 111.905 196.295 ;
        RECT 108.260 195.915 108.785 196.045 ;
        RECT 109.490 195.915 110.425 196.065 ;
        RECT 108.260 195.725 110.425 195.915 ;
        RECT 108.260 195.715 109.285 195.725 ;
        RECT 107.875 195.375 108.655 195.545 ;
        RECT 107.875 194.650 108.045 195.375 ;
        RECT 108.265 195.050 108.785 195.205 ;
        RECT 108.955 195.165 109.285 195.715 ;
        RECT 110.595 195.555 110.765 196.275 ;
        RECT 112.075 196.105 112.405 196.130 ;
        RECT 109.585 195.385 110.765 195.555 ;
        RECT 108.265 194.995 108.825 195.050 ;
        RECT 109.455 195.040 110.380 195.215 ;
        RECT 109.405 194.995 110.380 195.040 ;
        RECT 108.265 194.885 110.380 194.995 ;
        RECT 108.265 194.875 109.535 194.885 ;
        RECT 108.700 194.825 109.535 194.875 ;
        RECT 110.595 194.650 110.765 195.385 ;
        RECT 107.875 194.390 108.885 194.650 ;
        RECT 109.445 194.390 110.765 194.650 ;
        RECT 107.875 193.790 108.045 194.390 ;
        RECT 108.215 194.045 110.425 194.215 ;
        RECT 108.215 193.960 108.790 194.045 ;
        RECT 109.520 193.960 110.425 194.045 ;
        RECT 110.595 193.905 110.765 194.390 ;
        RECT 110.935 195.935 112.405 196.105 ;
        RECT 110.935 194.245 111.105 195.935 ;
        RECT 112.575 195.770 112.745 196.355 ;
        RECT 112.915 196.275 113.965 196.525 ;
        RECT 112.915 196.195 113.485 196.275 ;
        RECT 112.575 195.765 113.145 195.770 ;
        RECT 111.275 195.595 113.145 195.765 ;
        RECT 111.275 194.640 111.445 195.595 ;
        RECT 111.615 195.255 112.585 195.425 ;
        RECT 111.615 194.605 111.785 195.255 ;
        RECT 112.780 195.240 113.145 195.595 ;
        RECT 113.315 195.675 113.485 196.195 ;
        RECT 114.135 196.105 115.120 196.540 ;
        RECT 116.030 196.530 116.205 197.145 ;
        RECT 115.305 196.275 116.205 196.530 ;
        RECT 113.680 195.845 115.860 196.105 ;
        RECT 114.135 195.815 115.860 195.845 ;
        RECT 113.315 195.375 113.965 195.675 ;
        RECT 114.135 195.375 115.120 195.815 ;
        RECT 116.035 195.730 116.205 196.275 ;
        RECT 116.480 196.070 116.650 197.005 ;
        RECT 117.120 196.940 117.715 197.180 ;
        RECT 118.305 197.130 118.475 197.295 ;
        RECT 117.885 196.770 118.105 197.125 ;
        RECT 118.755 196.945 118.925 197.635 ;
        RECT 119.145 197.350 119.665 197.505 ;
        RECT 119.835 197.465 120.165 198.015 ;
        RECT 121.475 197.855 121.645 198.595 ;
        RECT 121.995 198.845 122.405 199.020 ;
        RECT 122.650 199.015 122.840 199.595 ;
        RECT 123.215 199.025 123.385 199.735 ;
        RECT 123.660 199.595 124.825 199.755 ;
        RECT 124.995 199.725 126.025 199.985 ;
        RECT 126.195 199.725 127.090 200.055 ;
        RECT 127.260 199.815 128.225 200.075 ;
        RECT 124.995 199.615 125.565 199.725 ;
        RECT 123.660 199.245 124.365 199.595 ;
        RECT 125.355 199.405 125.565 199.615 ;
        RECT 126.915 199.630 127.090 199.725 ;
        RECT 123.215 198.845 123.990 199.025 ;
        RECT 121.995 198.780 123.990 198.845 ;
        RECT 121.995 198.505 123.385 198.780 ;
        RECT 121.815 198.055 124.025 198.335 ;
        RECT 121.815 197.950 122.785 198.055 ;
        RECT 123.455 197.950 124.025 198.055 ;
        RECT 124.195 198.240 124.365 199.245 ;
        RECT 124.535 199.235 125.165 199.305 ;
        RECT 125.735 199.235 126.745 199.490 ;
        RECT 124.535 198.965 126.745 199.235 ;
        RECT 126.915 199.385 127.815 199.630 ;
        RECT 124.535 198.515 126.745 198.795 ;
        RECT 124.535 198.410 125.105 198.515 ;
        RECT 125.775 198.410 126.745 198.515 ;
        RECT 126.915 198.770 127.090 199.385 ;
        RECT 127.985 199.215 128.225 199.815 ;
        RECT 127.260 198.955 128.225 199.215 ;
        RECT 126.915 198.525 127.815 198.770 ;
        RECT 125.275 198.240 125.605 198.345 ;
        RECT 126.915 198.240 127.090 198.525 ;
        RECT 127.985 198.355 128.225 198.955 ;
        RECT 124.195 197.915 124.825 198.240 ;
        RECT 120.465 197.780 121.645 197.855 ;
        RECT 122.955 197.780 123.285 197.885 ;
        RECT 124.195 197.780 124.365 197.915 ;
        RECT 120.465 197.685 122.105 197.780 ;
        RECT 119.145 197.295 119.705 197.350 ;
        RECT 120.335 197.340 121.260 197.515 ;
        RECT 120.285 197.295 121.260 197.340 ;
        RECT 119.145 197.185 121.260 197.295 ;
        RECT 121.475 197.455 122.105 197.685 ;
        RECT 119.145 197.175 120.415 197.185 ;
        RECT 119.580 197.125 120.415 197.175 ;
        RECT 116.820 196.600 118.105 196.770 ;
        RECT 116.820 196.240 117.185 196.600 ;
        RECT 118.305 196.430 118.475 196.935 ;
        RECT 117.355 196.260 118.475 196.430 ;
        RECT 118.755 196.615 119.430 196.945 ;
        RECT 120.285 196.890 120.455 196.895 ;
        RECT 117.355 196.070 117.525 196.260 ;
        RECT 116.480 195.900 117.525 196.070 ;
        RECT 117.265 195.730 117.525 195.900 ;
        RECT 117.745 195.850 118.075 196.050 ;
        RECT 118.755 195.940 118.925 196.615 ;
        RECT 119.605 196.590 120.455 196.890 ;
        RECT 120.625 196.695 121.285 196.865 ;
        RECT 119.120 196.420 119.495 196.445 ;
        RECT 120.625 196.420 120.855 196.695 ;
        RECT 121.475 196.525 121.645 197.455 ;
        RECT 122.275 197.330 123.565 197.780 ;
        RECT 123.735 197.455 124.365 197.780 ;
        RECT 122.275 196.935 122.495 197.330 ;
        RECT 121.815 196.655 122.495 196.935 ;
        RECT 119.120 196.205 120.855 196.420 ;
        RECT 116.035 195.645 117.005 195.730 ;
        RECT 115.290 195.560 117.005 195.645 ;
        RECT 117.265 195.560 117.595 195.730 ;
        RECT 115.290 195.375 116.205 195.560 ;
        RECT 117.775 195.390 118.075 195.850 ;
        RECT 118.255 195.570 118.925 195.940 ;
        RECT 119.645 196.185 120.855 196.205 ;
        RECT 121.025 196.195 121.645 196.525 ;
        RECT 122.665 196.465 123.225 197.160 ;
        RECT 123.395 196.935 123.565 197.330 ;
        RECT 123.395 196.655 124.025 196.935 ;
        RECT 119.110 195.755 119.450 195.925 ;
        RECT 119.645 195.865 119.975 196.185 ;
        RECT 113.315 195.115 113.485 195.375 ;
        RECT 116.035 195.115 116.205 195.375 ;
        RECT 116.375 195.220 118.475 195.390 ;
        RECT 116.375 195.140 116.705 195.220 ;
        RECT 112.125 195.050 112.295 195.055 ;
        RECT 111.985 194.775 113.145 195.050 ;
        RECT 111.615 194.415 113.145 194.605 ;
        RECT 113.315 194.595 114.775 195.115 ;
        RECT 110.935 194.075 111.960 194.245 ;
        RECT 113.315 194.235 114.235 194.595 ;
        RECT 114.945 194.425 116.205 195.115 ;
        RECT 108.955 193.790 109.285 193.875 ;
        RECT 110.595 193.790 111.525 193.905 ;
        RECT 107.875 193.460 108.425 193.790 ;
        RECT 108.595 193.620 109.665 193.790 ;
        RECT 107.875 191.895 108.045 193.460 ;
        RECT 108.595 193.245 108.765 193.620 ;
        RECT 108.215 193.075 108.765 193.245 ;
        RECT 108.945 192.985 109.315 193.340 ;
        RECT 109.495 193.245 109.665 193.620 ;
        RECT 109.835 193.735 111.525 193.790 ;
        RECT 109.835 193.460 110.765 193.735 ;
        RECT 109.495 193.075 110.425 193.245 ;
        RECT 110.595 191.895 110.765 193.460 ;
        RECT 111.115 193.325 111.525 193.500 ;
        RECT 111.770 193.495 111.960 194.075 ;
        RECT 112.335 193.505 112.505 194.215 ;
        RECT 112.780 193.905 114.235 194.235 ;
        RECT 114.405 193.905 116.205 194.425 ;
        RECT 116.505 194.200 116.675 194.915 ;
        RECT 116.875 194.860 117.595 195.050 ;
        RECT 118.305 194.985 118.475 195.220 ;
        RECT 118.755 195.165 118.925 195.570 ;
        RECT 119.255 195.695 119.450 195.755 ;
        RECT 120.145 195.710 121.260 195.995 ;
        RECT 120.145 195.695 120.315 195.710 ;
        RECT 119.255 195.525 120.315 195.695 ;
        RECT 121.475 195.665 121.645 196.195 ;
        RECT 121.815 196.065 124.025 196.465 ;
        RECT 124.195 196.125 124.365 197.455 ;
        RECT 124.995 197.790 126.285 198.240 ;
        RECT 126.455 197.915 127.090 198.240 ;
        RECT 127.260 198.095 128.225 198.355 ;
        RECT 124.995 197.395 125.165 197.790 ;
        RECT 124.535 197.115 125.165 197.395 ;
        RECT 125.335 196.925 125.895 197.620 ;
        RECT 126.065 197.395 126.285 197.790 ;
        RECT 126.915 197.910 127.090 197.915 ;
        RECT 128.000 197.920 128.225 198.095 ;
        RECT 128.395 198.090 128.645 204.100 ;
        RECT 129.635 203.930 129.805 204.485 ;
        RECT 130.065 204.055 130.525 204.225 ;
        RECT 129.075 203.885 129.805 203.930 ;
        RECT 129.075 203.670 130.185 203.885 ;
        RECT 129.635 203.555 130.185 203.670 ;
        RECT 130.355 203.790 130.525 204.055 ;
        RECT 130.695 203.960 131.345 204.310 ;
        RECT 132.355 204.230 133.255 204.485 ;
        RECT 131.515 204.055 132.185 204.225 ;
        RECT 131.515 203.790 131.685 204.055 ;
        RECT 132.355 203.885 132.530 204.230 ;
        RECT 133.425 204.060 133.665 204.660 ;
        RECT 130.355 203.560 131.685 203.790 ;
        RECT 131.855 203.630 132.530 203.885 ;
        RECT 132.700 203.800 133.665 204.060 ;
        RECT 131.855 203.555 133.255 203.630 ;
        RECT 128.815 203.240 129.440 203.500 ;
        RECT 128.815 202.640 128.985 203.240 ;
        RECT 129.635 203.070 129.805 203.555 ;
        RECT 130.065 203.200 132.185 203.385 ;
        RECT 132.355 203.370 133.255 203.555 ;
        RECT 129.155 202.945 129.805 203.070 ;
        RECT 129.155 202.810 130.265 202.945 ;
        RECT 129.635 202.695 130.265 202.810 ;
        RECT 130.435 202.750 131.385 203.030 ;
        RECT 132.355 202.960 132.530 203.370 ;
        RECT 133.425 203.200 133.665 203.800 ;
        RECT 131.895 202.770 132.530 202.960 ;
        RECT 132.700 202.940 133.665 203.200 ;
        RECT 131.895 202.695 133.255 202.770 ;
        RECT 128.815 202.380 129.440 202.640 ;
        RECT 128.815 201.780 128.985 202.380 ;
        RECT 129.635 202.210 129.805 202.695 ;
        RECT 130.395 202.525 131.760 202.580 ;
        RECT 129.155 201.950 129.805 202.210 ;
        RECT 130.085 202.410 132.185 202.525 ;
        RECT 130.085 202.355 130.525 202.410 ;
        RECT 130.085 202.190 130.255 202.355 ;
        RECT 131.630 202.275 132.185 202.410 ;
        RECT 132.355 202.510 133.255 202.695 ;
        RECT 128.815 201.520 129.440 201.780 ;
        RECT 128.815 200.935 128.985 201.520 ;
        RECT 129.635 201.350 129.805 201.950 ;
        RECT 129.155 201.105 129.805 201.350 ;
        RECT 130.085 201.490 130.255 201.995 ;
        RECT 130.455 201.830 130.675 202.185 ;
        RECT 130.845 202.000 131.440 202.240 ;
        RECT 130.455 201.660 131.740 201.830 ;
        RECT 130.085 201.320 131.205 201.490 ;
        RECT 131.035 201.130 131.205 201.320 ;
        RECT 131.375 201.300 131.740 201.660 ;
        RECT 131.910 201.130 132.080 202.065 ;
        RECT 129.635 201.000 129.805 201.105 ;
        RECT 128.815 200.660 129.440 200.935 ;
        RECT 128.815 200.075 128.985 200.660 ;
        RECT 129.635 200.630 130.305 201.000 ;
        RECT 130.485 200.910 130.815 201.110 ;
        RECT 131.035 200.960 132.080 201.130 ;
        RECT 132.355 201.910 132.530 202.510 ;
        RECT 133.425 202.340 133.665 202.940 ;
        RECT 132.700 202.080 133.665 202.340 ;
        RECT 132.355 201.650 133.325 201.910 ;
        RECT 132.355 201.050 132.525 201.650 ;
        RECT 133.835 201.480 134.085 207.490 ;
        RECT 134.255 207.485 134.425 207.660 ;
        RECT 134.255 207.225 134.880 207.485 ;
        RECT 134.255 206.625 134.425 207.225 ;
        RECT 135.075 207.055 135.245 207.665 ;
        RECT 135.875 207.910 137.165 208.360 ;
        RECT 137.335 208.035 137.965 208.360 ;
        RECT 139.025 208.300 139.285 208.470 ;
        RECT 139.535 208.350 139.835 208.810 ;
        RECT 140.515 208.630 140.685 209.030 ;
        RECT 141.595 208.945 141.925 209.030 ;
        RECT 135.875 207.515 136.045 207.910 ;
        RECT 135.415 207.235 136.045 207.515 ;
        RECT 134.595 206.805 135.245 207.055 ;
        RECT 136.215 207.045 136.775 207.740 ;
        RECT 136.945 207.515 137.165 207.910 ;
        RECT 136.945 207.235 137.625 207.515 ;
        RECT 134.255 206.365 134.880 206.625 ;
        RECT 134.255 205.765 134.425 206.365 ;
        RECT 135.075 206.245 135.245 206.805 ;
        RECT 135.415 206.645 137.625 207.045 ;
        RECT 137.795 206.565 137.965 208.035 ;
        RECT 138.240 208.130 139.285 208.300 ;
        RECT 139.505 208.150 139.835 208.350 ;
        RECT 140.015 208.430 140.685 208.630 ;
        RECT 140.855 208.775 141.430 208.860 ;
        RECT 142.160 208.775 143.065 208.860 ;
        RECT 140.855 208.605 143.065 208.775 ;
        RECT 143.235 208.430 143.405 209.030 ;
        RECT 140.015 208.260 141.525 208.430 ;
        RECT 140.515 208.170 141.525 208.260 ;
        RECT 142.085 208.170 143.405 208.430 ;
        RECT 138.240 207.195 138.410 208.130 ;
        RECT 138.580 207.600 138.945 207.960 ;
        RECT 139.115 207.940 139.285 208.130 ;
        RECT 139.115 207.770 140.235 207.940 ;
        RECT 138.580 207.430 139.865 207.600 ;
        RECT 138.880 207.020 139.475 207.260 ;
        RECT 139.645 207.075 139.865 207.430 ;
        RECT 140.065 207.265 140.235 207.770 ;
        RECT 138.135 206.850 138.690 206.985 ;
        RECT 140.065 206.905 140.235 207.070 ;
        RECT 139.795 206.850 140.235 206.905 ;
        RECT 138.135 206.735 140.235 206.850 ;
        RECT 140.515 206.935 140.685 208.170 ;
        RECT 140.855 207.825 142.265 207.995 ;
        RECT 143.235 207.985 143.405 208.170 ;
        RECT 140.855 207.505 141.425 207.825 ;
        RECT 140.855 207.105 141.425 207.335 ;
        RECT 141.595 207.250 141.925 207.655 ;
        RECT 142.095 207.475 142.265 207.825 ;
        RECT 142.435 207.655 143.405 207.985 ;
        RECT 142.095 207.225 143.065 207.475 ;
        RECT 138.560 206.680 139.925 206.735 ;
        RECT 140.515 206.565 141.085 206.935 ;
        RECT 135.875 206.265 137.165 206.475 ;
        RECT 135.075 206.195 135.705 206.245 ;
        RECT 134.595 205.975 135.705 206.195 ;
        RECT 134.595 205.945 135.245 205.975 ;
        RECT 134.255 205.505 134.880 205.765 ;
        RECT 134.255 204.920 134.425 205.505 ;
        RECT 135.075 205.335 135.245 205.945 ;
        RECT 135.875 205.805 136.045 206.265 ;
        RECT 135.415 205.520 136.045 205.805 ;
        RECT 136.215 205.405 136.775 206.095 ;
        RECT 136.945 205.805 137.165 206.265 ;
        RECT 137.795 206.300 138.425 206.565 ;
        RECT 140.055 206.515 141.085 206.565 ;
        RECT 137.795 206.245 137.965 206.300 ;
        RECT 137.335 205.975 137.965 206.245 ;
        RECT 138.935 206.230 139.885 206.510 ;
        RECT 140.055 206.315 140.685 206.515 ;
        RECT 141.255 206.345 141.425 207.105 ;
        RECT 141.595 206.785 142.725 207.035 ;
        RECT 136.945 205.520 137.625 205.805 ;
        RECT 137.795 205.705 137.965 205.975 ;
        RECT 138.135 205.875 140.255 206.060 ;
        RECT 140.515 206.005 140.685 206.315 ;
        RECT 140.855 206.175 141.425 206.345 ;
        RECT 141.595 206.385 142.725 206.585 ;
        RECT 141.595 206.340 141.925 206.385 ;
        RECT 142.895 206.215 143.065 207.225 ;
        RECT 140.515 205.705 141.425 206.005 ;
        RECT 141.595 205.765 141.875 206.155 ;
        RECT 142.045 206.045 143.065 206.215 ;
        RECT 134.595 205.090 135.245 205.335 ;
        RECT 134.255 204.645 134.880 204.920 ;
        RECT 135.075 204.775 135.245 205.090 ;
        RECT 137.795 205.375 138.465 205.705 ;
        RECT 138.635 205.470 139.965 205.700 ;
        RECT 137.795 204.775 137.965 205.375 ;
        RECT 138.635 205.205 138.805 205.470 ;
        RECT 138.135 205.035 138.805 205.205 ;
        RECT 138.975 204.950 139.625 205.300 ;
        RECT 139.795 205.205 139.965 205.470 ;
        RECT 140.135 205.555 141.425 205.705 ;
        RECT 142.045 205.595 142.215 206.045 ;
        RECT 143.235 205.875 143.405 207.655 ;
        RECT 140.135 205.375 140.685 205.555 ;
        RECT 141.595 205.425 142.215 205.595 ;
        RECT 142.385 205.560 143.405 205.875 ;
        RECT 139.795 205.035 140.255 205.205 ;
        RECT 134.255 204.060 134.425 204.645 ;
        RECT 135.075 204.485 135.970 204.775 ;
        RECT 136.630 204.485 137.965 204.775 ;
        RECT 140.515 204.775 140.685 205.375 ;
        RECT 140.865 205.255 141.425 205.385 ;
        RECT 142.435 205.255 143.065 205.385 ;
        RECT 140.865 204.945 143.065 205.255 ;
        RECT 143.235 204.775 143.405 205.560 ;
        RECT 138.135 204.515 138.805 204.685 ;
        RECT 135.075 204.475 135.245 204.485 ;
        RECT 134.595 204.230 135.245 204.475 ;
        RECT 137.795 204.345 137.965 204.485 ;
        RECT 134.255 203.800 134.880 204.060 ;
        RECT 135.075 203.885 135.245 204.230 ;
        RECT 135.415 204.140 137.625 204.310 ;
        RECT 135.415 204.055 135.985 204.140 ;
        RECT 136.655 203.975 137.625 204.140 ;
        RECT 137.795 204.015 138.465 204.345 ;
        RECT 138.635 204.250 138.805 204.515 ;
        RECT 138.975 204.420 139.625 204.770 ;
        RECT 139.795 204.515 140.255 204.685 ;
        RECT 139.795 204.250 139.965 204.515 ;
        RECT 140.515 204.485 141.410 204.775 ;
        RECT 142.070 204.485 143.405 204.775 ;
        RECT 140.515 204.345 140.685 204.485 ;
        RECT 138.635 204.020 139.965 204.250 ;
        RECT 140.135 204.015 140.685 204.345 ;
        RECT 136.155 203.885 136.485 203.970 ;
        RECT 134.255 203.200 134.425 203.800 ;
        RECT 135.075 203.630 135.645 203.885 ;
        RECT 134.595 203.555 135.645 203.630 ;
        RECT 135.815 203.715 136.485 203.885 ;
        RECT 137.795 203.805 137.965 204.015 ;
        RECT 134.595 203.370 135.245 203.555 ;
        RECT 134.255 202.940 134.880 203.200 ;
        RECT 134.255 202.340 134.425 202.940 ;
        RECT 135.075 202.770 135.245 203.370 ;
        RECT 135.815 203.130 135.985 203.715 ;
        RECT 136.655 203.635 137.965 203.805 ;
        RECT 138.135 203.660 140.255 203.845 ;
        RECT 136.155 203.465 136.485 203.490 ;
        RECT 136.155 203.295 137.625 203.465 ;
        RECT 134.595 202.510 135.245 202.770 ;
        RECT 135.415 203.125 135.985 203.130 ;
        RECT 135.415 202.955 137.285 203.125 ;
        RECT 135.415 202.600 135.780 202.955 ;
        RECT 135.975 202.615 136.945 202.785 ;
        RECT 134.255 202.080 134.880 202.340 ;
        RECT 135.075 201.910 135.245 202.510 ;
        RECT 136.265 202.410 136.435 202.415 ;
        RECT 135.415 202.135 136.575 202.410 ;
        RECT 136.775 201.965 136.945 202.615 ;
        RECT 137.115 202.000 137.285 202.955 ;
        RECT 134.515 201.650 135.245 201.910 ;
        RECT 135.415 201.775 136.945 201.965 ;
        RECT 135.075 201.595 135.245 201.650 ;
        RECT 137.455 201.605 137.625 203.295 ;
        RECT 132.700 201.230 134.895 201.480 ;
        RECT 129.635 200.490 129.805 200.630 ;
        RECT 129.155 200.245 129.805 200.490 ;
        RECT 130.485 200.450 130.785 200.910 ;
        RECT 131.035 200.790 131.295 200.960 ;
        RECT 132.355 200.790 133.335 201.050 ;
        RECT 130.965 200.620 131.295 200.790 ;
        RECT 131.555 200.620 132.525 200.790 ;
        RECT 128.815 199.815 129.440 200.075 ;
        RECT 128.815 199.215 128.985 199.815 ;
        RECT 129.635 199.635 129.805 200.245 ;
        RECT 130.085 200.280 132.185 200.450 ;
        RECT 130.085 200.045 130.255 200.280 ;
        RECT 131.855 200.200 132.185 200.280 ;
        RECT 132.355 200.190 132.525 200.620 ;
        RECT 133.835 200.620 134.085 201.230 ;
        RECT 135.075 201.085 135.780 201.595 ;
        RECT 135.075 201.050 135.245 201.085 ;
        RECT 134.550 200.790 135.245 201.050 ;
        RECT 136.055 200.865 136.225 201.575 ;
        RECT 133.835 200.615 134.895 200.620 ;
        RECT 132.695 200.370 134.895 200.615 ;
        RECT 130.965 199.920 131.685 200.110 ;
        RECT 129.155 199.385 129.805 199.635 ;
        RECT 128.815 198.955 129.440 199.215 ;
        RECT 128.815 198.355 128.985 198.955 ;
        RECT 129.635 198.815 129.805 199.385 ;
        RECT 130.085 199.260 130.255 199.875 ;
        RECT 130.425 199.750 130.755 199.895 ;
        RECT 130.425 199.430 131.715 199.750 ;
        RECT 131.885 199.260 132.055 199.975 ;
        RECT 130.085 199.090 132.055 199.260 ;
        RECT 132.355 199.895 133.335 200.190 ;
        RECT 132.355 199.160 132.525 199.895 ;
        RECT 133.835 199.885 134.395 200.200 ;
        RECT 135.075 200.190 135.245 200.790 ;
        RECT 135.450 200.685 136.225 200.865 ;
        RECT 136.600 201.435 137.625 201.605 ;
        RECT 137.795 203.420 137.965 203.635 ;
        RECT 137.795 203.155 138.425 203.420 ;
        RECT 138.935 203.210 139.885 203.490 ;
        RECT 140.515 203.405 140.685 204.015 ;
        RECT 140.055 203.155 140.685 203.405 ;
        RECT 136.600 200.855 136.790 201.435 ;
        RECT 137.795 201.265 137.965 203.155 ;
        RECT 138.560 202.985 139.925 203.040 ;
        RECT 138.135 202.870 140.235 202.985 ;
        RECT 138.135 202.735 138.690 202.870 ;
        RECT 139.795 202.815 140.235 202.870 ;
        RECT 138.240 201.590 138.410 202.525 ;
        RECT 138.880 202.460 139.475 202.700 ;
        RECT 140.065 202.650 140.235 202.815 ;
        RECT 140.515 202.825 140.685 203.155 ;
        RECT 140.855 202.995 141.485 203.280 ;
        RECT 139.645 202.290 139.865 202.645 ;
        RECT 140.515 202.555 141.145 202.825 ;
        RECT 138.580 202.120 139.865 202.290 ;
        RECT 138.580 201.760 138.945 202.120 ;
        RECT 140.065 201.950 140.235 202.455 ;
        RECT 139.115 201.780 140.235 201.950 ;
        RECT 139.115 201.590 139.285 201.780 ;
        RECT 138.240 201.420 139.285 201.590 ;
        RECT 137.035 201.250 137.965 201.265 ;
        RECT 139.025 201.250 139.285 201.420 ;
        RECT 139.505 201.370 139.835 201.570 ;
        RECT 140.515 201.460 140.685 202.555 ;
        RECT 141.315 202.535 141.485 202.995 ;
        RECT 141.655 202.705 142.215 203.395 ;
        RECT 142.385 202.995 143.065 203.280 ;
        RECT 142.385 202.535 142.605 202.995 ;
        RECT 143.235 202.825 143.405 204.485 ;
        RECT 142.775 202.555 143.405 202.825 ;
        RECT 141.315 202.325 142.605 202.535 ;
        RECT 140.855 201.755 143.065 202.155 ;
        RECT 137.035 201.095 138.765 201.250 ;
        RECT 137.795 201.080 138.765 201.095 ;
        RECT 139.025 201.080 139.355 201.250 ;
        RECT 137.035 200.685 137.445 200.860 ;
        RECT 135.450 200.620 137.445 200.685 ;
        RECT 136.055 200.345 137.445 200.620 ;
        RECT 134.565 199.885 135.245 200.190 ;
        RECT 132.695 199.435 134.905 199.715 ;
        RECT 132.695 199.330 133.665 199.435 ;
        RECT 134.335 199.330 134.905 199.435 ;
        RECT 135.075 199.550 135.245 199.885 ;
        RECT 135.075 199.310 135.755 199.550 ;
        RECT 133.835 199.160 134.165 199.265 ;
        RECT 135.075 199.160 135.245 199.310 ;
        RECT 135.925 199.300 136.485 199.655 ;
        RECT 129.635 198.775 130.335 198.815 ;
        RECT 129.155 198.605 130.335 198.775 ;
        RECT 129.155 198.525 129.805 198.605 ;
        RECT 128.815 198.095 129.440 198.355 ;
        RECT 128.815 197.920 128.985 198.095 ;
        RECT 126.915 197.655 127.815 197.910 ;
        RECT 126.065 197.115 126.745 197.395 ;
        RECT 126.915 197.025 127.085 197.655 ;
        RECT 128.000 197.485 128.985 197.920 ;
        RECT 129.635 197.915 129.805 198.525 ;
        RECT 130.715 198.385 131.045 199.090 ;
        RECT 131.250 198.365 131.625 198.920 ;
        RECT 132.355 198.910 132.985 199.160 ;
        RECT 131.855 198.835 132.985 198.910 ;
        RECT 131.855 198.595 132.525 198.835 ;
        RECT 130.020 198.215 130.545 198.345 ;
        RECT 131.250 198.215 132.185 198.365 ;
        RECT 130.020 198.025 132.185 198.215 ;
        RECT 130.020 198.015 131.045 198.025 ;
        RECT 129.155 197.845 129.805 197.915 ;
        RECT 129.155 197.675 130.415 197.845 ;
        RECT 129.155 197.655 129.805 197.675 ;
        RECT 127.260 197.225 129.440 197.485 ;
        RECT 127.260 197.195 128.985 197.225 ;
        RECT 124.535 196.525 126.745 196.925 ;
        RECT 126.915 196.755 127.830 197.025 ;
        RECT 128.000 196.755 128.985 197.195 ;
        RECT 129.635 197.055 129.805 197.655 ;
        RECT 130.025 197.350 130.545 197.505 ;
        RECT 130.715 197.465 131.045 198.015 ;
        RECT 132.355 197.855 132.525 198.595 ;
        RECT 133.155 198.710 134.445 199.160 ;
        RECT 134.615 198.835 135.245 199.160 ;
        RECT 136.655 199.140 137.000 199.530 ;
        RECT 137.795 199.370 137.965 201.080 ;
        RECT 139.535 200.910 139.835 201.370 ;
        RECT 140.015 201.090 140.685 201.460 ;
        RECT 140.855 201.285 141.485 201.565 ;
        RECT 138.135 200.740 140.235 200.910 ;
        RECT 138.135 200.660 138.465 200.740 ;
        RECT 138.265 199.720 138.435 200.435 ;
        RECT 138.635 200.380 139.355 200.570 ;
        RECT 140.065 200.505 140.235 200.740 ;
        RECT 140.515 200.765 140.685 201.090 ;
        RECT 141.315 200.890 141.485 201.285 ;
        RECT 141.655 201.060 142.215 201.755 ;
        RECT 142.385 201.285 143.065 201.565 ;
        RECT 142.385 200.890 142.605 201.285 ;
        RECT 140.515 200.440 141.145 200.765 ;
        RECT 141.315 200.440 142.605 200.890 ;
        RECT 143.235 200.765 143.405 202.555 ;
        RECT 142.775 200.440 143.405 200.765 ;
        RECT 139.565 200.210 139.895 200.355 ;
        RECT 138.605 199.890 139.895 200.210 ;
        RECT 140.065 199.720 140.235 200.335 ;
        RECT 138.265 199.550 140.235 199.720 ;
        RECT 136.655 199.130 136.825 199.140 ;
        RECT 135.425 198.960 136.825 199.130 ;
        RECT 135.425 198.850 135.755 198.960 ;
        RECT 133.155 198.315 133.375 198.710 ;
        RECT 132.695 198.035 133.375 198.315 ;
        RECT 131.345 197.685 132.525 197.855 ;
        RECT 133.545 197.845 134.105 198.540 ;
        RECT 134.275 198.315 134.445 198.710 ;
        RECT 135.075 198.620 135.245 198.835 ;
        RECT 135.075 198.405 135.755 198.620 ;
        RECT 135.925 198.525 136.485 198.790 ;
        RECT 134.275 198.035 134.905 198.315 ;
        RECT 130.025 197.295 130.585 197.350 ;
        RECT 131.215 197.340 132.140 197.515 ;
        RECT 131.165 197.295 132.140 197.340 ;
        RECT 130.025 197.185 132.140 197.295 ;
        RECT 130.025 197.175 131.295 197.185 ;
        RECT 130.460 197.125 131.295 197.175 ;
        RECT 129.155 196.755 129.805 197.055 ;
        RECT 124.995 196.145 126.285 196.355 ;
        RECT 122.275 195.685 123.565 195.895 ;
        RECT 117.805 194.690 118.135 194.835 ;
        RECT 116.845 194.370 118.135 194.690 ;
        RECT 118.305 194.200 118.475 194.815 ;
        RECT 116.505 194.030 118.475 194.200 ;
        RECT 118.755 194.765 119.420 195.165 ;
        RECT 119.785 195.135 120.315 195.525 ;
        RECT 118.755 194.175 118.925 194.765 ;
        RECT 119.785 194.705 120.165 195.135 ;
        RECT 120.485 194.840 120.795 195.535 ;
        RECT 121.475 195.530 122.105 195.665 ;
        RECT 121.005 195.395 122.105 195.530 ;
        RECT 121.005 194.845 121.645 195.395 ;
        RECT 122.275 195.225 122.495 195.685 ;
        RECT 121.815 194.940 122.495 195.225 ;
        RECT 119.095 194.535 119.615 194.595 ;
        RECT 120.420 194.535 121.205 194.665 ;
        RECT 119.095 194.360 121.205 194.535 ;
        RECT 121.475 194.655 121.645 194.845 ;
        RECT 122.665 194.825 123.225 195.515 ;
        RECT 123.395 195.225 123.565 195.685 ;
        RECT 124.195 195.855 124.825 196.125 ;
        RECT 124.195 195.665 124.365 195.855 ;
        RECT 124.995 195.685 125.165 196.145 ;
        RECT 123.735 195.395 124.365 195.665 ;
        RECT 124.535 195.400 125.165 195.685 ;
        RECT 123.395 194.940 124.025 195.225 ;
        RECT 124.195 195.115 124.365 195.395 ;
        RECT 125.335 195.285 125.895 195.975 ;
        RECT 126.065 195.685 126.285 196.145 ;
        RECT 126.915 196.125 127.085 196.755 ;
        RECT 129.635 196.495 129.805 196.755 ;
        RECT 132.355 197.045 132.525 197.685 ;
        RECT 132.695 197.445 134.905 197.845 ;
        RECT 135.075 197.355 135.245 198.405 ;
        RECT 136.655 198.275 136.825 198.960 ;
        RECT 137.795 199.055 138.465 199.370 ;
        RECT 137.795 198.655 137.965 199.055 ;
        RECT 138.695 198.825 139.070 199.380 ;
        RECT 139.275 198.845 139.605 199.550 ;
        RECT 140.515 199.275 140.685 200.440 ;
        RECT 141.595 200.335 141.925 200.440 ;
        RECT 140.855 200.165 141.425 200.270 ;
        RECT 142.095 200.165 143.065 200.270 ;
        RECT 140.855 199.885 143.065 200.165 ;
        RECT 139.985 199.065 140.685 199.275 ;
        RECT 136.995 198.325 137.965 198.655 ;
        RECT 138.135 198.675 139.070 198.825 ;
        RECT 139.775 198.675 140.300 198.805 ;
        RECT 138.135 198.485 140.300 198.675 ;
        RECT 135.415 197.935 135.985 198.235 ;
        RECT 136.155 198.105 136.825 198.275 ;
        RECT 137.795 198.315 137.965 198.325 ;
        RECT 139.275 198.475 140.300 198.485 ;
        RECT 140.515 198.790 140.685 199.065 ;
        RECT 143.235 198.790 143.405 200.440 ;
        RECT 140.515 198.530 141.525 198.790 ;
        RECT 142.085 198.530 143.405 198.790 ;
        RECT 137.005 197.935 137.625 198.155 ;
        RECT 135.415 197.620 137.625 197.935 ;
        RECT 137.795 198.145 138.975 198.315 ;
        RECT 137.795 197.355 137.965 198.145 ;
        RECT 138.180 197.800 139.105 197.975 ;
        RECT 139.275 197.925 139.605 198.475 ;
        RECT 140.515 198.305 140.685 198.530 ;
        RECT 139.905 198.135 140.685 198.305 ;
        RECT 139.775 197.810 140.295 197.965 ;
        RECT 138.180 197.755 139.155 197.800 ;
        RECT 139.735 197.755 140.295 197.810 ;
        RECT 138.180 197.645 140.295 197.755 ;
        RECT 139.025 197.635 140.295 197.645 ;
        RECT 140.515 197.930 140.685 198.135 ;
        RECT 140.855 198.185 143.065 198.355 ;
        RECT 140.855 198.100 141.430 198.185 ;
        RECT 142.160 198.100 143.065 198.185 ;
        RECT 141.595 197.930 141.925 198.015 ;
        RECT 143.235 197.930 143.405 198.530 ;
        RECT 139.025 197.585 139.860 197.635 ;
        RECT 140.515 197.600 141.065 197.930 ;
        RECT 141.235 197.760 142.305 197.930 ;
        RECT 133.155 197.065 134.445 197.275 ;
        RECT 132.355 196.775 132.985 197.045 ;
        RECT 132.355 196.495 132.525 196.775 ;
        RECT 133.155 196.605 133.375 197.065 ;
        RECT 126.455 195.940 127.085 196.125 ;
        RECT 127.255 196.215 129.465 196.495 ;
        RECT 127.255 196.110 128.225 196.215 ;
        RECT 128.895 196.110 129.465 196.215 ;
        RECT 129.635 196.225 130.440 196.495 ;
        RECT 131.400 196.225 132.525 196.495 ;
        RECT 132.695 196.320 133.375 196.605 ;
        RECT 128.395 195.940 128.725 196.045 ;
        RECT 129.635 195.940 129.805 196.225 ;
        RECT 126.455 195.855 127.545 195.940 ;
        RECT 126.065 195.400 126.745 195.685 ;
        RECT 126.915 195.615 127.545 195.855 ;
        RECT 126.915 195.115 127.085 195.615 ;
        RECT 124.195 194.655 125.655 195.115 ;
        RECT 121.475 194.175 122.735 194.655 ;
        RECT 112.780 193.725 113.485 193.905 ;
        RECT 112.335 193.325 113.110 193.505 ;
        RECT 111.115 193.260 113.110 193.325 ;
        RECT 113.315 193.295 113.485 193.725 ;
        RECT 116.035 193.850 116.205 193.905 ;
        RECT 113.655 193.475 114.205 193.645 ;
        RECT 111.115 192.985 112.505 193.260 ;
        RECT 113.315 192.965 113.865 193.295 ;
        RECT 114.035 193.150 114.205 193.475 ;
        RECT 114.385 193.385 114.755 193.715 ;
        RECT 114.935 193.475 115.865 193.645 ;
        RECT 116.035 193.535 116.705 193.850 ;
        RECT 114.935 193.150 115.105 193.475 ;
        RECT 116.035 193.295 116.205 193.535 ;
        RECT 116.935 193.305 117.310 193.860 ;
        RECT 117.515 193.325 117.845 194.030 ;
        RECT 118.755 193.905 119.560 194.175 ;
        RECT 120.520 193.905 122.735 194.175 ;
        RECT 118.755 193.755 118.925 193.905 ;
        RECT 118.225 193.735 118.925 193.755 ;
        RECT 121.475 193.735 122.735 193.905 ;
        RECT 118.225 193.545 120.215 193.735 ;
        RECT 114.035 192.980 115.105 193.150 ;
        RECT 113.315 191.915 113.485 192.965 ;
        RECT 114.460 192.865 114.790 192.980 ;
        RECT 115.275 192.965 116.205 193.295 ;
        RECT 116.375 193.155 117.310 193.305 ;
        RECT 118.015 193.155 118.540 193.285 ;
        RECT 116.375 192.965 118.540 193.155 ;
        RECT 116.035 192.795 116.205 192.965 ;
        RECT 117.515 192.955 118.540 192.965 ;
        RECT 113.655 192.695 114.160 192.785 ;
        RECT 114.960 192.695 115.865 192.795 ;
        RECT 113.655 192.525 115.865 192.695 ;
        RECT 116.035 192.625 117.215 192.795 ;
        RECT 113.655 192.095 114.205 192.265 ;
        RECT 113.315 191.895 113.865 191.915 ;
        RECT 107.875 191.605 108.770 191.895 ;
        RECT 109.430 191.605 111.930 191.895 ;
        RECT 112.590 191.605 113.865 191.895 ;
        RECT 107.875 190.040 108.045 191.605 ;
        RECT 110.595 190.880 110.765 191.605 ;
        RECT 113.315 191.585 113.865 191.605 ;
        RECT 114.035 191.770 114.205 192.095 ;
        RECT 114.385 192.005 114.755 192.335 ;
        RECT 114.935 192.095 115.865 192.265 ;
        RECT 114.935 191.770 115.105 192.095 ;
        RECT 116.035 191.915 116.205 192.625 ;
        RECT 116.420 192.280 117.345 192.455 ;
        RECT 117.515 192.405 117.845 192.955 ;
        RECT 118.755 192.785 120.215 193.545 ;
        RECT 118.145 192.615 120.215 192.785 ;
        RECT 118.755 192.525 120.215 192.615 ;
        RECT 120.385 193.275 122.735 193.735 ;
        RECT 122.905 194.595 125.655 194.655 ;
        RECT 122.905 193.905 125.115 194.595 ;
        RECT 125.825 194.425 127.085 195.115 ;
        RECT 127.715 195.490 129.005 195.940 ;
        RECT 129.175 195.635 129.805 195.940 ;
        RECT 129.975 195.865 132.085 196.040 ;
        RECT 129.975 195.805 130.495 195.865 ;
        RECT 131.300 195.735 132.085 195.865 ;
        RECT 132.355 196.035 132.525 196.225 ;
        RECT 133.545 196.205 134.105 196.895 ;
        RECT 134.275 196.605 134.445 197.065 ;
        RECT 135.075 197.145 136.065 197.355 ;
        RECT 136.655 197.145 137.965 197.355 ;
        RECT 135.075 197.045 135.245 197.145 ;
        RECT 134.615 196.775 135.245 197.045 ;
        RECT 134.275 196.320 134.905 196.605 ;
        RECT 135.075 196.475 135.245 196.775 ;
        RECT 135.415 196.725 137.625 196.975 ;
        RECT 135.415 196.645 136.045 196.725 ;
        RECT 136.645 196.645 137.625 196.725 ;
        RECT 137.795 196.675 137.965 197.145 ;
        RECT 138.135 197.065 140.345 197.380 ;
        RECT 138.135 196.845 138.755 197.065 ;
        RECT 138.935 196.725 139.605 196.895 ;
        RECT 139.775 196.765 140.345 197.065 ;
        RECT 135.075 196.245 136.065 196.475 ;
        RECT 135.075 196.035 135.245 196.245 ;
        RECT 136.235 196.225 136.485 196.555 ;
        RECT 137.795 196.475 138.765 196.675 ;
        RECT 136.655 196.345 138.765 196.475 ;
        RECT 136.655 196.245 137.965 196.345 ;
        RECT 129.175 195.615 130.300 195.635 ;
        RECT 127.715 195.095 127.935 195.490 ;
        RECT 127.255 194.815 127.935 195.095 ;
        RECT 128.105 194.625 128.665 195.320 ;
        RECT 128.835 195.095 129.005 195.490 ;
        RECT 129.635 195.235 130.300 195.615 ;
        RECT 130.665 195.265 131.045 195.695 ;
        RECT 128.835 194.815 129.465 195.095 ;
        RECT 125.285 193.905 127.085 194.425 ;
        RECT 127.255 194.225 129.465 194.625 ;
        RECT 122.905 193.445 124.365 193.905 ;
        RECT 126.915 193.825 127.085 193.905 ;
        RECT 127.715 193.845 129.005 194.055 ;
        RECT 124.695 193.565 126.745 193.735 ;
        RECT 124.695 193.460 125.040 193.565 ;
        RECT 125.775 193.460 126.745 193.565 ;
        RECT 126.915 193.555 127.545 193.825 ;
        RECT 118.015 192.290 118.535 192.445 ;
        RECT 116.420 192.235 117.395 192.280 ;
        RECT 117.975 192.235 118.535 192.290 ;
        RECT 116.420 192.125 118.535 192.235 ;
        RECT 117.265 192.115 118.535 192.125 ;
        RECT 117.265 192.065 118.100 192.115 ;
        RECT 114.035 191.600 115.105 191.770 ;
        RECT 115.275 191.895 116.205 191.915 ;
        RECT 118.755 191.895 119.695 192.525 ;
        RECT 120.385 192.355 123.255 193.275 ;
        RECT 115.275 191.605 117.370 191.895 ;
        RECT 118.030 191.605 119.695 191.895 ;
        RECT 110.935 191.155 113.145 191.435 ;
        RECT 110.935 191.050 111.905 191.155 ;
        RECT 112.575 191.050 113.145 191.155 ;
        RECT 112.075 190.880 112.405 190.985 ;
        RECT 113.315 190.880 113.485 191.585 ;
        RECT 114.460 191.485 114.790 191.600 ;
        RECT 115.275 191.585 116.205 191.605 ;
        RECT 113.655 191.315 114.160 191.405 ;
        RECT 114.960 191.315 115.865 191.415 ;
        RECT 113.655 191.145 115.865 191.315 ;
        RECT 110.595 190.555 111.225 190.880 ;
        RECT 108.215 190.255 108.765 190.425 ;
        RECT 107.875 189.710 108.425 190.040 ;
        RECT 108.595 189.880 108.765 190.255 ;
        RECT 108.945 190.160 109.315 190.515 ;
        RECT 109.495 190.255 110.425 190.425 ;
        RECT 109.495 189.880 109.665 190.255 ;
        RECT 110.595 190.040 110.765 190.555 ;
        RECT 108.595 189.710 109.665 189.880 ;
        RECT 109.835 189.710 110.765 190.040 ;
        RECT 111.395 190.430 112.685 190.880 ;
        RECT 112.855 190.555 113.485 190.880 ;
        RECT 113.655 190.715 114.205 190.885 ;
        RECT 111.395 190.035 111.615 190.430 ;
        RECT 110.935 189.755 111.615 190.035 ;
        RECT 107.875 189.110 108.045 189.710 ;
        RECT 108.955 189.625 109.285 189.710 ;
        RECT 108.215 189.455 108.790 189.540 ;
        RECT 109.520 189.455 110.425 189.540 ;
        RECT 108.215 189.285 110.425 189.455 ;
        RECT 110.595 189.110 110.765 189.710 ;
        RECT 111.785 189.565 112.345 190.260 ;
        RECT 112.515 190.035 112.685 190.430 ;
        RECT 113.315 190.535 113.485 190.555 ;
        RECT 113.315 190.205 113.865 190.535 ;
        RECT 114.035 190.390 114.205 190.715 ;
        RECT 114.385 190.625 114.755 190.955 ;
        RECT 116.035 190.925 116.205 191.585 ;
        RECT 116.375 191.260 118.585 191.430 ;
        RECT 116.375 191.095 117.345 191.260 ;
        RECT 118.015 191.175 118.585 191.260 ;
        RECT 118.755 191.145 119.695 191.605 ;
        RECT 119.865 192.065 123.255 192.355 ;
        RECT 123.425 193.270 124.365 193.445 ;
        RECT 125.275 193.290 125.605 193.395 ;
        RECT 123.425 192.890 124.765 193.270 ;
        RECT 124.935 193.120 125.945 193.290 ;
        RECT 126.915 193.250 127.085 193.555 ;
        RECT 127.715 193.385 127.935 193.845 ;
        RECT 123.425 192.380 124.365 192.890 ;
        RECT 124.935 192.720 125.105 193.120 ;
        RECT 124.585 192.550 125.105 192.720 ;
        RECT 125.275 192.570 125.605 192.950 ;
        RECT 125.775 192.800 125.945 193.120 ;
        RECT 126.115 192.970 127.085 193.250 ;
        RECT 127.255 193.100 127.935 193.385 ;
        RECT 128.105 192.985 128.665 193.675 ;
        RECT 128.835 193.385 129.005 193.845 ;
        RECT 129.635 193.825 129.805 195.235 ;
        RECT 130.665 194.875 131.195 195.265 ;
        RECT 130.135 194.705 131.195 194.875 ;
        RECT 131.365 194.865 131.675 195.560 ;
        RECT 132.355 195.555 133.615 196.035 ;
        RECT 131.885 195.345 133.615 195.555 ;
        RECT 133.785 195.605 135.245 196.035 ;
        RECT 135.505 195.775 135.965 195.945 ;
        RECT 133.785 195.515 135.625 195.605 ;
        RECT 131.885 194.870 134.155 195.345 ;
        RECT 130.135 194.645 130.330 194.705 ;
        RECT 129.990 194.475 130.330 194.645 ;
        RECT 131.025 194.690 131.195 194.705 ;
        RECT 132.355 194.825 134.155 194.870 ;
        RECT 134.325 195.275 135.625 195.515 ;
        RECT 135.795 195.510 135.965 195.775 ;
        RECT 136.135 195.680 136.785 196.030 ;
        RECT 136.955 195.775 137.625 195.945 ;
        RECT 136.955 195.510 137.125 195.775 ;
        RECT 137.795 195.605 137.965 196.245 ;
        RECT 138.935 196.040 139.105 196.725 ;
        RECT 140.515 196.595 140.685 197.600 ;
        RECT 141.235 197.385 141.405 197.760 ;
        RECT 140.855 197.215 141.405 197.385 ;
        RECT 141.585 197.125 141.955 197.480 ;
        RECT 142.135 197.385 142.305 197.760 ;
        RECT 142.475 197.600 143.405 197.930 ;
        RECT 142.135 197.215 143.065 197.385 ;
        RECT 139.275 196.210 139.835 196.475 ;
        RECT 140.005 196.385 140.685 196.595 ;
        RECT 140.855 196.555 141.485 196.840 ;
        RECT 140.005 196.380 141.145 196.385 ;
        RECT 140.005 196.040 140.335 196.150 ;
        RECT 138.935 195.870 140.335 196.040 ;
        RECT 140.515 196.115 141.145 196.380 ;
        RECT 138.935 195.860 139.105 195.870 ;
        RECT 135.795 195.280 137.125 195.510 ;
        RECT 137.295 195.275 137.965 195.605 ;
        RECT 138.760 195.470 139.105 195.860 ;
        RECT 139.275 195.345 139.835 195.700 ;
        RECT 140.515 195.690 140.685 196.115 ;
        RECT 141.315 196.095 141.485 196.555 ;
        RECT 141.655 196.265 142.215 196.955 ;
        RECT 142.385 196.555 143.065 196.840 ;
        RECT 142.385 196.095 142.605 196.555 ;
        RECT 143.235 196.385 143.405 197.600 ;
        RECT 142.775 196.115 143.405 196.385 ;
        RECT 141.315 195.885 142.605 196.095 ;
        RECT 140.005 195.450 140.685 195.690 ;
        RECT 134.325 194.825 135.245 195.275 ;
        RECT 135.505 194.920 137.625 195.105 ;
        RECT 130.525 194.215 130.855 194.535 ;
        RECT 131.025 194.405 132.140 194.690 ;
        RECT 130.525 194.195 131.735 194.215 ;
        RECT 132.355 194.205 132.525 194.825 ;
        RECT 135.075 194.665 135.245 194.825 ;
        RECT 130.000 193.980 131.735 194.195 ;
        RECT 130.000 193.955 130.375 193.980 ;
        RECT 129.175 193.785 129.805 193.825 ;
        RECT 129.175 193.555 130.310 193.785 ;
        RECT 129.635 193.455 130.310 193.555 ;
        RECT 130.485 193.510 131.335 193.810 ;
        RECT 131.505 193.705 131.735 193.980 ;
        RECT 131.905 193.875 132.525 194.205 ;
        RECT 131.505 193.535 132.165 193.705 ;
        RECT 130.485 193.505 130.655 193.510 ;
        RECT 128.835 193.100 129.465 193.385 ;
        RECT 125.775 192.630 126.235 192.800 ;
        RECT 123.425 192.065 124.765 192.380 ;
        RECT 119.865 191.895 121.645 192.065 ;
        RECT 124.195 192.050 124.765 192.065 ;
        RECT 124.195 191.895 124.365 192.050 ;
        RECT 119.865 191.605 122.810 191.895 ;
        RECT 123.470 191.605 124.365 191.895 ;
        RECT 124.935 191.875 125.105 192.550 ;
        RECT 124.585 191.705 125.105 191.875 ;
        RECT 125.275 191.660 125.895 192.400 ;
        RECT 119.865 191.145 121.645 191.605 ;
        RECT 124.195 191.505 124.365 191.605 ;
        RECT 117.515 191.005 117.845 191.090 ;
        RECT 118.755 191.005 118.925 191.145 ;
        RECT 114.935 190.715 115.865 190.885 ;
        RECT 116.035 190.755 117.345 190.925 ;
        RECT 117.515 190.835 118.185 191.005 ;
        RECT 114.935 190.390 115.105 190.715 ;
        RECT 116.035 190.535 116.205 190.755 ;
        RECT 117.515 190.585 117.845 190.610 ;
        RECT 114.035 190.220 115.105 190.390 ;
        RECT 112.515 189.755 113.145 190.035 ;
        RECT 110.935 189.165 113.145 189.565 ;
        RECT 107.875 188.850 108.885 189.110 ;
        RECT 109.445 188.850 110.765 189.110 ;
        RECT 113.315 189.155 113.485 190.205 ;
        RECT 114.460 190.105 114.790 190.220 ;
        RECT 115.275 190.205 116.205 190.535 ;
        RECT 113.655 189.935 114.160 190.025 ;
        RECT 114.960 189.935 115.865 190.035 ;
        RECT 113.655 189.765 115.865 189.935 ;
        RECT 113.655 189.335 114.205 189.505 ;
        RECT 107.875 188.235 108.045 188.850 ;
        RECT 110.595 188.765 110.765 188.850 ;
        RECT 111.395 188.785 112.685 188.995 ;
        RECT 108.215 188.495 110.425 188.675 ;
        RECT 108.215 188.415 108.720 188.495 ;
        RECT 109.520 188.405 110.425 188.495 ;
        RECT 110.595 188.495 111.225 188.765 ;
        RECT 107.875 187.905 108.425 188.235 ;
        RECT 109.020 188.220 109.350 188.325 ;
        RECT 110.595 188.235 110.765 188.495 ;
        RECT 111.395 188.325 111.615 188.785 ;
        RECT 108.595 188.050 109.665 188.220 ;
        RECT 107.875 186.370 108.045 187.905 ;
        RECT 108.595 187.725 108.765 188.050 ;
        RECT 108.215 187.555 108.765 187.725 ;
        RECT 108.945 187.485 109.315 187.825 ;
        RECT 109.495 187.725 109.665 188.050 ;
        RECT 109.835 187.905 110.765 188.235 ;
        RECT 110.935 188.040 111.615 188.325 ;
        RECT 111.785 187.925 112.345 188.615 ;
        RECT 112.515 188.325 112.685 188.785 ;
        RECT 113.315 188.825 113.865 189.155 ;
        RECT 114.035 189.010 114.205 189.335 ;
        RECT 114.385 189.245 114.755 189.575 ;
        RECT 114.935 189.335 115.865 189.505 ;
        RECT 114.935 189.010 115.105 189.335 ;
        RECT 116.035 189.155 116.205 190.205 ;
        RECT 114.035 188.840 115.105 189.010 ;
        RECT 113.315 188.765 113.485 188.825 ;
        RECT 112.855 188.495 113.485 188.765 ;
        RECT 114.460 188.725 114.790 188.840 ;
        RECT 115.275 188.825 116.205 189.155 ;
        RECT 112.515 188.040 113.145 188.325 ;
        RECT 113.315 188.205 113.485 188.495 ;
        RECT 113.655 188.555 114.160 188.645 ;
        RECT 114.960 188.555 115.865 188.655 ;
        RECT 113.655 188.385 115.865 188.555 ;
        RECT 116.035 188.385 116.205 188.825 ;
        RECT 116.375 190.415 117.845 190.585 ;
        RECT 116.375 188.725 116.545 190.415 ;
        RECT 118.015 190.250 118.185 190.835 ;
        RECT 118.355 190.675 118.925 191.005 ;
        RECT 118.015 190.245 118.585 190.250 ;
        RECT 116.715 190.075 118.585 190.245 ;
        RECT 116.715 189.120 116.885 190.075 ;
        RECT 117.055 189.735 118.025 189.905 ;
        RECT 117.055 189.085 117.225 189.735 ;
        RECT 118.220 189.720 118.585 190.075 ;
        RECT 118.755 189.945 118.925 190.675 ;
        RECT 119.095 190.115 119.725 190.400 ;
        RECT 118.755 189.675 119.385 189.945 ;
        RECT 118.245 189.530 118.415 189.535 ;
        RECT 117.425 189.255 118.585 189.530 ;
        RECT 117.055 188.895 118.585 189.085 ;
        RECT 116.375 188.555 117.400 188.725 ;
        RECT 118.755 188.715 118.925 189.675 ;
        RECT 119.555 189.655 119.725 190.115 ;
        RECT 119.895 189.825 120.455 190.515 ;
        RECT 120.625 190.115 121.305 190.400 ;
        RECT 121.475 190.145 121.645 191.145 ;
        RECT 122.285 191.135 123.625 191.260 ;
        RECT 121.855 191.090 123.625 191.135 ;
        RECT 124.195 191.175 124.865 191.505 ;
        RECT 126.065 191.490 126.235 192.630 ;
        RECT 124.195 191.105 124.365 191.175 ;
        RECT 121.855 190.805 122.455 191.090 ;
        RECT 122.625 190.675 123.285 190.920 ;
        RECT 121.865 190.375 122.455 190.625 ;
        RECT 123.455 190.605 123.625 191.090 ;
        RECT 123.795 190.775 124.365 191.105 ;
        RECT 125.275 190.980 125.605 191.390 ;
        RECT 125.775 191.170 126.235 191.490 ;
        RECT 120.625 189.655 120.845 190.115 ;
        RECT 121.475 189.945 122.115 190.145 ;
        RECT 121.015 189.815 122.115 189.945 ;
        RECT 121.015 189.675 121.645 189.815 ;
        RECT 119.555 189.445 120.845 189.655 ;
        RECT 119.095 188.875 121.305 189.275 ;
        RECT 121.475 189.145 121.645 189.675 ;
        RECT 122.285 189.585 122.455 190.375 ;
        RECT 122.625 190.195 123.285 190.460 ;
        RECT 123.455 190.275 123.965 190.605 ;
        RECT 124.195 190.565 124.365 190.775 ;
        RECT 124.585 190.975 125.605 190.980 ;
        RECT 124.585 190.735 126.200 190.975 ;
        RECT 126.405 190.750 126.695 192.800 ;
        RECT 126.915 191.895 127.085 192.970 ;
        RECT 129.635 191.895 129.805 193.455 ;
        RECT 132.355 192.825 132.525 193.875 ;
        RECT 132.745 192.995 133.035 194.650 ;
        RECT 133.205 194.330 133.665 194.650 ;
        RECT 133.205 193.230 133.375 194.330 ;
        RECT 133.835 194.300 134.405 194.650 ;
        RECT 135.075 194.645 135.705 194.665 ;
        RECT 134.575 194.415 135.705 194.645 ;
        RECT 135.875 194.470 136.825 194.750 ;
        RECT 137.795 194.680 137.965 195.275 ;
        RECT 138.135 194.855 139.065 195.025 ;
        RECT 137.335 194.640 137.965 194.680 ;
        RECT 137.335 194.415 138.725 194.640 ;
        RECT 134.575 194.315 135.245 194.415 ;
        RECT 133.545 193.420 134.165 194.130 ;
        RECT 134.335 193.945 134.855 194.115 ;
        RECT 133.205 193.060 133.665 193.230 ;
        RECT 132.355 192.545 133.325 192.825 ;
        RECT 133.495 192.675 133.665 193.060 ;
        RECT 133.835 192.845 134.165 193.250 ;
        RECT 134.335 193.245 134.505 193.945 ;
        RECT 135.075 193.745 135.245 194.315 ;
        RECT 137.795 194.310 138.725 194.415 ;
        RECT 138.895 194.480 139.065 194.855 ;
        RECT 139.245 194.760 139.615 195.115 ;
        RECT 139.795 194.855 140.345 195.025 ;
        RECT 139.795 194.480 139.965 194.855 ;
        RECT 140.515 194.640 140.685 195.450 ;
        RECT 140.855 195.315 143.065 195.715 ;
        RECT 140.855 194.845 141.485 195.125 ;
        RECT 138.895 194.310 139.965 194.480 ;
        RECT 140.135 194.325 140.685 194.640 ;
        RECT 141.315 194.450 141.485 194.845 ;
        RECT 141.655 194.620 142.215 195.315 ;
        RECT 142.385 194.845 143.065 195.125 ;
        RECT 142.385 194.450 142.605 194.845 ;
        RECT 140.135 194.310 141.145 194.325 ;
        RECT 135.835 194.245 137.200 194.300 ;
        RECT 135.525 194.130 137.625 194.245 ;
        RECT 135.525 194.075 135.965 194.130 ;
        RECT 135.525 193.910 135.695 194.075 ;
        RECT 137.070 193.995 137.625 194.130 ;
        RECT 134.675 193.415 135.245 193.745 ;
        RECT 134.335 193.075 134.855 193.245 ;
        RECT 134.335 192.675 134.505 193.075 ;
        RECT 135.075 192.905 135.245 193.415 ;
        RECT 135.525 193.210 135.695 193.715 ;
        RECT 135.895 193.550 136.115 193.905 ;
        RECT 136.285 193.720 136.880 193.960 ;
        RECT 135.895 193.380 137.180 193.550 ;
        RECT 135.525 193.040 136.645 193.210 ;
        RECT 129.985 192.045 132.185 192.355 ;
        RECT 129.985 191.915 130.545 192.045 ;
        RECT 131.555 191.915 132.185 192.045 ;
        RECT 126.915 191.605 128.250 191.895 ;
        RECT 128.910 191.745 129.805 191.895 ;
        RECT 132.355 191.895 132.525 192.545 ;
        RECT 133.495 192.505 134.505 192.675 ;
        RECT 134.675 192.720 135.245 192.905 ;
        RECT 136.475 192.850 136.645 193.040 ;
        RECT 136.815 193.020 137.180 193.380 ;
        RECT 137.350 192.850 137.520 193.785 ;
        RECT 134.675 192.525 135.745 192.720 ;
        RECT 133.835 192.405 134.165 192.505 ;
        RECT 135.075 192.350 135.745 192.525 ;
        RECT 135.925 192.630 136.255 192.830 ;
        RECT 136.475 192.680 137.520 192.850 ;
        RECT 137.795 193.710 137.965 194.310 ;
        RECT 139.275 194.225 139.605 194.310 ;
        RECT 138.135 194.055 139.040 194.140 ;
        RECT 139.770 194.055 140.345 194.140 ;
        RECT 138.135 193.885 140.345 194.055 ;
        RECT 140.515 194.000 141.145 194.310 ;
        RECT 141.315 194.000 142.605 194.450 ;
        RECT 143.235 194.325 143.405 196.115 ;
        RECT 142.775 194.000 143.405 194.325 ;
        RECT 140.515 193.710 140.685 194.000 ;
        RECT 141.595 193.895 141.925 194.000 ;
        RECT 137.795 193.450 139.115 193.710 ;
        RECT 139.675 193.450 140.685 193.710 ;
        RECT 137.795 193.235 137.965 193.450 ;
        RECT 137.795 193.005 139.105 193.235 ;
        RECT 132.695 192.235 133.665 192.335 ;
        RECT 134.400 192.235 134.745 192.335 ;
        RECT 132.695 192.065 134.745 192.235 ;
        RECT 135.075 191.895 135.245 192.350 ;
        RECT 135.925 192.170 136.225 192.630 ;
        RECT 136.475 192.510 136.735 192.680 ;
        RECT 137.795 192.510 137.965 193.005 ;
        RECT 139.275 192.925 139.525 193.255 ;
        RECT 140.515 193.235 140.685 193.450 ;
        RECT 140.855 193.725 141.425 193.830 ;
        RECT 142.095 193.725 143.065 193.830 ;
        RECT 140.855 193.445 143.065 193.725 ;
        RECT 139.695 193.005 140.685 193.235 ;
        RECT 140.855 193.015 141.405 193.185 ;
        RECT 140.515 192.835 140.685 193.005 ;
        RECT 136.405 192.340 136.735 192.510 ;
        RECT 136.995 192.340 137.965 192.510 ;
        RECT 138.135 192.755 139.115 192.835 ;
        RECT 139.715 192.755 140.345 192.835 ;
        RECT 138.135 192.505 140.345 192.755 ;
        RECT 140.515 192.505 141.065 192.835 ;
        RECT 141.235 192.690 141.405 193.015 ;
        RECT 141.585 192.915 141.955 193.255 ;
        RECT 142.135 193.015 143.065 193.195 ;
        RECT 142.135 192.690 142.305 193.015 ;
        RECT 143.235 192.835 143.405 194.000 ;
        RECT 141.235 192.520 142.305 192.690 ;
        RECT 137.795 192.335 137.965 192.340 ;
        RECT 140.515 192.335 140.685 192.505 ;
        RECT 141.660 192.415 141.990 192.520 ;
        RECT 142.475 192.505 143.405 192.835 ;
        RECT 128.910 191.605 130.545 191.745 ;
        RECT 130.715 191.705 131.335 191.875 ;
        RECT 132.355 191.740 133.690 191.895 ;
        RECT 126.915 190.565 127.085 191.605 ;
        RECT 122.625 189.715 123.285 190.000 ;
        RECT 121.865 189.335 122.455 189.585 ;
        RECT 122.625 189.325 123.285 189.540 ;
        RECT 122.955 189.235 123.285 189.325 ;
        RECT 121.475 188.895 122.785 189.145 ;
        RECT 123.455 189.065 123.625 190.275 ;
        RECT 124.195 190.225 124.865 190.565 ;
        RECT 125.035 190.225 125.605 190.565 ;
        RECT 125.840 190.225 127.085 190.565 ;
        RECT 127.305 190.245 127.595 191.435 ;
        RECT 127.765 191.090 128.225 191.415 ;
        RECT 128.395 191.090 128.725 191.435 ;
        RECT 128.895 191.165 129.415 191.420 ;
        RECT 129.635 191.295 130.545 191.605 ;
        RECT 127.765 190.415 127.935 191.090 ;
        RECT 128.105 190.725 128.725 190.920 ;
        RECT 127.765 190.245 128.225 190.415 ;
        RECT 124.195 190.035 124.365 190.225 ;
        RECT 126.915 190.075 127.085 190.225 ;
        RECT 124.195 189.795 125.175 190.035 ;
        RECT 124.195 189.225 124.365 189.795 ;
        RECT 125.355 189.705 125.605 190.055 ;
        RECT 125.775 189.715 126.730 190.045 ;
        RECT 126.915 189.795 127.885 190.075 ;
        RECT 128.055 189.925 128.225 190.245 ;
        RECT 128.395 190.095 128.725 190.725 ;
        RECT 128.895 190.495 129.065 191.165 ;
        RECT 129.635 190.995 129.805 191.295 ;
        RECT 130.715 191.145 130.995 191.535 ;
        RECT 131.165 191.255 131.335 191.705 ;
        RECT 131.505 191.605 133.690 191.740 ;
        RECT 134.350 191.605 135.245 191.895 ;
        RECT 135.525 192.000 137.625 192.170 ;
        RECT 135.525 191.765 135.695 192.000 ;
        RECT 137.295 191.920 137.625 192.000 ;
        RECT 137.795 192.125 139.105 192.335 ;
        RECT 139.695 192.125 140.685 192.335 ;
        RECT 137.795 191.895 137.965 192.125 ;
        RECT 140.515 191.895 140.685 192.125 ;
        RECT 140.855 192.245 141.360 192.325 ;
        RECT 142.160 192.245 143.065 192.335 ;
        RECT 140.855 192.065 143.065 192.245 ;
        RECT 143.235 191.895 143.405 192.505 ;
        RECT 136.405 191.640 137.125 191.830 ;
        RECT 131.505 191.425 132.525 191.605 ;
        RECT 129.235 190.785 129.805 190.995 ;
        RECT 129.975 190.955 130.545 191.125 ;
        RECT 131.165 191.085 132.185 191.255 ;
        RECT 129.235 190.665 130.205 190.785 ;
        RECT 128.895 190.325 129.415 190.495 ;
        RECT 129.635 190.365 130.205 190.665 ;
        RECT 128.895 189.925 129.065 190.325 ;
        RECT 129.635 190.155 129.805 190.365 ;
        RECT 130.375 190.195 130.545 190.955 ;
        RECT 130.715 190.915 131.045 190.960 ;
        RECT 130.715 190.715 131.845 190.915 ;
        RECT 130.715 190.265 131.845 190.515 ;
        RECT 124.535 189.535 125.175 189.625 ;
        RECT 125.775 189.535 125.945 189.715 ;
        RECT 124.535 189.365 125.945 189.535 ;
        RECT 124.535 189.295 125.175 189.365 ;
        RECT 122.955 188.895 123.625 189.065 ;
        RECT 123.795 189.125 124.365 189.225 ;
        RECT 123.795 188.895 125.175 189.125 ;
        RECT 116.035 188.215 116.965 188.385 ;
        RECT 113.315 187.935 114.295 188.205 ;
        RECT 109.495 187.545 110.425 187.725 ;
        RECT 110.595 186.825 110.765 187.905 ;
        RECT 113.315 187.265 113.485 187.935 ;
        RECT 114.475 187.865 114.725 188.215 ;
        RECT 116.035 188.205 116.205 188.215 ;
        RECT 114.895 187.875 116.205 188.205 ;
        RECT 113.655 187.695 114.295 187.765 ;
        RECT 113.655 187.525 115.065 187.695 ;
        RECT 113.655 187.435 114.295 187.525 ;
        RECT 113.315 187.025 114.295 187.265 ;
        RECT 110.595 186.495 111.485 186.825 ;
        RECT 111.785 186.605 112.325 186.835 ;
        RECT 112.125 186.505 112.325 186.605 ;
        RECT 112.495 186.495 113.145 186.835 ;
        RECT 107.875 186.035 108.550 186.370 ;
        RECT 107.875 184.610 108.045 186.035 ;
        RECT 108.725 186.015 109.575 186.315 ;
        RECT 109.745 186.115 110.405 186.285 ;
        RECT 108.240 185.845 108.615 185.865 ;
        RECT 109.745 185.845 109.975 186.115 ;
        RECT 110.595 185.945 110.765 186.495 ;
        RECT 111.010 186.195 112.305 186.315 ;
        RECT 111.010 186.100 112.325 186.195 ;
        RECT 108.240 185.625 109.975 185.845 ;
        RECT 108.765 185.610 109.975 185.625 ;
        RECT 110.145 185.615 110.765 185.945 ;
        RECT 108.230 185.175 108.570 185.345 ;
        RECT 108.765 185.310 109.095 185.610 ;
        RECT 108.375 185.140 108.570 185.175 ;
        RECT 109.265 185.155 110.380 185.440 ;
        RECT 110.595 185.405 110.765 185.615 ;
        RECT 110.935 185.575 111.925 185.905 ;
        RECT 112.125 185.865 112.325 186.100 ;
        RECT 112.495 185.985 112.685 186.495 ;
        RECT 113.315 186.325 113.485 187.025 ;
        RECT 114.475 187.005 114.725 187.355 ;
        RECT 114.895 187.345 115.065 187.525 ;
        RECT 114.895 187.015 115.850 187.345 ;
        RECT 116.035 186.855 116.205 187.875 ;
        RECT 116.555 187.805 116.965 187.980 ;
        RECT 117.210 187.975 117.400 188.555 ;
        RECT 117.775 187.985 117.945 188.695 ;
        RECT 118.220 188.205 118.925 188.715 ;
        RECT 119.095 188.405 119.725 188.685 ;
        RECT 117.775 187.805 118.550 187.985 ;
        RECT 116.555 187.740 118.550 187.805 ;
        RECT 118.755 187.885 118.925 188.205 ;
        RECT 119.555 188.010 119.725 188.405 ;
        RECT 119.895 188.180 120.455 188.875 ;
        RECT 120.625 188.405 121.305 188.685 ;
        RECT 120.625 188.010 120.845 188.405 ;
        RECT 116.555 187.465 117.945 187.740 ;
        RECT 118.755 187.560 119.385 187.885 ;
        RECT 119.555 187.560 120.845 188.010 ;
        RECT 121.475 187.885 121.645 188.895 ;
        RECT 122.955 188.755 123.285 188.895 ;
        RECT 124.195 188.855 125.175 188.895 ;
        RECT 121.855 188.585 122.705 188.725 ;
        RECT 123.470 188.585 123.980 188.725 ;
        RECT 121.855 188.395 123.980 188.585 ;
        RECT 121.015 187.560 121.645 187.885 ;
        RECT 116.375 187.035 117.305 187.205 ;
        RECT 113.850 186.580 115.865 186.835 ;
        RECT 113.850 186.475 114.225 186.580 ;
        RECT 114.880 186.495 115.865 186.580 ;
        RECT 116.035 186.525 116.965 186.855 ;
        RECT 117.135 186.710 117.305 187.035 ;
        RECT 117.485 186.945 117.855 187.275 ;
        RECT 118.035 187.035 118.585 187.205 ;
        RECT 118.035 186.710 118.205 187.035 ;
        RECT 118.755 186.855 118.925 187.560 ;
        RECT 119.835 187.455 120.165 187.560 ;
        RECT 119.095 187.285 119.665 187.390 ;
        RECT 120.335 187.285 121.305 187.390 ;
        RECT 119.095 187.005 121.305 187.285 ;
        RECT 121.475 187.080 121.645 187.560 ;
        RECT 124.195 188.235 124.365 188.855 ;
        RECT 125.355 188.845 125.605 189.195 ;
        RECT 126.915 189.185 127.085 189.795 ;
        RECT 128.055 189.755 129.065 189.925 ;
        RECT 129.235 189.775 129.805 190.155 ;
        RECT 129.975 189.965 130.545 190.195 ;
        RECT 132.015 190.075 132.185 191.085 ;
        RECT 128.395 189.650 128.725 189.755 ;
        RECT 127.255 189.480 128.225 189.585 ;
        RECT 128.960 189.480 129.305 189.585 ;
        RECT 127.255 189.310 129.305 189.480 ;
        RECT 125.775 189.135 127.085 189.185 ;
        RECT 129.635 189.135 129.805 189.775 ;
        RECT 129.975 189.475 130.545 189.795 ;
        RECT 130.715 189.645 131.045 190.050 ;
        RECT 131.215 189.825 132.185 190.075 ;
        RECT 132.355 190.925 132.525 191.425 ;
        RECT 132.695 191.180 134.710 191.435 ;
        RECT 132.695 191.095 133.680 191.180 ;
        RECT 134.335 191.075 134.710 191.180 ;
        RECT 133.835 190.925 134.165 191.010 ;
        RECT 132.355 190.515 132.955 190.925 ;
        RECT 133.125 190.660 134.165 190.925 ;
        RECT 135.075 190.810 135.245 191.605 ;
        RECT 135.525 190.980 135.695 191.595 ;
        RECT 135.865 191.470 136.195 191.615 ;
        RECT 135.865 191.150 137.155 191.470 ;
        RECT 137.325 190.980 137.495 191.695 ;
        RECT 135.525 190.810 137.495 190.980 ;
        RECT 137.795 191.605 139.130 191.895 ;
        RECT 139.790 191.605 141.410 191.895 ;
        RECT 142.070 191.605 143.405 191.895 ;
        RECT 137.795 190.820 137.965 191.605 ;
        RECT 138.135 191.125 140.335 191.435 ;
        RECT 138.135 190.995 138.765 191.125 ;
        RECT 139.775 190.995 140.335 191.125 ;
        RECT 131.215 189.475 131.385 189.825 ;
        RECT 132.355 189.770 132.525 190.515 ;
        RECT 132.355 189.645 132.945 189.770 ;
        RECT 129.975 189.305 131.385 189.475 ;
        RECT 131.555 189.440 132.945 189.645 ;
        RECT 133.125 189.650 133.295 190.660 ;
        RECT 134.335 190.640 135.245 190.810 ;
        RECT 135.075 190.535 135.245 190.640 ;
        RECT 133.465 189.990 133.635 190.445 ;
        RECT 133.835 190.160 134.165 190.490 ;
        RECT 134.335 190.190 134.710 190.360 ;
        RECT 135.075 190.325 135.775 190.535 ;
        RECT 134.335 189.990 134.505 190.190 ;
        RECT 133.465 189.820 134.505 189.990 ;
        RECT 133.125 189.480 134.905 189.650 ;
        RECT 135.075 189.565 135.245 190.325 ;
        RECT 136.155 190.105 136.485 190.810 ;
        RECT 136.690 190.085 137.065 190.640 ;
        RECT 137.795 190.630 138.815 190.820 ;
        RECT 137.295 190.505 138.815 190.630 ;
        RECT 138.985 190.785 139.605 190.955 ;
        RECT 140.515 190.825 140.685 191.605 ;
        RECT 137.295 190.315 137.965 190.505 ;
        RECT 138.985 190.335 139.155 190.785 ;
        RECT 135.460 189.935 135.985 190.065 ;
        RECT 136.690 189.935 137.625 190.085 ;
        RECT 135.460 189.745 137.625 189.935 ;
        RECT 135.460 189.735 136.485 189.745 ;
        RECT 131.555 189.315 132.525 189.440 ;
        RECT 125.775 188.855 128.175 189.135 ;
        RECT 124.535 188.415 125.085 188.585 ;
        RECT 124.195 187.905 124.745 188.235 ;
        RECT 124.915 188.090 125.085 188.415 ;
        RECT 125.265 188.315 125.635 188.655 ;
        RECT 125.815 188.415 126.745 188.595 ;
        RECT 125.815 188.090 125.985 188.415 ;
        RECT 126.915 188.235 128.175 188.855 ;
        RECT 124.915 187.920 125.985 188.090 ;
        RECT 117.135 186.540 118.205 186.710 ;
        RECT 112.855 186.210 113.485 186.325 ;
        RECT 114.395 186.325 114.725 186.410 ;
        RECT 116.035 186.325 116.205 186.525 ;
        RECT 117.450 186.425 117.780 186.540 ;
        RECT 118.375 186.525 118.925 186.855 ;
        RECT 112.855 186.155 114.225 186.210 ;
        RECT 113.315 186.040 114.225 186.155 ;
        RECT 114.395 186.060 115.435 186.325 ;
        RECT 109.265 185.140 109.435 185.155 ;
        RECT 108.375 184.970 109.435 185.140 ;
        RECT 107.875 184.215 108.540 184.610 ;
        RECT 108.905 184.580 109.435 184.970 ;
        RECT 107.875 183.155 108.045 184.215 ;
        RECT 108.905 184.155 109.285 184.580 ;
        RECT 109.605 184.285 109.915 184.980 ;
        RECT 110.595 184.975 111.540 185.405 ;
        RECT 110.125 184.695 111.540 184.975 ;
        RECT 111.710 185.040 111.925 185.575 ;
        RECT 112.095 185.225 112.325 185.695 ;
        RECT 112.495 185.655 112.765 185.985 ;
        RECT 112.880 185.520 113.145 185.525 ;
        RECT 112.875 185.515 113.145 185.520 ;
        RECT 112.865 185.510 113.145 185.515 ;
        RECT 112.860 185.505 113.145 185.510 ;
        RECT 112.850 185.500 113.145 185.505 ;
        RECT 112.845 185.490 113.145 185.500 ;
        RECT 112.835 185.480 113.145 185.490 ;
        RECT 112.825 185.465 113.145 185.480 ;
        RECT 112.495 185.165 113.145 185.465 ;
        RECT 112.495 185.040 112.685 185.165 ;
        RECT 111.710 184.755 112.685 185.040 ;
        RECT 113.315 184.925 113.485 186.040 ;
        RECT 113.850 185.590 114.225 185.760 ;
        RECT 114.055 185.390 114.225 185.590 ;
        RECT 114.395 185.560 114.725 185.890 ;
        RECT 114.925 185.390 115.095 185.845 ;
        RECT 114.055 185.220 115.095 185.390 ;
        RECT 115.265 185.050 115.435 186.060 ;
        RECT 115.605 185.915 116.205 186.325 ;
        RECT 116.375 186.255 117.280 186.355 ;
        RECT 118.080 186.255 118.585 186.345 ;
        RECT 116.375 186.085 118.585 186.255 ;
        RECT 118.755 186.225 118.925 186.525 ;
        RECT 119.105 186.525 121.305 186.835 ;
        RECT 119.105 186.395 119.665 186.525 ;
        RECT 120.675 186.395 121.305 186.525 ;
        RECT 121.475 186.750 122.745 187.080 ;
        RECT 116.035 185.435 116.205 185.915 ;
        RECT 116.375 185.745 118.425 185.915 ;
        RECT 116.375 185.645 117.345 185.745 ;
        RECT 118.080 185.645 118.425 185.745 ;
        RECT 118.755 185.775 119.665 186.225 ;
        RECT 119.835 186.185 120.455 186.355 ;
        RECT 121.475 186.220 121.645 186.750 ;
        RECT 122.995 186.650 123.205 187.295 ;
        RECT 123.375 186.810 124.010 187.140 ;
        RECT 117.515 185.475 117.845 185.575 ;
        RECT 116.035 185.170 117.005 185.435 ;
        RECT 112.855 184.755 113.485 184.925 ;
        RECT 113.655 184.880 115.435 185.050 ;
        RECT 110.125 184.290 110.765 184.695 ;
        RECT 112.370 184.525 113.145 184.585 ;
        RECT 108.215 183.980 108.735 184.045 ;
        RECT 109.540 183.980 110.325 184.110 ;
        RECT 108.215 183.805 110.325 183.980 ;
        RECT 110.595 183.155 110.765 184.290 ;
        RECT 110.935 184.245 113.145 184.525 ;
        RECT 113.315 184.150 113.485 184.755 ;
        RECT 113.655 184.320 114.305 184.650 ;
        RECT 113.315 183.980 113.955 184.150 ;
        RECT 113.315 183.155 113.485 183.980 ;
        RECT 114.135 183.810 114.305 184.320 ;
        RECT 114.475 184.140 114.685 184.710 ;
        RECT 114.855 184.670 115.435 184.880 ;
        RECT 115.615 185.155 117.005 185.170 ;
        RECT 117.175 185.305 118.185 185.475 ;
        RECT 118.755 185.455 118.925 185.775 ;
        RECT 119.835 185.625 120.115 186.015 ;
        RECT 120.285 185.735 120.455 186.185 ;
        RECT 120.625 185.905 121.645 186.220 ;
        RECT 121.815 185.950 122.825 186.275 ;
        RECT 121.475 185.780 121.645 185.905 ;
        RECT 115.615 184.840 116.205 185.155 ;
        RECT 114.855 184.345 115.865 184.670 ;
        RECT 113.670 183.480 114.305 183.810 ;
        RECT 114.475 183.325 114.685 183.970 ;
        RECT 116.035 183.870 116.205 184.840 ;
        RECT 114.935 183.540 116.205 183.870 ;
        RECT 116.035 183.155 116.205 183.540 ;
        RECT 116.425 183.330 116.715 184.985 ;
        RECT 117.175 184.920 117.345 185.305 ;
        RECT 116.885 184.750 117.345 184.920 ;
        RECT 116.885 183.650 117.055 184.750 ;
        RECT 117.515 184.730 117.845 185.135 ;
        RECT 118.015 184.905 118.185 185.305 ;
        RECT 118.355 185.265 118.925 185.455 ;
        RECT 119.095 185.435 119.665 185.605 ;
        RECT 120.285 185.565 121.305 185.735 ;
        RECT 118.355 185.075 119.325 185.265 ;
        RECT 118.015 184.735 118.535 184.905 ;
        RECT 118.755 184.845 119.325 185.075 ;
        RECT 117.225 183.850 117.845 184.560 ;
        RECT 118.015 184.035 118.185 184.735 ;
        RECT 118.755 184.565 118.925 184.845 ;
        RECT 119.495 184.675 119.665 185.435 ;
        RECT 119.835 185.395 120.165 185.440 ;
        RECT 119.835 185.195 120.965 185.395 ;
        RECT 119.835 184.745 120.965 184.995 ;
        RECT 118.355 184.235 118.925 184.565 ;
        RECT 119.095 184.445 119.665 184.675 ;
        RECT 121.135 184.555 121.305 185.565 ;
        RECT 118.015 183.865 118.535 184.035 ;
        RECT 116.885 183.330 117.345 183.650 ;
        RECT 117.515 183.330 118.085 183.680 ;
        RECT 118.755 183.665 118.925 184.235 ;
        RECT 119.095 183.955 119.665 184.275 ;
        RECT 119.835 184.125 120.165 184.530 ;
        RECT 120.335 184.305 121.305 184.555 ;
        RECT 121.475 185.450 122.065 185.780 ;
        RECT 122.245 185.740 122.825 185.950 ;
        RECT 122.995 185.910 123.205 186.480 ;
        RECT 123.375 186.300 123.545 186.810 ;
        RECT 124.195 186.640 124.365 187.905 ;
        RECT 125.340 187.815 125.670 187.920 ;
        RECT 126.155 187.905 128.175 188.235 ;
        RECT 128.345 189.115 129.805 189.135 ;
        RECT 128.345 188.875 130.615 189.115 ;
        RECT 128.345 188.205 129.805 188.875 ;
        RECT 130.795 188.785 131.045 189.135 ;
        RECT 131.215 188.795 132.170 189.125 ;
        RECT 129.975 188.615 130.615 188.705 ;
        RECT 131.215 188.615 131.385 188.795 ;
        RECT 129.975 188.445 131.385 188.615 ;
        RECT 132.355 188.470 132.525 189.315 ;
        RECT 133.125 189.270 133.705 189.480 ;
        RECT 135.075 189.395 135.855 189.565 ;
        RECT 132.695 188.945 133.705 189.270 ;
        RECT 133.875 188.740 134.085 189.310 ;
        RECT 134.255 188.920 134.905 189.250 ;
        RECT 129.975 188.375 130.615 188.445 ;
        RECT 128.345 187.935 130.615 188.205 ;
        RECT 128.345 187.925 129.805 187.935 ;
        RECT 130.795 187.925 131.045 188.275 ;
        RECT 132.355 188.265 133.625 188.470 ;
        RECT 131.215 188.140 133.625 188.265 ;
        RECT 131.215 187.935 132.525 188.140 ;
        RECT 126.915 187.755 128.175 187.905 ;
        RECT 124.535 187.645 125.040 187.725 ;
        RECT 125.840 187.645 126.745 187.735 ;
        RECT 124.535 187.465 126.745 187.645 ;
        RECT 124.550 186.810 125.185 187.140 ;
        RECT 123.725 186.470 124.835 186.640 ;
        RECT 123.375 185.970 124.025 186.300 ;
        RECT 122.245 185.570 124.025 185.740 ;
        RECT 121.475 184.705 121.645 185.450 ;
        RECT 120.335 183.955 120.505 184.305 ;
        RECT 121.475 184.295 122.075 184.705 ;
        RECT 122.245 184.560 122.415 185.570 ;
        RECT 122.585 185.230 123.625 185.400 ;
        RECT 122.585 184.775 122.755 185.230 ;
        RECT 122.955 184.730 123.285 185.060 ;
        RECT 123.455 185.030 123.625 185.230 ;
        RECT 123.455 184.860 123.830 185.030 ;
        RECT 124.195 184.580 124.365 186.470 ;
        RECT 125.015 186.300 125.185 186.810 ;
        RECT 125.355 186.650 125.565 187.295 ;
        RECT 126.915 187.080 128.695 187.755 ;
        RECT 125.815 186.750 128.695 187.080 ;
        RECT 126.915 186.545 128.695 186.750 ;
        RECT 128.865 186.670 129.805 187.925 ;
        RECT 130.170 187.040 132.185 187.295 ;
        RECT 130.170 186.935 130.545 187.040 ;
        RECT 131.200 186.955 132.185 187.040 ;
        RECT 132.355 187.245 132.525 187.935 ;
        RECT 133.875 187.925 134.085 188.570 ;
        RECT 134.255 188.410 134.425 188.920 ;
        RECT 135.075 188.750 135.245 189.395 ;
        RECT 135.465 189.070 135.985 189.225 ;
        RECT 136.155 189.185 136.485 189.735 ;
        RECT 137.795 189.575 137.965 190.315 ;
        RECT 136.785 189.405 137.965 189.575 ;
        RECT 135.465 189.015 136.025 189.070 ;
        RECT 136.655 189.060 137.580 189.235 ;
        RECT 136.605 189.015 137.580 189.060 ;
        RECT 135.465 188.905 137.580 189.015 ;
        RECT 135.465 188.895 136.735 188.905 ;
        RECT 135.900 188.845 136.735 188.895 ;
        RECT 134.605 188.580 135.245 188.750 ;
        RECT 134.255 188.080 134.890 188.410 ;
        RECT 135.075 188.050 135.245 188.580 ;
        RECT 137.795 188.725 137.965 189.405 ;
        RECT 138.135 190.165 139.155 190.335 ;
        RECT 139.325 190.225 139.605 190.615 ;
        RECT 139.775 190.510 140.685 190.825 ;
        RECT 143.235 190.510 143.405 191.605 ;
        RECT 139.775 190.375 141.525 190.510 ;
        RECT 140.515 190.250 141.525 190.375 ;
        RECT 142.085 190.250 143.405 190.510 ;
        RECT 138.135 189.155 138.305 190.165 ;
        RECT 139.275 189.995 139.605 190.040 ;
        RECT 138.475 189.795 139.605 189.995 ;
        RECT 139.775 190.035 140.345 190.205 ;
        RECT 138.475 189.345 139.605 189.595 ;
        RECT 139.775 189.275 139.945 190.035 ;
        RECT 140.515 189.865 140.685 190.250 ;
        RECT 140.115 189.650 140.685 189.865 ;
        RECT 140.855 189.905 143.065 190.075 ;
        RECT 140.855 189.820 141.430 189.905 ;
        RECT 142.160 189.820 143.065 189.905 ;
        RECT 141.595 189.650 141.925 189.735 ;
        RECT 143.235 189.650 143.405 190.250 ;
        RECT 140.115 189.445 141.065 189.650 ;
        RECT 140.515 189.320 141.065 189.445 ;
        RECT 141.235 189.480 142.305 189.650 ;
        RECT 138.135 188.905 139.105 189.155 ;
        RECT 137.795 188.395 138.765 188.725 ;
        RECT 138.935 188.555 139.105 188.905 ;
        RECT 139.275 188.725 139.605 189.130 ;
        RECT 139.775 189.045 140.345 189.275 ;
        RECT 139.775 188.555 140.345 188.875 ;
        RECT 135.075 187.810 135.755 188.050 ;
        RECT 132.695 187.500 134.710 187.755 ;
        RECT 132.695 187.415 133.680 187.500 ;
        RECT 134.335 187.395 134.710 187.500 ;
        RECT 133.835 187.245 134.165 187.330 ;
        RECT 130.715 186.785 131.045 186.870 ;
        RECT 132.355 186.835 132.955 187.245 ;
        RECT 133.125 186.980 134.165 187.245 ;
        RECT 135.075 187.130 135.245 187.810 ;
        RECT 135.925 187.800 136.485 188.155 ;
        RECT 136.655 187.640 137.000 188.030 ;
        RECT 137.795 187.645 137.965 188.395 ;
        RECT 138.935 188.385 140.345 188.555 ;
        RECT 140.515 188.675 140.685 189.320 ;
        RECT 141.235 189.105 141.405 189.480 ;
        RECT 140.855 188.935 141.405 189.105 ;
        RECT 141.585 188.845 141.955 189.200 ;
        RECT 142.135 189.105 142.305 189.480 ;
        RECT 142.475 189.320 143.405 189.650 ;
        RECT 142.135 188.935 143.065 189.105 ;
        RECT 143.235 188.675 143.405 189.320 ;
        RECT 138.135 187.815 138.815 188.100 ;
        RECT 136.655 187.630 136.825 187.640 ;
        RECT 135.425 187.460 136.825 187.630 ;
        RECT 135.425 187.350 135.755 187.460 ;
        RECT 134.335 187.120 135.245 187.130 ;
        RECT 132.355 186.785 132.525 186.835 ;
        RECT 128.865 186.545 130.545 186.670 ;
        RECT 124.535 185.970 125.185 186.300 ;
        RECT 125.355 185.910 125.565 186.480 ;
        RECT 125.735 185.950 126.745 186.275 ;
        RECT 125.735 185.740 126.315 185.950 ;
        RECT 126.915 185.905 127.085 186.545 ;
        RECT 129.635 186.500 130.545 186.545 ;
        RECT 130.715 186.520 131.755 186.785 ;
        RECT 126.915 185.780 128.225 185.905 ;
        RECT 124.535 185.570 126.315 185.740 ;
        RECT 124.935 185.230 125.975 185.400 ;
        RECT 124.935 185.030 125.105 185.230 ;
        RECT 124.730 184.860 125.105 185.030 ;
        RECT 125.275 184.730 125.605 185.060 ;
        RECT 125.805 184.775 125.975 185.230 ;
        RECT 122.245 184.295 123.285 184.560 ;
        RECT 123.455 184.410 125.105 184.580 ;
        RECT 126.145 184.560 126.315 185.570 ;
        RECT 126.495 185.575 128.225 185.780 ;
        RECT 126.495 185.450 127.085 185.575 ;
        RECT 128.395 185.565 128.645 185.915 ;
        RECT 129.635 185.905 129.805 186.500 ;
        RECT 130.170 186.050 130.545 186.220 ;
        RECT 128.825 185.635 129.805 185.905 ;
        RECT 130.375 185.850 130.545 186.050 ;
        RECT 130.715 186.020 131.045 186.350 ;
        RECT 131.245 185.850 131.415 186.305 ;
        RECT 130.375 185.680 131.415 185.850 ;
        RECT 126.915 184.705 127.085 185.450 ;
        RECT 128.825 185.395 129.465 185.465 ;
        RECT 128.055 185.225 129.465 185.395 ;
        RECT 128.055 185.045 128.225 185.225 ;
        RECT 128.825 185.135 129.465 185.225 ;
        RECT 127.270 184.715 128.225 185.045 ;
        RECT 128.395 184.705 128.645 185.055 ;
        RECT 129.635 184.965 129.805 185.635 ;
        RECT 131.585 185.510 131.755 186.520 ;
        RECT 131.925 186.375 132.525 186.785 ;
        RECT 132.355 186.090 132.525 186.375 ;
        RECT 132.355 185.760 132.945 186.090 ;
        RECT 133.125 185.970 133.295 186.980 ;
        RECT 134.335 186.960 135.755 187.120 ;
        RECT 135.925 187.025 136.485 187.290 ;
        RECT 135.075 186.905 135.755 186.960 ;
        RECT 133.465 186.310 133.635 186.765 ;
        RECT 133.835 186.480 134.165 186.810 ;
        RECT 134.335 186.510 134.710 186.680 ;
        RECT 134.335 186.310 134.505 186.510 ;
        RECT 133.465 186.140 134.505 186.310 ;
        RECT 133.125 185.800 134.905 185.970 ;
        RECT 132.355 185.630 132.525 185.760 ;
        RECT 129.975 185.340 131.755 185.510 ;
        RECT 128.825 184.725 129.805 184.965 ;
        RECT 129.975 184.780 130.625 185.110 ;
        RECT 121.475 184.125 121.645 184.295 ;
        RECT 122.955 184.210 123.285 184.295 ;
        RECT 119.095 183.785 120.505 183.955 ;
        RECT 120.675 183.795 121.645 184.125 ;
        RECT 118.255 183.335 118.925 183.665 ;
        RECT 118.755 183.155 118.925 183.335 ;
        RECT 121.475 183.155 121.645 183.795 ;
        RECT 121.815 184.040 122.800 184.125 ;
        RECT 123.455 184.040 123.830 184.145 ;
        RECT 121.815 184.015 123.830 184.040 ;
        RECT 121.815 183.845 123.855 184.015 ;
        RECT 121.815 183.785 123.830 183.845 ;
        RECT 124.195 183.155 124.365 184.410 ;
        RECT 125.275 184.295 126.315 184.560 ;
        RECT 126.485 184.295 127.085 184.705 ;
        RECT 129.635 184.610 129.805 184.725 ;
        RECT 125.275 184.210 125.605 184.295 ;
        RECT 124.730 184.040 125.105 184.145 ;
        RECT 125.760 184.040 126.745 184.125 ;
        RECT 124.730 183.785 126.745 184.040 ;
        RECT 126.915 184.095 127.085 184.295 ;
        RECT 127.255 184.365 129.465 184.535 ;
        RECT 127.255 184.265 128.160 184.365 ;
        RECT 128.960 184.275 129.465 184.365 ;
        RECT 129.635 184.440 130.275 184.610 ;
        RECT 126.915 183.765 127.845 184.095 ;
        RECT 128.330 184.080 128.660 184.195 ;
        RECT 129.635 184.095 129.805 184.440 ;
        RECT 130.455 184.270 130.625 184.780 ;
        RECT 130.795 184.600 131.005 185.170 ;
        RECT 131.175 185.130 131.755 185.340 ;
        RECT 131.935 185.300 132.525 185.630 ;
        RECT 133.125 185.590 133.705 185.800 ;
        RECT 131.175 184.805 132.185 185.130 ;
        RECT 132.355 184.790 132.525 185.300 ;
        RECT 132.695 185.265 133.705 185.590 ;
        RECT 133.875 185.060 134.085 185.630 ;
        RECT 134.255 185.240 134.905 185.570 ;
        RECT 135.075 185.475 135.245 186.905 ;
        RECT 136.655 186.775 136.825 187.460 ;
        RECT 137.795 187.375 138.425 187.645 ;
        RECT 137.795 187.155 137.965 187.375 ;
        RECT 136.995 186.825 137.965 187.155 ;
        RECT 138.595 187.355 138.815 187.815 ;
        RECT 138.985 187.525 139.545 188.215 ;
        RECT 140.515 188.155 141.975 188.675 ;
        RECT 139.715 187.815 140.345 188.100 ;
        RECT 139.715 187.355 139.885 187.815 ;
        RECT 140.515 187.645 141.435 188.155 ;
        RECT 142.145 187.985 143.405 188.675 ;
        RECT 140.055 187.465 141.435 187.645 ;
        RECT 141.605 187.465 143.405 187.985 ;
        RECT 140.055 187.375 140.685 187.465 ;
        RECT 138.595 187.145 139.885 187.355 ;
        RECT 135.415 186.435 135.985 186.735 ;
        RECT 136.155 186.605 136.825 186.775 ;
        RECT 137.005 186.435 137.625 186.655 ;
        RECT 135.415 186.120 137.625 186.435 ;
        RECT 135.415 185.655 135.965 185.825 ;
        RECT 132.355 184.460 133.625 184.790 ;
        RECT 128.015 183.910 129.085 184.080 ;
        RECT 126.915 183.155 127.085 183.765 ;
        RECT 128.015 183.585 128.185 183.910 ;
        RECT 127.255 183.415 128.185 183.585 ;
        RECT 128.365 183.345 128.735 183.675 ;
        RECT 128.915 183.585 129.085 183.910 ;
        RECT 129.255 183.765 129.805 184.095 ;
        RECT 129.990 183.940 130.625 184.270 ;
        RECT 130.795 183.785 131.005 184.430 ;
        RECT 132.355 184.330 132.525 184.460 ;
        RECT 131.255 184.000 132.525 184.330 ;
        RECT 133.875 184.245 134.085 184.890 ;
        RECT 134.255 184.730 134.425 185.240 ;
        RECT 135.075 185.145 135.625 185.475 ;
        RECT 135.795 185.330 135.965 185.655 ;
        RECT 136.145 185.565 136.515 185.895 ;
        RECT 136.695 185.655 137.625 185.825 ;
        RECT 136.695 185.330 136.865 185.655 ;
        RECT 137.795 185.585 137.965 186.825 ;
        RECT 138.135 186.575 140.345 186.975 ;
        RECT 140.515 186.855 140.685 187.375 ;
        RECT 140.855 187.125 143.065 187.295 ;
        RECT 140.855 187.035 141.360 187.125 ;
        RECT 142.160 187.025 143.065 187.125 ;
        RECT 138.135 186.105 138.815 186.385 ;
        RECT 138.595 185.710 138.815 186.105 ;
        RECT 138.985 185.880 139.545 186.575 ;
        RECT 140.515 186.525 141.065 186.855 ;
        RECT 141.660 186.840 141.990 186.955 ;
        RECT 143.235 186.855 143.405 187.465 ;
        RECT 141.235 186.670 142.305 186.840 ;
        RECT 139.715 186.105 140.345 186.385 ;
        RECT 139.715 185.710 139.885 186.105 ;
        RECT 137.795 185.475 138.425 185.585 ;
        RECT 135.795 185.160 136.865 185.330 ;
        RECT 137.035 185.260 138.425 185.475 ;
        RECT 138.595 185.260 139.885 185.710 ;
        RECT 140.515 185.585 140.685 186.525 ;
        RECT 141.235 186.345 141.405 186.670 ;
        RECT 140.855 186.175 141.405 186.345 ;
        RECT 141.585 186.105 141.955 186.435 ;
        RECT 142.135 186.345 142.305 186.670 ;
        RECT 142.475 186.525 143.405 186.855 ;
        RECT 142.135 186.175 143.065 186.345 ;
        RECT 140.855 185.745 143.065 185.915 ;
        RECT 140.855 185.655 141.360 185.745 ;
        RECT 142.160 185.645 143.065 185.745 ;
        RECT 140.055 185.475 140.685 185.585 ;
        RECT 140.055 185.260 141.065 185.475 ;
        RECT 141.660 185.460 141.990 185.575 ;
        RECT 143.235 185.475 143.405 186.525 ;
        RECT 135.075 185.070 135.245 185.145 ;
        RECT 134.605 184.900 135.245 185.070 ;
        RECT 136.220 185.045 136.550 185.160 ;
        RECT 137.035 185.145 137.965 185.260 ;
        RECT 139.275 185.155 139.605 185.260 ;
        RECT 134.255 184.400 134.890 184.730 ;
        RECT 128.915 183.415 129.465 183.585 ;
        RECT 129.635 183.155 129.805 183.765 ;
        RECT 132.355 183.155 132.525 184.000 ;
        RECT 135.075 184.095 135.245 184.900 ;
        RECT 135.415 184.875 135.920 184.965 ;
        RECT 136.720 184.875 137.625 184.975 ;
        RECT 135.415 184.705 137.625 184.875 ;
        RECT 135.415 184.355 137.625 184.535 ;
        RECT 135.415 184.275 135.920 184.355 ;
        RECT 136.720 184.265 137.625 184.355 ;
        RECT 135.075 183.765 135.625 184.095 ;
        RECT 136.220 184.080 136.550 184.185 ;
        RECT 137.795 184.095 137.965 185.145 ;
        RECT 140.515 185.145 141.065 185.260 ;
        RECT 141.235 185.290 142.305 185.460 ;
        RECT 138.135 184.985 139.105 185.090 ;
        RECT 139.775 184.985 140.345 185.090 ;
        RECT 138.135 184.705 140.345 184.985 ;
        RECT 138.135 184.355 140.345 184.535 ;
        RECT 138.135 184.265 139.040 184.355 ;
        RECT 139.840 184.275 140.345 184.355 ;
        RECT 135.795 183.910 136.865 184.080 ;
        RECT 135.075 183.155 135.245 183.765 ;
        RECT 135.795 183.585 135.965 183.910 ;
        RECT 135.415 183.415 135.965 183.585 ;
        RECT 136.145 183.345 136.515 183.685 ;
        RECT 136.695 183.585 136.865 183.910 ;
        RECT 137.035 183.765 138.725 184.095 ;
        RECT 139.210 184.080 139.540 184.185 ;
        RECT 140.515 184.095 140.685 185.145 ;
        RECT 141.235 184.965 141.405 185.290 ;
        RECT 140.855 184.795 141.405 184.965 ;
        RECT 141.585 184.725 141.955 185.055 ;
        RECT 142.135 184.965 142.305 185.290 ;
        RECT 142.475 185.145 143.405 185.475 ;
        RECT 142.135 184.795 143.065 184.965 ;
        RECT 140.855 184.355 143.065 184.535 ;
        RECT 140.855 184.275 141.360 184.355 ;
        RECT 142.160 184.265 143.065 184.355 ;
        RECT 138.895 183.910 139.965 184.080 ;
        RECT 136.695 183.405 137.625 183.585 ;
        RECT 137.795 183.155 137.965 183.765 ;
        RECT 138.895 183.585 139.065 183.910 ;
        RECT 138.135 183.405 139.065 183.585 ;
        RECT 139.245 183.345 139.615 183.685 ;
        RECT 139.795 183.585 139.965 183.910 ;
        RECT 140.135 183.765 141.065 184.095 ;
        RECT 141.660 184.080 141.990 184.185 ;
        RECT 143.235 184.095 143.405 185.145 ;
        RECT 141.235 183.910 142.305 184.080 ;
        RECT 139.795 183.415 140.345 183.585 ;
        RECT 140.515 183.155 140.685 183.765 ;
        RECT 141.235 183.585 141.405 183.910 ;
        RECT 140.855 183.415 141.405 183.585 ;
        RECT 141.585 183.345 141.955 183.685 ;
        RECT 142.135 183.585 142.305 183.910 ;
        RECT 142.475 183.765 143.405 184.095 ;
        RECT 142.135 183.405 143.065 183.585 ;
        RECT 143.235 183.155 143.405 183.765 ;
        RECT 107.875 182.465 108.795 183.155 ;
        RECT 108.965 182.635 112.395 183.155 ;
        RECT 107.875 181.945 109.335 182.465 ;
        RECT 109.505 181.945 111.855 182.635 ;
        RECT 112.565 182.465 114.235 183.155 ;
        RECT 114.405 182.635 117.835 183.155 ;
        RECT 112.025 181.945 114.775 182.465 ;
        RECT 114.945 181.945 117.295 182.635 ;
        RECT 118.005 182.465 119.675 183.155 ;
        RECT 119.845 182.635 123.275 183.155 ;
        RECT 117.465 181.945 120.215 182.465 ;
        RECT 120.385 181.945 122.735 182.635 ;
        RECT 123.445 182.465 125.115 183.155 ;
        RECT 125.285 182.635 128.715 183.155 ;
        RECT 122.905 181.945 125.655 182.465 ;
        RECT 125.825 181.945 128.175 182.635 ;
        RECT 128.885 182.465 130.555 183.155 ;
        RECT 130.725 182.635 134.155 183.155 ;
        RECT 128.345 181.945 131.095 182.465 ;
        RECT 131.265 181.945 133.615 182.635 ;
        RECT 134.325 182.465 135.995 183.155 ;
        RECT 136.165 182.635 139.595 183.155 ;
        RECT 133.785 181.945 136.535 182.465 ;
        RECT 136.705 181.945 139.055 182.635 ;
        RECT 139.765 182.465 141.435 183.155 ;
        RECT 141.605 182.635 143.405 183.155 ;
        RECT 139.225 181.945 141.975 182.465 ;
        RECT 142.145 181.945 143.405 182.635 ;
        RECT 107.875 181.860 108.045 181.945 ;
        RECT 110.595 181.860 110.765 181.945 ;
        RECT 113.315 181.860 113.485 181.945 ;
        RECT 116.035 181.860 116.205 181.945 ;
        RECT 118.755 181.860 118.925 181.945 ;
        RECT 121.475 181.860 121.645 181.945 ;
        RECT 124.195 181.860 124.365 181.945 ;
        RECT 126.915 181.860 127.085 181.945 ;
        RECT 129.635 181.860 129.805 181.945 ;
        RECT 132.355 181.860 132.525 181.945 ;
        RECT 135.075 181.860 135.245 181.945 ;
        RECT 137.795 181.860 137.965 181.945 ;
        RECT 140.515 181.860 140.685 181.945 ;
        RECT 143.235 181.860 143.405 181.945 ;
        RECT 136.420 173.100 142.160 173.110 ;
        RECT 117.470 173.060 123.210 173.070 ;
        RECT 98.430 173.030 104.170 173.040 ;
        RECT 97.940 172.870 104.170 173.030 ;
        RECT 97.940 170.610 98.610 172.870 ;
        RECT 99.280 172.300 103.320 172.470 ;
        RECT 98.940 171.240 99.110 172.240 ;
        RECT 103.490 171.240 103.660 172.240 ;
        RECT 99.280 171.010 103.320 171.180 ;
        RECT 104.000 170.610 104.170 172.870 ;
        RECT 97.940 170.440 104.170 170.610 ;
        RECT 97.940 167.180 98.610 170.440 ;
        RECT 99.280 169.870 103.320 170.040 ;
        RECT 98.940 167.810 99.110 169.810 ;
        RECT 103.490 167.810 103.660 169.810 ;
        RECT 99.280 167.580 103.320 167.750 ;
        RECT 104.000 167.180 104.170 170.440 ;
        RECT 97.940 167.010 104.170 167.180 ;
        RECT 97.940 163.750 98.610 167.010 ;
        RECT 99.280 166.440 103.320 166.610 ;
        RECT 98.940 164.380 99.110 166.380 ;
        RECT 103.490 164.380 103.660 166.380 ;
        RECT 99.280 164.150 103.320 164.320 ;
        RECT 104.000 163.750 104.170 167.010 ;
        RECT 97.940 163.740 104.170 163.750 ;
        RECT 105.760 173.010 115.590 173.050 ;
        RECT 105.760 172.880 116.390 173.010 ;
        RECT 105.760 170.620 105.930 172.880 ;
        RECT 106.655 172.310 114.695 172.480 ;
        RECT 106.270 171.250 106.440 172.250 ;
        RECT 114.910 171.250 115.080 172.250 ;
        RECT 106.655 171.020 114.695 171.190 ;
        RECT 115.420 170.620 116.390 172.880 ;
        RECT 105.760 170.450 116.390 170.620 ;
        RECT 105.760 167.190 105.930 170.450 ;
        RECT 106.655 169.880 114.695 170.050 ;
        RECT 106.270 167.820 106.440 169.820 ;
        RECT 114.910 167.820 115.080 169.820 ;
        RECT 106.655 167.590 114.695 167.760 ;
        RECT 115.420 167.190 116.390 170.450 ;
        RECT 105.760 167.020 116.390 167.190 ;
        RECT 105.760 163.760 105.930 167.020 ;
        RECT 106.655 166.450 114.695 166.620 ;
        RECT 106.270 164.390 106.440 166.390 ;
        RECT 114.910 164.390 115.080 166.390 ;
        RECT 106.655 164.160 114.695 164.330 ;
        RECT 115.420 163.760 116.390 167.020 ;
        RECT 97.940 163.640 104.180 163.740 ;
        RECT 97.930 163.080 104.180 163.640 ;
        RECT 97.930 163.060 103.100 163.080 ;
        RECT 97.930 162.990 101.920 163.060 ;
        RECT 97.930 161.720 99.850 162.990 ;
        RECT 101.360 162.980 101.920 162.990 ;
        RECT 101.590 161.890 101.920 162.980 ;
        RECT 102.290 162.510 103.330 162.680 ;
        RECT 102.290 162.070 103.330 162.240 ;
        RECT 103.500 162.210 103.670 162.540 ;
        RECT 101.750 161.670 101.920 161.890 ;
        RECT 104.010 161.670 104.180 163.080 ;
        RECT 101.750 161.500 104.180 161.670 ;
        RECT 105.760 163.590 116.390 163.760 ;
        RECT 116.980 172.900 123.210 173.060 ;
        RECT 116.980 170.640 117.650 172.900 ;
        RECT 118.320 172.330 122.360 172.500 ;
        RECT 117.980 171.270 118.150 172.270 ;
        RECT 122.530 171.270 122.700 172.270 ;
        RECT 118.320 171.040 122.360 171.210 ;
        RECT 123.040 170.640 123.210 172.900 ;
        RECT 116.980 170.470 123.210 170.640 ;
        RECT 116.980 167.210 117.650 170.470 ;
        RECT 118.320 169.900 122.360 170.070 ;
        RECT 117.980 167.840 118.150 169.840 ;
        RECT 122.530 167.840 122.700 169.840 ;
        RECT 118.320 167.610 122.360 167.780 ;
        RECT 123.040 167.210 123.210 170.470 ;
        RECT 116.980 167.040 123.210 167.210 ;
        RECT 116.980 163.780 117.650 167.040 ;
        RECT 118.320 166.470 122.360 166.640 ;
        RECT 117.980 164.410 118.150 166.410 ;
        RECT 122.530 164.410 122.700 166.410 ;
        RECT 118.320 164.180 122.360 164.350 ;
        RECT 123.040 163.780 123.210 167.040 ;
        RECT 116.980 163.770 123.210 163.780 ;
        RECT 124.800 173.040 134.630 173.080 ;
        RECT 124.800 172.910 135.430 173.040 ;
        RECT 124.800 170.650 124.970 172.910 ;
        RECT 125.695 172.340 133.735 172.510 ;
        RECT 125.310 171.280 125.480 172.280 ;
        RECT 133.950 171.280 134.120 172.280 ;
        RECT 125.695 171.050 133.735 171.220 ;
        RECT 134.460 170.650 135.430 172.910 ;
        RECT 124.800 170.480 135.430 170.650 ;
        RECT 124.800 167.220 124.970 170.480 ;
        RECT 125.695 169.910 133.735 170.080 ;
        RECT 125.310 167.850 125.480 169.850 ;
        RECT 133.950 167.850 134.120 169.850 ;
        RECT 125.695 167.620 133.735 167.790 ;
        RECT 134.460 167.220 135.430 170.480 ;
        RECT 124.800 167.050 135.430 167.220 ;
        RECT 124.800 163.790 124.970 167.050 ;
        RECT 125.695 166.480 133.735 166.650 ;
        RECT 125.310 164.420 125.480 166.420 ;
        RECT 133.950 164.420 134.120 166.420 ;
        RECT 125.695 164.190 133.735 164.360 ;
        RECT 134.460 163.790 135.430 167.050 ;
        RECT 116.980 163.670 123.220 163.770 ;
        RECT 105.760 161.330 105.930 163.590 ;
        RECT 106.655 163.020 114.695 163.190 ;
        RECT 106.270 161.960 106.440 162.960 ;
        RECT 114.910 161.960 115.080 162.960 ;
        RECT 106.655 161.730 114.695 161.900 ;
        RECT 115.420 161.330 116.390 163.590 ;
        RECT 116.970 163.110 123.220 163.670 ;
        RECT 116.970 163.090 122.140 163.110 ;
        RECT 116.970 163.020 120.960 163.090 ;
        RECT 116.970 161.750 118.890 163.020 ;
        RECT 120.400 163.010 120.960 163.020 ;
        RECT 120.630 161.920 120.960 163.010 ;
        RECT 121.330 162.540 122.370 162.710 ;
        RECT 121.330 162.100 122.370 162.270 ;
        RECT 122.540 162.240 122.710 162.570 ;
        RECT 120.790 161.700 120.960 161.920 ;
        RECT 123.050 161.700 123.220 163.110 ;
        RECT 120.790 161.530 123.220 161.700 ;
        RECT 124.800 163.620 135.430 163.790 ;
        RECT 135.930 172.940 142.160 173.100 ;
        RECT 135.930 170.680 136.600 172.940 ;
        RECT 137.270 172.370 141.310 172.540 ;
        RECT 136.930 171.310 137.100 172.310 ;
        RECT 141.480 171.310 141.650 172.310 ;
        RECT 137.270 171.080 141.310 171.250 ;
        RECT 141.990 170.680 142.160 172.940 ;
        RECT 135.930 170.510 142.160 170.680 ;
        RECT 135.930 167.250 136.600 170.510 ;
        RECT 137.270 169.940 141.310 170.110 ;
        RECT 136.930 167.880 137.100 169.880 ;
        RECT 141.480 167.880 141.650 169.880 ;
        RECT 137.270 167.650 141.310 167.820 ;
        RECT 141.990 167.250 142.160 170.510 ;
        RECT 135.930 167.080 142.160 167.250 ;
        RECT 135.930 163.820 136.600 167.080 ;
        RECT 137.270 166.510 141.310 166.680 ;
        RECT 136.930 164.450 137.100 166.450 ;
        RECT 141.480 164.450 141.650 166.450 ;
        RECT 137.270 164.220 141.310 164.390 ;
        RECT 141.990 163.820 142.160 167.080 ;
        RECT 135.930 163.810 142.160 163.820 ;
        RECT 143.750 173.080 153.580 173.120 ;
        RECT 143.750 172.950 154.380 173.080 ;
        RECT 143.750 170.690 143.920 172.950 ;
        RECT 144.645 172.380 152.685 172.550 ;
        RECT 144.260 171.320 144.430 172.320 ;
        RECT 152.900 171.320 153.070 172.320 ;
        RECT 144.645 171.090 152.685 171.260 ;
        RECT 153.410 170.690 154.380 172.950 ;
        RECT 143.750 170.520 154.380 170.690 ;
        RECT 143.750 167.260 143.920 170.520 ;
        RECT 144.645 169.950 152.685 170.120 ;
        RECT 144.260 167.890 144.430 169.890 ;
        RECT 152.900 167.890 153.070 169.890 ;
        RECT 144.645 167.660 152.685 167.830 ;
        RECT 153.410 167.260 154.380 170.520 ;
        RECT 143.750 167.090 154.380 167.260 ;
        RECT 143.750 163.830 143.920 167.090 ;
        RECT 144.645 166.520 152.685 166.690 ;
        RECT 144.260 164.460 144.430 166.460 ;
        RECT 152.900 164.460 153.070 166.460 ;
        RECT 144.645 164.230 152.685 164.400 ;
        RECT 153.410 163.830 154.380 167.090 ;
        RECT 135.930 163.710 142.170 163.810 ;
        RECT 124.800 161.360 124.970 163.620 ;
        RECT 125.695 163.050 133.735 163.220 ;
        RECT 125.310 161.990 125.480 162.990 ;
        RECT 133.950 161.990 134.120 162.990 ;
        RECT 125.695 161.760 133.735 161.930 ;
        RECT 134.460 161.360 135.430 163.620 ;
        RECT 135.920 163.150 142.170 163.710 ;
        RECT 135.920 163.130 141.090 163.150 ;
        RECT 135.920 163.060 139.910 163.130 ;
        RECT 135.920 161.790 137.840 163.060 ;
        RECT 139.350 163.050 139.910 163.060 ;
        RECT 139.580 161.960 139.910 163.050 ;
        RECT 140.280 162.580 141.320 162.750 ;
        RECT 140.280 162.140 141.320 162.310 ;
        RECT 141.490 162.280 141.660 162.610 ;
        RECT 139.740 161.740 139.910 161.960 ;
        RECT 142.000 161.740 142.170 163.150 ;
        RECT 139.740 161.570 142.170 161.740 ;
        RECT 143.750 163.660 154.380 163.830 ;
        RECT 143.750 161.400 143.920 163.660 ;
        RECT 144.645 163.090 152.685 163.260 ;
        RECT 144.260 162.030 144.430 163.030 ;
        RECT 152.900 162.030 153.070 163.030 ;
        RECT 144.645 161.800 152.685 161.970 ;
        RECT 153.410 161.400 154.380 163.660 ;
        RECT 143.750 161.370 154.380 161.400 ;
        RECT 124.800 161.330 135.430 161.360 ;
        RECT 105.760 161.300 116.390 161.330 ;
        RECT 105.730 161.190 116.390 161.300 ;
        RECT 124.770 161.220 135.430 161.330 ;
        RECT 143.720 161.260 154.380 161.370 ;
        RECT 103.980 161.140 116.390 161.190 ;
        RECT 123.020 161.170 135.430 161.220 ;
        RECT 141.970 161.210 154.380 161.260 ;
        RECT 99.640 160.970 116.390 161.140 ;
        RECT 99.640 159.560 99.810 160.970 ;
        RECT 100.180 160.400 103.220 160.570 ;
        RECT 100.180 159.960 103.220 160.130 ;
        RECT 103.435 160.100 103.605 160.430 ;
        RECT 103.940 160.210 116.390 160.970 ;
        RECT 118.680 161.000 135.430 161.170 ;
        RECT 103.940 160.200 116.280 160.210 ;
        RECT 103.940 160.190 109.820 160.200 ;
        RECT 103.940 160.170 104.510 160.190 ;
        RECT 105.730 160.180 109.820 160.190 ;
        RECT 103.950 159.560 104.120 160.170 ;
        RECT 99.640 159.390 104.120 159.560 ;
        RECT 118.680 159.590 118.850 161.000 ;
        RECT 119.220 160.430 122.260 160.600 ;
        RECT 119.220 159.990 122.260 160.160 ;
        RECT 122.475 160.130 122.645 160.460 ;
        RECT 122.980 160.240 135.430 161.000 ;
        RECT 137.630 161.040 154.380 161.210 ;
        RECT 122.980 160.230 135.320 160.240 ;
        RECT 122.980 160.220 128.860 160.230 ;
        RECT 122.980 160.200 123.550 160.220 ;
        RECT 124.770 160.210 128.860 160.220 ;
        RECT 122.990 159.590 123.160 160.200 ;
        RECT 118.680 159.420 123.160 159.590 ;
        RECT 137.630 159.630 137.800 161.040 ;
        RECT 138.170 160.470 141.210 160.640 ;
        RECT 138.170 160.030 141.210 160.200 ;
        RECT 141.425 160.170 141.595 160.500 ;
        RECT 141.930 160.280 154.380 161.040 ;
        RECT 141.930 160.270 154.270 160.280 ;
        RECT 141.930 160.260 147.810 160.270 ;
        RECT 141.930 160.240 142.500 160.260 ;
        RECT 143.720 160.250 147.810 160.260 ;
        RECT 141.940 159.630 142.110 160.240 ;
        RECT 137.630 159.460 142.110 159.630 ;
        RECT 98.430 158.040 104.170 158.050 ;
        RECT 97.940 157.880 104.170 158.040 ;
        RECT 97.940 155.620 98.610 157.880 ;
        RECT 99.280 157.310 103.320 157.480 ;
        RECT 98.940 156.250 99.110 157.250 ;
        RECT 103.490 156.250 103.660 157.250 ;
        RECT 99.280 156.020 103.320 156.190 ;
        RECT 104.000 155.620 104.170 157.880 ;
        RECT 97.940 155.450 104.170 155.620 ;
        RECT 97.940 152.190 98.610 155.450 ;
        RECT 99.280 154.880 103.320 155.050 ;
        RECT 98.940 152.820 99.110 154.820 ;
        RECT 103.490 152.820 103.660 154.820 ;
        RECT 99.280 152.590 103.320 152.760 ;
        RECT 104.000 152.190 104.170 155.450 ;
        RECT 97.940 152.020 104.170 152.190 ;
        RECT 97.940 148.760 98.610 152.020 ;
        RECT 99.280 151.450 103.320 151.620 ;
        RECT 98.940 149.390 99.110 151.390 ;
        RECT 103.490 149.390 103.660 151.390 ;
        RECT 99.280 149.160 103.320 149.330 ;
        RECT 104.000 148.760 104.170 152.020 ;
        RECT 97.940 148.750 104.170 148.760 ;
        RECT 105.760 158.020 115.590 158.060 ;
        RECT 117.470 158.040 123.210 158.050 ;
        RECT 105.760 157.890 116.390 158.020 ;
        RECT 105.760 155.630 105.930 157.890 ;
        RECT 106.655 157.320 114.695 157.490 ;
        RECT 106.270 156.260 106.440 157.260 ;
        RECT 114.910 156.260 115.080 157.260 ;
        RECT 106.655 156.030 114.695 156.200 ;
        RECT 115.420 155.630 116.390 157.890 ;
        RECT 105.760 155.460 116.390 155.630 ;
        RECT 105.760 152.200 105.930 155.460 ;
        RECT 106.655 154.890 114.695 155.060 ;
        RECT 106.270 152.830 106.440 154.830 ;
        RECT 114.910 152.830 115.080 154.830 ;
        RECT 106.655 152.600 114.695 152.770 ;
        RECT 115.420 152.200 116.390 155.460 ;
        RECT 105.760 152.030 116.390 152.200 ;
        RECT 105.760 148.770 105.930 152.030 ;
        RECT 106.655 151.460 114.695 151.630 ;
        RECT 106.270 149.400 106.440 151.400 ;
        RECT 114.910 149.400 115.080 151.400 ;
        RECT 106.655 149.170 114.695 149.340 ;
        RECT 115.420 148.770 116.390 152.030 ;
        RECT 97.940 148.650 104.180 148.750 ;
        RECT 97.930 148.090 104.180 148.650 ;
        RECT 97.930 148.070 103.100 148.090 ;
        RECT 97.930 148.000 101.920 148.070 ;
        RECT 97.930 146.730 99.850 148.000 ;
        RECT 101.360 147.990 101.920 148.000 ;
        RECT 101.590 146.900 101.920 147.990 ;
        RECT 102.290 147.520 103.330 147.690 ;
        RECT 102.290 147.080 103.330 147.250 ;
        RECT 103.500 147.220 103.670 147.550 ;
        RECT 101.750 146.680 101.920 146.900 ;
        RECT 104.010 146.680 104.180 148.090 ;
        RECT 101.750 146.510 104.180 146.680 ;
        RECT 105.760 148.600 116.390 148.770 ;
        RECT 116.980 157.880 123.210 158.040 ;
        RECT 116.980 155.620 117.650 157.880 ;
        RECT 118.320 157.310 122.360 157.480 ;
        RECT 117.980 156.250 118.150 157.250 ;
        RECT 122.530 156.250 122.700 157.250 ;
        RECT 118.320 156.020 122.360 156.190 ;
        RECT 123.040 155.620 123.210 157.880 ;
        RECT 116.980 155.450 123.210 155.620 ;
        RECT 116.980 152.190 117.650 155.450 ;
        RECT 118.320 154.880 122.360 155.050 ;
        RECT 117.980 152.820 118.150 154.820 ;
        RECT 122.530 152.820 122.700 154.820 ;
        RECT 118.320 152.590 122.360 152.760 ;
        RECT 123.040 152.190 123.210 155.450 ;
        RECT 116.980 152.020 123.210 152.190 ;
        RECT 116.980 148.760 117.650 152.020 ;
        RECT 118.320 151.450 122.360 151.620 ;
        RECT 117.980 149.390 118.150 151.390 ;
        RECT 122.530 149.390 122.700 151.390 ;
        RECT 118.320 149.160 122.360 149.330 ;
        RECT 123.040 148.760 123.210 152.020 ;
        RECT 116.980 148.750 123.210 148.760 ;
        RECT 124.800 158.020 134.630 158.060 ;
        RECT 136.470 158.040 142.210 158.050 ;
        RECT 124.800 157.890 135.430 158.020 ;
        RECT 124.800 155.630 124.970 157.890 ;
        RECT 125.695 157.320 133.735 157.490 ;
        RECT 125.310 156.260 125.480 157.260 ;
        RECT 133.950 156.260 134.120 157.260 ;
        RECT 125.695 156.030 133.735 156.200 ;
        RECT 134.460 155.630 135.430 157.890 ;
        RECT 124.800 155.460 135.430 155.630 ;
        RECT 124.800 152.200 124.970 155.460 ;
        RECT 125.695 154.890 133.735 155.060 ;
        RECT 125.310 152.830 125.480 154.830 ;
        RECT 133.950 152.830 134.120 154.830 ;
        RECT 125.695 152.600 133.735 152.770 ;
        RECT 134.460 152.200 135.430 155.460 ;
        RECT 124.800 152.030 135.430 152.200 ;
        RECT 124.800 148.770 124.970 152.030 ;
        RECT 125.695 151.460 133.735 151.630 ;
        RECT 125.310 149.400 125.480 151.400 ;
        RECT 133.950 149.400 134.120 151.400 ;
        RECT 125.695 149.170 133.735 149.340 ;
        RECT 134.460 148.770 135.430 152.030 ;
        RECT 116.980 148.650 123.220 148.750 ;
        RECT 105.760 146.340 105.930 148.600 ;
        RECT 106.655 148.030 114.695 148.200 ;
        RECT 106.270 146.970 106.440 147.970 ;
        RECT 114.910 146.970 115.080 147.970 ;
        RECT 106.655 146.740 114.695 146.910 ;
        RECT 115.420 146.340 116.390 148.600 ;
        RECT 116.970 148.090 123.220 148.650 ;
        RECT 116.970 148.070 122.140 148.090 ;
        RECT 116.970 148.000 120.960 148.070 ;
        RECT 116.970 146.730 118.890 148.000 ;
        RECT 120.400 147.990 120.960 148.000 ;
        RECT 120.630 146.900 120.960 147.990 ;
        RECT 121.330 147.520 122.370 147.690 ;
        RECT 121.330 147.080 122.370 147.250 ;
        RECT 122.540 147.220 122.710 147.550 ;
        RECT 120.790 146.680 120.960 146.900 ;
        RECT 123.050 146.680 123.220 148.090 ;
        RECT 120.790 146.510 123.220 146.680 ;
        RECT 124.800 148.600 135.430 148.770 ;
        RECT 135.980 157.880 142.210 158.040 ;
        RECT 135.980 155.620 136.650 157.880 ;
        RECT 137.320 157.310 141.360 157.480 ;
        RECT 136.980 156.250 137.150 157.250 ;
        RECT 141.530 156.250 141.700 157.250 ;
        RECT 137.320 156.020 141.360 156.190 ;
        RECT 142.040 155.620 142.210 157.880 ;
        RECT 135.980 155.450 142.210 155.620 ;
        RECT 135.980 152.190 136.650 155.450 ;
        RECT 137.320 154.880 141.360 155.050 ;
        RECT 136.980 152.820 137.150 154.820 ;
        RECT 141.530 152.820 141.700 154.820 ;
        RECT 137.320 152.590 141.360 152.760 ;
        RECT 142.040 152.190 142.210 155.450 ;
        RECT 135.980 152.020 142.210 152.190 ;
        RECT 135.980 148.760 136.650 152.020 ;
        RECT 137.320 151.450 141.360 151.620 ;
        RECT 136.980 149.390 137.150 151.390 ;
        RECT 141.530 149.390 141.700 151.390 ;
        RECT 137.320 149.160 141.360 149.330 ;
        RECT 142.040 148.760 142.210 152.020 ;
        RECT 135.980 148.750 142.210 148.760 ;
        RECT 143.800 158.020 153.630 158.060 ;
        RECT 143.800 157.890 154.430 158.020 ;
        RECT 143.800 155.630 143.970 157.890 ;
        RECT 144.695 157.320 152.735 157.490 ;
        RECT 144.310 156.260 144.480 157.260 ;
        RECT 152.950 156.260 153.120 157.260 ;
        RECT 144.695 156.030 152.735 156.200 ;
        RECT 153.460 155.630 154.430 157.890 ;
        RECT 143.800 155.460 154.430 155.630 ;
        RECT 143.800 152.200 143.970 155.460 ;
        RECT 144.695 154.890 152.735 155.060 ;
        RECT 144.310 152.830 144.480 154.830 ;
        RECT 152.950 152.830 153.120 154.830 ;
        RECT 144.695 152.600 152.735 152.770 ;
        RECT 153.460 152.200 154.430 155.460 ;
        RECT 143.800 152.030 154.430 152.200 ;
        RECT 143.800 148.770 143.970 152.030 ;
        RECT 144.695 151.460 152.735 151.630 ;
        RECT 144.310 149.400 144.480 151.400 ;
        RECT 152.950 149.400 153.120 151.400 ;
        RECT 144.695 149.170 152.735 149.340 ;
        RECT 153.460 148.770 154.430 152.030 ;
        RECT 135.980 148.650 142.220 148.750 ;
        RECT 105.760 146.310 116.390 146.340 ;
        RECT 124.800 146.340 124.970 148.600 ;
        RECT 125.695 148.030 133.735 148.200 ;
        RECT 125.310 146.970 125.480 147.970 ;
        RECT 133.950 146.970 134.120 147.970 ;
        RECT 125.695 146.740 133.735 146.910 ;
        RECT 134.460 146.340 135.430 148.600 ;
        RECT 135.970 148.090 142.220 148.650 ;
        RECT 135.970 148.070 141.140 148.090 ;
        RECT 135.970 148.000 139.960 148.070 ;
        RECT 135.970 146.730 137.890 148.000 ;
        RECT 139.400 147.990 139.960 148.000 ;
        RECT 139.630 146.900 139.960 147.990 ;
        RECT 140.330 147.520 141.370 147.690 ;
        RECT 140.330 147.080 141.370 147.250 ;
        RECT 141.540 147.220 141.710 147.550 ;
        RECT 139.790 146.680 139.960 146.900 ;
        RECT 142.050 146.680 142.220 148.090 ;
        RECT 139.790 146.510 142.220 146.680 ;
        RECT 143.800 148.600 154.430 148.770 ;
        RECT 124.800 146.310 135.430 146.340 ;
        RECT 143.800 146.340 143.970 148.600 ;
        RECT 144.695 148.030 152.735 148.200 ;
        RECT 144.310 146.970 144.480 147.970 ;
        RECT 152.950 146.970 153.120 147.970 ;
        RECT 144.695 146.740 152.735 146.910 ;
        RECT 153.460 146.340 154.430 148.600 ;
        RECT 143.800 146.310 154.430 146.340 ;
        RECT 105.730 146.200 116.390 146.310 ;
        RECT 124.770 146.200 135.430 146.310 ;
        RECT 143.770 146.200 154.430 146.310 ;
        RECT 103.980 146.150 116.390 146.200 ;
        RECT 123.020 146.150 135.430 146.200 ;
        RECT 142.020 146.150 154.430 146.200 ;
        RECT 99.640 145.980 116.390 146.150 ;
        RECT 99.640 144.570 99.810 145.980 ;
        RECT 100.180 145.410 103.220 145.580 ;
        RECT 100.180 144.970 103.220 145.140 ;
        RECT 103.435 145.110 103.605 145.440 ;
        RECT 103.940 145.220 116.390 145.980 ;
        RECT 118.680 145.980 135.430 146.150 ;
        RECT 103.940 145.210 116.280 145.220 ;
        RECT 103.940 145.200 109.820 145.210 ;
        RECT 103.940 145.180 104.510 145.200 ;
        RECT 105.730 145.190 109.820 145.200 ;
        RECT 103.950 144.570 104.120 145.180 ;
        RECT 99.640 144.400 104.120 144.570 ;
        RECT 118.680 144.570 118.850 145.980 ;
        RECT 119.220 145.410 122.260 145.580 ;
        RECT 119.220 144.970 122.260 145.140 ;
        RECT 122.475 145.110 122.645 145.440 ;
        RECT 122.980 145.220 135.430 145.980 ;
        RECT 137.680 145.980 154.430 146.150 ;
        RECT 122.980 145.210 135.320 145.220 ;
        RECT 122.980 145.200 128.860 145.210 ;
        RECT 122.980 145.180 123.550 145.200 ;
        RECT 124.770 145.190 128.860 145.200 ;
        RECT 122.990 144.570 123.160 145.180 ;
        RECT 118.680 144.400 123.160 144.570 ;
        RECT 137.680 144.570 137.850 145.980 ;
        RECT 138.220 145.410 141.260 145.580 ;
        RECT 138.220 144.970 141.260 145.140 ;
        RECT 141.475 145.110 141.645 145.440 ;
        RECT 141.980 145.220 154.430 145.980 ;
        RECT 141.980 145.210 154.320 145.220 ;
        RECT 141.980 145.200 147.860 145.210 ;
        RECT 141.980 145.180 142.550 145.200 ;
        RECT 143.770 145.190 147.860 145.200 ;
        RECT 141.990 144.570 142.160 145.180 ;
        RECT 137.680 144.400 142.160 144.570 ;
        RECT 98.430 143.060 104.170 143.070 ;
        RECT 97.940 142.900 104.170 143.060 ;
        RECT 97.940 140.640 98.610 142.900 ;
        RECT 99.280 142.330 103.320 142.500 ;
        RECT 98.940 141.270 99.110 142.270 ;
        RECT 103.490 141.270 103.660 142.270 ;
        RECT 99.280 141.040 103.320 141.210 ;
        RECT 104.000 140.640 104.170 142.900 ;
        RECT 97.940 140.470 104.170 140.640 ;
        RECT 97.940 137.210 98.610 140.470 ;
        RECT 99.280 139.900 103.320 140.070 ;
        RECT 98.940 137.840 99.110 139.840 ;
        RECT 103.490 137.840 103.660 139.840 ;
        RECT 99.280 137.610 103.320 137.780 ;
        RECT 104.000 137.210 104.170 140.470 ;
        RECT 97.940 137.040 104.170 137.210 ;
        RECT 97.940 133.780 98.610 137.040 ;
        RECT 99.280 136.470 103.320 136.640 ;
        RECT 98.940 134.410 99.110 136.410 ;
        RECT 103.490 134.410 103.660 136.410 ;
        RECT 99.280 134.180 103.320 134.350 ;
        RECT 104.000 133.780 104.170 137.040 ;
        RECT 97.940 133.770 104.170 133.780 ;
        RECT 105.760 143.040 115.590 143.080 ;
        RECT 105.760 142.910 116.390 143.040 ;
        RECT 117.420 143.020 123.160 143.030 ;
        RECT 105.760 140.650 105.930 142.910 ;
        RECT 106.655 142.340 114.695 142.510 ;
        RECT 106.270 141.280 106.440 142.280 ;
        RECT 114.910 141.280 115.080 142.280 ;
        RECT 106.655 141.050 114.695 141.220 ;
        RECT 115.420 140.650 116.390 142.910 ;
        RECT 105.760 140.480 116.390 140.650 ;
        RECT 105.760 137.220 105.930 140.480 ;
        RECT 106.655 139.910 114.695 140.080 ;
        RECT 106.270 137.850 106.440 139.850 ;
        RECT 114.910 137.850 115.080 139.850 ;
        RECT 106.655 137.620 114.695 137.790 ;
        RECT 115.420 137.220 116.390 140.480 ;
        RECT 105.760 137.050 116.390 137.220 ;
        RECT 105.760 133.790 105.930 137.050 ;
        RECT 106.655 136.480 114.695 136.650 ;
        RECT 106.270 134.420 106.440 136.420 ;
        RECT 114.910 134.420 115.080 136.420 ;
        RECT 106.655 134.190 114.695 134.360 ;
        RECT 115.420 133.790 116.390 137.050 ;
        RECT 97.940 133.670 104.180 133.770 ;
        RECT 97.930 133.110 104.180 133.670 ;
        RECT 97.930 133.090 103.100 133.110 ;
        RECT 97.930 133.020 101.920 133.090 ;
        RECT 97.930 131.750 99.850 133.020 ;
        RECT 101.360 133.010 101.920 133.020 ;
        RECT 101.590 131.920 101.920 133.010 ;
        RECT 102.290 132.540 103.330 132.710 ;
        RECT 102.290 132.100 103.330 132.270 ;
        RECT 103.500 132.240 103.670 132.570 ;
        RECT 101.750 131.700 101.920 131.920 ;
        RECT 104.010 131.700 104.180 133.110 ;
        RECT 101.750 131.530 104.180 131.700 ;
        RECT 105.760 133.620 116.390 133.790 ;
        RECT 116.930 142.860 123.160 143.020 ;
        RECT 116.930 140.600 117.600 142.860 ;
        RECT 118.270 142.290 122.310 142.460 ;
        RECT 117.930 141.230 118.100 142.230 ;
        RECT 122.480 141.230 122.650 142.230 ;
        RECT 118.270 141.000 122.310 141.170 ;
        RECT 122.990 140.600 123.160 142.860 ;
        RECT 116.930 140.430 123.160 140.600 ;
        RECT 116.930 137.170 117.600 140.430 ;
        RECT 118.270 139.860 122.310 140.030 ;
        RECT 117.930 137.800 118.100 139.800 ;
        RECT 122.480 137.800 122.650 139.800 ;
        RECT 118.270 137.570 122.310 137.740 ;
        RECT 122.990 137.170 123.160 140.430 ;
        RECT 116.930 137.000 123.160 137.170 ;
        RECT 116.930 133.740 117.600 137.000 ;
        RECT 118.270 136.430 122.310 136.600 ;
        RECT 117.930 134.370 118.100 136.370 ;
        RECT 122.480 134.370 122.650 136.370 ;
        RECT 118.270 134.140 122.310 134.310 ;
        RECT 122.990 133.740 123.160 137.000 ;
        RECT 116.930 133.730 123.160 133.740 ;
        RECT 124.750 143.000 134.580 143.040 ;
        RECT 136.420 143.020 142.160 143.030 ;
        RECT 124.750 142.870 135.380 143.000 ;
        RECT 124.750 140.610 124.920 142.870 ;
        RECT 125.645 142.300 133.685 142.470 ;
        RECT 125.260 141.240 125.430 142.240 ;
        RECT 133.900 141.240 134.070 142.240 ;
        RECT 125.645 141.010 133.685 141.180 ;
        RECT 134.410 140.610 135.380 142.870 ;
        RECT 124.750 140.440 135.380 140.610 ;
        RECT 124.750 137.180 124.920 140.440 ;
        RECT 125.645 139.870 133.685 140.040 ;
        RECT 125.260 137.810 125.430 139.810 ;
        RECT 133.900 137.810 134.070 139.810 ;
        RECT 125.645 137.580 133.685 137.750 ;
        RECT 134.410 137.180 135.380 140.440 ;
        RECT 124.750 137.010 135.380 137.180 ;
        RECT 124.750 133.750 124.920 137.010 ;
        RECT 125.645 136.440 133.685 136.610 ;
        RECT 125.260 134.380 125.430 136.380 ;
        RECT 133.900 134.380 134.070 136.380 ;
        RECT 125.645 134.150 133.685 134.320 ;
        RECT 134.410 133.750 135.380 137.010 ;
        RECT 116.930 133.630 123.170 133.730 ;
        RECT 105.760 131.360 105.930 133.620 ;
        RECT 106.655 133.050 114.695 133.220 ;
        RECT 106.270 131.990 106.440 132.990 ;
        RECT 114.910 131.990 115.080 132.990 ;
        RECT 106.655 131.760 114.695 131.930 ;
        RECT 115.420 131.360 116.390 133.620 ;
        RECT 116.920 133.070 123.170 133.630 ;
        RECT 116.920 133.050 122.090 133.070 ;
        RECT 116.920 132.980 120.910 133.050 ;
        RECT 116.920 131.710 118.840 132.980 ;
        RECT 120.350 132.970 120.910 132.980 ;
        RECT 120.580 131.880 120.910 132.970 ;
        RECT 121.280 132.500 122.320 132.670 ;
        RECT 121.280 132.060 122.320 132.230 ;
        RECT 122.490 132.200 122.660 132.530 ;
        RECT 120.740 131.660 120.910 131.880 ;
        RECT 123.000 131.660 123.170 133.070 ;
        RECT 120.740 131.490 123.170 131.660 ;
        RECT 124.750 133.580 135.380 133.750 ;
        RECT 135.930 142.860 142.160 143.020 ;
        RECT 135.930 140.600 136.600 142.860 ;
        RECT 137.270 142.290 141.310 142.460 ;
        RECT 136.930 141.230 137.100 142.230 ;
        RECT 141.480 141.230 141.650 142.230 ;
        RECT 137.270 141.000 141.310 141.170 ;
        RECT 141.990 140.600 142.160 142.860 ;
        RECT 135.930 140.430 142.160 140.600 ;
        RECT 135.930 137.170 136.600 140.430 ;
        RECT 137.270 139.860 141.310 140.030 ;
        RECT 136.930 137.800 137.100 139.800 ;
        RECT 141.480 137.800 141.650 139.800 ;
        RECT 137.270 137.570 141.310 137.740 ;
        RECT 141.990 137.170 142.160 140.430 ;
        RECT 135.930 137.000 142.160 137.170 ;
        RECT 135.930 133.740 136.600 137.000 ;
        RECT 137.270 136.430 141.310 136.600 ;
        RECT 136.930 134.370 137.100 136.370 ;
        RECT 141.480 134.370 141.650 136.370 ;
        RECT 137.270 134.140 141.310 134.310 ;
        RECT 141.990 133.740 142.160 137.000 ;
        RECT 135.930 133.730 142.160 133.740 ;
        RECT 143.750 143.000 153.580 143.040 ;
        RECT 143.750 142.870 154.380 143.000 ;
        RECT 143.750 140.610 143.920 142.870 ;
        RECT 144.645 142.300 152.685 142.470 ;
        RECT 144.260 141.240 144.430 142.240 ;
        RECT 152.900 141.240 153.070 142.240 ;
        RECT 144.645 141.010 152.685 141.180 ;
        RECT 153.410 140.610 154.380 142.870 ;
        RECT 143.750 140.440 154.380 140.610 ;
        RECT 143.750 137.180 143.920 140.440 ;
        RECT 144.645 139.870 152.685 140.040 ;
        RECT 144.260 137.810 144.430 139.810 ;
        RECT 152.900 137.810 153.070 139.810 ;
        RECT 144.645 137.580 152.685 137.750 ;
        RECT 153.410 137.180 154.380 140.440 ;
        RECT 143.750 137.010 154.380 137.180 ;
        RECT 143.750 133.750 143.920 137.010 ;
        RECT 144.645 136.440 152.685 136.610 ;
        RECT 144.260 134.380 144.430 136.380 ;
        RECT 152.900 134.380 153.070 136.380 ;
        RECT 144.645 134.150 152.685 134.320 ;
        RECT 153.410 133.750 154.380 137.010 ;
        RECT 135.930 133.630 142.170 133.730 ;
        RECT 105.760 131.330 116.390 131.360 ;
        RECT 105.730 131.220 116.390 131.330 ;
        RECT 124.750 131.320 124.920 133.580 ;
        RECT 125.645 133.010 133.685 133.180 ;
        RECT 125.260 131.950 125.430 132.950 ;
        RECT 133.900 131.950 134.070 132.950 ;
        RECT 125.645 131.720 133.685 131.890 ;
        RECT 134.410 131.320 135.380 133.580 ;
        RECT 135.920 133.070 142.170 133.630 ;
        RECT 135.920 133.050 141.090 133.070 ;
        RECT 135.920 132.980 139.910 133.050 ;
        RECT 135.920 131.710 137.840 132.980 ;
        RECT 139.350 132.970 139.910 132.980 ;
        RECT 139.580 131.880 139.910 132.970 ;
        RECT 140.280 132.500 141.320 132.670 ;
        RECT 140.280 132.060 141.320 132.230 ;
        RECT 141.490 132.200 141.660 132.530 ;
        RECT 139.740 131.660 139.910 131.880 ;
        RECT 142.000 131.660 142.170 133.070 ;
        RECT 139.740 131.490 142.170 131.660 ;
        RECT 143.750 133.580 154.380 133.750 ;
        RECT 124.750 131.290 135.380 131.320 ;
        RECT 143.750 131.320 143.920 133.580 ;
        RECT 144.645 133.010 152.685 133.180 ;
        RECT 144.260 131.950 144.430 132.950 ;
        RECT 152.900 131.950 153.070 132.950 ;
        RECT 144.645 131.720 152.685 131.890 ;
        RECT 153.410 131.320 154.380 133.580 ;
        RECT 143.750 131.290 154.380 131.320 ;
        RECT 103.980 131.170 116.390 131.220 ;
        RECT 124.720 131.180 135.380 131.290 ;
        RECT 143.720 131.180 154.380 131.290 ;
        RECT 99.640 131.000 116.390 131.170 ;
        RECT 122.970 131.130 135.380 131.180 ;
        RECT 141.970 131.130 154.380 131.180 ;
        RECT 99.640 129.590 99.810 131.000 ;
        RECT 100.180 130.430 103.220 130.600 ;
        RECT 100.180 129.990 103.220 130.160 ;
        RECT 103.435 130.130 103.605 130.460 ;
        RECT 103.940 130.240 116.390 131.000 ;
        RECT 118.630 130.960 135.380 131.130 ;
        RECT 103.940 130.230 116.280 130.240 ;
        RECT 103.940 130.220 109.820 130.230 ;
        RECT 103.940 130.200 104.510 130.220 ;
        RECT 105.730 130.210 109.820 130.220 ;
        RECT 103.950 129.590 104.120 130.200 ;
        RECT 99.640 129.420 104.120 129.590 ;
        RECT 118.630 129.550 118.800 130.960 ;
        RECT 119.170 130.390 122.210 130.560 ;
        RECT 119.170 129.950 122.210 130.120 ;
        RECT 122.425 130.090 122.595 130.420 ;
        RECT 122.930 130.200 135.380 130.960 ;
        RECT 137.630 130.960 154.380 131.130 ;
        RECT 122.930 130.190 135.270 130.200 ;
        RECT 122.930 130.180 128.810 130.190 ;
        RECT 122.930 130.160 123.500 130.180 ;
        RECT 124.720 130.170 128.810 130.180 ;
        RECT 122.940 129.550 123.110 130.160 ;
        RECT 118.630 129.380 123.110 129.550 ;
        RECT 137.630 129.550 137.800 130.960 ;
        RECT 138.170 130.390 141.210 130.560 ;
        RECT 138.170 129.950 141.210 130.120 ;
        RECT 141.425 130.090 141.595 130.420 ;
        RECT 141.930 130.200 154.380 130.960 ;
        RECT 141.930 130.190 154.270 130.200 ;
        RECT 141.930 130.180 147.810 130.190 ;
        RECT 141.930 130.160 142.500 130.180 ;
        RECT 143.720 130.170 147.810 130.180 ;
        RECT 141.940 129.550 142.110 130.160 ;
        RECT 137.630 129.380 142.110 129.550 ;
        RECT 98.430 128.030 104.170 128.040 ;
        RECT 97.940 127.870 104.170 128.030 ;
        RECT 97.940 125.610 98.610 127.870 ;
        RECT 99.280 127.300 103.320 127.470 ;
        RECT 98.940 126.240 99.110 127.240 ;
        RECT 103.490 126.240 103.660 127.240 ;
        RECT 99.280 126.010 103.320 126.180 ;
        RECT 104.000 125.610 104.170 127.870 ;
        RECT 97.940 125.440 104.170 125.610 ;
        RECT 97.940 122.180 98.610 125.440 ;
        RECT 99.280 124.870 103.320 125.040 ;
        RECT 98.940 122.810 99.110 124.810 ;
        RECT 103.490 122.810 103.660 124.810 ;
        RECT 99.280 122.580 103.320 122.750 ;
        RECT 104.000 122.180 104.170 125.440 ;
        RECT 97.940 122.010 104.170 122.180 ;
        RECT 97.940 118.750 98.610 122.010 ;
        RECT 99.280 121.440 103.320 121.610 ;
        RECT 98.940 119.380 99.110 121.380 ;
        RECT 103.490 119.380 103.660 121.380 ;
        RECT 99.280 119.150 103.320 119.320 ;
        RECT 104.000 118.750 104.170 122.010 ;
        RECT 97.940 118.740 104.170 118.750 ;
        RECT 105.760 128.010 115.590 128.050 ;
        RECT 105.760 127.880 116.390 128.010 ;
        RECT 117.420 128.000 123.160 128.010 ;
        RECT 105.760 125.620 105.930 127.880 ;
        RECT 106.655 127.310 114.695 127.480 ;
        RECT 106.270 126.250 106.440 127.250 ;
        RECT 114.910 126.250 115.080 127.250 ;
        RECT 106.655 126.020 114.695 126.190 ;
        RECT 115.420 125.620 116.390 127.880 ;
        RECT 105.760 125.450 116.390 125.620 ;
        RECT 105.760 122.190 105.930 125.450 ;
        RECT 106.655 124.880 114.695 125.050 ;
        RECT 106.270 122.820 106.440 124.820 ;
        RECT 114.910 122.820 115.080 124.820 ;
        RECT 106.655 122.590 114.695 122.760 ;
        RECT 115.420 122.190 116.390 125.450 ;
        RECT 105.760 122.020 116.390 122.190 ;
        RECT 105.760 118.760 105.930 122.020 ;
        RECT 106.655 121.450 114.695 121.620 ;
        RECT 106.270 119.390 106.440 121.390 ;
        RECT 114.910 119.390 115.080 121.390 ;
        RECT 106.655 119.160 114.695 119.330 ;
        RECT 115.420 118.760 116.390 122.020 ;
        RECT 97.940 118.640 104.180 118.740 ;
        RECT 97.930 118.080 104.180 118.640 ;
        RECT 97.930 118.060 103.100 118.080 ;
        RECT 97.930 117.990 101.920 118.060 ;
        RECT 97.930 116.720 99.850 117.990 ;
        RECT 101.360 117.980 101.920 117.990 ;
        RECT 101.590 116.890 101.920 117.980 ;
        RECT 102.290 117.510 103.330 117.680 ;
        RECT 102.290 117.070 103.330 117.240 ;
        RECT 103.500 117.210 103.670 117.540 ;
        RECT 101.750 116.670 101.920 116.890 ;
        RECT 104.010 116.670 104.180 118.080 ;
        RECT 101.750 116.500 104.180 116.670 ;
        RECT 105.760 118.590 116.390 118.760 ;
        RECT 116.930 127.840 123.160 128.000 ;
        RECT 116.930 125.580 117.600 127.840 ;
        RECT 118.270 127.270 122.310 127.440 ;
        RECT 117.930 126.210 118.100 127.210 ;
        RECT 122.480 126.210 122.650 127.210 ;
        RECT 118.270 125.980 122.310 126.150 ;
        RECT 122.990 125.580 123.160 127.840 ;
        RECT 116.930 125.410 123.160 125.580 ;
        RECT 116.930 122.150 117.600 125.410 ;
        RECT 118.270 124.840 122.310 125.010 ;
        RECT 117.930 122.780 118.100 124.780 ;
        RECT 122.480 122.780 122.650 124.780 ;
        RECT 118.270 122.550 122.310 122.720 ;
        RECT 122.990 122.150 123.160 125.410 ;
        RECT 116.930 121.980 123.160 122.150 ;
        RECT 116.930 118.720 117.600 121.980 ;
        RECT 118.270 121.410 122.310 121.580 ;
        RECT 117.930 119.350 118.100 121.350 ;
        RECT 122.480 119.350 122.650 121.350 ;
        RECT 118.270 119.120 122.310 119.290 ;
        RECT 122.990 118.720 123.160 121.980 ;
        RECT 116.930 118.710 123.160 118.720 ;
        RECT 124.750 127.980 134.580 128.020 ;
        RECT 136.420 128.000 142.160 128.010 ;
        RECT 124.750 127.850 135.380 127.980 ;
        RECT 124.750 125.590 124.920 127.850 ;
        RECT 125.645 127.280 133.685 127.450 ;
        RECT 125.260 126.220 125.430 127.220 ;
        RECT 133.900 126.220 134.070 127.220 ;
        RECT 125.645 125.990 133.685 126.160 ;
        RECT 134.410 125.590 135.380 127.850 ;
        RECT 124.750 125.420 135.380 125.590 ;
        RECT 124.750 122.160 124.920 125.420 ;
        RECT 125.645 124.850 133.685 125.020 ;
        RECT 125.260 122.790 125.430 124.790 ;
        RECT 133.900 122.790 134.070 124.790 ;
        RECT 125.645 122.560 133.685 122.730 ;
        RECT 134.410 122.160 135.380 125.420 ;
        RECT 124.750 121.990 135.380 122.160 ;
        RECT 124.750 118.730 124.920 121.990 ;
        RECT 125.645 121.420 133.685 121.590 ;
        RECT 125.260 119.360 125.430 121.360 ;
        RECT 133.900 119.360 134.070 121.360 ;
        RECT 125.645 119.130 133.685 119.300 ;
        RECT 134.410 118.730 135.380 121.990 ;
        RECT 116.930 118.610 123.170 118.710 ;
        RECT 105.760 116.330 105.930 118.590 ;
        RECT 106.655 118.020 114.695 118.190 ;
        RECT 106.270 116.960 106.440 117.960 ;
        RECT 114.910 116.960 115.080 117.960 ;
        RECT 106.655 116.730 114.695 116.900 ;
        RECT 115.420 116.330 116.390 118.590 ;
        RECT 116.920 118.050 123.170 118.610 ;
        RECT 116.920 118.030 122.090 118.050 ;
        RECT 116.920 117.960 120.910 118.030 ;
        RECT 116.920 116.690 118.840 117.960 ;
        RECT 120.350 117.950 120.910 117.960 ;
        RECT 120.580 116.860 120.910 117.950 ;
        RECT 121.280 117.480 122.320 117.650 ;
        RECT 121.280 117.040 122.320 117.210 ;
        RECT 122.490 117.180 122.660 117.510 ;
        RECT 120.740 116.640 120.910 116.860 ;
        RECT 123.000 116.640 123.170 118.050 ;
        RECT 120.740 116.470 123.170 116.640 ;
        RECT 124.750 118.560 135.380 118.730 ;
        RECT 135.930 127.840 142.160 128.000 ;
        RECT 135.930 125.580 136.600 127.840 ;
        RECT 137.270 127.270 141.310 127.440 ;
        RECT 136.930 126.210 137.100 127.210 ;
        RECT 141.480 126.210 141.650 127.210 ;
        RECT 137.270 125.980 141.310 126.150 ;
        RECT 141.990 125.580 142.160 127.840 ;
        RECT 135.930 125.410 142.160 125.580 ;
        RECT 135.930 122.150 136.600 125.410 ;
        RECT 137.270 124.840 141.310 125.010 ;
        RECT 136.930 122.780 137.100 124.780 ;
        RECT 141.480 122.780 141.650 124.780 ;
        RECT 137.270 122.550 141.310 122.720 ;
        RECT 141.990 122.150 142.160 125.410 ;
        RECT 135.930 121.980 142.160 122.150 ;
        RECT 135.930 118.720 136.600 121.980 ;
        RECT 137.270 121.410 141.310 121.580 ;
        RECT 136.930 119.350 137.100 121.350 ;
        RECT 141.480 119.350 141.650 121.350 ;
        RECT 137.270 119.120 141.310 119.290 ;
        RECT 141.990 118.720 142.160 121.980 ;
        RECT 135.930 118.710 142.160 118.720 ;
        RECT 143.750 127.980 153.580 128.020 ;
        RECT 143.750 127.850 154.380 127.980 ;
        RECT 143.750 125.590 143.920 127.850 ;
        RECT 144.645 127.280 152.685 127.450 ;
        RECT 144.260 126.220 144.430 127.220 ;
        RECT 152.900 126.220 153.070 127.220 ;
        RECT 144.645 125.990 152.685 126.160 ;
        RECT 153.410 125.590 154.380 127.850 ;
        RECT 143.750 125.420 154.380 125.590 ;
        RECT 143.750 122.160 143.920 125.420 ;
        RECT 144.645 124.850 152.685 125.020 ;
        RECT 144.260 122.790 144.430 124.790 ;
        RECT 152.900 122.790 153.070 124.790 ;
        RECT 144.645 122.560 152.685 122.730 ;
        RECT 153.410 122.160 154.380 125.420 ;
        RECT 143.750 121.990 154.380 122.160 ;
        RECT 143.750 118.730 143.920 121.990 ;
        RECT 144.645 121.420 152.685 121.590 ;
        RECT 144.260 119.360 144.430 121.360 ;
        RECT 152.900 119.360 153.070 121.360 ;
        RECT 144.645 119.130 152.685 119.300 ;
        RECT 153.410 118.730 154.380 121.990 ;
        RECT 135.930 118.610 142.170 118.710 ;
        RECT 105.760 116.300 116.390 116.330 ;
        RECT 105.730 116.190 116.390 116.300 ;
        RECT 124.750 116.300 124.920 118.560 ;
        RECT 125.645 117.990 133.685 118.160 ;
        RECT 125.260 116.930 125.430 117.930 ;
        RECT 133.900 116.930 134.070 117.930 ;
        RECT 125.645 116.700 133.685 116.870 ;
        RECT 134.410 116.300 135.380 118.560 ;
        RECT 135.920 118.050 142.170 118.610 ;
        RECT 135.920 118.030 141.090 118.050 ;
        RECT 135.920 117.960 139.910 118.030 ;
        RECT 135.920 116.690 137.840 117.960 ;
        RECT 139.350 117.950 139.910 117.960 ;
        RECT 139.580 116.860 139.910 117.950 ;
        RECT 140.280 117.480 141.320 117.650 ;
        RECT 140.280 117.040 141.320 117.210 ;
        RECT 141.490 117.180 141.660 117.510 ;
        RECT 139.740 116.640 139.910 116.860 ;
        RECT 142.000 116.640 142.170 118.050 ;
        RECT 139.740 116.470 142.170 116.640 ;
        RECT 143.750 118.560 154.380 118.730 ;
        RECT 124.750 116.270 135.380 116.300 ;
        RECT 143.750 116.300 143.920 118.560 ;
        RECT 144.645 117.990 152.685 118.160 ;
        RECT 144.260 116.930 144.430 117.930 ;
        RECT 152.900 116.930 153.070 117.930 ;
        RECT 144.645 116.700 152.685 116.870 ;
        RECT 153.410 116.300 154.380 118.560 ;
        RECT 143.750 116.270 154.380 116.300 ;
        RECT 103.980 116.140 116.390 116.190 ;
        RECT 124.720 116.160 135.380 116.270 ;
        RECT 143.720 116.160 154.380 116.270 ;
        RECT 99.640 115.970 116.390 116.140 ;
        RECT 122.970 116.110 135.380 116.160 ;
        RECT 141.970 116.110 154.380 116.160 ;
        RECT 99.640 114.560 99.810 115.970 ;
        RECT 100.180 115.400 103.220 115.570 ;
        RECT 100.180 114.960 103.220 115.130 ;
        RECT 103.435 115.100 103.605 115.430 ;
        RECT 103.940 115.210 116.390 115.970 ;
        RECT 118.630 115.940 135.380 116.110 ;
        RECT 103.940 115.200 116.280 115.210 ;
        RECT 103.940 115.190 109.820 115.200 ;
        RECT 103.940 115.170 104.510 115.190 ;
        RECT 105.730 115.180 109.820 115.190 ;
        RECT 103.950 114.560 104.120 115.170 ;
        RECT 99.640 114.390 104.120 114.560 ;
        RECT 118.630 114.530 118.800 115.940 ;
        RECT 119.170 115.370 122.210 115.540 ;
        RECT 119.170 114.930 122.210 115.100 ;
        RECT 122.425 115.070 122.595 115.400 ;
        RECT 122.930 115.180 135.380 115.940 ;
        RECT 137.630 115.940 154.380 116.110 ;
        RECT 122.930 115.170 135.270 115.180 ;
        RECT 122.930 115.160 128.810 115.170 ;
        RECT 122.930 115.140 123.500 115.160 ;
        RECT 124.720 115.150 128.810 115.160 ;
        RECT 122.940 114.530 123.110 115.140 ;
        RECT 118.630 114.360 123.110 114.530 ;
        RECT 137.630 114.530 137.800 115.940 ;
        RECT 138.170 115.370 141.210 115.540 ;
        RECT 138.170 114.930 141.210 115.100 ;
        RECT 141.425 115.070 141.595 115.400 ;
        RECT 141.930 115.180 154.380 115.940 ;
        RECT 141.930 115.170 154.270 115.180 ;
        RECT 141.930 115.160 147.810 115.170 ;
        RECT 141.930 115.140 142.500 115.160 ;
        RECT 143.720 115.150 147.810 115.160 ;
        RECT 141.940 114.530 142.110 115.140 ;
        RECT 137.630 114.360 142.110 114.530 ;
        RECT 98.430 113.040 104.170 113.050 ;
        RECT 97.940 112.880 104.170 113.040 ;
        RECT 97.940 110.620 98.610 112.880 ;
        RECT 99.280 112.310 103.320 112.480 ;
        RECT 98.940 111.250 99.110 112.250 ;
        RECT 103.490 111.250 103.660 112.250 ;
        RECT 99.280 111.020 103.320 111.190 ;
        RECT 104.000 110.620 104.170 112.880 ;
        RECT 97.940 110.450 104.170 110.620 ;
        RECT 97.940 107.190 98.610 110.450 ;
        RECT 99.280 109.880 103.320 110.050 ;
        RECT 98.940 107.820 99.110 109.820 ;
        RECT 103.490 107.820 103.660 109.820 ;
        RECT 99.280 107.590 103.320 107.760 ;
        RECT 104.000 107.190 104.170 110.450 ;
        RECT 97.940 107.020 104.170 107.190 ;
        RECT 97.940 103.760 98.610 107.020 ;
        RECT 99.280 106.450 103.320 106.620 ;
        RECT 98.940 104.390 99.110 106.390 ;
        RECT 103.490 104.390 103.660 106.390 ;
        RECT 99.280 104.160 103.320 104.330 ;
        RECT 104.000 103.760 104.170 107.020 ;
        RECT 97.940 103.750 104.170 103.760 ;
        RECT 105.760 113.020 115.590 113.060 ;
        RECT 117.420 113.020 123.160 113.030 ;
        RECT 105.760 112.890 116.390 113.020 ;
        RECT 105.760 110.630 105.930 112.890 ;
        RECT 106.655 112.320 114.695 112.490 ;
        RECT 106.270 111.260 106.440 112.260 ;
        RECT 114.910 111.260 115.080 112.260 ;
        RECT 106.655 111.030 114.695 111.200 ;
        RECT 115.420 110.630 116.390 112.890 ;
        RECT 105.760 110.460 116.390 110.630 ;
        RECT 105.760 107.200 105.930 110.460 ;
        RECT 106.655 109.890 114.695 110.060 ;
        RECT 106.270 107.830 106.440 109.830 ;
        RECT 114.910 107.830 115.080 109.830 ;
        RECT 106.655 107.600 114.695 107.770 ;
        RECT 115.420 107.200 116.390 110.460 ;
        RECT 105.760 107.030 116.390 107.200 ;
        RECT 105.760 103.770 105.930 107.030 ;
        RECT 106.655 106.460 114.695 106.630 ;
        RECT 106.270 104.400 106.440 106.400 ;
        RECT 114.910 104.400 115.080 106.400 ;
        RECT 106.655 104.170 114.695 104.340 ;
        RECT 115.420 103.770 116.390 107.030 ;
        RECT 97.940 103.650 104.180 103.750 ;
        RECT 97.930 103.090 104.180 103.650 ;
        RECT 97.930 103.070 103.100 103.090 ;
        RECT 97.930 103.000 101.920 103.070 ;
        RECT 97.930 101.730 99.850 103.000 ;
        RECT 101.360 102.990 101.920 103.000 ;
        RECT 101.590 101.900 101.920 102.990 ;
        RECT 102.290 102.520 103.330 102.690 ;
        RECT 102.290 102.080 103.330 102.250 ;
        RECT 103.500 102.220 103.670 102.550 ;
        RECT 97.940 98.540 98.880 101.730 ;
        RECT 101.750 101.680 101.920 101.900 ;
        RECT 104.010 101.680 104.180 103.090 ;
        RECT 101.750 101.510 104.180 101.680 ;
        RECT 105.760 103.600 116.390 103.770 ;
        RECT 116.930 112.860 123.160 113.020 ;
        RECT 116.930 110.600 117.600 112.860 ;
        RECT 118.270 112.290 122.310 112.460 ;
        RECT 117.930 111.230 118.100 112.230 ;
        RECT 122.480 111.230 122.650 112.230 ;
        RECT 118.270 111.000 122.310 111.170 ;
        RECT 122.990 110.600 123.160 112.860 ;
        RECT 116.930 110.430 123.160 110.600 ;
        RECT 116.930 107.170 117.600 110.430 ;
        RECT 118.270 109.860 122.310 110.030 ;
        RECT 117.930 107.800 118.100 109.800 ;
        RECT 122.480 107.800 122.650 109.800 ;
        RECT 118.270 107.570 122.310 107.740 ;
        RECT 122.990 107.170 123.160 110.430 ;
        RECT 116.930 107.000 123.160 107.170 ;
        RECT 116.930 103.740 117.600 107.000 ;
        RECT 118.270 106.430 122.310 106.600 ;
        RECT 117.930 104.370 118.100 106.370 ;
        RECT 122.480 104.370 122.650 106.370 ;
        RECT 118.270 104.140 122.310 104.310 ;
        RECT 122.990 103.740 123.160 107.000 ;
        RECT 116.930 103.730 123.160 103.740 ;
        RECT 124.750 113.000 134.580 113.040 ;
        RECT 136.470 113.020 142.210 113.030 ;
        RECT 124.750 112.870 135.380 113.000 ;
        RECT 124.750 110.610 124.920 112.870 ;
        RECT 125.645 112.300 133.685 112.470 ;
        RECT 125.260 111.240 125.430 112.240 ;
        RECT 133.900 111.240 134.070 112.240 ;
        RECT 125.645 111.010 133.685 111.180 ;
        RECT 134.410 110.610 135.380 112.870 ;
        RECT 124.750 110.440 135.380 110.610 ;
        RECT 124.750 107.180 124.920 110.440 ;
        RECT 125.645 109.870 133.685 110.040 ;
        RECT 125.260 107.810 125.430 109.810 ;
        RECT 133.900 107.810 134.070 109.810 ;
        RECT 125.645 107.580 133.685 107.750 ;
        RECT 134.410 107.180 135.380 110.440 ;
        RECT 124.750 107.010 135.380 107.180 ;
        RECT 124.750 103.750 124.920 107.010 ;
        RECT 125.645 106.440 133.685 106.610 ;
        RECT 125.260 104.380 125.430 106.380 ;
        RECT 133.900 104.380 134.070 106.380 ;
        RECT 125.645 104.150 133.685 104.320 ;
        RECT 134.410 103.750 135.380 107.010 ;
        RECT 116.930 103.630 123.170 103.730 ;
        RECT 105.760 101.340 105.930 103.600 ;
        RECT 106.655 103.030 114.695 103.200 ;
        RECT 106.270 101.970 106.440 102.970 ;
        RECT 114.910 101.970 115.080 102.970 ;
        RECT 106.655 101.740 114.695 101.910 ;
        RECT 115.420 101.340 116.390 103.600 ;
        RECT 116.920 103.070 123.170 103.630 ;
        RECT 116.920 103.050 122.090 103.070 ;
        RECT 116.920 102.980 120.910 103.050 ;
        RECT 116.920 101.710 118.840 102.980 ;
        RECT 120.350 102.970 120.910 102.980 ;
        RECT 120.580 101.880 120.910 102.970 ;
        RECT 121.280 102.500 122.320 102.670 ;
        RECT 121.280 102.060 122.320 102.230 ;
        RECT 122.490 102.200 122.660 102.530 ;
        RECT 120.740 101.660 120.910 101.880 ;
        RECT 123.000 101.660 123.170 103.070 ;
        RECT 120.740 101.490 123.170 101.660 ;
        RECT 124.750 103.580 135.380 103.750 ;
        RECT 135.980 112.860 142.210 113.020 ;
        RECT 135.980 110.600 136.650 112.860 ;
        RECT 137.320 112.290 141.360 112.460 ;
        RECT 136.980 111.230 137.150 112.230 ;
        RECT 141.530 111.230 141.700 112.230 ;
        RECT 137.320 111.000 141.360 111.170 ;
        RECT 142.040 110.600 142.210 112.860 ;
        RECT 135.980 110.430 142.210 110.600 ;
        RECT 135.980 107.170 136.650 110.430 ;
        RECT 137.320 109.860 141.360 110.030 ;
        RECT 136.980 107.800 137.150 109.800 ;
        RECT 141.530 107.800 141.700 109.800 ;
        RECT 137.320 107.570 141.360 107.740 ;
        RECT 142.040 107.170 142.210 110.430 ;
        RECT 135.980 107.000 142.210 107.170 ;
        RECT 135.980 103.740 136.650 107.000 ;
        RECT 137.320 106.430 141.360 106.600 ;
        RECT 136.980 104.370 137.150 106.370 ;
        RECT 141.530 104.370 141.700 106.370 ;
        RECT 137.320 104.140 141.360 104.310 ;
        RECT 142.040 103.740 142.210 107.000 ;
        RECT 135.980 103.730 142.210 103.740 ;
        RECT 143.800 113.000 153.630 113.040 ;
        RECT 143.800 112.870 154.430 113.000 ;
        RECT 143.800 110.610 143.970 112.870 ;
        RECT 144.695 112.300 152.735 112.470 ;
        RECT 144.310 111.240 144.480 112.240 ;
        RECT 152.950 111.240 153.120 112.240 ;
        RECT 144.695 111.010 152.735 111.180 ;
        RECT 153.460 110.610 154.430 112.870 ;
        RECT 143.800 110.440 154.430 110.610 ;
        RECT 143.800 107.180 143.970 110.440 ;
        RECT 144.695 109.870 152.735 110.040 ;
        RECT 144.310 107.810 144.480 109.810 ;
        RECT 152.950 107.810 153.120 109.810 ;
        RECT 144.695 107.580 152.735 107.750 ;
        RECT 153.460 107.180 154.430 110.440 ;
        RECT 143.800 107.010 154.430 107.180 ;
        RECT 143.800 103.750 143.970 107.010 ;
        RECT 144.695 106.440 152.735 106.610 ;
        RECT 144.310 104.380 144.480 106.380 ;
        RECT 152.950 104.380 153.120 106.380 ;
        RECT 144.695 104.150 152.735 104.320 ;
        RECT 153.460 103.750 154.430 107.010 ;
        RECT 135.980 103.630 142.220 103.730 ;
        RECT 105.760 101.310 116.390 101.340 ;
        RECT 105.730 101.200 116.390 101.310 ;
        RECT 124.750 101.320 124.920 103.580 ;
        RECT 125.645 103.010 133.685 103.180 ;
        RECT 125.260 101.950 125.430 102.950 ;
        RECT 133.900 101.950 134.070 102.950 ;
        RECT 125.645 101.720 133.685 101.890 ;
        RECT 134.410 101.320 135.380 103.580 ;
        RECT 135.970 103.070 142.220 103.630 ;
        RECT 135.970 103.050 141.140 103.070 ;
        RECT 135.970 102.980 139.960 103.050 ;
        RECT 135.970 101.710 137.890 102.980 ;
        RECT 139.400 102.970 139.960 102.980 ;
        RECT 139.630 101.880 139.960 102.970 ;
        RECT 140.330 102.500 141.370 102.670 ;
        RECT 140.330 102.060 141.370 102.230 ;
        RECT 141.540 102.200 141.710 102.530 ;
        RECT 139.790 101.660 139.960 101.880 ;
        RECT 142.050 101.660 142.220 103.070 ;
        RECT 139.790 101.490 142.220 101.660 ;
        RECT 143.800 103.580 154.430 103.750 ;
        RECT 124.750 101.290 135.380 101.320 ;
        RECT 143.800 101.320 143.970 103.580 ;
        RECT 144.695 103.010 152.735 103.180 ;
        RECT 144.310 101.950 144.480 102.950 ;
        RECT 152.950 101.950 153.120 102.950 ;
        RECT 144.695 101.720 152.735 101.890 ;
        RECT 153.460 101.320 154.430 103.580 ;
        RECT 143.800 101.290 154.430 101.320 ;
        RECT 103.980 101.150 116.390 101.200 ;
        RECT 124.720 101.180 135.380 101.290 ;
        RECT 143.770 101.180 154.430 101.290 ;
        RECT 99.640 100.980 116.390 101.150 ;
        RECT 122.970 101.130 135.380 101.180 ;
        RECT 142.020 101.130 154.430 101.180 ;
        RECT 99.640 99.570 99.810 100.980 ;
        RECT 100.180 100.410 103.220 100.580 ;
        RECT 100.180 99.970 103.220 100.140 ;
        RECT 103.435 100.110 103.605 100.440 ;
        RECT 103.940 100.220 116.390 100.980 ;
        RECT 118.630 100.960 135.380 101.130 ;
        RECT 103.940 100.210 116.280 100.220 ;
        RECT 103.940 100.200 109.820 100.210 ;
        RECT 103.940 100.180 104.510 100.200 ;
        RECT 105.730 100.190 109.820 100.200 ;
        RECT 103.950 99.570 104.120 100.180 ;
        RECT 99.640 99.400 104.120 99.570 ;
        RECT 118.630 99.550 118.800 100.960 ;
        RECT 119.170 100.390 122.210 100.560 ;
        RECT 119.170 99.950 122.210 100.120 ;
        RECT 122.425 100.090 122.595 100.420 ;
        RECT 122.930 100.200 135.380 100.960 ;
        RECT 137.680 100.960 154.430 101.130 ;
        RECT 122.930 100.190 135.270 100.200 ;
        RECT 122.930 100.180 128.810 100.190 ;
        RECT 122.930 100.160 123.500 100.180 ;
        RECT 124.720 100.170 128.810 100.180 ;
        RECT 122.940 99.550 123.110 100.160 ;
        RECT 118.630 99.380 123.110 99.550 ;
        RECT 137.680 99.550 137.850 100.960 ;
        RECT 138.220 100.390 141.260 100.560 ;
        RECT 138.220 99.950 141.260 100.120 ;
        RECT 141.475 100.090 141.645 100.420 ;
        RECT 141.980 100.200 154.430 100.960 ;
        RECT 141.980 100.190 154.320 100.200 ;
        RECT 141.980 100.180 147.860 100.190 ;
        RECT 141.980 100.160 142.550 100.180 ;
        RECT 143.770 100.170 147.860 100.180 ;
        RECT 141.990 99.550 142.160 100.160 ;
        RECT 137.680 99.380 142.160 99.550 ;
        RECT 97.890 98.510 100.320 98.540 ;
        RECT 97.890 98.340 154.230 98.510 ;
        RECT 97.890 97.030 100.320 98.340 ;
        RECT 100.800 97.510 102.960 97.860 ;
        RECT 103.500 97.510 105.660 97.860 ;
        RECT 106.140 97.030 106.310 98.340 ;
        RECT 106.790 97.510 108.950 97.860 ;
        RECT 109.490 97.510 111.650 97.860 ;
        RECT 112.130 97.030 112.300 98.340 ;
        RECT 112.780 97.510 114.940 97.860 ;
        RECT 115.480 97.510 117.640 97.860 ;
        RECT 118.120 97.030 118.290 98.340 ;
        RECT 118.770 97.510 120.930 97.860 ;
        RECT 121.470 97.510 123.630 97.860 ;
        RECT 124.110 97.030 124.280 98.340 ;
        RECT 124.760 97.510 126.920 97.860 ;
        RECT 127.460 97.510 129.620 97.860 ;
        RECT 130.100 97.030 130.270 98.340 ;
        RECT 130.750 97.510 132.910 97.860 ;
        RECT 133.450 97.510 135.610 97.860 ;
        RECT 136.090 97.030 136.260 98.340 ;
        RECT 136.740 97.510 138.900 97.860 ;
        RECT 139.440 97.510 141.600 97.860 ;
        RECT 142.080 97.030 142.250 98.340 ;
        RECT 142.730 97.510 144.890 97.860 ;
        RECT 145.430 97.510 147.590 97.860 ;
        RECT 148.070 97.030 148.240 98.340 ;
        RECT 148.720 97.510 150.880 97.860 ;
        RECT 151.420 97.510 153.580 97.860 ;
        RECT 154.060 97.030 154.230 98.340 ;
        RECT 97.890 96.860 154.230 97.030 ;
        RECT 97.890 95.550 100.320 96.860 ;
        RECT 100.800 96.030 102.960 96.380 ;
        RECT 103.500 96.030 105.660 96.380 ;
        RECT 106.140 95.550 106.310 96.860 ;
        RECT 106.790 96.030 108.950 96.380 ;
        RECT 109.490 96.030 111.650 96.380 ;
        RECT 112.130 95.550 112.300 96.860 ;
        RECT 112.780 96.030 114.940 96.380 ;
        RECT 115.480 96.030 117.640 96.380 ;
        RECT 118.120 95.550 118.290 96.860 ;
        RECT 118.770 96.030 120.930 96.380 ;
        RECT 121.470 96.030 123.630 96.380 ;
        RECT 124.110 95.550 124.280 96.860 ;
        RECT 124.760 96.030 126.920 96.380 ;
        RECT 127.460 96.030 129.620 96.380 ;
        RECT 130.100 95.550 130.270 96.860 ;
        RECT 130.750 96.030 132.910 96.380 ;
        RECT 133.450 96.030 135.610 96.380 ;
        RECT 136.090 95.550 136.260 96.860 ;
        RECT 136.740 96.030 138.900 96.380 ;
        RECT 139.440 96.030 141.600 96.380 ;
        RECT 142.080 95.550 142.250 96.860 ;
        RECT 97.890 95.410 142.250 95.550 ;
        RECT 100.150 95.380 142.250 95.410 ;
      LAYER met1 ;
        RECT 145.380 221.200 145.700 221.460 ;
        RECT 144.980 220.260 145.240 220.580 ;
        RECT 111.400 218.730 111.660 219.050 ;
        RECT 144.360 218.920 144.620 219.240 ;
        RECT 105.460 205.520 105.720 205.840 ;
        RECT 105.520 191.010 105.660 205.520 ;
        RECT 106.150 205.120 106.470 205.180 ;
        RECT 106.150 204.920 106.540 205.120 ;
        RECT 106.400 197.030 106.540 204.920 ;
        RECT 106.760 204.060 107.020 204.370 ;
        RECT 106.760 204.050 107.130 204.060 ;
        RECT 106.820 203.920 107.130 204.050 ;
        RECT 106.990 201.080 107.130 203.920 ;
        RECT 106.900 200.820 107.220 201.080 ;
        RECT 106.300 196.640 106.700 197.030 ;
        RECT 105.390 190.620 105.790 191.010 ;
        RECT 107.720 181.860 108.200 217.740 ;
        RECT 109.020 206.310 109.280 206.630 ;
        RECT 108.355 205.405 108.585 205.695 ;
        RECT 108.400 203.870 108.540 205.405 ;
        RECT 108.340 203.550 108.600 203.870 ;
        RECT 108.355 203.105 108.585 203.395 ;
        RECT 108.400 201.110 108.540 203.105 ;
        RECT 109.035 202.400 109.265 202.475 ;
        RECT 109.035 202.260 110.240 202.400 ;
        RECT 109.035 202.185 109.265 202.260 ;
        RECT 109.035 201.725 109.265 202.015 ;
        RECT 109.080 201.570 109.220 201.725 ;
        RECT 109.020 201.250 109.280 201.570 ;
        RECT 109.715 201.240 109.945 201.530 ;
        RECT 108.340 200.790 108.600 201.110 ;
        RECT 109.375 200.845 109.605 201.135 ;
        RECT 108.695 200.390 108.925 200.680 ;
        RECT 108.740 199.270 108.880 200.390 ;
        RECT 109.420 199.945 109.560 200.845 ;
        RECT 109.375 199.655 109.605 199.945 ;
        RECT 108.680 198.950 108.940 199.270 ;
        RECT 109.420 197.425 109.560 199.655 ;
        RECT 109.760 199.430 109.900 201.240 ;
        RECT 109.715 199.140 109.945 199.430 ;
        RECT 109.760 197.860 109.900 199.140 ;
        RECT 109.715 197.570 109.945 197.860 ;
        RECT 109.375 197.135 109.605 197.425 ;
        RECT 108.340 196.880 108.600 196.970 ;
        RECT 108.340 196.740 108.880 196.880 ;
        RECT 108.340 196.650 108.600 196.740 ;
        RECT 108.355 194.120 108.585 194.195 ;
        RECT 108.740 194.120 108.880 196.740 ;
        RECT 110.100 196.510 110.240 202.260 ;
        RECT 110.040 196.190 110.300 196.510 ;
        RECT 109.715 194.825 109.945 195.115 ;
        RECT 108.355 193.980 108.880 194.120 ;
        RECT 108.355 193.905 108.585 193.980 ;
        RECT 109.760 193.290 109.900 194.825 ;
        RECT 109.020 192.970 109.280 193.290 ;
        RECT 109.700 192.970 109.960 193.290 ;
        RECT 108.340 190.670 108.600 190.990 ;
        RECT 108.400 189.595 108.540 190.670 ;
        RECT 109.020 190.210 109.280 190.530 ;
        RECT 108.355 189.305 108.585 189.595 ;
        RECT 110.055 188.385 110.285 188.675 ;
        RECT 109.360 187.910 109.620 188.230 ;
        RECT 109.020 187.450 109.280 187.770 ;
        RECT 109.420 186.375 109.560 187.910 ;
        RECT 109.700 186.990 109.960 187.310 ;
        RECT 109.375 186.085 109.605 186.375 ;
        RECT 109.760 184.995 109.900 186.990 ;
        RECT 110.100 186.850 110.240 188.385 ;
        RECT 110.040 186.530 110.300 186.850 ;
        RECT 109.715 184.705 109.945 184.995 ;
        RECT 110.040 184.230 110.300 184.550 ;
        RECT 110.100 184.075 110.240 184.230 ;
        RECT 110.055 183.785 110.285 184.075 ;
        RECT 110.440 181.860 110.920 217.740 ;
        RECT 111.460 215.815 111.600 218.730 ;
        RECT 143.850 217.960 144.110 218.280 ;
        RECT 112.080 215.970 112.340 216.290 ;
        RECT 111.415 215.525 111.645 215.815 ;
        RECT 112.140 214.895 112.280 215.970 ;
        RECT 112.095 214.605 112.325 214.895 ;
        RECT 112.760 213.210 113.020 213.530 ;
        RECT 112.760 211.370 113.020 211.690 ;
        RECT 112.760 210.910 113.020 211.230 ;
        RECT 111.755 210.005 111.985 210.295 ;
        RECT 111.800 204.790 111.940 210.005 ;
        RECT 112.760 208.610 113.020 208.930 ;
        RECT 112.820 206.630 112.960 208.610 ;
        RECT 112.760 206.310 113.020 206.630 ;
        RECT 111.740 204.470 112.000 204.790 ;
        RECT 112.820 204.315 112.960 206.310 ;
        RECT 112.775 204.025 113.005 204.315 ;
        RECT 111.755 201.715 111.985 202.005 ;
        RECT 111.415 201.280 111.645 201.570 ;
        RECT 111.460 200.000 111.600 201.280 ;
        RECT 111.415 199.710 111.645 200.000 ;
        RECT 111.060 198.950 111.320 199.270 ;
        RECT 111.120 196.955 111.260 198.950 ;
        RECT 111.460 197.900 111.600 199.710 ;
        RECT 111.800 199.485 111.940 201.715 ;
        RECT 112.760 200.100 113.020 200.190 ;
        RECT 112.140 199.960 113.020 200.100 ;
        RECT 111.755 199.195 111.985 199.485 ;
        RECT 111.800 198.295 111.940 199.195 ;
        RECT 112.140 198.750 112.280 199.960 ;
        RECT 112.760 199.870 113.020 199.960 ;
        RECT 112.420 198.950 112.680 199.270 ;
        RECT 112.095 198.460 112.325 198.750 ;
        RECT 111.755 198.005 111.985 198.295 ;
        RECT 111.415 197.610 111.645 197.900 ;
        RECT 112.095 197.340 112.325 197.415 ;
        RECT 112.480 197.340 112.620 198.950 ;
        RECT 112.095 197.200 112.620 197.340 ;
        RECT 112.095 197.125 112.325 197.200 ;
        RECT 111.075 196.665 111.305 196.955 ;
        RECT 112.095 194.825 112.325 195.115 ;
        RECT 111.740 193.430 112.000 193.750 ;
        RECT 111.740 192.970 112.000 193.290 ;
        RECT 111.800 188.675 111.940 192.970 ;
        RECT 112.140 191.435 112.280 194.825 ;
        RECT 112.760 194.350 113.020 194.670 ;
        RECT 112.095 191.145 112.325 191.435 ;
        RECT 111.755 188.385 111.985 188.675 ;
        RECT 111.740 187.910 112.000 188.230 ;
        RECT 111.800 186.835 111.940 187.910 ;
        RECT 112.080 187.450 112.340 187.770 ;
        RECT 111.755 186.545 111.985 186.835 ;
        RECT 111.755 186.085 111.985 186.375 ;
        RECT 111.800 183.630 111.940 186.085 ;
        RECT 112.140 185.455 112.280 187.450 ;
        RECT 112.095 185.165 112.325 185.455 ;
        RECT 112.760 184.690 113.020 185.010 ;
        RECT 112.820 184.535 112.960 184.690 ;
        RECT 112.775 184.245 113.005 184.535 ;
        RECT 111.740 183.310 112.000 183.630 ;
        RECT 113.160 181.860 113.640 217.740 ;
        RECT 115.480 215.970 115.740 216.290 ;
        RECT 114.815 213.675 115.045 213.965 ;
        RECT 114.120 213.210 114.380 213.530 ;
        RECT 114.180 210.710 114.320 213.210 ;
        RECT 114.860 211.445 115.000 213.675 ;
        RECT 115.155 213.240 115.385 213.530 ;
        RECT 115.200 211.960 115.340 213.240 ;
        RECT 115.155 211.670 115.385 211.960 ;
        RECT 114.815 211.155 115.045 211.445 ;
        RECT 114.135 210.420 114.365 210.710 ;
        RECT 114.860 210.255 115.000 211.155 ;
        RECT 114.815 209.965 115.045 210.255 ;
        RECT 115.200 209.860 115.340 211.670 ;
        RECT 115.155 209.570 115.385 209.860 ;
        RECT 114.800 209.070 115.060 209.390 ;
        RECT 114.475 204.025 114.705 204.315 ;
        RECT 114.520 199.730 114.660 204.025 ;
        RECT 114.460 199.410 114.720 199.730 ;
        RECT 115.480 198.950 115.740 199.270 ;
        RECT 115.540 197.875 115.680 198.950 ;
        RECT 115.495 197.585 115.725 197.875 ;
        RECT 114.475 193.660 114.705 193.735 ;
        RECT 114.475 193.520 115.000 193.660 ;
        RECT 114.475 193.445 114.705 193.520 ;
        RECT 114.460 192.050 114.720 192.370 ;
        RECT 113.795 191.360 114.025 191.435 ;
        RECT 113.795 191.220 114.320 191.360 ;
        RECT 113.795 191.145 114.025 191.220 ;
        RECT 113.795 188.385 114.025 188.675 ;
        RECT 113.840 188.230 113.980 188.385 ;
        RECT 113.780 187.910 114.040 188.230 ;
        RECT 114.180 188.140 114.320 191.220 ;
        RECT 114.460 190.670 114.720 190.990 ;
        RECT 114.460 189.290 114.720 189.610 ;
        RECT 114.475 188.140 114.705 188.215 ;
        RECT 114.180 188.000 114.705 188.140 ;
        RECT 113.780 187.450 114.040 187.770 ;
        RECT 114.180 185.840 114.320 188.000 ;
        RECT 114.475 187.925 114.705 188.000 ;
        RECT 114.475 187.005 114.705 187.295 ;
        RECT 114.520 186.850 114.660 187.005 ;
        RECT 114.460 186.530 114.720 186.850 ;
        RECT 114.460 185.840 114.720 185.930 ;
        RECT 114.180 185.700 114.720 185.840 ;
        RECT 114.460 185.610 114.720 185.700 ;
        RECT 114.460 184.230 114.720 184.550 ;
        RECT 114.860 184.090 115.000 193.520 ;
        RECT 115.155 192.525 115.385 192.815 ;
        RECT 115.200 187.310 115.340 192.525 ;
        RECT 115.495 189.765 115.725 190.055 ;
        RECT 115.540 187.770 115.680 189.765 ;
        RECT 115.480 187.450 115.740 187.770 ;
        RECT 115.140 186.990 115.400 187.310 ;
        RECT 115.495 186.545 115.725 186.835 ;
        RECT 115.540 186.390 115.680 186.545 ;
        RECT 115.480 186.070 115.740 186.390 ;
        RECT 114.800 183.770 115.060 184.090 ;
        RECT 114.460 183.310 114.720 183.630 ;
        RECT 115.880 181.860 116.360 217.740 ;
        RECT 116.840 216.430 117.100 216.750 ;
        RECT 116.900 215.815 117.040 216.430 ;
        RECT 117.180 215.970 117.440 216.290 ;
        RECT 116.855 215.525 117.085 215.815 ;
        RECT 117.240 213.515 117.380 215.970 ;
        RECT 117.535 214.605 117.765 214.895 ;
        RECT 117.195 213.225 117.425 213.515 ;
        RECT 116.500 211.370 116.760 211.690 ;
        RECT 116.560 210.295 116.700 211.370 ;
        RECT 116.840 210.910 117.100 211.230 ;
        RECT 116.515 210.005 116.745 210.295 ;
        RECT 116.515 201.265 116.745 201.555 ;
        RECT 116.560 200.190 116.700 201.265 ;
        RECT 116.500 199.870 116.760 200.190 ;
        RECT 116.900 199.180 117.040 210.910 ;
        RECT 117.180 208.610 117.440 208.930 ;
        RECT 117.580 208.470 117.720 214.605 ;
        RECT 117.520 208.150 117.780 208.470 ;
        RECT 117.535 205.405 117.765 205.695 ;
        RECT 117.180 204.470 117.440 204.790 ;
        RECT 117.195 203.565 117.425 203.855 ;
        RECT 117.240 199.640 117.380 203.565 ;
        RECT 117.580 203.395 117.720 205.405 ;
        RECT 117.535 203.105 117.765 203.395 ;
        RECT 117.240 199.500 118.060 199.640 ;
        RECT 116.560 199.040 117.040 199.180 ;
        RECT 116.560 192.830 116.700 199.040 ;
        RECT 117.520 198.950 117.780 199.270 ;
        RECT 116.855 198.480 117.085 198.770 ;
        RECT 116.900 196.670 117.040 198.480 ;
        RECT 117.195 198.085 117.425 198.375 ;
        RECT 117.240 197.185 117.380 198.085 ;
        RECT 117.535 197.630 117.765 197.920 ;
        RECT 117.195 196.895 117.425 197.185 ;
        RECT 116.855 196.380 117.085 196.670 ;
        RECT 116.900 195.100 117.040 196.380 ;
        RECT 116.855 194.810 117.085 195.100 ;
        RECT 117.240 194.665 117.380 196.895 ;
        RECT 117.195 194.375 117.425 194.665 ;
        RECT 117.580 194.120 117.720 197.630 ;
        RECT 117.920 194.670 118.060 199.500 ;
        RECT 117.860 194.350 118.120 194.670 ;
        RECT 116.900 193.980 117.720 194.120 ;
        RECT 116.500 192.510 116.760 192.830 ;
        RECT 116.515 192.065 116.745 192.355 ;
        RECT 116.560 190.530 116.700 192.065 ;
        RECT 116.900 191.435 117.040 193.980 ;
        RECT 117.520 193.430 117.780 193.750 ;
        RECT 117.180 192.510 117.440 192.830 ;
        RECT 116.855 191.145 117.085 191.435 ;
        RECT 116.500 190.210 116.760 190.530 ;
        RECT 117.240 189.135 117.380 192.510 ;
        RECT 117.195 188.845 117.425 189.135 ;
        RECT 117.195 188.600 117.425 188.675 ;
        RECT 117.580 188.600 117.720 193.430 ;
        RECT 118.200 189.290 118.460 189.610 ;
        RECT 117.195 188.460 117.720 188.600 ;
        RECT 117.195 188.385 117.425 188.460 ;
        RECT 117.180 187.450 117.440 187.770 ;
        RECT 116.500 186.530 116.760 186.850 ;
        RECT 116.560 184.995 116.700 186.530 ;
        RECT 116.855 186.085 117.085 186.375 ;
        RECT 116.515 184.705 116.745 184.995 ;
        RECT 116.900 183.630 117.040 186.085 ;
        RECT 117.240 184.550 117.380 187.450 ;
        RECT 117.520 186.990 117.780 187.310 ;
        RECT 117.520 185.610 117.780 185.930 ;
        RECT 118.200 185.610 118.460 185.930 ;
        RECT 117.580 184.995 117.720 185.610 ;
        RECT 117.860 185.150 118.120 185.470 ;
        RECT 117.535 184.705 117.765 184.995 ;
        RECT 117.180 184.230 117.440 184.550 ;
        RECT 116.840 183.310 117.100 183.630 ;
        RECT 117.920 183.615 118.060 185.150 ;
        RECT 117.875 183.325 118.105 183.615 ;
        RECT 118.600 181.860 119.080 217.740 ;
        RECT 120.240 216.200 120.500 216.290 ;
        RECT 119.960 216.060 120.500 216.200 ;
        RECT 119.575 214.650 119.805 214.940 ;
        RECT 119.620 213.990 119.760 214.650 ;
        RECT 119.560 213.670 119.820 213.990 ;
        RECT 119.960 209.390 120.100 216.060 ;
        RECT 120.240 215.970 120.500 216.060 ;
        RECT 120.595 215.500 120.825 215.790 ;
        RECT 120.255 215.105 120.485 215.395 ;
        RECT 120.300 214.205 120.440 215.105 ;
        RECT 120.255 213.915 120.485 214.205 ;
        RECT 120.300 211.685 120.440 213.915 ;
        RECT 120.640 213.690 120.780 215.500 ;
        RECT 120.595 213.400 120.825 213.690 ;
        RECT 120.640 212.120 120.780 213.400 ;
        RECT 120.595 211.830 120.825 212.120 ;
        RECT 120.255 211.395 120.485 211.685 ;
        RECT 119.900 209.070 120.160 209.390 ;
        RECT 120.935 209.085 121.165 209.375 ;
        RECT 119.960 204.315 120.100 209.070 ;
        RECT 120.980 208.470 121.120 209.085 ;
        RECT 120.920 208.150 121.180 208.470 ;
        RECT 119.915 204.240 120.145 204.315 ;
        RECT 119.280 204.100 120.145 204.240 ;
        RECT 119.280 199.270 119.420 204.100 ;
        RECT 119.915 204.025 120.145 204.100 ;
        RECT 120.595 203.540 120.825 203.830 ;
        RECT 119.560 203.090 119.820 203.410 ;
        RECT 120.255 203.145 120.485 203.435 ;
        RECT 119.620 202.860 119.760 203.090 ;
        RECT 119.915 202.860 120.145 202.980 ;
        RECT 119.620 202.720 120.145 202.860 ;
        RECT 119.915 202.690 120.145 202.720 ;
        RECT 120.300 202.245 120.440 203.145 ;
        RECT 120.255 201.955 120.485 202.245 ;
        RECT 120.300 199.725 120.440 201.955 ;
        RECT 120.640 201.730 120.780 203.540 ;
        RECT 120.595 201.440 120.825 201.730 ;
        RECT 120.640 200.160 120.780 201.440 ;
        RECT 120.595 199.870 120.825 200.160 ;
        RECT 120.255 199.435 120.485 199.725 ;
        RECT 119.220 198.950 119.480 199.270 ;
        RECT 119.235 197.125 119.465 197.415 ;
        RECT 119.280 196.510 119.420 197.125 ;
        RECT 120.255 196.665 120.485 196.955 ;
        RECT 119.220 196.190 119.480 196.510 ;
        RECT 120.300 196.050 120.440 196.665 ;
        RECT 120.240 195.730 120.500 196.050 ;
        RECT 120.580 194.810 120.840 195.130 ;
        RECT 120.935 194.365 121.165 194.655 ;
        RECT 120.980 193.750 121.120 194.365 ;
        RECT 120.920 193.430 121.180 193.750 ;
        RECT 119.900 190.210 120.160 190.530 ;
        RECT 119.220 189.290 119.480 189.610 ;
        RECT 119.280 187.295 119.420 189.290 ;
        RECT 120.240 187.910 120.500 188.230 ;
        RECT 119.900 187.450 120.160 187.770 ;
        RECT 119.235 187.005 119.465 187.295 ;
        RECT 119.960 185.915 120.100 187.450 ;
        RECT 119.915 185.625 120.145 185.915 ;
        RECT 119.900 185.150 120.160 185.470 ;
        RECT 119.900 184.690 120.160 185.010 ;
        RECT 119.915 184.460 120.145 184.535 ;
        RECT 120.300 184.460 120.440 187.910 ;
        RECT 120.920 187.450 121.180 187.770 ;
        RECT 120.980 186.835 121.120 187.450 ;
        RECT 120.935 186.545 121.165 186.835 ;
        RECT 119.915 184.320 120.440 184.460 ;
        RECT 119.915 184.245 120.145 184.320 ;
        RECT 121.320 181.860 121.800 217.740 ;
        RECT 123.640 216.430 123.900 216.750 ;
        RECT 122.280 215.970 122.540 216.290 ;
        RECT 122.960 215.970 123.220 216.290 ;
        RECT 121.940 213.670 122.200 213.990 ;
        RECT 122.340 209.760 122.480 215.970 ;
        RECT 123.020 214.895 123.160 215.970 ;
        RECT 123.700 215.815 123.840 216.430 ;
        RECT 123.655 215.525 123.885 215.815 ;
        RECT 122.975 214.605 123.205 214.895 ;
        RECT 123.655 211.845 123.885 212.135 ;
        RECT 122.635 211.385 122.865 211.675 ;
        RECT 122.680 211.230 122.820 211.385 ;
        RECT 123.700 211.230 123.840 211.845 ;
        RECT 122.620 210.910 122.880 211.230 ;
        RECT 123.640 210.910 123.900 211.230 ;
        RECT 122.620 210.450 122.880 210.770 ;
        RECT 122.635 209.760 122.865 209.835 ;
        RECT 122.340 209.620 122.865 209.760 ;
        RECT 122.635 209.545 122.865 209.620 ;
        RECT 122.295 209.060 122.525 209.350 ;
        RECT 122.340 207.250 122.480 209.060 ;
        RECT 122.635 208.665 122.865 208.955 ;
        RECT 122.680 207.765 122.820 208.665 ;
        RECT 123.315 208.210 123.545 208.500 ;
        RECT 122.635 207.475 122.865 207.765 ;
        RECT 122.295 206.960 122.525 207.250 ;
        RECT 122.340 205.680 122.480 206.960 ;
        RECT 122.295 205.390 122.525 205.680 ;
        RECT 122.680 205.245 122.820 207.475 ;
        RECT 122.635 204.955 122.865 205.245 ;
        RECT 123.360 204.790 123.500 208.210 ;
        RECT 123.300 204.470 123.560 204.790 ;
        RECT 123.360 203.410 123.500 204.470 ;
        RECT 122.280 203.090 122.540 203.410 ;
        RECT 123.300 203.090 123.560 203.410 ;
        RECT 122.340 202.475 122.480 203.090 ;
        RECT 123.640 202.630 123.900 202.950 ;
        RECT 122.295 202.185 122.525 202.475 ;
        RECT 122.975 200.345 123.205 200.635 ;
        RECT 122.635 200.100 122.865 200.175 ;
        RECT 122.340 199.960 122.865 200.100 ;
        RECT 122.340 194.670 122.480 199.960 ;
        RECT 122.635 199.885 122.865 199.960 ;
        RECT 122.635 198.965 122.865 199.255 ;
        RECT 122.680 196.970 122.820 198.965 ;
        RECT 123.020 198.335 123.160 200.345 ;
        RECT 122.975 198.045 123.205 198.335 ;
        RECT 122.620 196.650 122.880 196.970 ;
        RECT 122.620 196.190 122.880 196.510 ;
        RECT 122.680 195.575 122.820 196.190 ;
        RECT 123.700 196.050 123.840 202.630 ;
        RECT 123.640 195.730 123.900 196.050 ;
        RECT 122.635 195.285 122.865 195.575 ;
        RECT 122.280 194.350 122.540 194.670 ;
        RECT 122.340 188.675 122.480 194.350 ;
        RECT 122.960 192.050 123.220 192.370 ;
        RECT 123.020 190.975 123.160 192.050 ;
        RECT 122.975 190.685 123.205 190.975 ;
        RECT 122.975 190.440 123.205 190.515 ;
        RECT 122.975 190.300 123.500 190.440 ;
        RECT 122.975 190.225 123.205 190.300 ;
        RECT 122.960 189.750 123.220 190.070 ;
        RECT 122.635 189.305 122.865 189.595 ;
        RECT 122.295 188.385 122.525 188.675 ;
        RECT 122.680 185.930 122.820 189.305 ;
        RECT 123.360 188.230 123.500 190.300 ;
        RECT 123.300 187.910 123.560 188.230 ;
        RECT 122.975 187.005 123.205 187.295 ;
        RECT 123.020 186.850 123.160 187.005 ;
        RECT 122.960 186.530 123.220 186.850 ;
        RECT 122.960 186.070 123.220 186.390 ;
        RECT 123.640 186.070 123.900 186.390 ;
        RECT 122.620 185.610 122.880 185.930 ;
        RECT 122.975 184.705 123.205 184.995 ;
        RECT 123.020 184.550 123.160 184.705 ;
        RECT 122.960 184.230 123.220 184.550 ;
        RECT 123.700 184.075 123.840 186.070 ;
        RECT 123.655 183.785 123.885 184.075 ;
        RECT 124.040 181.860 124.520 217.740 ;
        RECT 125.680 215.970 125.940 216.290 ;
        RECT 125.740 214.895 125.880 215.970 ;
        RECT 125.695 214.605 125.925 214.895 ;
        RECT 126.360 211.370 126.620 211.690 ;
        RECT 124.660 210.910 124.920 211.230 ;
        RECT 125.340 208.150 125.600 208.470 ;
        RECT 125.355 204.240 125.585 204.315 ;
        RECT 125.060 204.100 125.585 204.240 ;
        RECT 125.060 198.795 125.200 204.100 ;
        RECT 125.355 204.025 125.585 204.100 ;
        RECT 125.355 203.320 125.585 203.395 ;
        RECT 125.355 203.180 125.880 203.320 ;
        RECT 125.355 203.105 125.585 203.180 ;
        RECT 125.340 202.630 125.600 202.950 ;
        RECT 125.740 201.940 125.880 203.180 ;
        RECT 126.360 203.090 126.620 203.410 ;
        RECT 126.360 202.630 126.620 202.950 ;
        RECT 126.035 201.940 126.265 202.015 ;
        RECT 125.740 201.800 126.265 201.940 ;
        RECT 126.035 201.725 126.265 201.800 ;
        RECT 125.695 201.265 125.925 201.555 ;
        RECT 125.355 200.345 125.585 200.635 ;
        RECT 125.400 200.190 125.540 200.345 ;
        RECT 125.340 199.870 125.600 200.190 ;
        RECT 125.340 198.950 125.600 199.270 ;
        RECT 125.015 198.505 125.245 198.795 ;
        RECT 125.740 195.960 125.880 201.265 ;
        RECT 126.080 198.810 126.220 201.725 ;
        RECT 126.420 201.095 126.560 202.630 ;
        RECT 126.375 200.805 126.605 201.095 ;
        RECT 126.020 198.490 126.280 198.810 ;
        RECT 125.740 195.820 126.220 195.960 ;
        RECT 125.680 195.270 125.940 195.590 ;
        RECT 126.080 194.670 126.220 195.820 ;
        RECT 126.020 194.350 126.280 194.670 ;
        RECT 124.675 193.445 124.905 193.735 ;
        RECT 124.720 192.830 124.860 193.445 ;
        RECT 124.660 192.510 124.920 192.830 ;
        RECT 125.355 192.740 125.585 192.815 ;
        RECT 125.355 192.600 125.880 192.740 ;
        RECT 125.355 192.525 125.585 192.600 ;
        RECT 125.355 191.605 125.585 191.895 ;
        RECT 125.015 190.225 125.245 190.515 ;
        RECT 124.660 189.750 124.920 190.070 ;
        RECT 124.720 189.595 124.860 189.750 ;
        RECT 124.675 189.305 124.905 189.595 ;
        RECT 125.060 188.230 125.200 190.225 ;
        RECT 125.400 190.055 125.540 191.605 ;
        RECT 125.355 189.765 125.585 190.055 ;
        RECT 125.400 189.610 125.540 189.765 ;
        RECT 125.340 189.290 125.600 189.610 ;
        RECT 125.355 189.060 125.585 189.135 ;
        RECT 125.740 189.060 125.880 192.600 ;
        RECT 126.360 192.050 126.620 192.370 ;
        RECT 125.355 188.920 125.880 189.060 ;
        RECT 125.355 188.845 125.585 188.920 ;
        RECT 125.340 188.370 125.600 188.690 ;
        RECT 125.000 187.910 125.260 188.230 ;
        RECT 124.675 187.680 124.905 187.755 ;
        RECT 124.675 187.540 125.200 187.680 ;
        RECT 124.675 187.465 124.905 187.540 ;
        RECT 125.060 187.220 125.200 187.540 ;
        RECT 125.355 187.220 125.585 187.295 ;
        RECT 125.060 187.080 125.585 187.220 ;
        RECT 125.060 185.470 125.200 187.080 ;
        RECT 125.355 187.005 125.585 187.080 ;
        RECT 125.340 186.070 125.600 186.390 ;
        RECT 125.740 186.300 125.880 188.920 ;
        RECT 126.020 186.300 126.280 186.390 ;
        RECT 125.740 186.160 126.280 186.300 ;
        RECT 126.020 186.070 126.280 186.160 ;
        RECT 125.340 185.610 125.600 185.930 ;
        RECT 125.000 185.150 125.260 185.470 ;
        RECT 125.400 184.995 125.540 185.610 ;
        RECT 125.355 184.705 125.585 184.995 ;
        RECT 126.360 184.690 126.620 185.010 ;
        RECT 126.420 184.075 126.560 184.690 ;
        RECT 126.375 183.785 126.605 184.075 ;
        RECT 126.760 181.860 127.240 217.740 ;
        RECT 127.380 215.970 127.640 216.290 ;
        RECT 128.740 215.970 129.000 216.290 ;
        RECT 128.075 213.675 128.305 213.965 ;
        RECT 127.735 213.240 127.965 213.530 ;
        RECT 127.780 211.960 127.920 213.240 ;
        RECT 127.735 211.670 127.965 211.960 ;
        RECT 127.780 209.860 127.920 211.670 ;
        RECT 128.120 211.445 128.260 213.675 ;
        RECT 128.075 211.155 128.305 211.445 ;
        RECT 128.120 210.255 128.260 211.155 ;
        RECT 128.800 210.710 128.940 215.970 ;
        RECT 128.755 210.420 128.985 210.710 ;
        RECT 128.075 209.965 128.305 210.255 ;
        RECT 127.735 209.570 127.965 209.860 ;
        RECT 128.400 209.070 128.660 209.390 ;
        RECT 128.740 205.390 129.000 205.710 ;
        RECT 127.380 199.410 127.640 199.730 ;
        RECT 127.440 199.255 127.580 199.410 ;
        RECT 127.395 198.965 127.625 199.255 ;
        RECT 128.060 198.950 128.320 199.270 ;
        RECT 127.380 194.350 127.640 194.670 ;
        RECT 127.440 191.435 127.580 194.350 ;
        RECT 128.120 193.735 128.260 198.950 ;
        RECT 129.080 196.190 129.340 196.510 ;
        RECT 129.080 193.890 129.340 194.210 ;
        RECT 128.075 193.445 128.305 193.735 ;
        RECT 127.395 191.145 127.625 191.435 ;
        RECT 128.400 191.130 128.660 191.450 ;
        RECT 128.400 190.210 128.660 190.530 ;
        RECT 129.140 189.595 129.280 193.890 ;
        RECT 129.095 189.305 129.325 189.595 ;
        RECT 127.380 187.910 127.640 188.230 ;
        RECT 127.440 184.995 127.580 187.910 ;
        RECT 128.400 185.840 128.660 185.930 ;
        RECT 128.400 185.700 128.940 185.840 ;
        RECT 128.400 185.610 128.660 185.700 ;
        RECT 127.395 184.705 127.625 184.995 ;
        RECT 128.415 184.705 128.645 184.995 ;
        RECT 128.460 184.550 128.600 184.705 ;
        RECT 128.400 184.230 128.660 184.550 ;
        RECT 128.800 184.460 128.940 185.700 ;
        RECT 129.095 184.460 129.325 184.535 ;
        RECT 128.800 184.320 129.325 184.460 ;
        RECT 129.095 184.245 129.325 184.320 ;
        RECT 128.400 183.310 128.660 183.630 ;
        RECT 129.480 181.860 129.960 217.740 ;
        RECT 130.100 215.970 130.360 216.290 ;
        RECT 130.115 214.145 130.345 214.435 ;
        RECT 130.160 211.690 130.300 214.145 ;
        RECT 131.120 213.670 131.380 213.990 ;
        RECT 131.135 212.765 131.365 213.055 ;
        RECT 130.795 211.845 131.025 212.135 ;
        RECT 131.180 212.060 131.320 212.765 ;
        RECT 131.180 211.920 132.000 212.060 ;
        RECT 130.100 211.370 130.360 211.690 ;
        RECT 130.500 210.800 130.640 211.205 ;
        RECT 130.455 210.770 130.685 210.800 ;
        RECT 130.440 210.450 130.700 210.770 ;
        RECT 130.500 203.320 130.640 210.450 ;
        RECT 130.840 209.390 130.980 211.845 ;
        RECT 131.475 211.360 131.705 211.650 ;
        RECT 131.135 210.965 131.365 211.255 ;
        RECT 131.180 210.065 131.320 210.965 ;
        RECT 131.135 209.775 131.365 210.065 ;
        RECT 130.780 209.070 131.040 209.390 ;
        RECT 130.840 206.630 130.980 209.070 ;
        RECT 131.180 207.545 131.320 209.775 ;
        RECT 131.520 209.550 131.660 211.360 ;
        RECT 131.475 209.260 131.705 209.550 ;
        RECT 131.520 207.980 131.660 209.260 ;
        RECT 131.475 207.690 131.705 207.980 ;
        RECT 131.135 207.255 131.365 207.545 ;
        RECT 130.780 206.310 131.040 206.630 ;
        RECT 131.475 205.160 131.705 205.235 ;
        RECT 130.160 203.180 130.640 203.320 ;
        RECT 130.840 205.020 131.705 205.160 ;
        RECT 130.160 196.970 130.300 203.180 ;
        RECT 130.455 202.690 130.685 202.980 ;
        RECT 130.100 196.650 130.360 196.970 ;
        RECT 130.160 196.035 130.300 196.650 ;
        RECT 130.500 196.510 130.640 202.690 ;
        RECT 130.440 196.190 130.700 196.510 ;
        RECT 130.840 196.050 130.980 205.020 ;
        RECT 131.475 204.945 131.705 205.020 ;
        RECT 131.120 204.010 131.380 204.330 ;
        RECT 131.475 203.540 131.705 203.830 ;
        RECT 131.135 203.145 131.365 203.435 ;
        RECT 131.180 202.245 131.320 203.145 ;
        RECT 131.135 201.955 131.365 202.245 ;
        RECT 131.180 199.725 131.320 201.955 ;
        RECT 131.520 201.730 131.660 203.540 ;
        RECT 131.860 203.410 132.000 211.920 ;
        RECT 131.800 203.090 132.060 203.410 ;
        RECT 131.475 201.440 131.705 201.730 ;
        RECT 131.520 200.160 131.660 201.440 ;
        RECT 131.475 199.870 131.705 200.160 ;
        RECT 131.135 199.435 131.365 199.725 ;
        RECT 131.815 197.125 132.045 197.415 ;
        RECT 131.860 196.970 132.000 197.125 ;
        RECT 131.800 196.650 132.060 196.970 ;
        RECT 130.115 195.745 130.345 196.035 ;
        RECT 130.780 195.730 131.040 196.050 ;
        RECT 130.440 195.040 130.700 195.130 ;
        RECT 130.840 195.040 130.980 195.730 ;
        RECT 131.460 195.270 131.720 195.590 ;
        RECT 130.440 194.900 130.980 195.040 ;
        RECT 130.440 194.810 130.700 194.900 ;
        RECT 130.500 193.735 130.640 194.810 ;
        RECT 130.455 193.445 130.685 193.735 ;
        RECT 130.115 192.065 130.345 192.355 ;
        RECT 130.160 191.450 130.300 192.065 ;
        RECT 130.100 191.130 130.360 191.450 ;
        RECT 130.795 191.360 131.025 191.435 ;
        RECT 130.500 191.220 131.025 191.360 ;
        RECT 130.500 190.900 130.640 191.220 ;
        RECT 130.795 191.145 131.025 191.220 ;
        RECT 130.160 190.760 130.640 190.900 ;
        RECT 131.135 190.900 131.365 190.975 ;
        RECT 131.135 190.760 131.660 190.900 ;
        RECT 130.160 186.300 130.300 190.760 ;
        RECT 131.135 190.685 131.365 190.760 ;
        RECT 131.135 190.225 131.365 190.515 ;
        RECT 130.795 189.980 131.025 190.055 ;
        RECT 130.500 189.840 131.025 189.980 ;
        RECT 130.500 188.675 130.640 189.840 ;
        RECT 130.795 189.765 131.025 189.840 ;
        RECT 130.780 189.290 131.040 189.610 ;
        RECT 130.840 189.135 130.980 189.290 ;
        RECT 130.795 188.845 131.025 189.135 ;
        RECT 130.455 188.385 130.685 188.675 ;
        RECT 130.795 187.925 131.025 188.215 ;
        RECT 130.840 186.850 130.980 187.925 ;
        RECT 131.180 187.770 131.320 190.225 ;
        RECT 131.520 188.690 131.660 190.760 ;
        RECT 131.460 188.370 131.720 188.690 ;
        RECT 131.120 187.450 131.380 187.770 ;
        RECT 130.780 186.530 131.040 186.850 ;
        RECT 130.780 186.300 131.040 186.390 ;
        RECT 130.160 186.160 131.040 186.300 ;
        RECT 130.780 186.070 131.040 186.160 ;
        RECT 130.780 184.690 131.040 185.010 ;
        RECT 130.780 184.230 131.040 184.550 ;
        RECT 130.840 184.075 130.980 184.230 ;
        RECT 131.520 184.090 131.660 188.370 ;
        RECT 131.815 187.005 132.045 187.295 ;
        RECT 131.860 185.470 132.000 187.005 ;
        RECT 131.800 185.150 132.060 185.470 ;
        RECT 130.795 183.785 131.025 184.075 ;
        RECT 131.460 183.770 131.720 184.090 ;
        RECT 132.200 181.860 132.680 217.740 ;
        RECT 134.520 216.430 134.780 216.750 ;
        RECT 134.580 215.815 134.720 216.430 ;
        RECT 134.535 215.525 134.765 215.815 ;
        RECT 133.855 214.605 134.085 214.895 ;
        RECT 133.160 213.670 133.420 213.990 ;
        RECT 133.220 212.060 133.360 213.670 ;
        RECT 133.515 212.060 133.745 212.135 ;
        RECT 133.220 211.920 133.745 212.060 ;
        RECT 132.835 199.425 133.065 199.715 ;
        RECT 132.880 199.270 133.020 199.425 ;
        RECT 132.820 198.950 133.080 199.270 ;
        RECT 133.220 194.210 133.360 211.920 ;
        RECT 133.515 211.845 133.745 211.920 ;
        RECT 133.515 210.925 133.745 211.215 ;
        RECT 133.560 210.770 133.700 210.925 ;
        RECT 133.500 210.450 133.760 210.770 ;
        RECT 133.900 209.390 134.040 214.605 ;
        RECT 134.520 214.130 134.780 214.450 ;
        RECT 134.535 212.305 134.765 212.595 ;
        RECT 133.840 209.070 134.100 209.390 ;
        RECT 134.580 208.930 134.720 212.305 ;
        RECT 134.520 208.610 134.780 208.930 ;
        RECT 134.520 206.310 134.780 206.630 ;
        RECT 134.580 204.330 134.720 206.310 ;
        RECT 134.520 204.010 134.780 204.330 ;
        RECT 134.520 203.090 134.780 203.410 ;
        RECT 133.855 199.885 134.085 200.175 ;
        RECT 133.900 199.730 134.040 199.885 ;
        RECT 134.580 199.730 134.720 203.090 ;
        RECT 133.840 199.410 134.100 199.730 ;
        RECT 134.520 199.410 134.780 199.730 ;
        RECT 133.515 196.205 133.745 196.495 ;
        RECT 133.560 196.050 133.700 196.205 ;
        RECT 133.500 195.730 133.760 196.050 ;
        RECT 134.180 194.350 134.440 194.670 ;
        RECT 133.160 193.890 133.420 194.210 ;
        RECT 133.515 193.445 133.745 193.735 ;
        RECT 132.835 193.200 133.065 193.275 ;
        RECT 132.835 193.060 133.360 193.200 ;
        RECT 132.835 192.985 133.065 193.060 ;
        RECT 132.820 192.050 133.080 192.370 ;
        RECT 133.220 189.610 133.360 193.060 ;
        RECT 133.560 190.440 133.700 193.445 ;
        RECT 133.855 193.200 134.085 193.275 ;
        RECT 133.855 193.060 134.720 193.200 ;
        RECT 133.855 192.985 134.085 193.060 ;
        RECT 134.195 191.145 134.425 191.435 ;
        RECT 133.840 190.440 134.100 190.530 ;
        RECT 133.560 190.300 134.100 190.440 ;
        RECT 133.840 190.210 134.100 190.300 ;
        RECT 134.240 190.070 134.380 191.145 ;
        RECT 134.180 189.750 134.440 190.070 ;
        RECT 133.160 189.290 133.420 189.610 ;
        RECT 134.180 189.290 134.440 189.610 ;
        RECT 133.855 189.060 134.085 189.135 ;
        RECT 133.560 188.920 134.085 189.060 ;
        RECT 133.560 187.755 133.700 188.920 ;
        RECT 133.855 188.845 134.085 188.920 ;
        RECT 133.855 188.140 134.085 188.215 ;
        RECT 134.240 188.140 134.380 189.290 ;
        RECT 133.855 188.000 134.380 188.140 ;
        RECT 133.855 187.925 134.085 188.000 ;
        RECT 133.515 187.465 133.745 187.755 ;
        RECT 133.840 186.530 134.100 186.850 ;
        RECT 133.840 185.150 134.100 185.470 ;
        RECT 133.855 184.245 134.085 184.535 ;
        RECT 134.240 184.460 134.380 188.000 ;
        RECT 134.580 186.850 134.720 193.060 ;
        RECT 134.520 186.530 134.780 186.850 ;
        RECT 134.520 184.460 134.780 184.550 ;
        RECT 134.240 184.320 134.780 184.460 ;
        RECT 133.900 184.090 134.040 184.245 ;
        RECT 134.520 184.230 134.780 184.320 ;
        RECT 133.840 183.770 134.100 184.090 ;
        RECT 134.920 181.860 135.400 217.740 ;
        RECT 136.235 215.985 136.465 216.275 ;
        RECT 135.895 214.650 136.125 214.940 ;
        RECT 135.940 214.450 136.080 214.650 ;
        RECT 135.880 214.130 136.140 214.450 ;
        RECT 135.540 209.300 135.800 209.390 ;
        RECT 135.540 209.160 136.080 209.300 ;
        RECT 135.540 209.070 135.800 209.160 ;
        RECT 135.540 208.610 135.800 208.930 ;
        RECT 135.940 206.080 136.080 209.160 ;
        RECT 136.280 206.630 136.420 215.985 ;
        RECT 136.915 215.500 137.145 215.790 ;
        RECT 136.575 215.105 136.805 215.395 ;
        RECT 136.620 214.205 136.760 215.105 ;
        RECT 136.575 213.915 136.805 214.205 ;
        RECT 136.620 211.685 136.760 213.915 ;
        RECT 136.960 213.690 137.100 215.500 ;
        RECT 136.915 213.400 137.145 213.690 ;
        RECT 136.960 212.120 137.100 213.400 ;
        RECT 136.915 211.830 137.145 212.120 ;
        RECT 136.575 211.395 136.805 211.685 ;
        RECT 136.220 206.310 136.480 206.630 ;
        RECT 136.235 206.080 136.465 206.155 ;
        RECT 135.940 205.940 136.465 206.080 ;
        RECT 136.235 205.865 136.465 205.940 ;
        RECT 137.240 204.010 137.500 204.330 ;
        RECT 136.235 202.185 136.465 202.475 ;
        RECT 135.895 201.725 136.125 202.015 ;
        RECT 135.540 199.870 135.800 200.190 ;
        RECT 135.600 197.875 135.740 199.870 ;
        RECT 135.555 197.585 135.785 197.875 ;
        RECT 135.940 194.210 136.080 201.725 ;
        RECT 136.280 200.190 136.420 202.185 ;
        RECT 136.575 201.020 136.805 201.095 ;
        RECT 136.575 200.880 137.100 201.020 ;
        RECT 136.575 200.805 136.805 200.880 ;
        RECT 136.220 199.870 136.480 200.190 ;
        RECT 136.220 199.410 136.480 199.730 ;
        RECT 136.220 198.490 136.480 198.810 ;
        RECT 136.280 196.970 136.420 198.490 ;
        RECT 136.220 196.650 136.480 196.970 ;
        RECT 136.220 196.190 136.480 196.510 ;
        RECT 136.280 195.590 136.420 196.190 ;
        RECT 136.560 195.730 136.820 196.050 ;
        RECT 136.960 195.960 137.100 200.880 ;
        RECT 137.240 198.950 137.500 199.270 ;
        RECT 137.300 196.955 137.440 198.950 ;
        RECT 137.255 196.665 137.485 196.955 ;
        RECT 136.960 195.820 137.440 195.960 ;
        RECT 136.220 195.270 136.480 195.590 ;
        RECT 136.915 195.260 137.145 195.550 ;
        RECT 136.575 194.865 136.805 195.155 ;
        RECT 136.235 194.410 136.465 194.700 ;
        RECT 135.880 193.890 136.140 194.210 ;
        RECT 136.280 193.290 136.420 194.410 ;
        RECT 136.620 193.965 136.760 194.865 ;
        RECT 136.575 193.675 136.805 193.965 ;
        RECT 136.220 192.970 136.480 193.290 ;
        RECT 136.620 191.445 136.760 193.675 ;
        RECT 136.960 193.450 137.100 195.260 ;
        RECT 137.300 194.210 137.440 195.820 ;
        RECT 137.240 193.890 137.500 194.210 ;
        RECT 136.915 193.160 137.145 193.450 ;
        RECT 136.960 191.880 137.100 193.160 ;
        RECT 136.915 191.590 137.145 191.880 ;
        RECT 136.575 191.155 136.805 191.445 ;
        RECT 137.300 190.900 137.440 193.890 ;
        RECT 136.280 190.760 137.440 190.900 ;
        RECT 136.280 188.215 136.420 190.760 ;
        RECT 137.240 188.830 137.500 189.150 ;
        RECT 136.235 187.925 136.465 188.215 ;
        RECT 136.220 186.990 136.480 187.310 ;
        RECT 137.240 186.070 137.500 186.390 ;
        RECT 136.220 185.610 136.480 185.930 ;
        RECT 135.540 184.690 135.800 185.010 ;
        RECT 135.540 184.230 135.800 184.550 ;
        RECT 136.220 183.310 136.480 183.630 ;
        RECT 137.640 181.860 138.120 217.740 ;
        RECT 139.960 211.830 140.220 212.150 ;
        RECT 138.955 209.535 139.185 209.825 ;
        RECT 138.615 209.100 138.845 209.390 ;
        RECT 138.660 207.820 138.800 209.100 ;
        RECT 138.615 207.530 138.845 207.820 ;
        RECT 138.260 206.310 138.520 206.630 ;
        RECT 138.320 204.700 138.460 206.310 ;
        RECT 138.660 205.720 138.800 207.530 ;
        RECT 139.000 207.305 139.140 209.535 ;
        RECT 138.955 207.015 139.185 207.305 ;
        RECT 139.960 207.230 140.220 207.550 ;
        RECT 139.000 206.115 139.140 207.015 ;
        RECT 139.295 206.225 139.525 206.515 ;
        RECT 138.955 205.825 139.185 206.115 ;
        RECT 138.615 205.430 138.845 205.720 ;
        RECT 138.955 204.945 139.185 205.235 ;
        RECT 139.000 204.775 139.140 204.945 ;
        RECT 138.955 204.700 139.185 204.775 ;
        RECT 138.320 204.560 139.185 204.700 ;
        RECT 138.320 196.050 138.460 204.560 ;
        RECT 138.955 204.485 139.185 204.560 ;
        RECT 139.340 204.330 139.480 206.225 ;
        RECT 139.620 204.930 139.880 205.250 ;
        RECT 138.615 204.000 138.845 204.290 ;
        RECT 139.280 204.010 139.540 204.330 ;
        RECT 138.660 202.190 138.800 204.000 ;
        RECT 138.955 203.605 139.185 203.895 ;
        RECT 139.000 202.705 139.140 203.605 ;
        RECT 139.680 203.550 139.820 204.930 ;
        RECT 139.635 203.260 139.865 203.550 ;
        RECT 138.955 202.415 139.185 202.705 ;
        RECT 138.615 201.900 138.845 202.190 ;
        RECT 138.660 200.620 138.800 201.900 ;
        RECT 138.615 200.330 138.845 200.620 ;
        RECT 139.000 200.185 139.140 202.415 ;
        RECT 140.020 202.400 140.160 207.230 ;
        RECT 139.680 202.260 140.160 202.400 ;
        RECT 138.955 199.895 139.185 200.185 ;
        RECT 138.600 199.410 138.860 199.730 ;
        RECT 138.260 195.730 138.520 196.050 ;
        RECT 138.660 194.195 138.800 199.410 ;
        RECT 138.940 198.490 139.200 198.810 ;
        RECT 139.000 195.040 139.140 198.490 ;
        RECT 139.680 197.415 139.820 202.260 ;
        RECT 139.975 197.585 140.205 197.875 ;
        RECT 139.635 197.125 139.865 197.415 ;
        RECT 140.020 196.970 140.160 197.585 ;
        RECT 139.960 196.650 140.220 196.970 ;
        RECT 139.620 196.190 139.880 196.510 ;
        RECT 139.280 195.270 139.540 195.590 ;
        RECT 139.295 195.040 139.525 195.115 ;
        RECT 139.000 194.900 139.525 195.040 ;
        RECT 139.295 194.825 139.525 194.900 ;
        RECT 138.940 194.350 139.200 194.670 ;
        RECT 138.615 193.905 138.845 194.195 ;
        RECT 138.260 192.970 138.520 193.290 ;
        RECT 138.320 191.435 138.460 192.970 ;
        RECT 138.615 192.525 138.845 192.815 ;
        RECT 138.275 191.145 138.505 191.435 ;
        RECT 138.660 190.055 138.800 192.525 ;
        RECT 139.000 192.280 139.140 194.350 ;
        RECT 139.280 193.890 139.540 194.210 ;
        RECT 139.340 193.275 139.480 193.890 ;
        RECT 139.295 192.985 139.525 193.275 ;
        RECT 139.280 192.280 139.540 192.370 ;
        RECT 139.000 192.140 139.540 192.280 ;
        RECT 139.280 192.050 139.540 192.140 ;
        RECT 139.340 190.515 139.480 192.050 ;
        RECT 139.295 190.225 139.525 190.515 ;
        RECT 138.615 189.765 138.845 190.055 ;
        RECT 139.280 189.290 139.540 189.610 ;
        RECT 138.600 188.830 138.860 189.150 ;
        RECT 139.295 188.845 139.525 189.135 ;
        RECT 138.660 188.140 138.800 188.830 ;
        RECT 138.955 188.140 139.185 188.215 ;
        RECT 138.660 188.000 139.185 188.140 ;
        RECT 138.955 187.925 139.185 188.000 ;
        RECT 138.260 186.990 138.520 187.310 ;
        RECT 138.320 184.995 138.460 186.990 ;
        RECT 139.340 186.390 139.480 188.845 ;
        RECT 139.280 186.070 139.540 186.390 ;
        RECT 138.600 185.610 138.860 185.930 ;
        RECT 138.275 184.705 138.505 184.995 ;
        RECT 138.660 184.535 138.800 185.610 ;
        RECT 138.615 184.245 138.845 184.535 ;
        RECT 139.280 183.310 139.540 183.630 ;
        RECT 140.360 181.860 140.840 217.740 ;
        RECT 141.660 211.830 141.920 212.150 ;
        RECT 141.720 209.835 141.860 211.830 ;
        RECT 141.675 209.760 141.905 209.835 ;
        RECT 141.675 209.620 142.200 209.760 ;
        RECT 141.675 209.545 141.905 209.620 ;
        RECT 141.660 207.230 141.920 207.550 ;
        RECT 141.660 206.770 141.920 207.090 ;
        RECT 141.675 205.865 141.905 206.155 ;
        RECT 140.980 204.930 141.240 205.250 ;
        RECT 140.980 199.870 141.240 200.190 ;
        RECT 141.720 197.800 141.860 205.865 ;
        RECT 142.060 203.395 142.200 209.620 ;
        RECT 142.695 208.625 142.925 208.915 ;
        RECT 142.355 206.325 142.585 206.615 ;
        RECT 142.015 203.105 142.245 203.395 ;
        RECT 142.400 199.270 142.540 206.325 ;
        RECT 142.740 203.870 142.880 208.625 ;
        RECT 142.680 203.550 142.940 203.870 ;
        RECT 142.340 198.950 142.600 199.270 ;
        RECT 142.695 198.045 142.925 198.335 ;
        RECT 141.720 197.660 142.540 197.800 ;
        RECT 141.675 197.125 141.905 197.415 ;
        RECT 141.720 196.970 141.860 197.125 ;
        RECT 141.660 196.650 141.920 196.970 ;
        RECT 140.980 196.190 141.240 196.510 ;
        RECT 141.040 193.735 141.180 196.190 ;
        RECT 141.660 193.890 141.920 194.210 ;
        RECT 140.995 193.445 141.225 193.735 ;
        RECT 141.720 193.275 141.860 193.890 ;
        RECT 141.675 192.985 141.905 193.275 ;
        RECT 142.400 192.370 142.540 197.660 ;
        RECT 142.740 197.430 142.880 198.045 ;
        RECT 142.680 197.110 142.940 197.430 ;
        RECT 142.340 192.050 142.600 192.370 ;
        RECT 142.680 190.670 142.940 190.990 ;
        RECT 140.980 190.210 141.240 190.530 ;
        RECT 141.040 187.295 141.180 190.210 ;
        RECT 142.740 190.055 142.880 190.670 ;
        RECT 142.695 189.765 142.925 190.055 ;
        RECT 141.660 188.830 141.920 189.150 ;
        RECT 140.995 187.005 141.225 187.295 ;
        RECT 140.980 186.530 141.240 186.850 ;
        RECT 141.040 185.915 141.180 186.530 ;
        RECT 141.660 186.070 141.920 186.390 ;
        RECT 140.995 185.625 141.225 185.915 ;
        RECT 141.660 184.690 141.920 185.010 ;
        RECT 140.995 184.245 141.225 184.535 ;
        RECT 141.040 184.090 141.180 184.245 ;
        RECT 140.980 183.770 141.240 184.090 ;
        RECT 141.660 183.310 141.920 183.630 ;
        RECT 143.080 181.860 143.560 217.740 ;
        RECT 143.905 201.705 144.055 217.960 ;
        RECT 143.910 199.760 144.050 201.705 ;
        RECT 143.810 199.370 144.160 199.760 ;
        RECT 144.420 197.400 144.560 218.920 ;
        RECT 144.330 197.140 144.650 197.400 ;
        RECT 145.040 191.000 145.180 220.260 ;
        RECT 145.470 203.870 145.610 221.200 ;
        RECT 145.380 203.550 145.700 203.870 ;
        RECT 144.940 190.660 145.270 191.000 ;
        RECT 115.310 173.480 117.720 174.140 ;
        RECT 97.850 173.010 98.110 173.040 ;
        RECT 97.850 170.910 98.680 173.010 ;
        RECT 104.350 172.620 105.600 173.060 ;
        RECT 102.290 172.610 107.530 172.620 ;
        RECT 99.340 172.510 114.640 172.610 ;
        RECT 99.340 172.500 114.675 172.510 ;
        RECT 99.300 172.380 114.675 172.500 ;
        RECT 99.300 172.270 103.300 172.380 ;
        RECT 104.350 172.300 106.090 172.380 ;
        RECT 106.670 172.300 114.675 172.380 ;
        RECT 104.350 172.220 105.600 172.300 ;
        RECT 106.675 172.280 114.675 172.300 ;
        RECT 98.910 171.970 99.140 172.220 ;
        RECT 103.460 172.080 103.690 172.220 ;
        RECT 106.240 172.080 106.470 172.230 ;
        RECT 103.460 171.970 106.470 172.080 ;
        RECT 114.880 171.970 115.110 172.230 ;
        RECT 98.910 171.530 115.110 171.970 ;
        RECT 98.910 171.260 99.140 171.530 ;
        RECT 103.460 171.500 115.110 171.530 ;
        RECT 103.460 171.410 106.470 171.500 ;
        RECT 103.460 171.260 103.690 171.410 ;
        RECT 106.240 171.270 106.470 171.410 ;
        RECT 114.880 171.270 115.110 171.500 ;
        RECT 99.300 170.980 103.300 171.210 ;
        RECT 106.675 171.000 114.675 171.220 ;
        RECT 115.440 171.000 116.400 173.040 ;
        RECT 116.870 172.350 117.720 173.480 ;
        RECT 123.390 172.650 124.640 173.090 ;
        RECT 135.840 173.080 136.100 173.110 ;
        RECT 121.330 172.640 126.570 172.650 ;
        RECT 118.380 172.540 133.680 172.640 ;
        RECT 118.380 172.530 133.715 172.540 ;
        RECT 106.675 170.990 116.400 171.000 ;
        RECT 99.300 170.910 103.290 170.980 ;
        RECT 97.850 170.800 103.290 170.910 ;
        RECT 106.730 170.830 116.400 170.990 ;
        RECT 97.850 170.710 100.980 170.800 ;
        RECT 114.470 170.780 116.400 170.830 ;
        RECT 97.850 167.440 98.680 170.710 ;
        RECT 102.330 170.250 107.580 170.260 ;
        RECT 102.330 170.140 114.640 170.250 ;
        RECT 99.360 170.080 114.640 170.140 ;
        RECT 99.360 170.070 114.675 170.080 ;
        RECT 99.300 169.940 114.675 170.070 ;
        RECT 99.300 169.930 104.460 169.940 ;
        RECT 99.300 169.840 103.300 169.930 ;
        RECT 106.675 169.850 114.675 169.940 ;
        RECT 106.760 169.840 114.650 169.850 ;
        RECT 98.910 169.480 99.140 169.790 ;
        RECT 99.360 169.480 103.260 169.840 ;
        RECT 103.460 169.480 103.690 169.790 ;
        RECT 98.910 168.140 103.690 169.480 ;
        RECT 98.910 167.830 99.140 168.140 ;
        RECT 103.460 167.830 103.690 168.140 ;
        RECT 106.240 169.260 106.470 169.800 ;
        RECT 107.280 169.260 108.290 169.290 ;
        RECT 114.880 169.260 115.110 169.800 ;
        RECT 106.240 168.360 115.110 169.260 ;
        RECT 106.240 167.840 106.470 168.360 ;
        RECT 107.280 168.290 108.290 168.360 ;
        RECT 114.880 167.840 115.110 168.360 ;
        RECT 99.300 167.550 103.300 167.780 ;
        RECT 106.675 167.560 114.675 167.790 ;
        RECT 97.850 167.400 98.980 167.440 ;
        RECT 97.850 167.320 99.220 167.400 ;
        RECT 99.590 167.330 103.250 167.550 ;
        RECT 99.590 167.320 101.030 167.330 ;
        RECT 97.850 167.280 101.030 167.320 ;
        RECT 97.850 167.190 100.540 167.280 ;
        RECT 106.740 167.270 114.630 167.560 ;
        RECT 97.850 167.130 99.870 167.190 ;
        RECT 97.850 167.080 99.620 167.130 ;
        RECT 97.850 163.740 98.680 167.080 ;
        RECT 106.730 166.780 114.650 166.790 ;
        RECT 102.960 166.770 114.650 166.780 ;
        RECT 99.340 166.650 114.650 166.770 ;
        RECT 99.340 166.640 114.675 166.650 ;
        RECT 99.300 166.520 114.675 166.640 ;
        RECT 99.300 166.410 103.300 166.520 ;
        RECT 98.910 166.070 99.140 166.360 ;
        RECT 99.360 166.070 103.250 166.410 ;
        RECT 103.460 166.070 103.690 166.360 ;
        RECT 98.910 164.700 103.690 166.070 ;
        RECT 98.910 164.400 99.140 164.700 ;
        RECT 103.460 164.400 103.690 164.700 ;
        RECT 99.300 164.120 103.300 164.350 ;
        RECT 99.550 163.890 103.120 164.120 ;
        RECT 99.550 163.740 103.240 163.890 ;
        RECT 97.850 163.460 103.240 163.740 ;
        RECT 104.490 163.570 105.110 166.520 ;
        RECT 106.675 166.420 114.675 166.520 ;
        RECT 106.730 166.410 114.650 166.420 ;
        RECT 106.240 165.710 106.470 166.370 ;
        RECT 107.250 165.710 108.250 165.800 ;
        RECT 114.880 165.710 115.110 166.370 ;
        RECT 106.240 164.890 115.110 165.710 ;
        RECT 106.240 164.410 106.470 164.890 ;
        RECT 107.250 164.800 108.250 164.890 ;
        RECT 114.880 164.410 115.110 164.890 ;
        RECT 106.675 164.130 114.675 164.360 ;
        RECT 97.850 163.000 103.250 163.460 ;
        RECT 97.850 161.660 99.850 163.000 ;
        RECT 101.600 162.990 103.250 163.000 ;
        RECT 100.290 161.720 101.290 162.440 ;
        RECT 101.600 162.180 101.910 162.990 ;
        RECT 102.370 162.710 103.250 162.990 ;
        RECT 103.490 163.170 105.110 163.570 ;
        RECT 106.760 163.220 114.630 164.130 ;
        RECT 102.310 162.480 103.310 162.710 ;
        RECT 103.490 162.520 103.840 163.170 ;
        RECT 104.490 163.160 105.110 163.170 ;
        RECT 106.675 162.990 114.675 163.220 ;
        RECT 106.760 162.980 114.630 162.990 ;
        RECT 102.370 162.270 103.250 162.290 ;
        RECT 101.640 161.890 101.910 162.180 ;
        RECT 102.310 162.040 103.310 162.270 ;
        RECT 103.470 162.230 103.840 162.520 ;
        RECT 103.500 162.170 103.840 162.230 ;
        RECT 104.600 162.840 105.360 162.890 ;
        RECT 106.240 162.840 106.470 162.940 ;
        RECT 104.600 162.630 106.470 162.840 ;
        RECT 114.880 162.630 115.110 162.940 ;
        RECT 104.600 162.210 107.140 162.630 ;
        RECT 114.510 162.210 115.110 162.630 ;
        RECT 102.370 161.890 103.250 162.040 ;
        RECT 102.380 161.720 103.110 161.890 ;
        RECT 97.860 161.650 99.850 161.660 ;
        RECT 97.860 158.050 98.640 161.650 ;
        RECT 100.260 160.600 103.110 161.720 ;
        RECT 103.500 161.420 103.850 162.170 ;
        RECT 104.600 162.050 106.470 162.210 ;
        RECT 104.600 162.000 105.360 162.050 ;
        RECT 106.240 161.980 106.470 162.050 ;
        RECT 114.880 161.980 115.110 162.210 ;
        RECT 106.675 161.700 114.675 161.930 ;
        RECT 103.500 161.360 103.790 161.420 ;
        RECT 103.410 161.240 103.790 161.360 ;
        RECT 106.770 161.300 114.630 161.700 ;
        RECT 115.440 161.400 116.400 170.780 ;
        RECT 116.890 170.940 117.720 172.350 ;
        RECT 118.340 172.410 133.715 172.530 ;
        RECT 118.340 172.300 122.340 172.410 ;
        RECT 123.390 172.330 125.130 172.410 ;
        RECT 125.710 172.330 133.715 172.410 ;
        RECT 123.390 172.250 124.640 172.330 ;
        RECT 125.715 172.310 133.715 172.330 ;
        RECT 117.950 172.000 118.180 172.250 ;
        RECT 122.500 172.110 122.730 172.250 ;
        RECT 125.280 172.110 125.510 172.260 ;
        RECT 122.500 172.000 125.510 172.110 ;
        RECT 133.920 172.000 134.150 172.260 ;
        RECT 117.950 171.560 134.150 172.000 ;
        RECT 117.950 171.290 118.180 171.560 ;
        RECT 122.500 171.530 134.150 171.560 ;
        RECT 122.500 171.440 125.510 171.530 ;
        RECT 122.500 171.290 122.730 171.440 ;
        RECT 125.280 171.300 125.510 171.440 ;
        RECT 133.920 171.300 134.150 171.530 ;
        RECT 118.340 171.010 122.340 171.240 ;
        RECT 125.715 171.030 133.715 171.250 ;
        RECT 134.480 171.030 135.440 173.070 ;
        RECT 125.715 171.020 135.440 171.030 ;
        RECT 118.340 170.940 122.330 171.010 ;
        RECT 116.890 170.830 122.330 170.940 ;
        RECT 125.770 170.860 135.440 171.020 ;
        RECT 116.890 170.740 120.020 170.830 ;
        RECT 133.510 170.810 135.440 170.860 ;
        RECT 116.890 167.480 117.720 170.740 ;
        RECT 121.370 170.280 126.620 170.290 ;
        RECT 121.370 170.170 133.680 170.280 ;
        RECT 118.400 170.110 133.680 170.170 ;
        RECT 118.400 170.100 133.715 170.110 ;
        RECT 118.340 169.970 133.715 170.100 ;
        RECT 118.340 169.960 123.500 169.970 ;
        RECT 118.340 169.870 122.340 169.960 ;
        RECT 125.715 169.880 133.715 169.970 ;
        RECT 125.800 169.870 133.690 169.880 ;
        RECT 117.950 169.510 118.180 169.820 ;
        RECT 118.400 169.510 122.300 169.870 ;
        RECT 122.500 169.510 122.730 169.820 ;
        RECT 117.950 168.170 122.730 169.510 ;
        RECT 117.950 167.860 118.180 168.170 ;
        RECT 122.500 167.860 122.730 168.170 ;
        RECT 125.280 169.290 125.510 169.830 ;
        RECT 126.320 169.290 127.330 169.320 ;
        RECT 133.920 169.290 134.150 169.830 ;
        RECT 125.280 168.390 134.150 169.290 ;
        RECT 125.280 167.870 125.510 168.390 ;
        RECT 126.320 168.320 127.330 168.390 ;
        RECT 133.920 167.870 134.150 168.390 ;
        RECT 118.340 167.580 122.340 167.810 ;
        RECT 125.715 167.590 133.715 167.820 ;
        RECT 115.430 161.300 116.400 161.400 ;
        RECT 100.200 160.370 103.200 160.600 ;
        RECT 103.410 160.410 103.750 161.240 ;
        RECT 105.760 161.230 116.400 161.300 ;
        RECT 100.250 160.340 103.110 160.370 ;
        RECT 100.250 160.320 101.420 160.340 ;
        RECT 102.380 160.330 103.110 160.340 ;
        RECT 100.200 159.930 103.200 160.160 ;
        RECT 103.405 160.120 103.750 160.410 ;
        RECT 103.940 160.190 116.400 161.230 ;
        RECT 116.860 167.470 117.720 167.480 ;
        RECT 116.860 167.430 118.020 167.470 ;
        RECT 116.860 167.350 118.260 167.430 ;
        RECT 118.630 167.360 122.290 167.580 ;
        RECT 118.630 167.350 120.070 167.360 ;
        RECT 116.860 167.310 120.070 167.350 ;
        RECT 116.860 167.220 119.580 167.310 ;
        RECT 125.780 167.300 133.670 167.590 ;
        RECT 116.860 167.160 118.910 167.220 ;
        RECT 116.860 167.110 118.660 167.160 ;
        RECT 116.860 163.770 117.720 167.110 ;
        RECT 125.770 166.810 133.690 166.820 ;
        RECT 122.000 166.800 133.690 166.810 ;
        RECT 118.380 166.680 133.690 166.800 ;
        RECT 118.380 166.670 133.715 166.680 ;
        RECT 118.340 166.550 133.715 166.670 ;
        RECT 118.340 166.440 122.340 166.550 ;
        RECT 117.950 166.100 118.180 166.390 ;
        RECT 118.400 166.100 122.290 166.440 ;
        RECT 122.500 166.100 122.730 166.390 ;
        RECT 117.950 164.730 122.730 166.100 ;
        RECT 117.950 164.430 118.180 164.730 ;
        RECT 122.500 164.430 122.730 164.730 ;
        RECT 118.340 164.150 122.340 164.380 ;
        RECT 118.590 163.920 122.160 164.150 ;
        RECT 118.590 163.770 122.280 163.920 ;
        RECT 116.860 163.490 122.280 163.770 ;
        RECT 123.530 163.600 124.150 166.550 ;
        RECT 125.715 166.450 133.715 166.550 ;
        RECT 125.770 166.440 133.690 166.450 ;
        RECT 125.280 165.740 125.510 166.400 ;
        RECT 126.290 165.740 127.290 165.830 ;
        RECT 133.920 165.740 134.150 166.400 ;
        RECT 125.280 164.920 134.150 165.740 ;
        RECT 125.280 164.440 125.510 164.920 ;
        RECT 126.290 164.830 127.290 164.920 ;
        RECT 133.920 164.440 134.150 164.920 ;
        RECT 125.715 164.160 133.715 164.390 ;
        RECT 116.860 163.030 122.290 163.490 ;
        RECT 116.860 161.680 118.890 163.030 ;
        RECT 120.640 163.020 122.290 163.030 ;
        RECT 119.330 161.750 120.330 162.470 ;
        RECT 120.640 162.210 120.950 163.020 ;
        RECT 121.410 162.740 122.290 163.020 ;
        RECT 122.530 163.200 124.150 163.600 ;
        RECT 125.800 163.250 133.670 164.160 ;
        RECT 121.350 162.510 122.350 162.740 ;
        RECT 122.530 162.550 122.880 163.200 ;
        RECT 123.530 163.190 124.150 163.200 ;
        RECT 125.715 163.020 133.715 163.250 ;
        RECT 125.800 163.010 133.670 163.020 ;
        RECT 121.410 162.300 122.290 162.320 ;
        RECT 120.680 161.920 120.950 162.210 ;
        RECT 121.350 162.070 122.350 162.300 ;
        RECT 122.510 162.260 122.880 162.550 ;
        RECT 122.540 162.200 122.880 162.260 ;
        RECT 123.640 162.870 124.400 162.920 ;
        RECT 125.280 162.870 125.510 162.970 ;
        RECT 123.640 162.660 125.510 162.870 ;
        RECT 133.920 162.660 134.150 162.970 ;
        RECT 123.640 162.240 126.180 162.660 ;
        RECT 133.550 162.240 134.150 162.660 ;
        RECT 121.410 161.920 122.290 162.070 ;
        RECT 121.420 161.750 122.150 161.920 ;
        RECT 103.940 160.170 116.370 160.190 ;
        RECT 104.210 160.160 109.650 160.170 ;
        RECT 110.650 160.160 116.370 160.170 ;
        RECT 103.410 160.010 103.750 160.120 ;
        RECT 97.850 158.020 98.640 158.050 ;
        RECT 97.850 155.920 98.680 158.020 ;
        RECT 104.350 157.630 105.600 158.070 ;
        RECT 115.430 158.050 116.370 160.160 ;
        RECT 102.290 157.620 107.530 157.630 ;
        RECT 99.340 157.520 114.640 157.620 ;
        RECT 99.340 157.510 114.675 157.520 ;
        RECT 99.300 157.390 114.675 157.510 ;
        RECT 99.300 157.280 103.300 157.390 ;
        RECT 104.350 157.310 106.090 157.390 ;
        RECT 106.670 157.310 114.675 157.390 ;
        RECT 104.350 157.230 105.600 157.310 ;
        RECT 106.675 157.290 114.675 157.310 ;
        RECT 98.910 156.980 99.140 157.230 ;
        RECT 103.460 157.090 103.690 157.230 ;
        RECT 106.240 157.090 106.470 157.240 ;
        RECT 103.460 156.980 106.470 157.090 ;
        RECT 114.880 156.980 115.110 157.240 ;
        RECT 98.910 156.540 115.110 156.980 ;
        RECT 98.910 156.270 99.140 156.540 ;
        RECT 103.460 156.510 115.110 156.540 ;
        RECT 103.460 156.420 106.470 156.510 ;
        RECT 103.460 156.270 103.690 156.420 ;
        RECT 106.240 156.280 106.470 156.420 ;
        RECT 114.880 156.280 115.110 156.510 ;
        RECT 115.430 156.420 116.400 158.050 ;
        RECT 99.300 155.990 103.300 156.220 ;
        RECT 106.675 156.010 114.675 156.230 ;
        RECT 115.440 156.010 116.400 156.420 ;
        RECT 106.675 156.000 116.400 156.010 ;
        RECT 99.300 155.920 103.290 155.990 ;
        RECT 97.850 155.810 103.290 155.920 ;
        RECT 106.730 155.840 116.400 156.000 ;
        RECT 97.850 155.720 100.980 155.810 ;
        RECT 114.470 155.790 116.400 155.840 ;
        RECT 97.850 152.450 98.680 155.720 ;
        RECT 102.330 155.260 107.580 155.270 ;
        RECT 102.330 155.150 114.640 155.260 ;
        RECT 99.360 155.090 114.640 155.150 ;
        RECT 99.360 155.080 114.675 155.090 ;
        RECT 99.300 154.950 114.675 155.080 ;
        RECT 99.300 154.940 104.460 154.950 ;
        RECT 99.300 154.850 103.300 154.940 ;
        RECT 106.675 154.860 114.675 154.950 ;
        RECT 106.760 154.850 114.650 154.860 ;
        RECT 98.910 154.490 99.140 154.800 ;
        RECT 99.360 154.490 103.260 154.850 ;
        RECT 103.460 154.490 103.690 154.800 ;
        RECT 98.910 153.150 103.690 154.490 ;
        RECT 98.910 152.840 99.140 153.150 ;
        RECT 103.460 152.840 103.690 153.150 ;
        RECT 106.240 154.270 106.470 154.810 ;
        RECT 107.280 154.270 108.290 154.300 ;
        RECT 114.880 154.270 115.110 154.810 ;
        RECT 106.240 153.370 115.110 154.270 ;
        RECT 106.240 152.850 106.470 153.370 ;
        RECT 107.280 153.300 108.290 153.370 ;
        RECT 114.880 152.850 115.110 153.370 ;
        RECT 99.300 152.560 103.300 152.790 ;
        RECT 106.675 152.570 114.675 152.800 ;
        RECT 97.850 152.410 98.980 152.450 ;
        RECT 97.850 152.330 99.220 152.410 ;
        RECT 99.590 152.340 103.250 152.560 ;
        RECT 99.590 152.330 101.030 152.340 ;
        RECT 97.850 152.290 101.030 152.330 ;
        RECT 97.850 152.200 100.540 152.290 ;
        RECT 106.740 152.280 114.630 152.570 ;
        RECT 97.850 152.140 99.870 152.200 ;
        RECT 97.850 152.090 99.620 152.140 ;
        RECT 97.850 148.750 98.680 152.090 ;
        RECT 106.730 151.790 114.650 151.800 ;
        RECT 102.960 151.780 114.650 151.790 ;
        RECT 99.340 151.660 114.650 151.780 ;
        RECT 99.340 151.650 114.675 151.660 ;
        RECT 99.300 151.530 114.675 151.650 ;
        RECT 99.300 151.420 103.300 151.530 ;
        RECT 98.910 151.080 99.140 151.370 ;
        RECT 99.360 151.080 103.250 151.420 ;
        RECT 103.460 151.080 103.690 151.370 ;
        RECT 98.910 149.710 103.690 151.080 ;
        RECT 98.910 149.410 99.140 149.710 ;
        RECT 103.460 149.410 103.690 149.710 ;
        RECT 99.300 149.130 103.300 149.360 ;
        RECT 99.550 148.900 103.120 149.130 ;
        RECT 99.550 148.750 103.240 148.900 ;
        RECT 97.850 148.470 103.240 148.750 ;
        RECT 104.490 148.580 105.110 151.530 ;
        RECT 106.675 151.430 114.675 151.530 ;
        RECT 106.730 151.420 114.650 151.430 ;
        RECT 106.240 150.720 106.470 151.380 ;
        RECT 107.250 150.720 108.250 150.810 ;
        RECT 114.880 150.720 115.110 151.380 ;
        RECT 106.240 149.900 115.110 150.720 ;
        RECT 106.240 149.420 106.470 149.900 ;
        RECT 107.250 149.810 108.250 149.900 ;
        RECT 114.880 149.420 115.110 149.900 ;
        RECT 106.675 149.140 114.675 149.370 ;
        RECT 97.850 148.010 103.250 148.470 ;
        RECT 97.850 146.670 99.850 148.010 ;
        RECT 101.600 148.000 103.250 148.010 ;
        RECT 100.290 146.730 101.290 147.450 ;
        RECT 101.600 147.190 101.910 148.000 ;
        RECT 102.370 147.720 103.250 148.000 ;
        RECT 103.490 148.180 105.110 148.580 ;
        RECT 106.760 148.230 114.630 149.140 ;
        RECT 102.310 147.490 103.310 147.720 ;
        RECT 103.490 147.530 103.840 148.180 ;
        RECT 104.490 148.170 105.110 148.180 ;
        RECT 106.675 148.000 114.675 148.230 ;
        RECT 106.760 147.990 114.630 148.000 ;
        RECT 102.370 147.280 103.250 147.300 ;
        RECT 101.640 146.900 101.910 147.190 ;
        RECT 102.310 147.050 103.310 147.280 ;
        RECT 103.470 147.240 103.840 147.530 ;
        RECT 103.500 147.180 103.840 147.240 ;
        RECT 104.600 147.850 105.360 147.900 ;
        RECT 106.240 147.850 106.470 147.950 ;
        RECT 104.600 147.640 106.470 147.850 ;
        RECT 114.880 147.640 115.110 147.950 ;
        RECT 104.600 147.220 107.140 147.640 ;
        RECT 114.510 147.220 115.110 147.640 ;
        RECT 102.370 146.900 103.250 147.050 ;
        RECT 102.380 146.730 103.110 146.900 ;
        RECT 97.860 146.660 99.850 146.670 ;
        RECT 97.860 143.070 98.640 146.660 ;
        RECT 100.260 145.610 103.110 146.730 ;
        RECT 103.500 146.430 103.850 147.180 ;
        RECT 104.600 147.060 106.470 147.220 ;
        RECT 104.600 147.010 105.360 147.060 ;
        RECT 106.240 146.990 106.470 147.060 ;
        RECT 114.880 146.990 115.110 147.220 ;
        RECT 106.675 146.710 114.675 146.940 ;
        RECT 103.500 146.370 103.790 146.430 ;
        RECT 103.410 146.250 103.790 146.370 ;
        RECT 106.770 146.310 114.630 146.710 ;
        RECT 115.440 146.500 116.400 155.790 ;
        RECT 115.390 146.310 116.400 146.500 ;
        RECT 100.200 145.380 103.200 145.610 ;
        RECT 103.410 145.420 103.750 146.250 ;
        RECT 105.760 146.240 116.400 146.310 ;
        RECT 100.250 145.350 103.110 145.380 ;
        RECT 100.250 145.330 101.420 145.350 ;
        RECT 102.380 145.340 103.110 145.350 ;
        RECT 100.200 144.940 103.200 145.170 ;
        RECT 103.405 145.130 103.750 145.420 ;
        RECT 103.940 145.200 116.400 146.240 ;
        RECT 116.860 158.020 117.620 161.680 ;
        RECT 119.300 160.630 122.150 161.750 ;
        RECT 122.540 161.450 122.890 162.200 ;
        RECT 123.640 162.080 125.510 162.240 ;
        RECT 123.640 162.030 124.400 162.080 ;
        RECT 125.280 162.010 125.510 162.080 ;
        RECT 133.920 162.010 134.150 162.240 ;
        RECT 125.715 161.730 133.715 161.960 ;
        RECT 122.540 161.390 122.830 161.450 ;
        RECT 122.450 161.270 122.830 161.390 ;
        RECT 125.810 161.330 133.670 161.730 ;
        RECT 134.480 161.330 135.440 170.810 ;
        RECT 135.840 170.980 136.670 173.080 ;
        RECT 142.340 172.690 143.590 173.130 ;
        RECT 140.280 172.680 145.520 172.690 ;
        RECT 137.330 172.580 152.630 172.680 ;
        RECT 137.330 172.570 152.665 172.580 ;
        RECT 137.290 172.450 152.665 172.570 ;
        RECT 137.290 172.340 141.290 172.450 ;
        RECT 142.340 172.370 144.080 172.450 ;
        RECT 144.660 172.370 152.665 172.450 ;
        RECT 142.340 172.290 143.590 172.370 ;
        RECT 144.665 172.350 152.665 172.370 ;
        RECT 136.900 172.040 137.130 172.290 ;
        RECT 141.450 172.150 141.680 172.290 ;
        RECT 144.230 172.150 144.460 172.300 ;
        RECT 141.450 172.040 144.460 172.150 ;
        RECT 152.870 172.040 153.100 172.300 ;
        RECT 136.900 171.600 153.100 172.040 ;
        RECT 136.900 171.330 137.130 171.600 ;
        RECT 141.450 171.570 153.100 171.600 ;
        RECT 141.450 171.480 144.460 171.570 ;
        RECT 141.450 171.330 141.680 171.480 ;
        RECT 144.230 171.340 144.460 171.480 ;
        RECT 152.870 171.340 153.100 171.570 ;
        RECT 137.290 171.050 141.290 171.280 ;
        RECT 144.665 171.070 152.665 171.290 ;
        RECT 153.430 171.070 154.390 173.110 ;
        RECT 144.665 171.060 154.390 171.070 ;
        RECT 137.290 170.980 141.280 171.050 ;
        RECT 135.840 170.870 141.280 170.980 ;
        RECT 144.720 170.900 154.390 171.060 ;
        RECT 135.840 170.780 138.970 170.870 ;
        RECT 152.460 170.850 154.390 170.900 ;
        RECT 135.840 170.640 136.670 170.780 ;
        RECT 135.590 169.180 136.670 170.640 ;
        RECT 140.320 170.320 145.570 170.330 ;
        RECT 140.320 170.210 152.630 170.320 ;
        RECT 137.350 170.150 152.630 170.210 ;
        RECT 137.350 170.140 152.665 170.150 ;
        RECT 137.290 170.010 152.665 170.140 ;
        RECT 137.290 170.000 142.450 170.010 ;
        RECT 137.290 169.910 141.290 170.000 ;
        RECT 144.665 169.920 152.665 170.010 ;
        RECT 144.750 169.910 152.640 169.920 ;
        RECT 135.840 167.510 136.670 169.180 ;
        RECT 136.900 169.550 137.130 169.860 ;
        RECT 137.350 169.550 141.250 169.910 ;
        RECT 141.450 169.550 141.680 169.860 ;
        RECT 136.900 168.210 141.680 169.550 ;
        RECT 136.900 167.900 137.130 168.210 ;
        RECT 141.450 167.900 141.680 168.210 ;
        RECT 144.230 169.330 144.460 169.870 ;
        RECT 145.270 169.330 146.280 169.360 ;
        RECT 152.870 169.330 153.100 169.870 ;
        RECT 144.230 168.430 153.100 169.330 ;
        RECT 144.230 167.910 144.460 168.430 ;
        RECT 145.270 168.360 146.280 168.430 ;
        RECT 152.870 167.910 153.100 168.430 ;
        RECT 137.290 167.620 141.290 167.850 ;
        RECT 144.665 167.630 152.665 167.860 ;
        RECT 135.840 167.470 136.970 167.510 ;
        RECT 135.840 167.390 137.210 167.470 ;
        RECT 137.580 167.400 141.240 167.620 ;
        RECT 137.580 167.390 139.020 167.400 ;
        RECT 135.840 167.350 139.020 167.390 ;
        RECT 135.840 167.260 138.530 167.350 ;
        RECT 144.730 167.340 152.620 167.630 ;
        RECT 135.840 167.200 137.860 167.260 ;
        RECT 135.840 167.150 137.610 167.200 ;
        RECT 135.840 163.810 136.670 167.150 ;
        RECT 144.720 166.850 152.640 166.860 ;
        RECT 140.950 166.840 152.640 166.850 ;
        RECT 137.330 166.720 152.640 166.840 ;
        RECT 137.330 166.710 152.665 166.720 ;
        RECT 137.290 166.590 152.665 166.710 ;
        RECT 137.290 166.480 141.290 166.590 ;
        RECT 136.900 166.140 137.130 166.430 ;
        RECT 137.350 166.140 141.240 166.480 ;
        RECT 141.450 166.140 141.680 166.430 ;
        RECT 136.900 164.770 141.680 166.140 ;
        RECT 136.900 164.470 137.130 164.770 ;
        RECT 141.450 164.470 141.680 164.770 ;
        RECT 137.290 164.190 141.290 164.420 ;
        RECT 137.540 163.960 141.110 164.190 ;
        RECT 137.540 163.810 141.230 163.960 ;
        RECT 135.840 163.530 141.230 163.810 ;
        RECT 142.480 163.640 143.100 166.590 ;
        RECT 144.665 166.490 152.665 166.590 ;
        RECT 144.720 166.480 152.640 166.490 ;
        RECT 144.230 165.780 144.460 166.440 ;
        RECT 145.240 165.780 146.240 165.870 ;
        RECT 152.870 165.780 153.100 166.440 ;
        RECT 144.230 164.960 153.100 165.780 ;
        RECT 144.230 164.480 144.460 164.960 ;
        RECT 145.240 164.870 146.240 164.960 ;
        RECT 152.870 164.480 153.100 164.960 ;
        RECT 144.665 164.200 152.665 164.430 ;
        RECT 135.840 163.070 141.240 163.530 ;
        RECT 135.840 161.730 137.840 163.070 ;
        RECT 139.590 163.060 141.240 163.070 ;
        RECT 138.280 161.790 139.280 162.510 ;
        RECT 139.590 162.250 139.900 163.060 ;
        RECT 140.360 162.780 141.240 163.060 ;
        RECT 141.480 163.240 143.100 163.640 ;
        RECT 144.750 163.290 152.620 164.200 ;
        RECT 140.300 162.550 141.300 162.780 ;
        RECT 141.480 162.590 141.830 163.240 ;
        RECT 142.480 163.230 143.100 163.240 ;
        RECT 144.665 163.060 152.665 163.290 ;
        RECT 144.750 163.050 152.620 163.060 ;
        RECT 140.360 162.340 141.240 162.360 ;
        RECT 139.630 161.960 139.900 162.250 ;
        RECT 140.300 162.110 141.300 162.340 ;
        RECT 141.460 162.300 141.830 162.590 ;
        RECT 141.490 162.240 141.830 162.300 ;
        RECT 142.590 162.910 143.350 162.960 ;
        RECT 144.230 162.910 144.460 163.010 ;
        RECT 142.590 162.700 144.460 162.910 ;
        RECT 152.870 162.700 153.100 163.010 ;
        RECT 142.590 162.280 145.130 162.700 ;
        RECT 152.500 162.280 153.100 162.700 ;
        RECT 140.360 161.960 141.240 162.110 ;
        RECT 140.370 161.790 141.100 161.960 ;
        RECT 119.240 160.400 122.240 160.630 ;
        RECT 122.450 160.440 122.790 161.270 ;
        RECT 124.800 161.260 135.440 161.330 ;
        RECT 119.290 160.370 122.150 160.400 ;
        RECT 119.290 160.350 120.460 160.370 ;
        RECT 121.420 160.360 122.150 160.370 ;
        RECT 119.240 159.960 122.240 160.190 ;
        RECT 122.445 160.150 122.790 160.440 ;
        RECT 122.980 160.200 135.440 161.260 ;
        RECT 123.250 160.190 128.690 160.200 ;
        RECT 129.690 160.190 135.440 160.200 ;
        RECT 122.450 160.040 122.790 160.150 ;
        RECT 116.860 155.920 117.720 158.020 ;
        RECT 123.390 157.630 124.640 158.070 ;
        RECT 134.500 158.050 135.440 160.190 ;
        RECT 135.920 161.720 137.840 161.730 ;
        RECT 135.920 158.050 136.640 161.720 ;
        RECT 138.250 160.670 141.100 161.790 ;
        RECT 141.490 161.490 141.840 162.240 ;
        RECT 142.590 162.120 144.460 162.280 ;
        RECT 142.590 162.070 143.350 162.120 ;
        RECT 144.230 162.050 144.460 162.120 ;
        RECT 152.870 162.050 153.100 162.280 ;
        RECT 144.665 161.770 152.665 162.000 ;
        RECT 141.490 161.430 141.780 161.490 ;
        RECT 141.400 161.310 141.780 161.430 ;
        RECT 144.760 161.370 152.620 161.770 ;
        RECT 153.430 161.370 154.390 170.850 ;
        RECT 138.190 160.440 141.190 160.670 ;
        RECT 141.400 160.480 141.740 161.310 ;
        RECT 143.750 161.300 154.390 161.370 ;
        RECT 138.240 160.410 141.100 160.440 ;
        RECT 138.240 160.390 139.410 160.410 ;
        RECT 140.370 160.400 141.100 160.410 ;
        RECT 138.190 160.000 141.190 160.230 ;
        RECT 141.395 160.190 141.740 160.480 ;
        RECT 141.930 161.220 154.390 161.300 ;
        RECT 141.930 160.240 154.420 161.220 ;
        RECT 142.200 160.230 147.640 160.240 ;
        RECT 148.640 160.230 154.420 160.240 ;
        RECT 141.400 160.080 141.740 160.190 ;
        RECT 153.480 159.710 154.420 160.230 ;
        RECT 152.180 158.420 154.420 159.710 ;
        RECT 121.330 157.620 126.570 157.630 ;
        RECT 118.380 157.520 133.680 157.620 ;
        RECT 118.380 157.510 133.715 157.520 ;
        RECT 118.340 157.390 133.715 157.510 ;
        RECT 118.340 157.280 122.340 157.390 ;
        RECT 123.390 157.310 125.130 157.390 ;
        RECT 125.710 157.310 133.715 157.390 ;
        RECT 123.390 157.230 124.640 157.310 ;
        RECT 125.715 157.290 133.715 157.310 ;
        RECT 117.950 156.980 118.180 157.230 ;
        RECT 122.500 157.090 122.730 157.230 ;
        RECT 125.280 157.090 125.510 157.240 ;
        RECT 122.500 156.980 125.510 157.090 ;
        RECT 133.920 156.980 134.150 157.240 ;
        RECT 117.950 156.540 134.150 156.980 ;
        RECT 117.950 156.270 118.180 156.540 ;
        RECT 122.500 156.510 134.150 156.540 ;
        RECT 122.500 156.420 125.510 156.510 ;
        RECT 122.500 156.270 122.730 156.420 ;
        RECT 125.280 156.280 125.510 156.420 ;
        RECT 133.920 156.280 134.150 156.510 ;
        RECT 118.340 155.990 122.340 156.220 ;
        RECT 125.715 156.010 133.715 156.230 ;
        RECT 134.480 156.010 135.440 158.050 ;
        RECT 125.715 156.000 135.440 156.010 ;
        RECT 118.340 155.920 122.330 155.990 ;
        RECT 116.860 155.810 122.330 155.920 ;
        RECT 125.770 155.840 135.440 156.000 ;
        RECT 116.860 155.720 120.020 155.810 ;
        RECT 133.510 155.790 135.440 155.840 ;
        RECT 116.860 152.450 117.720 155.720 ;
        RECT 121.370 155.260 126.620 155.270 ;
        RECT 121.370 155.150 133.680 155.260 ;
        RECT 118.400 155.090 133.680 155.150 ;
        RECT 118.400 155.080 133.715 155.090 ;
        RECT 118.340 154.950 133.715 155.080 ;
        RECT 118.340 154.940 123.500 154.950 ;
        RECT 118.340 154.850 122.340 154.940 ;
        RECT 125.715 154.860 133.715 154.950 ;
        RECT 125.800 154.850 133.690 154.860 ;
        RECT 117.950 154.490 118.180 154.800 ;
        RECT 118.400 154.490 122.300 154.850 ;
        RECT 122.500 154.490 122.730 154.800 ;
        RECT 117.950 153.150 122.730 154.490 ;
        RECT 117.950 152.840 118.180 153.150 ;
        RECT 122.500 152.840 122.730 153.150 ;
        RECT 125.280 154.270 125.510 154.810 ;
        RECT 126.320 154.270 127.330 154.300 ;
        RECT 133.920 154.270 134.150 154.810 ;
        RECT 125.280 153.370 134.150 154.270 ;
        RECT 125.280 152.850 125.510 153.370 ;
        RECT 126.320 153.300 127.330 153.370 ;
        RECT 133.920 152.850 134.150 153.370 ;
        RECT 118.340 152.560 122.340 152.790 ;
        RECT 125.715 152.570 133.715 152.800 ;
        RECT 116.860 152.410 118.020 152.450 ;
        RECT 116.860 152.330 118.260 152.410 ;
        RECT 118.630 152.340 122.290 152.560 ;
        RECT 118.630 152.330 120.070 152.340 ;
        RECT 116.860 152.290 120.070 152.330 ;
        RECT 116.860 152.200 119.580 152.290 ;
        RECT 125.780 152.280 133.670 152.570 ;
        RECT 116.860 152.140 118.910 152.200 ;
        RECT 116.860 152.090 118.660 152.140 ;
        RECT 116.860 148.750 117.720 152.090 ;
        RECT 125.770 151.790 133.690 151.800 ;
        RECT 122.000 151.780 133.690 151.790 ;
        RECT 118.380 151.660 133.690 151.780 ;
        RECT 118.380 151.650 133.715 151.660 ;
        RECT 118.340 151.530 133.715 151.650 ;
        RECT 118.340 151.420 122.340 151.530 ;
        RECT 117.950 151.080 118.180 151.370 ;
        RECT 118.400 151.080 122.290 151.420 ;
        RECT 122.500 151.080 122.730 151.370 ;
        RECT 117.950 149.710 122.730 151.080 ;
        RECT 117.950 149.410 118.180 149.710 ;
        RECT 122.500 149.410 122.730 149.710 ;
        RECT 118.340 149.130 122.340 149.360 ;
        RECT 118.590 148.900 122.160 149.130 ;
        RECT 118.590 148.750 122.280 148.900 ;
        RECT 116.860 148.470 122.280 148.750 ;
        RECT 123.530 148.580 124.150 151.530 ;
        RECT 125.715 151.430 133.715 151.530 ;
        RECT 125.770 151.420 133.690 151.430 ;
        RECT 125.280 150.720 125.510 151.380 ;
        RECT 126.290 150.720 127.290 150.810 ;
        RECT 133.920 150.720 134.150 151.380 ;
        RECT 125.280 149.900 134.150 150.720 ;
        RECT 125.280 149.420 125.510 149.900 ;
        RECT 126.290 149.810 127.290 149.900 ;
        RECT 133.920 149.420 134.150 149.900 ;
        RECT 125.715 149.140 133.715 149.370 ;
        RECT 116.860 148.010 122.290 148.470 ;
        RECT 116.860 146.660 118.890 148.010 ;
        RECT 120.640 148.000 122.290 148.010 ;
        RECT 119.330 146.730 120.330 147.450 ;
        RECT 120.640 147.190 120.950 148.000 ;
        RECT 121.410 147.720 122.290 148.000 ;
        RECT 122.530 148.180 124.150 148.580 ;
        RECT 125.800 148.230 133.670 149.140 ;
        RECT 121.350 147.490 122.350 147.720 ;
        RECT 122.530 147.530 122.880 148.180 ;
        RECT 123.530 148.170 124.150 148.180 ;
        RECT 125.715 148.000 133.715 148.230 ;
        RECT 125.800 147.990 133.670 148.000 ;
        RECT 121.410 147.280 122.290 147.300 ;
        RECT 120.680 146.900 120.950 147.190 ;
        RECT 121.350 147.050 122.350 147.280 ;
        RECT 122.510 147.240 122.880 147.530 ;
        RECT 122.540 147.180 122.880 147.240 ;
        RECT 123.640 147.850 124.400 147.900 ;
        RECT 125.280 147.850 125.510 147.950 ;
        RECT 123.640 147.640 125.510 147.850 ;
        RECT 133.920 147.640 134.150 147.950 ;
        RECT 123.640 147.220 126.180 147.640 ;
        RECT 133.550 147.220 134.150 147.640 ;
        RECT 121.410 146.900 122.290 147.050 ;
        RECT 121.420 146.730 122.150 146.900 ;
        RECT 103.940 145.180 116.330 145.200 ;
        RECT 104.210 145.170 109.650 145.180 ;
        RECT 110.650 145.170 116.330 145.180 ;
        RECT 103.410 145.020 103.750 145.130 ;
        RECT 97.850 143.040 98.640 143.070 ;
        RECT 97.850 140.940 98.680 143.040 ;
        RECT 104.350 142.650 105.600 143.090 ;
        RECT 115.390 143.070 116.330 145.170 ;
        RECT 102.290 142.640 107.530 142.650 ;
        RECT 99.340 142.540 114.640 142.640 ;
        RECT 99.340 142.530 114.675 142.540 ;
        RECT 99.300 142.410 114.675 142.530 ;
        RECT 99.300 142.300 103.300 142.410 ;
        RECT 104.350 142.330 106.090 142.410 ;
        RECT 106.670 142.330 114.675 142.410 ;
        RECT 104.350 142.250 105.600 142.330 ;
        RECT 106.675 142.310 114.675 142.330 ;
        RECT 98.910 142.000 99.140 142.250 ;
        RECT 103.460 142.110 103.690 142.250 ;
        RECT 106.240 142.110 106.470 142.260 ;
        RECT 103.460 142.000 106.470 142.110 ;
        RECT 114.880 142.000 115.110 142.260 ;
        RECT 98.910 141.560 115.110 142.000 ;
        RECT 98.910 141.290 99.140 141.560 ;
        RECT 103.460 141.530 115.110 141.560 ;
        RECT 103.460 141.440 106.470 141.530 ;
        RECT 103.460 141.290 103.690 141.440 ;
        RECT 106.240 141.300 106.470 141.440 ;
        RECT 114.880 141.300 115.110 141.530 ;
        RECT 115.390 141.520 116.400 143.070 ;
        RECT 116.860 143.030 117.620 146.660 ;
        RECT 119.300 145.610 122.150 146.730 ;
        RECT 122.540 146.430 122.890 147.180 ;
        RECT 123.640 147.060 125.510 147.220 ;
        RECT 123.640 147.010 124.400 147.060 ;
        RECT 125.280 146.990 125.510 147.060 ;
        RECT 133.920 146.990 134.150 147.220 ;
        RECT 125.715 146.710 133.715 146.940 ;
        RECT 122.540 146.370 122.830 146.430 ;
        RECT 122.450 146.250 122.830 146.370 ;
        RECT 125.810 146.310 133.670 146.710 ;
        RECT 134.480 146.310 135.440 155.790 ;
        RECT 135.890 158.020 136.640 158.050 ;
        RECT 135.890 155.920 136.720 158.020 ;
        RECT 142.390 157.630 143.640 158.070 ;
        RECT 153.480 158.050 154.420 158.420 ;
        RECT 140.330 157.620 145.570 157.630 ;
        RECT 137.380 157.520 152.680 157.620 ;
        RECT 137.380 157.510 152.715 157.520 ;
        RECT 137.340 157.390 152.715 157.510 ;
        RECT 137.340 157.280 141.340 157.390 ;
        RECT 142.390 157.310 144.130 157.390 ;
        RECT 144.710 157.310 152.715 157.390 ;
        RECT 142.390 157.230 143.640 157.310 ;
        RECT 144.715 157.290 152.715 157.310 ;
        RECT 136.950 156.980 137.180 157.230 ;
        RECT 141.500 157.090 141.730 157.230 ;
        RECT 144.280 157.090 144.510 157.240 ;
        RECT 141.500 156.980 144.510 157.090 ;
        RECT 152.920 156.980 153.150 157.240 ;
        RECT 136.950 156.540 153.150 156.980 ;
        RECT 136.950 156.270 137.180 156.540 ;
        RECT 141.500 156.510 153.150 156.540 ;
        RECT 141.500 156.420 144.510 156.510 ;
        RECT 141.500 156.270 141.730 156.420 ;
        RECT 144.280 156.280 144.510 156.420 ;
        RECT 152.920 156.280 153.150 156.510 ;
        RECT 137.340 155.990 141.340 156.220 ;
        RECT 144.715 156.010 152.715 156.230 ;
        RECT 153.480 156.010 154.440 158.050 ;
        RECT 144.715 156.000 154.440 156.010 ;
        RECT 137.340 155.920 141.330 155.990 ;
        RECT 135.890 155.810 141.330 155.920 ;
        RECT 144.770 155.840 154.440 156.000 ;
        RECT 135.890 155.720 139.020 155.810 ;
        RECT 152.510 155.790 154.440 155.840 ;
        RECT 135.890 152.450 136.720 155.720 ;
        RECT 140.370 155.260 145.620 155.270 ;
        RECT 140.370 155.150 152.680 155.260 ;
        RECT 137.400 155.090 152.680 155.150 ;
        RECT 137.400 155.080 152.715 155.090 ;
        RECT 137.340 154.950 152.715 155.080 ;
        RECT 137.340 154.940 142.500 154.950 ;
        RECT 137.340 154.850 141.340 154.940 ;
        RECT 144.715 154.860 152.715 154.950 ;
        RECT 144.800 154.850 152.690 154.860 ;
        RECT 136.950 154.490 137.180 154.800 ;
        RECT 137.400 154.490 141.300 154.850 ;
        RECT 141.500 154.490 141.730 154.800 ;
        RECT 136.950 153.150 141.730 154.490 ;
        RECT 136.950 152.840 137.180 153.150 ;
        RECT 141.500 152.840 141.730 153.150 ;
        RECT 144.280 154.270 144.510 154.810 ;
        RECT 145.320 154.270 146.330 154.300 ;
        RECT 152.920 154.270 153.150 154.810 ;
        RECT 144.280 153.370 153.150 154.270 ;
        RECT 144.280 152.850 144.510 153.370 ;
        RECT 145.320 153.300 146.330 153.370 ;
        RECT 152.920 152.850 153.150 153.370 ;
        RECT 137.340 152.560 141.340 152.790 ;
        RECT 144.715 152.570 152.715 152.800 ;
        RECT 135.890 152.410 137.020 152.450 ;
        RECT 135.890 152.330 137.260 152.410 ;
        RECT 137.630 152.340 141.290 152.560 ;
        RECT 137.630 152.330 139.070 152.340 ;
        RECT 135.890 152.290 139.070 152.330 ;
        RECT 135.890 152.200 138.580 152.290 ;
        RECT 144.780 152.280 152.670 152.570 ;
        RECT 135.890 152.140 137.910 152.200 ;
        RECT 135.890 152.090 137.660 152.140 ;
        RECT 135.890 148.750 136.720 152.090 ;
        RECT 144.770 151.790 152.690 151.800 ;
        RECT 141.000 151.780 152.690 151.790 ;
        RECT 137.380 151.660 152.690 151.780 ;
        RECT 137.380 151.650 152.715 151.660 ;
        RECT 137.340 151.530 152.715 151.650 ;
        RECT 137.340 151.420 141.340 151.530 ;
        RECT 136.950 151.080 137.180 151.370 ;
        RECT 137.400 151.080 141.290 151.420 ;
        RECT 141.500 151.080 141.730 151.370 ;
        RECT 136.950 149.710 141.730 151.080 ;
        RECT 136.950 149.410 137.180 149.710 ;
        RECT 141.500 149.410 141.730 149.710 ;
        RECT 137.340 149.130 141.340 149.360 ;
        RECT 137.590 148.900 141.160 149.130 ;
        RECT 137.590 148.750 141.280 148.900 ;
        RECT 135.890 148.470 141.280 148.750 ;
        RECT 142.530 148.580 143.150 151.530 ;
        RECT 144.715 151.430 152.715 151.530 ;
        RECT 144.770 151.420 152.690 151.430 ;
        RECT 144.280 150.720 144.510 151.380 ;
        RECT 145.290 150.720 146.290 150.810 ;
        RECT 152.920 150.720 153.150 151.380 ;
        RECT 144.280 149.900 153.150 150.720 ;
        RECT 144.280 149.420 144.510 149.900 ;
        RECT 145.290 149.810 146.290 149.900 ;
        RECT 152.920 149.420 153.150 149.900 ;
        RECT 144.715 149.140 152.715 149.370 ;
        RECT 135.890 148.010 141.290 148.470 ;
        RECT 135.890 146.670 137.890 148.010 ;
        RECT 139.640 148.000 141.290 148.010 ;
        RECT 138.330 146.730 139.330 147.450 ;
        RECT 139.640 147.190 139.950 148.000 ;
        RECT 140.410 147.720 141.290 148.000 ;
        RECT 141.530 148.180 143.150 148.580 ;
        RECT 144.800 148.230 152.670 149.140 ;
        RECT 140.350 147.490 141.350 147.720 ;
        RECT 141.530 147.530 141.880 148.180 ;
        RECT 142.530 148.170 143.150 148.180 ;
        RECT 144.715 148.000 152.715 148.230 ;
        RECT 144.800 147.990 152.670 148.000 ;
        RECT 140.410 147.280 141.290 147.300 ;
        RECT 139.680 146.900 139.950 147.190 ;
        RECT 140.350 147.050 141.350 147.280 ;
        RECT 141.510 147.240 141.880 147.530 ;
        RECT 141.540 147.180 141.880 147.240 ;
        RECT 142.640 147.850 143.400 147.900 ;
        RECT 144.280 147.850 144.510 147.950 ;
        RECT 142.640 147.640 144.510 147.850 ;
        RECT 152.920 147.640 153.150 147.950 ;
        RECT 142.640 147.220 145.180 147.640 ;
        RECT 152.550 147.220 153.150 147.640 ;
        RECT 140.410 146.900 141.290 147.050 ;
        RECT 140.420 146.730 141.150 146.900 ;
        RECT 119.240 145.380 122.240 145.610 ;
        RECT 122.450 145.420 122.790 146.250 ;
        RECT 124.800 146.240 135.440 146.310 ;
        RECT 119.290 145.350 122.150 145.380 ;
        RECT 119.290 145.330 120.460 145.350 ;
        RECT 121.420 145.340 122.150 145.350 ;
        RECT 119.240 144.940 122.240 145.170 ;
        RECT 122.445 145.130 122.790 145.420 ;
        RECT 122.980 145.200 135.440 146.240 ;
        RECT 135.910 146.660 137.890 146.670 ;
        RECT 122.980 145.180 135.380 145.200 ;
        RECT 123.250 145.170 128.690 145.180 ;
        RECT 129.690 145.170 135.380 145.180 ;
        RECT 122.450 145.020 122.790 145.130 ;
        RECT 99.300 141.010 103.300 141.240 ;
        RECT 106.675 141.030 114.675 141.250 ;
        RECT 115.440 141.030 116.400 141.520 ;
        RECT 106.675 141.020 116.400 141.030 ;
        RECT 99.300 140.940 103.290 141.010 ;
        RECT 97.850 140.830 103.290 140.940 ;
        RECT 106.730 140.860 116.400 141.020 ;
        RECT 97.850 140.740 100.980 140.830 ;
        RECT 114.470 140.810 116.400 140.860 ;
        RECT 97.850 137.470 98.680 140.740 ;
        RECT 102.330 140.280 107.580 140.290 ;
        RECT 102.330 140.170 114.640 140.280 ;
        RECT 99.360 140.110 114.640 140.170 ;
        RECT 99.360 140.100 114.675 140.110 ;
        RECT 99.300 139.970 114.675 140.100 ;
        RECT 99.300 139.960 104.460 139.970 ;
        RECT 99.300 139.870 103.300 139.960 ;
        RECT 106.675 139.880 114.675 139.970 ;
        RECT 106.760 139.870 114.650 139.880 ;
        RECT 98.910 139.510 99.140 139.820 ;
        RECT 99.360 139.510 103.260 139.870 ;
        RECT 103.460 139.510 103.690 139.820 ;
        RECT 98.910 138.170 103.690 139.510 ;
        RECT 98.910 137.860 99.140 138.170 ;
        RECT 103.460 137.860 103.690 138.170 ;
        RECT 106.240 139.290 106.470 139.830 ;
        RECT 107.280 139.290 108.290 139.320 ;
        RECT 114.880 139.290 115.110 139.830 ;
        RECT 106.240 138.390 115.110 139.290 ;
        RECT 106.240 137.870 106.470 138.390 ;
        RECT 107.280 138.320 108.290 138.390 ;
        RECT 114.880 137.870 115.110 138.390 ;
        RECT 99.300 137.580 103.300 137.810 ;
        RECT 106.675 137.590 114.675 137.820 ;
        RECT 97.850 137.430 98.980 137.470 ;
        RECT 97.850 137.350 99.220 137.430 ;
        RECT 99.590 137.360 103.250 137.580 ;
        RECT 99.590 137.350 101.030 137.360 ;
        RECT 97.850 137.310 101.030 137.350 ;
        RECT 97.850 137.220 100.540 137.310 ;
        RECT 106.740 137.300 114.630 137.590 ;
        RECT 97.850 137.160 99.870 137.220 ;
        RECT 97.850 137.110 99.620 137.160 ;
        RECT 97.850 133.770 98.680 137.110 ;
        RECT 106.730 136.810 114.650 136.820 ;
        RECT 102.960 136.800 114.650 136.810 ;
        RECT 99.340 136.680 114.650 136.800 ;
        RECT 99.340 136.670 114.675 136.680 ;
        RECT 99.300 136.550 114.675 136.670 ;
        RECT 99.300 136.440 103.300 136.550 ;
        RECT 98.910 136.100 99.140 136.390 ;
        RECT 99.360 136.100 103.250 136.440 ;
        RECT 103.460 136.100 103.690 136.390 ;
        RECT 98.910 134.730 103.690 136.100 ;
        RECT 98.910 134.430 99.140 134.730 ;
        RECT 103.460 134.430 103.690 134.730 ;
        RECT 99.300 134.150 103.300 134.380 ;
        RECT 99.550 133.920 103.120 134.150 ;
        RECT 99.550 133.770 103.240 133.920 ;
        RECT 97.850 133.490 103.240 133.770 ;
        RECT 104.490 133.600 105.110 136.550 ;
        RECT 106.675 136.450 114.675 136.550 ;
        RECT 106.730 136.440 114.650 136.450 ;
        RECT 106.240 135.740 106.470 136.400 ;
        RECT 107.250 135.740 108.250 135.830 ;
        RECT 114.880 135.740 115.110 136.400 ;
        RECT 106.240 134.920 115.110 135.740 ;
        RECT 106.240 134.440 106.470 134.920 ;
        RECT 107.250 134.830 108.250 134.920 ;
        RECT 114.880 134.440 115.110 134.920 ;
        RECT 106.675 134.160 114.675 134.390 ;
        RECT 97.850 133.030 103.250 133.490 ;
        RECT 97.850 131.690 99.850 133.030 ;
        RECT 101.600 133.020 103.250 133.030 ;
        RECT 100.290 131.750 101.290 132.470 ;
        RECT 101.600 132.210 101.910 133.020 ;
        RECT 102.370 132.740 103.250 133.020 ;
        RECT 103.490 133.200 105.110 133.600 ;
        RECT 106.760 133.250 114.630 134.160 ;
        RECT 102.310 132.510 103.310 132.740 ;
        RECT 103.490 132.550 103.840 133.200 ;
        RECT 104.490 133.190 105.110 133.200 ;
        RECT 106.675 133.020 114.675 133.250 ;
        RECT 106.760 133.010 114.630 133.020 ;
        RECT 102.370 132.300 103.250 132.320 ;
        RECT 101.640 131.920 101.910 132.210 ;
        RECT 102.310 132.070 103.310 132.300 ;
        RECT 103.470 132.260 103.840 132.550 ;
        RECT 103.500 132.200 103.840 132.260 ;
        RECT 104.600 132.870 105.360 132.920 ;
        RECT 106.240 132.870 106.470 132.970 ;
        RECT 104.600 132.660 106.470 132.870 ;
        RECT 114.880 132.660 115.110 132.970 ;
        RECT 104.600 132.240 107.140 132.660 ;
        RECT 114.510 132.240 115.110 132.660 ;
        RECT 102.370 131.920 103.250 132.070 ;
        RECT 102.380 131.750 103.110 131.920 ;
        RECT 97.860 131.680 99.850 131.690 ;
        RECT 97.860 128.040 98.640 131.680 ;
        RECT 100.260 130.630 103.110 131.750 ;
        RECT 103.500 131.450 103.850 132.200 ;
        RECT 104.600 132.080 106.470 132.240 ;
        RECT 104.600 132.030 105.360 132.080 ;
        RECT 106.240 132.010 106.470 132.080 ;
        RECT 114.880 132.010 115.110 132.240 ;
        RECT 106.675 131.730 114.675 131.960 ;
        RECT 103.500 131.390 103.790 131.450 ;
        RECT 103.410 131.270 103.790 131.390 ;
        RECT 106.770 131.330 114.630 131.730 ;
        RECT 115.440 131.510 116.400 140.810 ;
        RECT 116.840 143.000 117.620 143.030 ;
        RECT 116.840 140.900 117.670 143.000 ;
        RECT 123.340 142.610 124.590 143.050 ;
        RECT 134.440 143.030 135.380 145.170 ;
        RECT 135.910 143.030 136.610 146.660 ;
        RECT 138.300 145.610 141.150 146.730 ;
        RECT 141.540 146.430 141.890 147.180 ;
        RECT 142.640 147.060 144.510 147.220 ;
        RECT 142.640 147.010 143.400 147.060 ;
        RECT 144.280 146.990 144.510 147.060 ;
        RECT 152.920 146.990 153.150 147.220 ;
        RECT 144.715 146.710 152.715 146.940 ;
        RECT 141.540 146.370 141.830 146.430 ;
        RECT 141.450 146.250 141.830 146.370 ;
        RECT 144.810 146.310 152.670 146.710 ;
        RECT 153.480 146.310 154.440 155.790 ;
        RECT 138.240 145.380 141.240 145.610 ;
        RECT 141.450 145.420 141.790 146.250 ;
        RECT 143.800 146.240 154.440 146.310 ;
        RECT 138.290 145.350 141.150 145.380 ;
        RECT 138.290 145.330 139.460 145.350 ;
        RECT 140.420 145.340 141.150 145.350 ;
        RECT 138.240 144.940 141.240 145.170 ;
        RECT 141.445 145.130 141.790 145.420 ;
        RECT 141.980 145.200 154.440 146.240 ;
        RECT 141.980 145.180 154.360 145.200 ;
        RECT 142.250 145.170 147.690 145.180 ;
        RECT 148.690 145.170 154.360 145.180 ;
        RECT 141.450 145.020 141.790 145.130 ;
        RECT 121.280 142.600 126.520 142.610 ;
        RECT 118.330 142.500 133.630 142.600 ;
        RECT 118.330 142.490 133.665 142.500 ;
        RECT 118.290 142.370 133.665 142.490 ;
        RECT 118.290 142.260 122.290 142.370 ;
        RECT 123.340 142.290 125.080 142.370 ;
        RECT 125.660 142.290 133.665 142.370 ;
        RECT 123.340 142.210 124.590 142.290 ;
        RECT 125.665 142.270 133.665 142.290 ;
        RECT 117.900 141.960 118.130 142.210 ;
        RECT 122.450 142.070 122.680 142.210 ;
        RECT 125.230 142.070 125.460 142.220 ;
        RECT 122.450 141.960 125.460 142.070 ;
        RECT 133.870 141.960 134.100 142.220 ;
        RECT 117.900 141.520 134.100 141.960 ;
        RECT 117.900 141.250 118.130 141.520 ;
        RECT 122.450 141.490 134.100 141.520 ;
        RECT 122.450 141.400 125.460 141.490 ;
        RECT 122.450 141.250 122.680 141.400 ;
        RECT 125.230 141.260 125.460 141.400 ;
        RECT 133.870 141.260 134.100 141.490 ;
        RECT 118.290 140.970 122.290 141.200 ;
        RECT 125.665 140.990 133.665 141.210 ;
        RECT 134.430 140.990 135.390 143.030 ;
        RECT 125.665 140.980 135.390 140.990 ;
        RECT 118.290 140.900 122.280 140.970 ;
        RECT 116.840 140.790 122.280 140.900 ;
        RECT 125.720 140.820 135.390 140.980 ;
        RECT 116.840 140.700 119.970 140.790 ;
        RECT 133.460 140.770 135.390 140.820 ;
        RECT 116.840 137.430 117.670 140.700 ;
        RECT 121.320 140.240 126.570 140.250 ;
        RECT 121.320 140.130 133.630 140.240 ;
        RECT 118.350 140.070 133.630 140.130 ;
        RECT 118.350 140.060 133.665 140.070 ;
        RECT 118.290 139.930 133.665 140.060 ;
        RECT 118.290 139.920 123.450 139.930 ;
        RECT 118.290 139.830 122.290 139.920 ;
        RECT 125.665 139.840 133.665 139.930 ;
        RECT 125.750 139.830 133.640 139.840 ;
        RECT 117.900 139.470 118.130 139.780 ;
        RECT 118.350 139.470 122.250 139.830 ;
        RECT 122.450 139.470 122.680 139.780 ;
        RECT 117.900 138.130 122.680 139.470 ;
        RECT 117.900 137.820 118.130 138.130 ;
        RECT 122.450 137.820 122.680 138.130 ;
        RECT 125.230 139.250 125.460 139.790 ;
        RECT 126.270 139.250 127.280 139.280 ;
        RECT 133.870 139.250 134.100 139.790 ;
        RECT 125.230 138.350 134.100 139.250 ;
        RECT 125.230 137.830 125.460 138.350 ;
        RECT 126.270 138.280 127.280 138.350 ;
        RECT 133.870 137.830 134.100 138.350 ;
        RECT 118.290 137.540 122.290 137.770 ;
        RECT 125.665 137.550 133.665 137.780 ;
        RECT 116.840 137.390 117.970 137.430 ;
        RECT 116.840 137.310 118.210 137.390 ;
        RECT 118.580 137.320 122.240 137.540 ;
        RECT 118.580 137.310 120.020 137.320 ;
        RECT 116.840 137.270 120.020 137.310 ;
        RECT 116.840 137.180 119.530 137.270 ;
        RECT 125.730 137.260 133.620 137.550 ;
        RECT 116.840 137.120 118.860 137.180 ;
        RECT 116.840 137.070 118.610 137.120 ;
        RECT 116.840 133.730 117.670 137.070 ;
        RECT 125.720 136.770 133.640 136.780 ;
        RECT 121.950 136.760 133.640 136.770 ;
        RECT 118.330 136.640 133.640 136.760 ;
        RECT 118.330 136.630 133.665 136.640 ;
        RECT 118.290 136.510 133.665 136.630 ;
        RECT 118.290 136.400 122.290 136.510 ;
        RECT 117.900 136.060 118.130 136.350 ;
        RECT 118.350 136.060 122.240 136.400 ;
        RECT 122.450 136.060 122.680 136.350 ;
        RECT 117.900 134.690 122.680 136.060 ;
        RECT 117.900 134.390 118.130 134.690 ;
        RECT 122.450 134.390 122.680 134.690 ;
        RECT 118.290 134.110 122.290 134.340 ;
        RECT 118.540 133.880 122.110 134.110 ;
        RECT 118.540 133.730 122.230 133.880 ;
        RECT 116.840 133.450 122.230 133.730 ;
        RECT 123.480 133.560 124.100 136.510 ;
        RECT 125.665 136.410 133.665 136.510 ;
        RECT 125.720 136.400 133.640 136.410 ;
        RECT 125.230 135.700 125.460 136.360 ;
        RECT 126.240 135.700 127.240 135.790 ;
        RECT 133.870 135.700 134.100 136.360 ;
        RECT 125.230 134.880 134.100 135.700 ;
        RECT 125.230 134.400 125.460 134.880 ;
        RECT 126.240 134.790 127.240 134.880 ;
        RECT 133.870 134.400 134.100 134.880 ;
        RECT 125.665 134.120 133.665 134.350 ;
        RECT 116.840 132.990 122.240 133.450 ;
        RECT 116.840 131.650 118.840 132.990 ;
        RECT 120.590 132.980 122.240 132.990 ;
        RECT 119.280 131.710 120.280 132.430 ;
        RECT 120.590 132.170 120.900 132.980 ;
        RECT 121.360 132.700 122.240 132.980 ;
        RECT 122.480 133.160 124.100 133.560 ;
        RECT 125.750 133.210 133.620 134.120 ;
        RECT 121.300 132.470 122.300 132.700 ;
        RECT 122.480 132.510 122.830 133.160 ;
        RECT 123.480 133.150 124.100 133.160 ;
        RECT 125.665 132.980 133.665 133.210 ;
        RECT 125.750 132.970 133.620 132.980 ;
        RECT 121.360 132.260 122.240 132.280 ;
        RECT 120.630 131.880 120.900 132.170 ;
        RECT 121.300 132.030 122.300 132.260 ;
        RECT 122.460 132.220 122.830 132.510 ;
        RECT 122.490 132.160 122.830 132.220 ;
        RECT 123.590 132.830 124.350 132.880 ;
        RECT 125.230 132.830 125.460 132.930 ;
        RECT 123.590 132.620 125.460 132.830 ;
        RECT 133.870 132.620 134.100 132.930 ;
        RECT 123.590 132.200 126.130 132.620 ;
        RECT 133.500 132.200 134.100 132.620 ;
        RECT 121.360 131.880 122.240 132.030 ;
        RECT 121.370 131.710 122.100 131.880 ;
        RECT 115.430 131.330 116.400 131.510 ;
        RECT 100.200 130.400 103.200 130.630 ;
        RECT 103.410 130.440 103.750 131.270 ;
        RECT 105.760 131.260 116.400 131.330 ;
        RECT 100.250 130.370 103.110 130.400 ;
        RECT 100.250 130.350 101.420 130.370 ;
        RECT 102.380 130.360 103.110 130.370 ;
        RECT 100.200 129.960 103.200 130.190 ;
        RECT 103.405 130.150 103.750 130.440 ;
        RECT 103.940 130.220 116.400 131.260 ;
        RECT 116.860 131.640 118.840 131.650 ;
        RECT 103.940 130.200 116.370 130.220 ;
        RECT 104.210 130.190 109.650 130.200 ;
        RECT 110.650 130.190 116.370 130.200 ;
        RECT 103.410 130.040 103.750 130.150 ;
        RECT 97.850 128.010 98.640 128.040 ;
        RECT 97.850 125.910 98.680 128.010 ;
        RECT 104.350 127.620 105.600 128.060 ;
        RECT 115.430 128.040 116.370 130.190 ;
        RECT 102.290 127.610 107.530 127.620 ;
        RECT 99.340 127.510 114.640 127.610 ;
        RECT 99.340 127.500 114.675 127.510 ;
        RECT 99.300 127.380 114.675 127.500 ;
        RECT 99.300 127.270 103.300 127.380 ;
        RECT 104.350 127.300 106.090 127.380 ;
        RECT 106.670 127.300 114.675 127.380 ;
        RECT 104.350 127.220 105.600 127.300 ;
        RECT 106.675 127.280 114.675 127.300 ;
        RECT 98.910 126.970 99.140 127.220 ;
        RECT 103.460 127.080 103.690 127.220 ;
        RECT 106.240 127.080 106.470 127.230 ;
        RECT 103.460 126.970 106.470 127.080 ;
        RECT 114.880 126.970 115.110 127.230 ;
        RECT 98.910 126.530 115.110 126.970 ;
        RECT 115.430 126.530 116.400 128.040 ;
        RECT 116.860 128.010 117.620 131.640 ;
        RECT 119.250 130.590 122.100 131.710 ;
        RECT 122.490 131.410 122.840 132.160 ;
        RECT 123.590 132.040 125.460 132.200 ;
        RECT 123.590 131.990 124.350 132.040 ;
        RECT 125.230 131.970 125.460 132.040 ;
        RECT 133.870 131.970 134.100 132.200 ;
        RECT 125.665 131.690 133.665 131.920 ;
        RECT 122.490 131.350 122.780 131.410 ;
        RECT 122.400 131.230 122.780 131.350 ;
        RECT 125.760 131.290 133.620 131.690 ;
        RECT 134.430 131.290 135.390 140.770 ;
        RECT 135.840 143.000 136.610 143.030 ;
        RECT 135.840 140.900 136.670 143.000 ;
        RECT 142.340 142.610 143.590 143.050 ;
        RECT 153.420 143.030 154.360 145.170 ;
        RECT 140.280 142.600 145.520 142.610 ;
        RECT 137.330 142.500 152.630 142.600 ;
        RECT 137.330 142.490 152.665 142.500 ;
        RECT 137.290 142.370 152.665 142.490 ;
        RECT 137.290 142.260 141.290 142.370 ;
        RECT 142.340 142.290 144.080 142.370 ;
        RECT 144.660 142.290 152.665 142.370 ;
        RECT 142.340 142.210 143.590 142.290 ;
        RECT 144.665 142.270 152.665 142.290 ;
        RECT 136.900 141.960 137.130 142.210 ;
        RECT 141.450 142.070 141.680 142.210 ;
        RECT 144.230 142.070 144.460 142.220 ;
        RECT 141.450 141.960 144.460 142.070 ;
        RECT 152.870 141.960 153.100 142.220 ;
        RECT 136.900 141.520 153.100 141.960 ;
        RECT 136.900 141.250 137.130 141.520 ;
        RECT 141.450 141.490 153.100 141.520 ;
        RECT 141.450 141.400 144.460 141.490 ;
        RECT 141.450 141.250 141.680 141.400 ;
        RECT 144.230 141.260 144.460 141.400 ;
        RECT 152.870 141.260 153.100 141.490 ;
        RECT 153.420 141.260 154.390 143.030 ;
        RECT 137.290 140.970 141.290 141.200 ;
        RECT 144.665 140.990 152.665 141.210 ;
        RECT 153.430 140.990 154.390 141.260 ;
        RECT 144.665 140.980 154.390 140.990 ;
        RECT 137.290 140.900 141.280 140.970 ;
        RECT 135.840 140.790 141.280 140.900 ;
        RECT 144.720 140.820 154.390 140.980 ;
        RECT 135.840 140.700 138.970 140.790 ;
        RECT 152.460 140.770 154.390 140.820 ;
        RECT 135.840 137.430 136.670 140.700 ;
        RECT 140.320 140.240 145.570 140.250 ;
        RECT 140.320 140.130 152.630 140.240 ;
        RECT 137.350 140.070 152.630 140.130 ;
        RECT 137.350 140.060 152.665 140.070 ;
        RECT 137.290 139.930 152.665 140.060 ;
        RECT 137.290 139.920 142.450 139.930 ;
        RECT 137.290 139.830 141.290 139.920 ;
        RECT 144.665 139.840 152.665 139.930 ;
        RECT 144.750 139.830 152.640 139.840 ;
        RECT 136.900 139.470 137.130 139.780 ;
        RECT 137.350 139.470 141.250 139.830 ;
        RECT 141.450 139.470 141.680 139.780 ;
        RECT 136.900 138.130 141.680 139.470 ;
        RECT 136.900 137.820 137.130 138.130 ;
        RECT 141.450 137.820 141.680 138.130 ;
        RECT 144.230 139.250 144.460 139.790 ;
        RECT 145.270 139.250 146.280 139.280 ;
        RECT 152.870 139.250 153.100 139.790 ;
        RECT 144.230 138.350 153.100 139.250 ;
        RECT 144.230 137.830 144.460 138.350 ;
        RECT 145.270 138.280 146.280 138.350 ;
        RECT 152.870 137.830 153.100 138.350 ;
        RECT 137.290 137.540 141.290 137.770 ;
        RECT 144.665 137.550 152.665 137.780 ;
        RECT 135.840 137.390 136.970 137.430 ;
        RECT 135.840 137.310 137.210 137.390 ;
        RECT 137.580 137.320 141.240 137.540 ;
        RECT 137.580 137.310 139.020 137.320 ;
        RECT 135.840 137.270 139.020 137.310 ;
        RECT 135.840 137.180 138.530 137.270 ;
        RECT 144.730 137.260 152.620 137.550 ;
        RECT 135.840 137.120 137.860 137.180 ;
        RECT 135.840 137.070 137.610 137.120 ;
        RECT 135.840 133.730 136.670 137.070 ;
        RECT 144.720 136.770 152.640 136.780 ;
        RECT 140.950 136.760 152.640 136.770 ;
        RECT 137.330 136.640 152.640 136.760 ;
        RECT 137.330 136.630 152.665 136.640 ;
        RECT 137.290 136.510 152.665 136.630 ;
        RECT 137.290 136.400 141.290 136.510 ;
        RECT 136.900 136.060 137.130 136.350 ;
        RECT 137.350 136.060 141.240 136.400 ;
        RECT 141.450 136.060 141.680 136.350 ;
        RECT 136.900 134.690 141.680 136.060 ;
        RECT 136.900 134.390 137.130 134.690 ;
        RECT 141.450 134.390 141.680 134.690 ;
        RECT 137.290 134.110 141.290 134.340 ;
        RECT 137.540 133.880 141.110 134.110 ;
        RECT 137.540 133.730 141.230 133.880 ;
        RECT 135.840 133.450 141.230 133.730 ;
        RECT 142.480 133.560 143.100 136.510 ;
        RECT 144.665 136.410 152.665 136.510 ;
        RECT 144.720 136.400 152.640 136.410 ;
        RECT 144.230 135.700 144.460 136.360 ;
        RECT 145.240 135.700 146.240 135.790 ;
        RECT 152.870 135.700 153.100 136.360 ;
        RECT 144.230 134.880 153.100 135.700 ;
        RECT 144.230 134.400 144.460 134.880 ;
        RECT 145.240 134.790 146.240 134.880 ;
        RECT 152.870 134.400 153.100 134.880 ;
        RECT 144.665 134.120 152.665 134.350 ;
        RECT 135.840 132.990 141.240 133.450 ;
        RECT 135.840 131.650 137.840 132.990 ;
        RECT 139.590 132.980 141.240 132.990 ;
        RECT 138.280 131.710 139.280 132.430 ;
        RECT 139.590 132.170 139.900 132.980 ;
        RECT 140.360 132.700 141.240 132.980 ;
        RECT 141.480 133.160 143.100 133.560 ;
        RECT 144.750 133.210 152.620 134.120 ;
        RECT 140.300 132.470 141.300 132.700 ;
        RECT 141.480 132.510 141.830 133.160 ;
        RECT 142.480 133.150 143.100 133.160 ;
        RECT 144.665 132.980 152.665 133.210 ;
        RECT 144.750 132.970 152.620 132.980 ;
        RECT 140.360 132.260 141.240 132.280 ;
        RECT 139.630 131.880 139.900 132.170 ;
        RECT 140.300 132.030 141.300 132.260 ;
        RECT 141.460 132.220 141.830 132.510 ;
        RECT 141.490 132.160 141.830 132.220 ;
        RECT 142.590 132.830 143.350 132.880 ;
        RECT 144.230 132.830 144.460 132.930 ;
        RECT 142.590 132.620 144.460 132.830 ;
        RECT 152.870 132.620 153.100 132.930 ;
        RECT 142.590 132.200 145.130 132.620 ;
        RECT 152.500 132.200 153.100 132.620 ;
        RECT 140.360 131.880 141.240 132.030 ;
        RECT 140.370 131.710 141.100 131.880 ;
        RECT 119.190 130.360 122.190 130.590 ;
        RECT 122.400 130.400 122.740 131.230 ;
        RECT 124.750 131.220 135.390 131.290 ;
        RECT 119.240 130.330 122.100 130.360 ;
        RECT 119.240 130.310 120.410 130.330 ;
        RECT 121.370 130.320 122.100 130.330 ;
        RECT 119.190 129.920 122.190 130.150 ;
        RECT 122.395 130.110 122.740 130.400 ;
        RECT 122.930 130.180 135.390 131.220 ;
        RECT 135.910 131.640 137.840 131.650 ;
        RECT 122.930 130.160 135.380 130.180 ;
        RECT 123.200 130.150 128.640 130.160 ;
        RECT 129.640 130.150 135.380 130.160 ;
        RECT 122.400 130.000 122.740 130.110 ;
        RECT 98.910 126.260 99.140 126.530 ;
        RECT 103.460 126.500 115.110 126.530 ;
        RECT 103.460 126.410 106.470 126.500 ;
        RECT 103.460 126.260 103.690 126.410 ;
        RECT 106.240 126.270 106.470 126.410 ;
        RECT 114.880 126.270 115.110 126.500 ;
        RECT 99.300 125.980 103.300 126.210 ;
        RECT 106.675 126.000 114.675 126.220 ;
        RECT 115.440 126.000 116.400 126.530 ;
        RECT 106.675 125.990 116.400 126.000 ;
        RECT 99.300 125.910 103.290 125.980 ;
        RECT 97.850 125.800 103.290 125.910 ;
        RECT 106.730 125.830 116.400 125.990 ;
        RECT 97.850 125.710 100.980 125.800 ;
        RECT 114.470 125.780 116.400 125.830 ;
        RECT 97.850 122.440 98.680 125.710 ;
        RECT 102.330 125.250 107.580 125.260 ;
        RECT 102.330 125.140 114.640 125.250 ;
        RECT 99.360 125.080 114.640 125.140 ;
        RECT 99.360 125.070 114.675 125.080 ;
        RECT 99.300 124.940 114.675 125.070 ;
        RECT 99.300 124.930 104.460 124.940 ;
        RECT 99.300 124.840 103.300 124.930 ;
        RECT 106.675 124.850 114.675 124.940 ;
        RECT 106.760 124.840 114.650 124.850 ;
        RECT 98.910 124.480 99.140 124.790 ;
        RECT 99.360 124.480 103.260 124.840 ;
        RECT 103.460 124.480 103.690 124.790 ;
        RECT 98.910 123.140 103.690 124.480 ;
        RECT 98.910 122.830 99.140 123.140 ;
        RECT 103.460 122.830 103.690 123.140 ;
        RECT 106.240 124.260 106.470 124.800 ;
        RECT 107.280 124.260 108.290 124.290 ;
        RECT 114.880 124.260 115.110 124.800 ;
        RECT 106.240 123.360 115.110 124.260 ;
        RECT 106.240 122.840 106.470 123.360 ;
        RECT 107.280 123.290 108.290 123.360 ;
        RECT 114.880 122.840 115.110 123.360 ;
        RECT 99.300 122.550 103.300 122.780 ;
        RECT 106.675 122.560 114.675 122.790 ;
        RECT 97.850 122.400 98.980 122.440 ;
        RECT 97.850 122.320 99.220 122.400 ;
        RECT 99.590 122.330 103.250 122.550 ;
        RECT 99.590 122.320 101.030 122.330 ;
        RECT 97.850 122.280 101.030 122.320 ;
        RECT 97.850 122.190 100.540 122.280 ;
        RECT 106.740 122.270 114.630 122.560 ;
        RECT 97.850 122.130 99.870 122.190 ;
        RECT 97.850 122.080 99.620 122.130 ;
        RECT 97.850 118.740 98.680 122.080 ;
        RECT 106.730 121.780 114.650 121.790 ;
        RECT 102.960 121.770 114.650 121.780 ;
        RECT 99.340 121.650 114.650 121.770 ;
        RECT 99.340 121.640 114.675 121.650 ;
        RECT 99.300 121.520 114.675 121.640 ;
        RECT 99.300 121.410 103.300 121.520 ;
        RECT 98.910 121.070 99.140 121.360 ;
        RECT 99.360 121.070 103.250 121.410 ;
        RECT 103.460 121.070 103.690 121.360 ;
        RECT 98.910 119.700 103.690 121.070 ;
        RECT 98.910 119.400 99.140 119.700 ;
        RECT 103.460 119.400 103.690 119.700 ;
        RECT 99.300 119.120 103.300 119.350 ;
        RECT 99.550 118.890 103.120 119.120 ;
        RECT 99.550 118.740 103.240 118.890 ;
        RECT 97.850 118.460 103.240 118.740 ;
        RECT 104.490 118.570 105.110 121.520 ;
        RECT 106.675 121.420 114.675 121.520 ;
        RECT 106.730 121.410 114.650 121.420 ;
        RECT 106.240 120.710 106.470 121.370 ;
        RECT 107.250 120.710 108.250 120.800 ;
        RECT 114.880 120.710 115.110 121.370 ;
        RECT 106.240 119.890 115.110 120.710 ;
        RECT 106.240 119.410 106.470 119.890 ;
        RECT 107.250 119.800 108.250 119.890 ;
        RECT 114.880 119.410 115.110 119.890 ;
        RECT 106.675 119.130 114.675 119.360 ;
        RECT 97.850 118.000 103.250 118.460 ;
        RECT 97.850 116.660 99.850 118.000 ;
        RECT 101.600 117.990 103.250 118.000 ;
        RECT 100.290 116.720 101.290 117.440 ;
        RECT 101.600 117.180 101.910 117.990 ;
        RECT 102.370 117.710 103.250 117.990 ;
        RECT 103.490 118.170 105.110 118.570 ;
        RECT 106.760 118.220 114.630 119.130 ;
        RECT 102.310 117.480 103.310 117.710 ;
        RECT 103.490 117.520 103.840 118.170 ;
        RECT 104.490 118.160 105.110 118.170 ;
        RECT 106.675 117.990 114.675 118.220 ;
        RECT 106.760 117.980 114.630 117.990 ;
        RECT 102.370 117.270 103.250 117.290 ;
        RECT 101.640 116.890 101.910 117.180 ;
        RECT 102.310 117.040 103.310 117.270 ;
        RECT 103.470 117.230 103.840 117.520 ;
        RECT 103.500 117.170 103.840 117.230 ;
        RECT 104.600 117.840 105.360 117.890 ;
        RECT 106.240 117.840 106.470 117.940 ;
        RECT 104.600 117.630 106.470 117.840 ;
        RECT 114.880 117.630 115.110 117.940 ;
        RECT 104.600 117.210 107.140 117.630 ;
        RECT 114.510 117.210 115.110 117.630 ;
        RECT 102.370 116.890 103.250 117.040 ;
        RECT 102.380 116.720 103.110 116.890 ;
        RECT 97.860 116.650 99.850 116.660 ;
        RECT 97.860 113.050 98.640 116.650 ;
        RECT 100.260 115.600 103.110 116.720 ;
        RECT 103.500 116.420 103.850 117.170 ;
        RECT 104.600 117.050 106.470 117.210 ;
        RECT 104.600 117.000 105.360 117.050 ;
        RECT 106.240 116.980 106.470 117.050 ;
        RECT 114.880 116.980 115.110 117.210 ;
        RECT 106.675 116.700 114.675 116.930 ;
        RECT 103.500 116.360 103.790 116.420 ;
        RECT 103.410 116.240 103.790 116.360 ;
        RECT 106.770 116.300 114.630 116.700 ;
        RECT 115.440 116.520 116.400 125.780 ;
        RECT 116.840 127.980 117.620 128.010 ;
        RECT 116.840 125.880 117.670 127.980 ;
        RECT 123.340 127.590 124.590 128.030 ;
        RECT 134.440 128.010 135.380 130.150 ;
        RECT 135.910 128.010 136.610 131.640 ;
        RECT 138.250 130.590 141.100 131.710 ;
        RECT 141.490 131.410 141.840 132.160 ;
        RECT 142.590 132.040 144.460 132.200 ;
        RECT 142.590 131.990 143.350 132.040 ;
        RECT 144.230 131.970 144.460 132.040 ;
        RECT 152.870 131.970 153.100 132.200 ;
        RECT 144.665 131.690 152.665 131.920 ;
        RECT 141.490 131.350 141.780 131.410 ;
        RECT 141.400 131.230 141.780 131.350 ;
        RECT 144.760 131.290 152.620 131.690 ;
        RECT 153.430 131.290 154.390 140.770 ;
        RECT 138.190 130.360 141.190 130.590 ;
        RECT 141.400 130.400 141.740 131.230 ;
        RECT 143.750 131.220 154.390 131.290 ;
        RECT 138.240 130.330 141.100 130.360 ;
        RECT 138.240 130.310 139.410 130.330 ;
        RECT 140.370 130.320 141.100 130.330 ;
        RECT 138.190 129.920 141.190 130.150 ;
        RECT 141.395 130.110 141.740 130.400 ;
        RECT 141.930 130.180 154.390 131.220 ;
        RECT 141.930 130.160 154.380 130.180 ;
        RECT 142.200 130.150 147.640 130.160 ;
        RECT 148.640 130.150 154.380 130.160 ;
        RECT 141.400 130.000 141.740 130.110 ;
        RECT 121.280 127.580 126.520 127.590 ;
        RECT 118.330 127.480 133.630 127.580 ;
        RECT 118.330 127.470 133.665 127.480 ;
        RECT 118.290 127.350 133.665 127.470 ;
        RECT 118.290 127.240 122.290 127.350 ;
        RECT 123.340 127.270 125.080 127.350 ;
        RECT 125.660 127.270 133.665 127.350 ;
        RECT 123.340 127.190 124.590 127.270 ;
        RECT 125.665 127.250 133.665 127.270 ;
        RECT 117.900 126.940 118.130 127.190 ;
        RECT 122.450 127.050 122.680 127.190 ;
        RECT 125.230 127.050 125.460 127.200 ;
        RECT 122.450 126.940 125.460 127.050 ;
        RECT 133.870 126.940 134.100 127.200 ;
        RECT 117.900 126.500 134.100 126.940 ;
        RECT 117.900 126.230 118.130 126.500 ;
        RECT 122.450 126.470 134.100 126.500 ;
        RECT 122.450 126.380 125.460 126.470 ;
        RECT 122.450 126.230 122.680 126.380 ;
        RECT 125.230 126.240 125.460 126.380 ;
        RECT 133.870 126.240 134.100 126.470 ;
        RECT 118.290 125.950 122.290 126.180 ;
        RECT 125.665 125.970 133.665 126.190 ;
        RECT 134.430 125.970 135.390 128.010 ;
        RECT 125.665 125.960 135.390 125.970 ;
        RECT 118.290 125.880 122.280 125.950 ;
        RECT 116.840 125.770 122.280 125.880 ;
        RECT 125.720 125.800 135.390 125.960 ;
        RECT 116.840 125.680 119.970 125.770 ;
        RECT 133.460 125.750 135.390 125.800 ;
        RECT 116.840 122.410 117.670 125.680 ;
        RECT 121.320 125.220 126.570 125.230 ;
        RECT 121.320 125.110 133.630 125.220 ;
        RECT 118.350 125.050 133.630 125.110 ;
        RECT 118.350 125.040 133.665 125.050 ;
        RECT 118.290 124.910 133.665 125.040 ;
        RECT 118.290 124.900 123.450 124.910 ;
        RECT 118.290 124.810 122.290 124.900 ;
        RECT 125.665 124.820 133.665 124.910 ;
        RECT 125.750 124.810 133.640 124.820 ;
        RECT 117.900 124.450 118.130 124.760 ;
        RECT 118.350 124.450 122.250 124.810 ;
        RECT 122.450 124.450 122.680 124.760 ;
        RECT 117.900 123.110 122.680 124.450 ;
        RECT 117.900 122.800 118.130 123.110 ;
        RECT 122.450 122.800 122.680 123.110 ;
        RECT 125.230 124.230 125.460 124.770 ;
        RECT 126.270 124.230 127.280 124.260 ;
        RECT 133.870 124.230 134.100 124.770 ;
        RECT 125.230 123.330 134.100 124.230 ;
        RECT 125.230 122.810 125.460 123.330 ;
        RECT 126.270 123.260 127.280 123.330 ;
        RECT 133.870 122.810 134.100 123.330 ;
        RECT 118.290 122.520 122.290 122.750 ;
        RECT 125.665 122.530 133.665 122.760 ;
        RECT 116.840 122.370 117.970 122.410 ;
        RECT 116.840 122.290 118.210 122.370 ;
        RECT 118.580 122.300 122.240 122.520 ;
        RECT 118.580 122.290 120.020 122.300 ;
        RECT 116.840 122.250 120.020 122.290 ;
        RECT 116.840 122.160 119.530 122.250 ;
        RECT 125.730 122.240 133.620 122.530 ;
        RECT 116.840 122.100 118.860 122.160 ;
        RECT 116.840 122.050 118.610 122.100 ;
        RECT 116.840 118.710 117.670 122.050 ;
        RECT 125.720 121.750 133.640 121.760 ;
        RECT 121.950 121.740 133.640 121.750 ;
        RECT 118.330 121.620 133.640 121.740 ;
        RECT 118.330 121.610 133.665 121.620 ;
        RECT 118.290 121.490 133.665 121.610 ;
        RECT 118.290 121.380 122.290 121.490 ;
        RECT 117.900 121.040 118.130 121.330 ;
        RECT 118.350 121.040 122.240 121.380 ;
        RECT 122.450 121.040 122.680 121.330 ;
        RECT 117.900 119.670 122.680 121.040 ;
        RECT 117.900 119.370 118.130 119.670 ;
        RECT 122.450 119.370 122.680 119.670 ;
        RECT 118.290 119.090 122.290 119.320 ;
        RECT 118.540 118.860 122.110 119.090 ;
        RECT 118.540 118.710 122.230 118.860 ;
        RECT 116.840 118.430 122.230 118.710 ;
        RECT 123.480 118.540 124.100 121.490 ;
        RECT 125.665 121.390 133.665 121.490 ;
        RECT 125.720 121.380 133.640 121.390 ;
        RECT 125.230 120.680 125.460 121.340 ;
        RECT 126.240 120.680 127.240 120.770 ;
        RECT 133.870 120.680 134.100 121.340 ;
        RECT 125.230 119.860 134.100 120.680 ;
        RECT 125.230 119.380 125.460 119.860 ;
        RECT 126.240 119.770 127.240 119.860 ;
        RECT 133.870 119.380 134.100 119.860 ;
        RECT 125.665 119.100 133.665 119.330 ;
        RECT 116.840 117.970 122.240 118.430 ;
        RECT 116.840 116.630 118.840 117.970 ;
        RECT 120.590 117.960 122.240 117.970 ;
        RECT 119.280 116.690 120.280 117.410 ;
        RECT 120.590 117.150 120.900 117.960 ;
        RECT 121.360 117.680 122.240 117.960 ;
        RECT 122.480 118.140 124.100 118.540 ;
        RECT 125.750 118.190 133.620 119.100 ;
        RECT 121.300 117.450 122.300 117.680 ;
        RECT 122.480 117.490 122.830 118.140 ;
        RECT 123.480 118.130 124.100 118.140 ;
        RECT 125.665 117.960 133.665 118.190 ;
        RECT 125.750 117.950 133.620 117.960 ;
        RECT 121.360 117.240 122.240 117.260 ;
        RECT 120.630 116.860 120.900 117.150 ;
        RECT 121.300 117.010 122.300 117.240 ;
        RECT 122.460 117.200 122.830 117.490 ;
        RECT 122.490 117.140 122.830 117.200 ;
        RECT 123.590 117.810 124.350 117.860 ;
        RECT 125.230 117.810 125.460 117.910 ;
        RECT 123.590 117.600 125.460 117.810 ;
        RECT 133.870 117.600 134.100 117.910 ;
        RECT 123.590 117.180 126.130 117.600 ;
        RECT 133.500 117.180 134.100 117.600 ;
        RECT 121.360 116.860 122.240 117.010 ;
        RECT 121.370 116.690 122.100 116.860 ;
        RECT 115.420 116.300 116.400 116.520 ;
        RECT 100.200 115.370 103.200 115.600 ;
        RECT 103.410 115.410 103.750 116.240 ;
        RECT 105.760 116.230 116.400 116.300 ;
        RECT 100.250 115.340 103.110 115.370 ;
        RECT 100.250 115.320 101.420 115.340 ;
        RECT 102.380 115.330 103.110 115.340 ;
        RECT 100.200 114.930 103.200 115.160 ;
        RECT 103.405 115.120 103.750 115.410 ;
        RECT 103.940 115.190 116.400 116.230 ;
        RECT 116.860 116.620 118.840 116.630 ;
        RECT 103.940 115.170 116.360 115.190 ;
        RECT 104.210 115.160 109.650 115.170 ;
        RECT 110.650 115.160 116.360 115.170 ;
        RECT 103.410 115.010 103.750 115.120 ;
        RECT 97.850 113.020 98.640 113.050 ;
        RECT 97.850 110.920 98.680 113.020 ;
        RECT 104.350 112.630 105.600 113.070 ;
        RECT 115.420 113.050 116.360 115.160 ;
        RECT 102.290 112.620 107.530 112.630 ;
        RECT 99.340 112.520 114.640 112.620 ;
        RECT 99.340 112.510 114.675 112.520 ;
        RECT 99.300 112.390 114.675 112.510 ;
        RECT 99.300 112.280 103.300 112.390 ;
        RECT 104.350 112.310 106.090 112.390 ;
        RECT 106.670 112.310 114.675 112.390 ;
        RECT 104.350 112.230 105.600 112.310 ;
        RECT 106.675 112.290 114.675 112.310 ;
        RECT 98.910 111.980 99.140 112.230 ;
        RECT 103.460 112.090 103.690 112.230 ;
        RECT 106.240 112.090 106.470 112.240 ;
        RECT 103.460 111.980 106.470 112.090 ;
        RECT 114.880 111.980 115.110 112.240 ;
        RECT 98.910 111.540 115.110 111.980 ;
        RECT 115.420 111.540 116.400 113.050 ;
        RECT 116.860 113.030 117.620 116.620 ;
        RECT 119.250 115.570 122.100 116.690 ;
        RECT 122.490 116.390 122.840 117.140 ;
        RECT 123.590 117.020 125.460 117.180 ;
        RECT 123.590 116.970 124.350 117.020 ;
        RECT 125.230 116.950 125.460 117.020 ;
        RECT 133.870 116.950 134.100 117.180 ;
        RECT 125.665 116.670 133.665 116.900 ;
        RECT 122.490 116.330 122.780 116.390 ;
        RECT 122.400 116.210 122.780 116.330 ;
        RECT 125.760 116.270 133.620 116.670 ;
        RECT 134.430 116.270 135.390 125.750 ;
        RECT 135.840 127.980 136.610 128.010 ;
        RECT 135.840 125.880 136.670 127.980 ;
        RECT 142.340 127.590 143.590 128.030 ;
        RECT 153.440 128.010 154.380 130.150 ;
        RECT 140.280 127.580 145.520 127.590 ;
        RECT 137.330 127.480 152.630 127.580 ;
        RECT 137.330 127.470 152.665 127.480 ;
        RECT 137.290 127.350 152.665 127.470 ;
        RECT 137.290 127.240 141.290 127.350 ;
        RECT 142.340 127.270 144.080 127.350 ;
        RECT 144.660 127.270 152.665 127.350 ;
        RECT 142.340 127.190 143.590 127.270 ;
        RECT 144.665 127.250 152.665 127.270 ;
        RECT 136.900 126.940 137.130 127.190 ;
        RECT 141.450 127.050 141.680 127.190 ;
        RECT 144.230 127.050 144.460 127.200 ;
        RECT 141.450 126.940 144.460 127.050 ;
        RECT 152.870 126.940 153.100 127.200 ;
        RECT 136.900 126.500 153.100 126.940 ;
        RECT 136.900 126.230 137.130 126.500 ;
        RECT 141.450 126.470 153.100 126.500 ;
        RECT 141.450 126.380 144.460 126.470 ;
        RECT 141.450 126.230 141.680 126.380 ;
        RECT 144.230 126.240 144.460 126.380 ;
        RECT 152.870 126.240 153.100 126.470 ;
        RECT 137.290 125.950 141.290 126.180 ;
        RECT 144.665 125.970 152.665 126.190 ;
        RECT 153.430 125.970 154.390 128.010 ;
        RECT 144.665 125.960 154.390 125.970 ;
        RECT 137.290 125.880 141.280 125.950 ;
        RECT 135.840 125.770 141.280 125.880 ;
        RECT 144.720 125.800 154.390 125.960 ;
        RECT 135.840 125.680 138.970 125.770 ;
        RECT 152.460 125.750 154.390 125.800 ;
        RECT 135.840 122.410 136.670 125.680 ;
        RECT 140.320 125.220 145.570 125.230 ;
        RECT 140.320 125.110 152.630 125.220 ;
        RECT 137.350 125.050 152.630 125.110 ;
        RECT 137.350 125.040 152.665 125.050 ;
        RECT 137.290 124.910 152.665 125.040 ;
        RECT 137.290 124.900 142.450 124.910 ;
        RECT 137.290 124.810 141.290 124.900 ;
        RECT 144.665 124.820 152.665 124.910 ;
        RECT 144.750 124.810 152.640 124.820 ;
        RECT 136.900 124.450 137.130 124.760 ;
        RECT 137.350 124.450 141.250 124.810 ;
        RECT 141.450 124.450 141.680 124.760 ;
        RECT 136.900 123.110 141.680 124.450 ;
        RECT 136.900 122.800 137.130 123.110 ;
        RECT 141.450 122.800 141.680 123.110 ;
        RECT 144.230 124.230 144.460 124.770 ;
        RECT 145.270 124.230 146.280 124.260 ;
        RECT 152.870 124.230 153.100 124.770 ;
        RECT 144.230 123.330 153.100 124.230 ;
        RECT 144.230 122.810 144.460 123.330 ;
        RECT 145.270 123.260 146.280 123.330 ;
        RECT 152.870 122.810 153.100 123.330 ;
        RECT 137.290 122.520 141.290 122.750 ;
        RECT 144.665 122.530 152.665 122.760 ;
        RECT 135.840 122.370 136.970 122.410 ;
        RECT 135.840 122.290 137.210 122.370 ;
        RECT 137.580 122.300 141.240 122.520 ;
        RECT 137.580 122.290 139.020 122.300 ;
        RECT 135.840 122.250 139.020 122.290 ;
        RECT 135.840 122.160 138.530 122.250 ;
        RECT 144.730 122.240 152.620 122.530 ;
        RECT 135.840 122.100 137.860 122.160 ;
        RECT 135.840 122.050 137.610 122.100 ;
        RECT 135.840 118.710 136.670 122.050 ;
        RECT 144.720 121.750 152.640 121.760 ;
        RECT 140.950 121.740 152.640 121.750 ;
        RECT 137.330 121.620 152.640 121.740 ;
        RECT 137.330 121.610 152.665 121.620 ;
        RECT 137.290 121.490 152.665 121.610 ;
        RECT 137.290 121.380 141.290 121.490 ;
        RECT 136.900 121.040 137.130 121.330 ;
        RECT 137.350 121.040 141.240 121.380 ;
        RECT 141.450 121.040 141.680 121.330 ;
        RECT 136.900 119.670 141.680 121.040 ;
        RECT 136.900 119.370 137.130 119.670 ;
        RECT 141.450 119.370 141.680 119.670 ;
        RECT 137.290 119.090 141.290 119.320 ;
        RECT 137.540 118.860 141.110 119.090 ;
        RECT 137.540 118.710 141.230 118.860 ;
        RECT 135.840 118.430 141.230 118.710 ;
        RECT 142.480 118.540 143.100 121.490 ;
        RECT 144.665 121.390 152.665 121.490 ;
        RECT 144.720 121.380 152.640 121.390 ;
        RECT 144.230 120.680 144.460 121.340 ;
        RECT 145.240 120.680 146.240 120.770 ;
        RECT 152.870 120.680 153.100 121.340 ;
        RECT 144.230 119.860 153.100 120.680 ;
        RECT 144.230 119.380 144.460 119.860 ;
        RECT 145.240 119.770 146.240 119.860 ;
        RECT 152.870 119.380 153.100 119.860 ;
        RECT 144.665 119.100 152.665 119.330 ;
        RECT 135.840 117.970 141.240 118.430 ;
        RECT 135.840 116.630 137.840 117.970 ;
        RECT 139.590 117.960 141.240 117.970 ;
        RECT 138.280 116.690 139.280 117.410 ;
        RECT 139.590 117.150 139.900 117.960 ;
        RECT 140.360 117.680 141.240 117.960 ;
        RECT 141.480 118.140 143.100 118.540 ;
        RECT 144.750 118.190 152.620 119.100 ;
        RECT 140.300 117.450 141.300 117.680 ;
        RECT 141.480 117.490 141.830 118.140 ;
        RECT 142.480 118.130 143.100 118.140 ;
        RECT 144.665 117.960 152.665 118.190 ;
        RECT 144.750 117.950 152.620 117.960 ;
        RECT 140.360 117.240 141.240 117.260 ;
        RECT 139.630 116.860 139.900 117.150 ;
        RECT 140.300 117.010 141.300 117.240 ;
        RECT 141.460 117.200 141.830 117.490 ;
        RECT 141.490 117.140 141.830 117.200 ;
        RECT 142.590 117.810 143.350 117.860 ;
        RECT 144.230 117.810 144.460 117.910 ;
        RECT 142.590 117.600 144.460 117.810 ;
        RECT 152.870 117.600 153.100 117.910 ;
        RECT 142.590 117.180 145.130 117.600 ;
        RECT 152.500 117.180 153.100 117.600 ;
        RECT 140.360 116.860 141.240 117.010 ;
        RECT 140.370 116.690 141.100 116.860 ;
        RECT 119.190 115.340 122.190 115.570 ;
        RECT 122.400 115.380 122.740 116.210 ;
        RECT 124.750 116.200 135.390 116.270 ;
        RECT 119.240 115.310 122.100 115.340 ;
        RECT 119.240 115.290 120.410 115.310 ;
        RECT 121.370 115.300 122.100 115.310 ;
        RECT 119.190 114.900 122.190 115.130 ;
        RECT 122.395 115.090 122.740 115.380 ;
        RECT 122.930 115.160 135.390 116.200 ;
        RECT 135.910 116.620 137.840 116.630 ;
        RECT 122.930 115.140 135.330 115.160 ;
        RECT 123.200 115.130 128.640 115.140 ;
        RECT 129.640 115.130 135.330 115.140 ;
        RECT 122.400 114.980 122.740 115.090 ;
        RECT 98.910 111.270 99.140 111.540 ;
        RECT 103.460 111.510 115.110 111.540 ;
        RECT 103.460 111.420 106.470 111.510 ;
        RECT 103.460 111.270 103.690 111.420 ;
        RECT 106.240 111.280 106.470 111.420 ;
        RECT 114.880 111.280 115.110 111.510 ;
        RECT 99.300 110.990 103.300 111.220 ;
        RECT 106.675 111.010 114.675 111.230 ;
        RECT 115.440 111.010 116.400 111.540 ;
        RECT 106.675 111.000 116.400 111.010 ;
        RECT 99.300 110.920 103.290 110.990 ;
        RECT 97.850 110.810 103.290 110.920 ;
        RECT 106.730 110.840 116.400 111.000 ;
        RECT 97.850 110.720 100.980 110.810 ;
        RECT 114.470 110.790 116.400 110.840 ;
        RECT 97.850 107.450 98.680 110.720 ;
        RECT 102.330 110.260 107.580 110.270 ;
        RECT 102.330 110.150 114.640 110.260 ;
        RECT 99.360 110.090 114.640 110.150 ;
        RECT 99.360 110.080 114.675 110.090 ;
        RECT 99.300 109.950 114.675 110.080 ;
        RECT 99.300 109.940 104.460 109.950 ;
        RECT 99.300 109.850 103.300 109.940 ;
        RECT 106.675 109.860 114.675 109.950 ;
        RECT 106.760 109.850 114.650 109.860 ;
        RECT 98.910 109.490 99.140 109.800 ;
        RECT 99.360 109.490 103.260 109.850 ;
        RECT 103.460 109.490 103.690 109.800 ;
        RECT 98.910 108.150 103.690 109.490 ;
        RECT 98.910 107.840 99.140 108.150 ;
        RECT 103.460 107.840 103.690 108.150 ;
        RECT 106.240 109.270 106.470 109.810 ;
        RECT 107.280 109.270 108.290 109.300 ;
        RECT 114.880 109.270 115.110 109.810 ;
        RECT 106.240 108.370 115.110 109.270 ;
        RECT 106.240 107.850 106.470 108.370 ;
        RECT 107.280 108.300 108.290 108.370 ;
        RECT 114.880 107.850 115.110 108.370 ;
        RECT 99.300 107.560 103.300 107.790 ;
        RECT 106.675 107.570 114.675 107.800 ;
        RECT 97.850 107.410 98.980 107.450 ;
        RECT 97.850 107.330 99.220 107.410 ;
        RECT 99.590 107.340 103.250 107.560 ;
        RECT 99.590 107.330 101.030 107.340 ;
        RECT 97.850 107.290 101.030 107.330 ;
        RECT 97.850 107.200 100.540 107.290 ;
        RECT 106.740 107.280 114.630 107.570 ;
        RECT 97.850 107.140 99.870 107.200 ;
        RECT 97.850 107.090 99.620 107.140 ;
        RECT 97.850 103.750 98.680 107.090 ;
        RECT 106.730 106.790 114.650 106.800 ;
        RECT 102.960 106.780 114.650 106.790 ;
        RECT 99.340 106.660 114.650 106.780 ;
        RECT 99.340 106.650 114.675 106.660 ;
        RECT 99.300 106.530 114.675 106.650 ;
        RECT 99.300 106.420 103.300 106.530 ;
        RECT 98.910 106.080 99.140 106.370 ;
        RECT 99.360 106.080 103.250 106.420 ;
        RECT 103.460 106.080 103.690 106.370 ;
        RECT 98.910 104.710 103.690 106.080 ;
        RECT 98.910 104.410 99.140 104.710 ;
        RECT 103.460 104.410 103.690 104.710 ;
        RECT 99.300 104.130 103.300 104.360 ;
        RECT 99.550 103.900 103.120 104.130 ;
        RECT 99.550 103.750 103.240 103.900 ;
        RECT 97.850 103.470 103.240 103.750 ;
        RECT 104.490 103.580 105.110 106.530 ;
        RECT 106.675 106.430 114.675 106.530 ;
        RECT 106.730 106.420 114.650 106.430 ;
        RECT 106.240 105.720 106.470 106.380 ;
        RECT 107.250 105.720 108.250 105.810 ;
        RECT 114.880 105.720 115.110 106.380 ;
        RECT 106.240 104.900 115.110 105.720 ;
        RECT 106.240 104.420 106.470 104.900 ;
        RECT 107.250 104.810 108.250 104.900 ;
        RECT 114.880 104.420 115.110 104.900 ;
        RECT 106.675 104.140 114.675 104.370 ;
        RECT 97.850 103.010 103.250 103.470 ;
        RECT 97.850 101.670 99.850 103.010 ;
        RECT 101.600 103.000 103.250 103.010 ;
        RECT 100.290 102.330 101.290 102.450 ;
        RECT 97.870 101.660 99.850 101.670 ;
        RECT 100.260 101.730 101.290 102.330 ;
        RECT 101.600 102.190 101.910 103.000 ;
        RECT 102.370 102.720 103.250 103.000 ;
        RECT 103.490 103.180 105.110 103.580 ;
        RECT 106.760 103.230 114.630 104.140 ;
        RECT 102.310 102.490 103.310 102.720 ;
        RECT 103.490 102.530 103.840 103.180 ;
        RECT 104.490 103.170 105.110 103.180 ;
        RECT 106.675 103.000 114.675 103.230 ;
        RECT 106.760 102.990 114.630 103.000 ;
        RECT 102.370 102.280 103.250 102.300 ;
        RECT 101.640 101.900 101.910 102.190 ;
        RECT 102.310 102.050 103.310 102.280 ;
        RECT 103.470 102.240 103.840 102.530 ;
        RECT 103.500 102.180 103.840 102.240 ;
        RECT 104.600 102.850 105.360 102.900 ;
        RECT 106.240 102.850 106.470 102.950 ;
        RECT 104.600 102.640 106.470 102.850 ;
        RECT 114.880 102.640 115.110 102.950 ;
        RECT 104.600 102.220 107.140 102.640 ;
        RECT 114.510 102.220 115.110 102.640 ;
        RECT 102.370 101.900 103.250 102.050 ;
        RECT 102.380 101.730 103.110 101.900 ;
        RECT 97.870 98.540 98.920 101.660 ;
        RECT 100.260 100.610 103.110 101.730 ;
        RECT 103.500 101.430 103.850 102.180 ;
        RECT 104.600 102.060 106.470 102.220 ;
        RECT 104.600 102.010 105.360 102.060 ;
        RECT 106.240 101.990 106.470 102.060 ;
        RECT 114.880 101.990 115.110 102.220 ;
        RECT 106.675 101.710 114.675 101.940 ;
        RECT 103.500 101.370 103.790 101.430 ;
        RECT 103.410 101.250 103.790 101.370 ;
        RECT 106.770 101.310 114.630 101.710 ;
        RECT 115.440 101.310 116.400 110.790 ;
        RECT 116.840 113.000 117.620 113.030 ;
        RECT 116.840 110.900 117.670 113.000 ;
        RECT 123.340 112.610 124.590 113.050 ;
        RECT 134.390 113.030 135.330 115.130 ;
        RECT 135.910 113.030 136.610 116.620 ;
        RECT 138.250 115.570 141.100 116.690 ;
        RECT 141.490 116.390 141.840 117.140 ;
        RECT 142.590 117.020 144.460 117.180 ;
        RECT 142.590 116.970 143.350 117.020 ;
        RECT 144.230 116.950 144.460 117.020 ;
        RECT 152.870 116.950 153.100 117.180 ;
        RECT 144.665 116.670 152.665 116.900 ;
        RECT 141.490 116.330 141.780 116.390 ;
        RECT 141.400 116.210 141.780 116.330 ;
        RECT 144.760 116.270 152.620 116.670 ;
        RECT 153.430 116.270 154.390 125.750 ;
        RECT 138.190 115.340 141.190 115.570 ;
        RECT 141.400 115.380 141.740 116.210 ;
        RECT 143.750 116.200 154.390 116.270 ;
        RECT 138.240 115.310 141.100 115.340 ;
        RECT 138.240 115.290 139.410 115.310 ;
        RECT 140.370 115.300 141.100 115.310 ;
        RECT 138.190 114.900 141.190 115.130 ;
        RECT 141.395 115.090 141.740 115.380 ;
        RECT 141.930 116.180 154.390 116.200 ;
        RECT 141.930 115.140 154.420 116.180 ;
        RECT 142.200 115.130 147.640 115.140 ;
        RECT 148.640 115.130 154.420 115.140 ;
        RECT 141.400 114.980 141.740 115.090 ;
        RECT 121.280 112.600 126.520 112.610 ;
        RECT 118.330 112.500 133.630 112.600 ;
        RECT 118.330 112.490 133.665 112.500 ;
        RECT 118.290 112.370 133.665 112.490 ;
        RECT 118.290 112.260 122.290 112.370 ;
        RECT 123.340 112.290 125.080 112.370 ;
        RECT 125.660 112.290 133.665 112.370 ;
        RECT 123.340 112.210 124.590 112.290 ;
        RECT 125.665 112.270 133.665 112.290 ;
        RECT 117.900 111.960 118.130 112.210 ;
        RECT 122.450 112.070 122.680 112.210 ;
        RECT 125.230 112.070 125.460 112.220 ;
        RECT 122.450 111.960 125.460 112.070 ;
        RECT 133.870 111.960 134.100 112.220 ;
        RECT 117.900 111.520 134.100 111.960 ;
        RECT 117.900 111.250 118.130 111.520 ;
        RECT 122.450 111.490 134.100 111.520 ;
        RECT 122.450 111.400 125.460 111.490 ;
        RECT 122.450 111.250 122.680 111.400 ;
        RECT 125.230 111.260 125.460 111.400 ;
        RECT 133.870 111.260 134.100 111.490 ;
        RECT 134.390 111.240 135.390 113.030 ;
        RECT 118.290 110.970 122.290 111.200 ;
        RECT 125.665 110.990 133.665 111.210 ;
        RECT 134.430 110.990 135.390 111.240 ;
        RECT 125.665 110.980 135.390 110.990 ;
        RECT 118.290 110.900 122.280 110.970 ;
        RECT 116.840 110.790 122.280 110.900 ;
        RECT 125.720 110.820 135.390 110.980 ;
        RECT 116.840 110.700 119.970 110.790 ;
        RECT 133.460 110.770 135.390 110.820 ;
        RECT 116.840 107.430 117.670 110.700 ;
        RECT 121.320 110.240 126.570 110.250 ;
        RECT 121.320 110.130 133.630 110.240 ;
        RECT 118.350 110.070 133.630 110.130 ;
        RECT 118.350 110.060 133.665 110.070 ;
        RECT 118.290 109.930 133.665 110.060 ;
        RECT 118.290 109.920 123.450 109.930 ;
        RECT 118.290 109.830 122.290 109.920 ;
        RECT 125.665 109.840 133.665 109.930 ;
        RECT 125.750 109.830 133.640 109.840 ;
        RECT 117.900 109.470 118.130 109.780 ;
        RECT 118.350 109.470 122.250 109.830 ;
        RECT 122.450 109.470 122.680 109.780 ;
        RECT 117.900 108.130 122.680 109.470 ;
        RECT 117.900 107.820 118.130 108.130 ;
        RECT 122.450 107.820 122.680 108.130 ;
        RECT 125.230 109.250 125.460 109.790 ;
        RECT 126.270 109.250 127.280 109.280 ;
        RECT 133.870 109.250 134.100 109.790 ;
        RECT 125.230 108.350 134.100 109.250 ;
        RECT 125.230 107.830 125.460 108.350 ;
        RECT 126.270 108.280 127.280 108.350 ;
        RECT 133.870 107.830 134.100 108.350 ;
        RECT 118.290 107.540 122.290 107.770 ;
        RECT 125.665 107.550 133.665 107.780 ;
        RECT 116.840 107.390 117.970 107.430 ;
        RECT 116.840 107.310 118.210 107.390 ;
        RECT 118.580 107.320 122.240 107.540 ;
        RECT 118.580 107.310 120.020 107.320 ;
        RECT 116.840 107.270 120.020 107.310 ;
        RECT 116.840 107.180 119.530 107.270 ;
        RECT 125.730 107.260 133.620 107.550 ;
        RECT 116.840 107.120 118.860 107.180 ;
        RECT 116.840 107.070 118.610 107.120 ;
        RECT 116.840 103.730 117.670 107.070 ;
        RECT 125.720 106.770 133.640 106.780 ;
        RECT 121.950 106.760 133.640 106.770 ;
        RECT 118.330 106.640 133.640 106.760 ;
        RECT 118.330 106.630 133.665 106.640 ;
        RECT 118.290 106.510 133.665 106.630 ;
        RECT 118.290 106.400 122.290 106.510 ;
        RECT 117.900 106.060 118.130 106.350 ;
        RECT 118.350 106.060 122.240 106.400 ;
        RECT 122.450 106.060 122.680 106.350 ;
        RECT 117.900 104.690 122.680 106.060 ;
        RECT 117.900 104.390 118.130 104.690 ;
        RECT 122.450 104.390 122.680 104.690 ;
        RECT 118.290 104.110 122.290 104.340 ;
        RECT 118.540 103.880 122.110 104.110 ;
        RECT 118.540 103.730 122.230 103.880 ;
        RECT 116.840 103.450 122.230 103.730 ;
        RECT 123.480 103.560 124.100 106.510 ;
        RECT 125.665 106.410 133.665 106.510 ;
        RECT 125.720 106.400 133.640 106.410 ;
        RECT 125.230 105.700 125.460 106.360 ;
        RECT 126.240 105.700 127.240 105.790 ;
        RECT 133.870 105.700 134.100 106.360 ;
        RECT 125.230 104.880 134.100 105.700 ;
        RECT 125.230 104.400 125.460 104.880 ;
        RECT 126.240 104.790 127.240 104.880 ;
        RECT 133.870 104.400 134.100 104.880 ;
        RECT 125.665 104.120 133.665 104.350 ;
        RECT 116.840 102.990 122.240 103.450 ;
        RECT 116.840 101.650 118.840 102.990 ;
        RECT 120.590 102.980 122.240 102.990 ;
        RECT 119.280 101.710 120.280 102.430 ;
        RECT 120.590 102.170 120.900 102.980 ;
        RECT 121.360 102.700 122.240 102.980 ;
        RECT 122.480 103.160 124.100 103.560 ;
        RECT 125.750 103.210 133.620 104.120 ;
        RECT 121.300 102.470 122.300 102.700 ;
        RECT 122.480 102.510 122.830 103.160 ;
        RECT 123.480 103.150 124.100 103.160 ;
        RECT 125.665 102.980 133.665 103.210 ;
        RECT 125.750 102.970 133.620 102.980 ;
        RECT 121.360 102.260 122.240 102.280 ;
        RECT 120.630 101.880 120.900 102.170 ;
        RECT 121.300 102.030 122.300 102.260 ;
        RECT 122.460 102.220 122.830 102.510 ;
        RECT 122.490 102.160 122.830 102.220 ;
        RECT 123.590 102.830 124.350 102.880 ;
        RECT 125.230 102.830 125.460 102.930 ;
        RECT 123.590 102.620 125.460 102.830 ;
        RECT 133.870 102.620 134.100 102.930 ;
        RECT 123.590 102.200 126.130 102.620 ;
        RECT 133.500 102.200 134.100 102.620 ;
        RECT 121.360 101.880 122.240 102.030 ;
        RECT 121.370 101.710 122.100 101.880 ;
        RECT 116.920 101.640 118.840 101.650 ;
        RECT 100.200 100.380 103.200 100.610 ;
        RECT 103.410 100.420 103.750 101.250 ;
        RECT 105.760 101.240 116.400 101.310 ;
        RECT 100.250 100.350 103.110 100.380 ;
        RECT 100.250 100.330 101.420 100.350 ;
        RECT 102.380 100.340 103.110 100.350 ;
        RECT 100.200 99.940 103.200 100.170 ;
        RECT 103.405 100.130 103.750 100.420 ;
        RECT 103.940 100.200 116.400 101.240 ;
        RECT 119.250 100.590 122.100 101.710 ;
        RECT 122.490 101.410 122.840 102.160 ;
        RECT 123.590 102.040 125.460 102.200 ;
        RECT 123.590 101.990 124.350 102.040 ;
        RECT 125.230 101.970 125.460 102.040 ;
        RECT 133.870 101.970 134.100 102.200 ;
        RECT 125.665 101.690 133.665 101.920 ;
        RECT 122.490 101.350 122.780 101.410 ;
        RECT 122.400 101.230 122.780 101.350 ;
        RECT 125.760 101.290 133.620 101.690 ;
        RECT 134.430 101.290 135.390 110.770 ;
        RECT 135.890 113.000 136.610 113.030 ;
        RECT 135.890 110.900 136.720 113.000 ;
        RECT 142.390 112.610 143.640 113.050 ;
        RECT 153.480 113.030 154.420 115.130 ;
        RECT 140.330 112.600 145.570 112.610 ;
        RECT 137.380 112.500 152.680 112.600 ;
        RECT 137.380 112.490 152.715 112.500 ;
        RECT 137.340 112.370 152.715 112.490 ;
        RECT 137.340 112.260 141.340 112.370 ;
        RECT 142.390 112.290 144.130 112.370 ;
        RECT 144.710 112.290 152.715 112.370 ;
        RECT 142.390 112.210 143.640 112.290 ;
        RECT 144.715 112.270 152.715 112.290 ;
        RECT 136.950 111.960 137.180 112.210 ;
        RECT 141.500 112.070 141.730 112.210 ;
        RECT 144.280 112.070 144.510 112.220 ;
        RECT 141.500 111.960 144.510 112.070 ;
        RECT 152.920 111.960 153.150 112.220 ;
        RECT 136.950 111.520 153.150 111.960 ;
        RECT 136.950 111.250 137.180 111.520 ;
        RECT 141.500 111.490 153.150 111.520 ;
        RECT 141.500 111.400 144.510 111.490 ;
        RECT 141.500 111.250 141.730 111.400 ;
        RECT 144.280 111.260 144.510 111.400 ;
        RECT 152.920 111.260 153.150 111.490 ;
        RECT 137.340 110.970 141.340 111.200 ;
        RECT 144.715 110.990 152.715 111.210 ;
        RECT 153.480 110.990 154.440 113.030 ;
        RECT 144.715 110.980 154.440 110.990 ;
        RECT 137.340 110.900 141.330 110.970 ;
        RECT 135.890 110.790 141.330 110.900 ;
        RECT 144.770 110.820 154.440 110.980 ;
        RECT 135.890 110.700 139.020 110.790 ;
        RECT 152.510 110.770 154.440 110.820 ;
        RECT 135.890 107.430 136.720 110.700 ;
        RECT 140.370 110.240 145.620 110.250 ;
        RECT 140.370 110.130 152.680 110.240 ;
        RECT 137.400 110.070 152.680 110.130 ;
        RECT 137.400 110.060 152.715 110.070 ;
        RECT 137.340 109.930 152.715 110.060 ;
        RECT 137.340 109.920 142.500 109.930 ;
        RECT 137.340 109.830 141.340 109.920 ;
        RECT 144.715 109.840 152.715 109.930 ;
        RECT 144.800 109.830 152.690 109.840 ;
        RECT 136.950 109.470 137.180 109.780 ;
        RECT 137.400 109.470 141.300 109.830 ;
        RECT 141.500 109.470 141.730 109.780 ;
        RECT 136.950 108.130 141.730 109.470 ;
        RECT 136.950 107.820 137.180 108.130 ;
        RECT 141.500 107.820 141.730 108.130 ;
        RECT 144.280 109.250 144.510 109.790 ;
        RECT 145.320 109.250 146.330 109.280 ;
        RECT 152.920 109.250 153.150 109.790 ;
        RECT 144.280 108.350 153.150 109.250 ;
        RECT 144.280 107.830 144.510 108.350 ;
        RECT 145.320 108.280 146.330 108.350 ;
        RECT 152.920 107.830 153.150 108.350 ;
        RECT 137.340 107.540 141.340 107.770 ;
        RECT 144.715 107.550 152.715 107.780 ;
        RECT 135.890 107.390 137.020 107.430 ;
        RECT 135.890 107.310 137.260 107.390 ;
        RECT 137.630 107.320 141.290 107.540 ;
        RECT 137.630 107.310 139.070 107.320 ;
        RECT 135.890 107.270 139.070 107.310 ;
        RECT 135.890 107.180 138.580 107.270 ;
        RECT 144.780 107.260 152.670 107.550 ;
        RECT 135.890 107.120 137.910 107.180 ;
        RECT 135.890 107.070 137.660 107.120 ;
        RECT 135.890 103.730 136.720 107.070 ;
        RECT 144.770 106.770 152.690 106.780 ;
        RECT 141.000 106.760 152.690 106.770 ;
        RECT 137.380 106.640 152.690 106.760 ;
        RECT 137.380 106.630 152.715 106.640 ;
        RECT 137.340 106.510 152.715 106.630 ;
        RECT 137.340 106.400 141.340 106.510 ;
        RECT 136.950 106.060 137.180 106.350 ;
        RECT 137.400 106.060 141.290 106.400 ;
        RECT 141.500 106.060 141.730 106.350 ;
        RECT 136.950 104.690 141.730 106.060 ;
        RECT 136.950 104.390 137.180 104.690 ;
        RECT 141.500 104.390 141.730 104.690 ;
        RECT 137.340 104.110 141.340 104.340 ;
        RECT 137.590 103.880 141.160 104.110 ;
        RECT 137.590 103.730 141.280 103.880 ;
        RECT 135.890 103.450 141.280 103.730 ;
        RECT 142.530 103.560 143.150 106.510 ;
        RECT 144.715 106.410 152.715 106.510 ;
        RECT 144.770 106.400 152.690 106.410 ;
        RECT 144.280 105.700 144.510 106.360 ;
        RECT 145.290 105.700 146.290 105.790 ;
        RECT 152.920 105.700 153.150 106.360 ;
        RECT 144.280 104.880 153.150 105.700 ;
        RECT 144.280 104.400 144.510 104.880 ;
        RECT 145.290 104.790 146.290 104.880 ;
        RECT 152.920 104.400 153.150 104.880 ;
        RECT 144.715 104.120 152.715 104.350 ;
        RECT 135.890 102.990 141.290 103.450 ;
        RECT 135.890 101.650 137.890 102.990 ;
        RECT 139.640 102.980 141.290 102.990 ;
        RECT 138.330 101.710 139.330 102.430 ;
        RECT 139.640 102.170 139.950 102.980 ;
        RECT 140.410 102.700 141.290 102.980 ;
        RECT 141.530 103.160 143.150 103.560 ;
        RECT 144.800 103.210 152.670 104.120 ;
        RECT 140.350 102.470 141.350 102.700 ;
        RECT 141.530 102.510 141.880 103.160 ;
        RECT 142.530 103.150 143.150 103.160 ;
        RECT 144.715 102.980 152.715 103.210 ;
        RECT 144.800 102.970 152.670 102.980 ;
        RECT 140.410 102.260 141.290 102.280 ;
        RECT 139.680 101.880 139.950 102.170 ;
        RECT 140.350 102.030 141.350 102.260 ;
        RECT 141.510 102.220 141.880 102.510 ;
        RECT 141.540 102.160 141.880 102.220 ;
        RECT 142.640 102.830 143.400 102.880 ;
        RECT 144.280 102.830 144.510 102.930 ;
        RECT 142.640 102.620 144.510 102.830 ;
        RECT 152.920 102.620 153.150 102.930 ;
        RECT 142.640 102.200 145.180 102.620 ;
        RECT 152.550 102.200 153.150 102.620 ;
        RECT 140.410 101.880 141.290 102.030 ;
        RECT 140.420 101.710 141.150 101.880 ;
        RECT 135.970 101.640 137.890 101.650 ;
        RECT 119.190 100.360 122.190 100.590 ;
        RECT 122.400 100.400 122.740 101.230 ;
        RECT 124.750 101.220 135.390 101.290 ;
        RECT 119.240 100.330 122.100 100.360 ;
        RECT 119.240 100.310 120.410 100.330 ;
        RECT 121.370 100.320 122.100 100.330 ;
        RECT 103.940 100.180 116.270 100.200 ;
        RECT 104.210 100.170 109.650 100.180 ;
        RECT 110.650 100.170 116.270 100.180 ;
        RECT 103.410 100.020 103.750 100.130 ;
        RECT 119.190 99.920 122.190 100.150 ;
        RECT 122.395 100.110 122.740 100.400 ;
        RECT 122.930 100.180 135.390 101.220 ;
        RECT 138.300 100.590 141.150 101.710 ;
        RECT 141.540 101.410 141.890 102.160 ;
        RECT 142.640 102.040 144.510 102.200 ;
        RECT 142.640 101.990 143.400 102.040 ;
        RECT 144.280 101.970 144.510 102.040 ;
        RECT 152.920 101.970 153.150 102.200 ;
        RECT 144.715 101.690 152.715 101.920 ;
        RECT 141.540 101.350 141.830 101.410 ;
        RECT 141.450 101.230 141.830 101.350 ;
        RECT 144.810 101.290 152.670 101.690 ;
        RECT 153.480 101.290 154.440 110.770 ;
        RECT 138.240 100.360 141.240 100.590 ;
        RECT 141.450 100.400 141.790 101.230 ;
        RECT 143.800 101.220 154.440 101.290 ;
        RECT 138.290 100.330 141.150 100.360 ;
        RECT 138.290 100.310 139.460 100.330 ;
        RECT 140.420 100.320 141.150 100.330 ;
        RECT 122.930 100.160 135.260 100.180 ;
        RECT 123.200 100.150 128.640 100.160 ;
        RECT 129.640 100.150 135.260 100.160 ;
        RECT 122.400 100.000 122.740 100.110 ;
        RECT 138.240 99.920 141.240 100.150 ;
        RECT 141.445 100.110 141.790 100.400 ;
        RECT 141.980 100.180 154.440 101.220 ;
        RECT 141.980 100.160 154.400 100.180 ;
        RECT 142.250 100.150 147.690 100.160 ;
        RECT 148.690 100.150 154.400 100.160 ;
        RECT 141.450 100.000 141.790 100.110 ;
        RECT 97.870 96.610 100.320 98.540 ;
        RECT 102.200 97.840 102.900 97.860 ;
        RECT 100.500 97.810 102.900 97.840 ;
        RECT 100.500 97.560 102.935 97.810 ;
        RECT 100.500 97.540 102.900 97.560 ;
        RECT 103.520 97.550 105.890 97.850 ;
        RECT 106.550 97.810 108.920 97.850 ;
        RECT 111.000 97.820 111.700 97.860 ;
        RECT 114.160 97.820 114.860 97.830 ;
        RECT 109.530 97.810 111.900 97.820 ;
        RECT 106.550 97.560 108.925 97.810 ;
        RECT 109.515 97.560 111.900 97.810 ;
        RECT 106.550 97.550 108.920 97.560 ;
        RECT 102.200 97.170 102.900 97.540 ;
        RECT 104.780 97.210 105.480 97.550 ;
        RECT 108.180 97.210 108.880 97.550 ;
        RECT 109.530 97.520 111.900 97.560 ;
        RECT 112.460 97.810 114.860 97.820 ;
        RECT 112.460 97.560 114.915 97.810 ;
        RECT 112.460 97.520 114.860 97.560 ;
        RECT 115.480 97.530 117.850 97.830 ;
        RECT 118.480 97.810 120.850 97.840 ;
        RECT 121.540 97.810 123.910 97.870 ;
        RECT 126.110 97.810 126.810 97.830 ;
        RECT 127.490 97.810 129.860 97.850 ;
        RECT 118.480 97.560 120.905 97.810 ;
        RECT 121.495 97.570 123.910 97.810 ;
        RECT 121.495 97.560 123.600 97.570 ;
        RECT 124.460 97.560 126.895 97.810 ;
        RECT 127.485 97.560 129.860 97.810 ;
        RECT 130.780 97.790 132.885 97.810 ;
        RECT 118.480 97.540 120.850 97.560 ;
        RECT 102.200 97.040 103.890 97.170 ;
        RECT 104.780 97.050 107.070 97.210 ;
        RECT 102.200 96.900 104.230 97.040 ;
        RECT 102.640 96.860 104.230 96.900 ;
        RECT 104.780 96.870 107.490 97.050 ;
        RECT 108.180 97.020 110.100 97.210 ;
        RECT 111.000 97.110 111.700 97.520 ;
        RECT 114.160 97.180 114.860 97.520 ;
        RECT 108.180 96.890 110.210 97.020 ;
        RECT 111.000 96.980 112.950 97.110 ;
        RECT 114.160 97.000 116.110 97.180 ;
        RECT 117.020 97.130 117.720 97.530 ;
        RECT 120.020 97.190 120.720 97.540 ;
        RECT 111.000 96.900 113.320 96.980 ;
        RECT 97.870 96.340 101.310 96.610 ;
        RECT 103.530 96.370 104.230 96.860 ;
        RECT 105.250 96.800 107.490 96.870 ;
        RECT 97.870 96.330 102.910 96.340 ;
        RECT 97.870 96.080 102.935 96.330 ;
        RECT 97.870 96.040 102.910 96.080 ;
        RECT 103.520 96.070 105.890 96.370 ;
        RECT 106.790 96.330 107.490 96.800 ;
        RECT 108.590 96.790 110.210 96.890 ;
        RECT 109.510 96.350 110.210 96.790 ;
        RECT 111.440 96.690 113.320 96.900 ;
        RECT 114.160 96.870 116.270 97.000 ;
        RECT 114.600 96.760 116.270 96.870 ;
        RECT 117.020 96.940 118.930 97.130 ;
        RECT 120.020 96.990 122.020 97.190 ;
        RECT 122.720 97.140 123.420 97.560 ;
        RECT 124.460 97.510 126.830 97.560 ;
        RECT 127.490 97.550 129.860 97.560 ;
        RECT 130.470 97.560 132.885 97.790 ;
        RECT 126.110 97.240 126.810 97.510 ;
        RECT 122.720 97.010 125.250 97.140 ;
        RECT 126.110 97.050 128.120 97.240 ;
        RECT 128.960 97.160 129.660 97.550 ;
        RECT 130.470 97.490 132.840 97.560 ;
        RECT 133.460 97.510 135.900 97.860 ;
        RECT 138.120 97.850 138.820 97.880 ;
        RECT 141.380 97.850 142.700 97.860 ;
        RECT 117.020 96.840 119.350 96.940 ;
        RECT 112.620 96.370 113.320 96.690 ;
        RECT 115.570 96.370 116.270 96.760 ;
        RECT 117.420 96.710 119.350 96.840 ;
        RECT 120.020 96.820 122.200 96.990 ;
        RECT 122.720 96.880 125.460 97.010 ;
        RECT 120.510 96.770 122.200 96.820 ;
        RECT 106.540 96.080 108.925 96.330 ;
        RECT 97.870 95.760 101.310 96.040 ;
        RECT 106.540 96.030 108.910 96.080 ;
        RECT 109.510 96.050 111.880 96.350 ;
        RECT 112.540 96.330 114.910 96.370 ;
        RECT 112.540 96.080 114.915 96.330 ;
        RECT 112.540 96.070 114.910 96.080 ;
        RECT 115.500 96.070 117.870 96.370 ;
        RECT 118.650 96.350 119.350 96.710 ;
        RECT 118.490 96.330 120.860 96.350 ;
        RECT 121.500 96.330 122.200 96.770 ;
        RECT 123.080 96.740 125.460 96.880 ;
        RECT 126.110 96.870 128.200 97.050 ;
        RECT 128.960 96.960 130.970 97.160 ;
        RECT 132.140 97.090 132.780 97.490 ;
        RECT 132.140 97.000 133.730 97.090 ;
        RECT 128.960 96.880 131.200 96.960 ;
        RECT 132.140 96.930 134.260 97.000 ;
        RECT 134.580 96.970 135.900 97.510 ;
        RECT 136.740 97.330 138.880 97.850 ;
        RECT 139.460 97.500 144.890 97.850 ;
        RECT 145.460 97.810 150.860 97.850 ;
        RECT 145.455 97.560 150.860 97.810 ;
        RECT 145.460 97.510 150.860 97.560 ;
        RECT 151.440 97.510 154.400 100.150 ;
        RECT 141.380 97.490 142.700 97.500 ;
        RECT 138.240 97.090 138.840 97.330 ;
        RECT 141.780 97.310 142.290 97.490 ;
        RECT 147.900 97.340 148.410 97.510 ;
        RECT 134.580 96.950 136.860 96.970 ;
        RECT 138.240 96.950 139.850 97.090 ;
        RECT 126.200 96.820 128.200 96.870 ;
        RECT 124.760 96.340 125.460 96.740 ;
        RECT 127.500 96.360 128.200 96.820 ;
        RECT 129.050 96.740 131.200 96.880 ;
        RECT 132.670 96.800 134.260 96.930 ;
        RECT 124.460 96.330 126.830 96.340 ;
        RECT 127.490 96.330 129.860 96.360 ;
        RECT 130.500 96.350 131.200 96.740 ;
        RECT 133.520 96.380 134.260 96.800 ;
        RECT 135.430 96.860 136.860 96.950 ;
        RECT 135.430 96.730 137.610 96.860 ;
        RECT 118.490 96.080 120.905 96.330 ;
        RECT 121.495 96.320 123.600 96.330 ;
        RECT 121.495 96.080 123.870 96.320 ;
        RECT 112.620 96.020 113.320 96.070 ;
        RECT 115.570 96.040 116.270 96.070 ;
        RECT 118.490 96.050 120.860 96.080 ;
        RECT 118.650 95.980 119.350 96.050 ;
        RECT 121.500 96.020 123.870 96.080 ;
        RECT 124.460 96.080 126.895 96.330 ;
        RECT 127.485 96.080 129.860 96.330 ;
        RECT 124.460 96.040 126.830 96.080 ;
        RECT 127.490 96.060 129.860 96.080 ;
        RECT 130.490 96.330 132.860 96.350 ;
        RECT 133.480 96.330 135.920 96.380 ;
        RECT 136.560 96.370 137.610 96.730 ;
        RECT 138.330 96.790 139.850 96.950 ;
        RECT 138.330 96.690 141.580 96.790 ;
        RECT 130.490 96.080 132.885 96.330 ;
        RECT 133.475 96.080 135.920 96.330 ;
        RECT 130.490 96.050 132.860 96.080 ;
        RECT 130.500 96.000 131.200 96.050 ;
        RECT 133.480 96.030 135.920 96.080 ;
        RECT 136.440 96.020 138.880 96.370 ;
        RECT 139.440 96.360 141.580 96.690 ;
        RECT 139.440 96.270 141.900 96.360 ;
        RECT 139.460 96.010 141.900 96.270 ;
        RECT 97.870 95.410 100.320 95.760 ;
        RECT 97.870 95.390 98.920 95.410 ;
      LAYER met2 ;
        RECT 69.245 221.580 69.635 221.660 ;
        RECT 69.245 221.440 73.040 221.580 ;
        RECT 69.245 221.360 69.635 221.440 ;
        RECT 72.900 221.400 73.040 221.440 ;
        RECT 145.410 221.400 145.670 221.490 ;
        RECT 72.900 221.260 145.670 221.400 ;
        RECT 72.015 221.110 72.405 221.190 ;
        RECT 145.410 221.170 145.670 221.260 ;
        RECT 72.015 220.970 122.420 221.110 ;
        RECT 72.015 220.890 72.405 220.970 ;
        RECT 74.825 220.540 75.125 220.640 ;
        RECT 121.035 220.540 121.405 220.580 ;
        RECT 74.825 220.345 121.405 220.540 ;
        RECT 122.280 220.490 122.420 220.970 ;
        RECT 144.950 220.490 145.270 220.550 ;
        RECT 122.280 220.350 145.270 220.490 ;
        RECT 74.825 220.250 75.125 220.345 ;
        RECT 121.035 220.300 121.405 220.345 ;
        RECT 144.950 220.290 145.270 220.350 ;
        RECT 80.315 219.955 80.615 220.070 ;
        RECT 134.635 219.975 135.005 220.010 ;
        RECT 131.280 219.955 135.005 219.975 ;
        RECT 80.315 219.790 135.005 219.955 ;
        RECT 80.315 219.680 80.615 219.790 ;
        RECT 131.280 219.770 135.005 219.790 ;
        RECT 134.635 219.730 135.005 219.770 ;
        RECT 83.035 219.550 83.425 219.630 ;
        RECT 83.035 219.410 96.240 219.550 ;
        RECT 83.035 219.330 83.425 219.410 ;
        RECT 96.100 219.270 112.640 219.410 ;
        RECT 85.775 219.155 86.165 219.190 ;
        RECT 85.775 219.000 95.545 219.155 ;
        RECT 112.500 219.150 112.640 219.270 ;
        RECT 144.330 219.150 144.650 219.210 ;
        RECT 111.515 219.020 111.885 219.030 ;
        RECT 111.100 219.000 111.885 219.020 ;
        RECT 112.500 219.010 144.650 219.150 ;
        RECT 85.775 218.925 111.885 219.000 ;
        RECT 144.330 218.950 144.650 219.010 ;
        RECT 85.775 218.890 86.165 218.925 ;
        RECT 95.315 218.770 111.885 218.925 ;
        RECT 111.100 218.750 111.885 218.770 ;
        RECT 91.355 218.655 91.745 218.720 ;
        RECT 91.355 218.545 94.915 218.655 ;
        RECT 127.830 218.545 128.220 218.820 ;
        RECT 91.355 218.485 128.220 218.545 ;
        RECT 91.355 218.420 91.745 218.485 ;
        RECT 94.745 218.440 128.220 218.485 ;
        RECT 94.745 218.375 128.105 218.440 ;
        RECT 94.045 218.195 94.435 218.270 ;
        RECT 143.820 218.195 144.140 218.250 ;
        RECT 94.045 218.045 144.140 218.195 ;
        RECT 94.045 217.970 94.435 218.045 ;
        RECT 143.820 217.990 144.140 218.045 ;
        RECT 88.575 217.860 88.965 217.940 ;
        RECT 88.575 217.820 93.900 217.860 ;
        RECT 94.590 217.820 107.450 217.860 ;
        RECT 88.575 217.720 107.450 217.820 ;
        RECT 88.575 217.640 88.965 217.720 ;
        RECT 93.740 217.680 94.720 217.720 ;
        RECT 77.555 217.490 77.945 217.570 ;
        RECT 77.555 217.350 106.960 217.490 ;
        RECT 77.555 217.270 77.945 217.350 ;
        RECT 66.475 217.090 66.865 217.170 ;
        RECT 66.475 216.950 106.380 217.090 ;
        RECT 66.475 216.870 66.865 216.950 ;
        RECT 63.665 216.550 64.055 216.630 ;
        RECT 63.665 216.410 105.660 216.550 ;
        RECT 63.665 216.330 64.055 216.410 ;
        RECT 105.520 205.810 105.660 216.410 ;
        RECT 105.430 205.550 105.750 205.810 ;
        RECT 106.240 205.210 106.380 216.950 ;
        RECT 106.180 204.890 106.440 205.210 ;
        RECT 106.820 204.340 106.960 217.350 ;
        RECT 106.730 204.080 107.050 204.340 ;
        RECT 97.080 203.780 101.080 203.850 ;
        RECT 107.310 203.780 107.450 217.720 ;
        RECT 116.810 216.660 117.130 216.720 ;
        RECT 121.035 216.660 121.405 216.730 ;
        RECT 116.810 216.520 121.405 216.660 ;
        RECT 116.810 216.460 117.130 216.520 ;
        RECT 121.035 216.450 121.405 216.520 ;
        RECT 123.610 216.660 123.930 216.720 ;
        RECT 127.835 216.660 128.205 216.730 ;
        RECT 134.635 216.720 135.005 216.730 ;
        RECT 123.610 216.520 128.205 216.660 ;
        RECT 123.610 216.460 123.930 216.520 ;
        RECT 127.835 216.450 128.205 216.520 ;
        RECT 134.490 216.460 135.005 216.720 ;
        RECT 134.635 216.450 135.005 216.460 ;
        RECT 112.050 216.200 112.370 216.260 ;
        RECT 115.450 216.200 115.770 216.260 ;
        RECT 117.150 216.200 117.470 216.260 ;
        RECT 112.050 216.060 117.470 216.200 ;
        RECT 112.050 216.000 112.370 216.060 ;
        RECT 115.450 216.000 115.770 216.060 ;
        RECT 117.150 216.000 117.470 216.060 ;
        RECT 120.210 216.200 120.530 216.260 ;
        RECT 122.250 216.200 122.570 216.260 ;
        RECT 120.210 216.060 122.570 216.200 ;
        RECT 120.210 216.000 120.530 216.060 ;
        RECT 122.250 216.000 122.570 216.060 ;
        RECT 122.930 216.200 123.250 216.260 ;
        RECT 125.650 216.200 125.970 216.260 ;
        RECT 127.350 216.200 127.670 216.260 ;
        RECT 122.930 216.060 127.670 216.200 ;
        RECT 122.930 216.000 123.250 216.060 ;
        RECT 125.650 216.000 125.970 216.060 ;
        RECT 127.350 216.000 127.670 216.060 ;
        RECT 128.710 216.200 129.030 216.260 ;
        RECT 130.070 216.200 130.390 216.260 ;
        RECT 128.710 216.060 130.390 216.200 ;
        RECT 128.710 216.000 129.030 216.060 ;
        RECT 130.070 216.000 130.390 216.060 ;
        RECT 134.490 214.360 134.810 214.420 ;
        RECT 135.850 214.360 136.170 214.420 ;
        RECT 134.490 214.220 136.170 214.360 ;
        RECT 134.490 214.160 134.810 214.220 ;
        RECT 135.850 214.160 136.170 214.220 ;
        RECT 119.530 213.900 119.850 213.960 ;
        RECT 121.910 213.900 122.230 213.960 ;
        RECT 119.530 213.760 122.230 213.900 ;
        RECT 119.530 213.700 119.850 213.760 ;
        RECT 121.910 213.700 122.230 213.760 ;
        RECT 131.090 213.900 131.410 213.960 ;
        RECT 133.130 213.900 133.450 213.960 ;
        RECT 131.090 213.760 133.450 213.900 ;
        RECT 131.090 213.700 131.410 213.760 ;
        RECT 133.130 213.700 133.450 213.760 ;
        RECT 112.730 213.440 113.050 213.500 ;
        RECT 114.090 213.440 114.410 213.500 ;
        RECT 112.730 213.300 114.410 213.440 ;
        RECT 112.730 213.240 113.050 213.300 ;
        RECT 114.090 213.240 114.410 213.300 ;
        RECT 139.930 212.060 140.250 212.120 ;
        RECT 141.630 212.060 141.950 212.120 ;
        RECT 139.930 211.920 141.950 212.060 ;
        RECT 139.930 211.860 140.250 211.920 ;
        RECT 141.630 211.860 141.950 211.920 ;
        RECT 112.730 211.600 113.050 211.660 ;
        RECT 116.470 211.600 116.790 211.660 ;
        RECT 112.730 211.460 116.790 211.600 ;
        RECT 112.730 211.400 113.050 211.460 ;
        RECT 116.470 211.400 116.790 211.460 ;
        RECT 126.330 211.600 126.650 211.660 ;
        RECT 130.070 211.600 130.390 211.660 ;
        RECT 126.330 211.460 130.390 211.600 ;
        RECT 126.330 211.400 126.650 211.460 ;
        RECT 130.070 211.400 130.390 211.460 ;
        RECT 112.730 211.140 113.050 211.200 ;
        RECT 116.810 211.140 117.130 211.200 ;
        RECT 122.590 211.140 122.910 211.200 ;
        RECT 112.730 211.000 122.910 211.140 ;
        RECT 112.730 210.940 113.050 211.000 ;
        RECT 116.810 210.940 117.130 211.000 ;
        RECT 122.590 210.940 122.910 211.000 ;
        RECT 123.610 211.140 123.930 211.200 ;
        RECT 124.630 211.140 124.950 211.200 ;
        RECT 123.610 211.000 124.950 211.140 ;
        RECT 123.610 210.940 123.930 211.000 ;
        RECT 124.630 210.940 124.950 211.000 ;
        RECT 122.590 210.680 122.910 210.740 ;
        RECT 130.410 210.680 130.730 210.740 ;
        RECT 133.470 210.680 133.790 210.740 ;
        RECT 122.590 210.540 133.790 210.680 ;
        RECT 122.590 210.480 122.910 210.540 ;
        RECT 130.410 210.480 130.730 210.540 ;
        RECT 133.470 210.480 133.790 210.540 ;
        RECT 114.770 209.300 115.090 209.360 ;
        RECT 119.870 209.300 120.190 209.360 ;
        RECT 114.770 209.160 120.190 209.300 ;
        RECT 114.770 209.100 115.090 209.160 ;
        RECT 119.870 209.100 120.190 209.160 ;
        RECT 128.370 209.300 128.690 209.360 ;
        RECT 130.750 209.300 131.070 209.360 ;
        RECT 128.370 209.160 131.070 209.300 ;
        RECT 128.370 209.100 128.690 209.160 ;
        RECT 130.750 209.100 131.070 209.160 ;
        RECT 133.810 209.300 134.130 209.360 ;
        RECT 135.510 209.300 135.830 209.360 ;
        RECT 133.810 209.160 135.830 209.300 ;
        RECT 133.810 209.100 134.130 209.160 ;
        RECT 135.510 209.100 135.830 209.160 ;
        RECT 112.730 208.840 113.050 208.900 ;
        RECT 117.150 208.840 117.470 208.900 ;
        RECT 112.730 208.700 117.470 208.840 ;
        RECT 112.730 208.640 113.050 208.700 ;
        RECT 117.150 208.640 117.470 208.700 ;
        RECT 134.490 208.840 134.810 208.900 ;
        RECT 135.510 208.840 135.830 208.900 ;
        RECT 134.490 208.700 135.830 208.840 ;
        RECT 134.490 208.640 134.810 208.700 ;
        RECT 135.510 208.640 135.830 208.700 ;
        RECT 117.490 208.380 117.810 208.440 ;
        RECT 120.890 208.380 121.210 208.440 ;
        RECT 125.310 208.380 125.630 208.440 ;
        RECT 117.490 208.240 125.630 208.380 ;
        RECT 117.490 208.180 117.810 208.240 ;
        RECT 120.890 208.180 121.210 208.240 ;
        RECT 125.310 208.180 125.630 208.240 ;
        RECT 139.930 207.460 140.250 207.520 ;
        RECT 141.630 207.460 141.950 207.520 ;
        RECT 139.930 207.320 141.950 207.460 ;
        RECT 139.930 207.260 140.250 207.320 ;
        RECT 141.630 207.260 141.950 207.320 ;
        RECT 139.395 207.000 139.765 207.070 ;
        RECT 141.630 207.000 141.950 207.060 ;
        RECT 139.395 206.860 141.950 207.000 ;
        RECT 139.395 206.790 139.765 206.860 ;
        RECT 141.630 206.800 141.950 206.860 ;
        RECT 108.990 206.540 109.310 206.600 ;
        RECT 112.730 206.540 113.050 206.600 ;
        RECT 108.990 206.400 113.050 206.540 ;
        RECT 108.990 206.340 109.310 206.400 ;
        RECT 112.730 206.340 113.050 206.400 ;
        RECT 130.750 206.540 131.070 206.600 ;
        RECT 134.490 206.540 134.810 206.600 ;
        RECT 136.190 206.540 136.510 206.600 ;
        RECT 138.230 206.540 138.550 206.600 ;
        RECT 130.750 206.400 138.550 206.540 ;
        RECT 130.750 206.340 131.070 206.400 ;
        RECT 134.490 206.340 134.810 206.400 ;
        RECT 136.190 206.340 136.510 206.400 ;
        RECT 138.230 206.340 138.550 206.400 ;
        RECT 128.710 205.620 129.030 205.680 ;
        RECT 138.035 205.620 138.405 205.690 ;
        RECT 128.710 205.480 138.405 205.620 ;
        RECT 128.710 205.420 129.030 205.480 ;
        RECT 138.035 205.410 138.405 205.480 ;
        RECT 139.590 205.160 139.910 205.220 ;
        RECT 140.950 205.160 141.270 205.220 ;
        RECT 139.590 205.020 141.270 205.160 ;
        RECT 139.590 204.960 139.910 205.020 ;
        RECT 140.950 204.960 141.270 205.020 ;
        RECT 111.710 204.700 112.030 204.760 ;
        RECT 117.150 204.700 117.470 204.760 ;
        RECT 123.270 204.700 123.590 204.760 ;
        RECT 111.710 204.560 123.590 204.700 ;
        RECT 111.710 204.500 112.030 204.560 ;
        RECT 117.150 204.500 117.470 204.560 ;
        RECT 123.270 204.500 123.590 204.560 ;
        RECT 131.090 204.240 131.410 204.300 ;
        RECT 134.490 204.240 134.810 204.300 ;
        RECT 131.090 204.100 134.810 204.240 ;
        RECT 131.090 204.040 131.410 204.100 ;
        RECT 134.490 204.040 134.810 204.100 ;
        RECT 137.210 204.240 137.530 204.300 ;
        RECT 139.250 204.240 139.570 204.300 ;
        RECT 137.210 204.100 139.570 204.240 ;
        RECT 137.210 204.040 137.530 204.100 ;
        RECT 139.250 204.040 139.570 204.100 ;
        RECT 108.310 203.780 108.630 203.840 ;
        RECT 97.080 203.640 108.630 203.780 ;
        RECT 97.080 203.570 101.080 203.640 ;
        RECT 108.310 203.580 108.630 203.640 ;
        RECT 142.650 203.780 142.970 203.840 ;
        RECT 145.380 203.780 145.700 203.870 ;
        RECT 150.845 203.780 154.845 203.850 ;
        RECT 142.650 203.640 154.845 203.780 ;
        RECT 142.650 203.580 142.970 203.640 ;
        RECT 145.380 203.550 145.700 203.640 ;
        RECT 150.845 203.570 154.845 203.640 ;
        RECT 119.530 203.320 119.850 203.380 ;
        RECT 122.250 203.320 122.570 203.380 ;
        RECT 119.530 203.180 122.570 203.320 ;
        RECT 119.530 203.120 119.850 203.180 ;
        RECT 122.250 203.120 122.570 203.180 ;
        RECT 123.270 203.320 123.590 203.380 ;
        RECT 126.330 203.320 126.650 203.380 ;
        RECT 131.770 203.320 132.090 203.380 ;
        RECT 134.490 203.320 134.810 203.380 ;
        RECT 123.270 203.180 134.810 203.320 ;
        RECT 123.270 203.120 123.590 203.180 ;
        RECT 126.330 203.120 126.650 203.180 ;
        RECT 131.770 203.120 132.090 203.180 ;
        RECT 134.490 203.120 134.810 203.180 ;
        RECT 123.610 202.860 123.930 202.920 ;
        RECT 125.310 202.860 125.630 202.920 ;
        RECT 123.610 202.720 125.630 202.860 ;
        RECT 123.610 202.660 123.930 202.720 ;
        RECT 125.310 202.660 125.630 202.720 ;
        RECT 126.330 202.860 126.650 202.920 ;
        RECT 139.395 202.860 139.765 202.930 ;
        RECT 126.330 202.720 139.765 202.860 ;
        RECT 126.330 202.660 126.650 202.720 ;
        RECT 139.395 202.650 139.765 202.720 ;
        RECT 108.990 201.280 109.310 201.540 ;
        RECT 106.930 201.020 107.190 201.110 ;
        RECT 108.310 201.020 108.630 201.080 ;
        RECT 102.790 200.880 108.630 201.020 ;
        RECT 97.080 200.560 101.080 200.630 ;
        RECT 102.790 200.560 102.930 200.880 ;
        RECT 106.930 200.790 107.190 200.880 ;
        RECT 108.310 200.820 108.630 200.880 ;
        RECT 97.080 200.420 102.930 200.560 ;
        RECT 97.080 200.350 101.080 200.420 ;
        RECT 109.080 200.100 109.220 201.280 ;
        RECT 110.495 200.650 110.865 202.190 ;
        RECT 115.935 200.650 116.305 202.190 ;
        RECT 121.375 200.650 121.745 202.190 ;
        RECT 126.815 200.650 127.185 202.190 ;
        RECT 132.255 200.650 132.625 202.190 ;
        RECT 137.695 200.650 138.065 202.190 ;
        RECT 143.135 200.650 143.505 202.190 ;
        RECT 150.845 200.560 154.845 200.630 ;
        RECT 144.270 200.420 154.845 200.560 ;
        RECT 112.730 200.100 113.050 200.160 ;
        RECT 116.470 200.100 116.790 200.160 ;
        RECT 109.080 199.960 112.450 200.100 ;
        RECT 112.310 199.240 112.450 199.960 ;
        RECT 112.730 199.960 116.790 200.100 ;
        RECT 112.730 199.900 113.050 199.960 ;
        RECT 116.470 199.900 116.790 199.960 ;
        RECT 125.310 200.100 125.630 200.160 ;
        RECT 135.510 200.100 135.830 200.160 ;
        RECT 125.310 199.960 135.830 200.100 ;
        RECT 125.310 199.900 125.630 199.960 ;
        RECT 135.510 199.900 135.830 199.960 ;
        RECT 136.190 200.100 136.510 200.160 ;
        RECT 140.950 200.100 141.270 200.160 ;
        RECT 136.190 199.960 141.270 200.100 ;
        RECT 136.190 199.900 136.510 199.960 ;
        RECT 140.950 199.900 141.270 199.960 ;
        RECT 144.270 199.770 144.410 200.420 ;
        RECT 150.845 200.350 154.845 200.420 ;
        RECT 144.020 199.760 144.410 199.770 ;
        RECT 114.430 199.640 114.750 199.700 ;
        RECT 127.350 199.640 127.670 199.700 ;
        RECT 133.810 199.640 134.130 199.700 ;
        RECT 114.430 199.500 134.130 199.640 ;
        RECT 114.430 199.440 114.750 199.500 ;
        RECT 127.350 199.440 127.670 199.500 ;
        RECT 133.810 199.440 134.130 199.500 ;
        RECT 134.490 199.640 134.810 199.700 ;
        RECT 136.190 199.640 136.510 199.700 ;
        RECT 134.490 199.500 136.510 199.640 ;
        RECT 134.490 199.440 134.810 199.500 ;
        RECT 136.190 199.440 136.510 199.500 ;
        RECT 138.570 199.640 138.890 199.700 ;
        RECT 143.810 199.640 144.410 199.760 ;
        RECT 138.570 199.500 144.410 199.640 ;
        RECT 138.570 199.440 138.890 199.500 ;
        RECT 143.810 199.370 144.160 199.500 ;
        RECT 108.650 199.180 108.970 199.240 ;
        RECT 111.030 199.180 111.350 199.240 ;
        RECT 108.650 199.040 111.350 199.180 ;
        RECT 112.310 199.180 112.710 199.240 ;
        RECT 115.450 199.180 115.770 199.240 ;
        RECT 117.490 199.180 117.810 199.240 ;
        RECT 119.190 199.180 119.510 199.240 ;
        RECT 112.310 199.040 119.510 199.180 ;
        RECT 108.650 198.980 108.970 199.040 ;
        RECT 111.030 198.980 111.350 199.040 ;
        RECT 112.390 198.980 112.710 199.040 ;
        RECT 115.450 198.980 115.770 199.040 ;
        RECT 117.490 198.980 117.810 199.040 ;
        RECT 119.190 198.980 119.510 199.040 ;
        RECT 125.310 199.180 125.630 199.240 ;
        RECT 128.030 199.180 128.350 199.240 ;
        RECT 132.790 199.180 133.110 199.240 ;
        RECT 125.310 199.040 128.350 199.180 ;
        RECT 125.310 198.980 125.630 199.040 ;
        RECT 128.030 198.980 128.350 199.040 ;
        RECT 128.630 199.040 133.110 199.180 ;
        RECT 97.080 197.340 101.080 197.410 ;
        RECT 107.775 197.350 108.145 198.890 ;
        RECT 113.215 197.350 113.585 198.890 ;
        RECT 118.655 197.350 119.025 198.890 ;
        RECT 124.095 197.350 124.465 198.890 ;
        RECT 125.990 198.720 126.310 198.780 ;
        RECT 128.630 198.720 128.770 199.040 ;
        RECT 132.790 198.980 133.110 199.040 ;
        RECT 137.210 199.180 137.530 199.240 ;
        RECT 142.310 199.180 142.630 199.240 ;
        RECT 137.210 199.040 142.630 199.180 ;
        RECT 137.210 198.980 137.530 199.040 ;
        RECT 142.310 198.980 142.630 199.040 ;
        RECT 125.990 198.580 128.770 198.720 ;
        RECT 125.990 198.520 126.310 198.580 ;
        RECT 129.535 197.350 129.905 198.890 ;
        RECT 134.975 197.350 135.345 198.890 ;
        RECT 136.190 198.720 136.510 198.780 ;
        RECT 138.910 198.720 139.230 198.780 ;
        RECT 136.190 198.580 139.230 198.720 ;
        RECT 136.190 198.520 136.510 198.580 ;
        RECT 138.910 198.520 139.230 198.580 ;
        RECT 140.415 197.350 140.785 198.890 ;
        RECT 142.650 197.340 142.970 197.400 ;
        RECT 144.360 197.340 144.620 197.430 ;
        RECT 150.845 197.340 154.845 197.410 ;
        RECT 97.080 197.200 102.930 197.340 ;
        RECT 97.080 197.130 101.080 197.200 ;
        RECT 102.790 196.880 102.930 197.200 ;
        RECT 142.650 197.200 154.845 197.340 ;
        RECT 142.650 197.140 142.970 197.200 ;
        RECT 144.360 197.110 144.620 197.200 ;
        RECT 150.845 197.130 154.845 197.200 ;
        RECT 106.300 196.880 106.700 197.030 ;
        RECT 108.310 196.880 108.630 196.940 ;
        RECT 102.790 196.740 108.630 196.880 ;
        RECT 106.300 196.640 106.700 196.740 ;
        RECT 108.310 196.680 108.630 196.740 ;
        RECT 122.590 196.880 122.910 196.940 ;
        RECT 130.070 196.880 130.390 196.940 ;
        RECT 131.770 196.880 132.090 196.940 ;
        RECT 136.190 196.880 136.510 196.940 ;
        RECT 122.590 196.740 131.490 196.880 ;
        RECT 122.590 196.680 122.910 196.740 ;
        RECT 130.070 196.680 130.390 196.740 ;
        RECT 110.010 196.420 110.330 196.480 ;
        RECT 119.190 196.420 119.510 196.480 ;
        RECT 122.590 196.420 122.910 196.480 ;
        RECT 110.010 196.280 122.910 196.420 ;
        RECT 110.010 196.220 110.330 196.280 ;
        RECT 119.190 196.220 119.510 196.280 ;
        RECT 122.590 196.220 122.910 196.280 ;
        RECT 129.050 196.420 129.370 196.480 ;
        RECT 130.410 196.420 130.730 196.480 ;
        RECT 129.050 196.280 130.730 196.420 ;
        RECT 131.350 196.420 131.490 196.740 ;
        RECT 131.770 196.740 136.510 196.880 ;
        RECT 131.770 196.680 132.090 196.740 ;
        RECT 136.190 196.680 136.510 196.740 ;
        RECT 139.930 196.880 140.250 196.940 ;
        RECT 141.630 196.880 141.950 196.940 ;
        RECT 139.930 196.740 141.950 196.880 ;
        RECT 139.930 196.680 140.250 196.740 ;
        RECT 141.630 196.680 141.950 196.740 ;
        RECT 136.190 196.420 136.510 196.480 ;
        RECT 131.350 196.280 136.510 196.420 ;
        RECT 129.050 196.220 129.370 196.280 ;
        RECT 130.410 196.220 130.730 196.280 ;
        RECT 136.190 196.220 136.510 196.280 ;
        RECT 139.590 196.420 139.910 196.480 ;
        RECT 140.950 196.420 141.270 196.480 ;
        RECT 139.590 196.280 141.270 196.420 ;
        RECT 139.590 196.220 139.910 196.280 ;
        RECT 140.950 196.220 141.270 196.280 ;
        RECT 120.210 195.960 120.530 196.020 ;
        RECT 120.210 195.760 120.610 195.960 ;
        RECT 123.610 195.760 123.930 196.020 ;
        RECT 130.750 195.960 131.070 196.020 ;
        RECT 133.470 195.960 133.790 196.020 ;
        RECT 130.750 195.820 133.790 195.960 ;
        RECT 130.750 195.760 131.070 195.820 ;
        RECT 133.470 195.760 133.790 195.820 ;
        RECT 136.530 195.960 136.850 196.020 ;
        RECT 138.230 195.960 138.550 196.020 ;
        RECT 136.530 195.820 138.550 195.960 ;
        RECT 136.530 195.760 136.850 195.820 ;
        RECT 138.230 195.760 138.550 195.820 ;
        RECT 120.470 195.500 120.610 195.760 ;
        RECT 123.700 195.500 123.840 195.760 ;
        RECT 125.650 195.500 125.970 195.560 ;
        RECT 131.430 195.500 131.750 195.560 ;
        RECT 120.470 195.360 131.750 195.500 ;
        RECT 125.650 195.300 125.970 195.360 ;
        RECT 131.430 195.300 131.750 195.360 ;
        RECT 136.190 195.500 136.510 195.560 ;
        RECT 139.250 195.500 139.570 195.560 ;
        RECT 136.190 195.360 139.570 195.500 ;
        RECT 136.190 195.300 136.510 195.360 ;
        RECT 139.250 195.300 139.570 195.360 ;
        RECT 120.550 195.040 120.870 195.100 ;
        RECT 130.410 195.040 130.730 195.100 ;
        RECT 120.550 194.900 130.730 195.040 ;
        RECT 120.550 194.840 120.870 194.900 ;
        RECT 130.410 194.840 130.730 194.900 ;
        RECT 112.730 194.580 113.050 194.640 ;
        RECT 117.830 194.580 118.150 194.640 ;
        RECT 122.250 194.580 122.570 194.640 ;
        RECT 112.730 194.440 122.570 194.580 ;
        RECT 112.730 194.380 113.050 194.440 ;
        RECT 117.830 194.380 118.150 194.440 ;
        RECT 122.250 194.380 122.570 194.440 ;
        RECT 125.990 194.580 126.310 194.640 ;
        RECT 127.350 194.580 127.670 194.640 ;
        RECT 134.150 194.580 134.470 194.640 ;
        RECT 138.910 194.580 139.230 194.640 ;
        RECT 125.990 194.440 139.230 194.580 ;
        RECT 125.990 194.380 126.310 194.440 ;
        RECT 127.350 194.380 127.670 194.440 ;
        RECT 134.150 194.380 134.470 194.440 ;
        RECT 138.910 194.380 139.230 194.440 ;
        RECT 129.050 194.120 129.370 194.180 ;
        RECT 133.130 194.120 133.450 194.180 ;
        RECT 135.850 194.120 136.170 194.180 ;
        RECT 137.210 194.120 137.530 194.180 ;
        RECT 139.250 194.120 139.570 194.180 ;
        RECT 129.050 193.980 136.170 194.120 ;
        RECT 129.050 193.920 129.370 193.980 ;
        RECT 133.130 193.920 133.450 193.980 ;
        RECT 135.850 193.920 136.170 193.980 ;
        RECT 136.790 193.980 139.570 194.120 ;
        RECT 111.710 193.660 112.030 193.720 ;
        RECT 117.490 193.660 117.810 193.720 ;
        RECT 120.890 193.660 121.210 193.720 ;
        RECT 136.790 193.660 136.930 193.980 ;
        RECT 137.210 193.920 137.530 193.980 ;
        RECT 139.250 193.920 139.570 193.980 ;
        RECT 141.630 194.120 141.950 194.180 ;
        RECT 143.775 194.120 144.165 194.200 ;
        RECT 150.845 194.120 154.845 194.190 ;
        RECT 141.630 193.980 154.845 194.120 ;
        RECT 141.630 193.920 141.950 193.980 ;
        RECT 143.775 193.900 144.165 193.980 ;
        RECT 150.845 193.910 154.845 193.980 ;
        RECT 111.710 193.520 136.930 193.660 ;
        RECT 111.710 193.460 112.030 193.520 ;
        RECT 117.490 193.460 117.810 193.520 ;
        RECT 120.890 193.460 121.210 193.520 ;
        RECT 108.990 193.200 109.310 193.260 ;
        RECT 109.670 193.200 109.990 193.260 ;
        RECT 111.710 193.200 112.030 193.260 ;
        RECT 108.990 193.060 112.030 193.200 ;
        RECT 108.990 193.000 109.310 193.060 ;
        RECT 109.670 193.000 109.990 193.060 ;
        RECT 111.710 193.000 112.030 193.060 ;
        RECT 136.190 193.200 136.510 193.260 ;
        RECT 138.230 193.200 138.550 193.260 ;
        RECT 136.190 193.060 138.550 193.200 ;
        RECT 136.190 193.000 136.510 193.060 ;
        RECT 138.230 193.000 138.550 193.060 ;
        RECT 116.470 192.740 116.790 192.800 ;
        RECT 117.150 192.740 117.470 192.800 ;
        RECT 124.630 192.740 124.950 192.800 ;
        RECT 116.470 192.600 124.950 192.740 ;
        RECT 116.470 192.540 116.790 192.600 ;
        RECT 117.150 192.540 117.470 192.600 ;
        RECT 124.630 192.540 124.950 192.600 ;
        RECT 110.835 192.280 111.205 192.350 ;
        RECT 114.430 192.280 114.750 192.340 ;
        RECT 110.835 192.140 114.750 192.280 ;
        RECT 110.835 192.070 111.205 192.140 ;
        RECT 114.430 192.080 114.750 192.140 ;
        RECT 122.930 192.280 123.250 192.340 ;
        RECT 126.330 192.280 126.650 192.340 ;
        RECT 132.790 192.280 133.110 192.340 ;
        RECT 122.930 192.140 133.110 192.280 ;
        RECT 122.930 192.080 123.250 192.140 ;
        RECT 126.330 192.080 126.650 192.140 ;
        RECT 132.790 192.080 133.110 192.140 ;
        RECT 139.250 192.280 139.570 192.340 ;
        RECT 142.310 192.280 142.630 192.340 ;
        RECT 139.250 192.140 142.630 192.280 ;
        RECT 139.250 192.080 139.570 192.140 ;
        RECT 142.310 192.080 142.630 192.140 ;
        RECT 128.370 191.360 128.690 191.420 ;
        RECT 130.070 191.360 130.390 191.420 ;
        RECT 128.370 191.220 130.390 191.360 ;
        RECT 128.370 191.160 128.690 191.220 ;
        RECT 130.070 191.160 130.390 191.220 ;
        RECT 97.080 190.900 101.080 190.970 ;
        RECT 105.390 190.900 105.790 191.010 ;
        RECT 108.310 190.900 108.630 190.960 ;
        RECT 97.080 190.760 108.630 190.900 ;
        RECT 97.080 190.690 101.080 190.760 ;
        RECT 105.390 190.620 105.790 190.760 ;
        RECT 108.310 190.700 108.630 190.760 ;
        RECT 114.430 190.900 114.750 190.960 ;
        RECT 121.035 190.900 121.405 190.970 ;
        RECT 114.430 190.760 121.405 190.900 ;
        RECT 114.430 190.700 114.750 190.760 ;
        RECT 121.035 190.690 121.405 190.760 ;
        RECT 142.650 190.900 142.970 190.960 ;
        RECT 144.940 190.900 145.270 191.000 ;
        RECT 150.845 190.900 154.845 190.970 ;
        RECT 142.650 190.760 154.845 190.900 ;
        RECT 142.650 190.700 142.970 190.760 ;
        RECT 144.940 190.660 145.270 190.760 ;
        RECT 150.845 190.690 154.845 190.760 ;
        RECT 108.990 190.440 109.310 190.500 ;
        RECT 116.470 190.440 116.790 190.500 ;
        RECT 119.870 190.440 120.190 190.500 ;
        RECT 108.990 190.300 120.190 190.440 ;
        RECT 108.990 190.240 109.310 190.300 ;
        RECT 116.470 190.240 116.790 190.300 ;
        RECT 119.870 190.240 120.190 190.300 ;
        RECT 128.370 190.440 128.690 190.500 ;
        RECT 133.810 190.440 134.130 190.500 ;
        RECT 140.950 190.440 141.270 190.500 ;
        RECT 128.370 190.300 141.270 190.440 ;
        RECT 128.370 190.240 128.690 190.300 ;
        RECT 133.810 190.240 134.130 190.300 ;
        RECT 140.950 190.240 141.270 190.300 ;
        RECT 122.930 189.980 123.250 190.040 ;
        RECT 124.630 189.980 124.950 190.040 ;
        RECT 122.930 189.840 124.950 189.980 ;
        RECT 122.930 189.780 123.250 189.840 ;
        RECT 124.630 189.780 124.950 189.840 ;
        RECT 134.150 189.980 134.470 190.040 ;
        RECT 134.150 189.840 139.480 189.980 ;
        RECT 134.150 189.780 134.470 189.840 ;
        RECT 139.340 189.590 139.480 189.840 ;
        RECT 114.235 189.580 114.605 189.590 ;
        RECT 139.340 189.580 139.765 189.590 ;
        RECT 114.235 189.320 114.750 189.580 ;
        RECT 118.170 189.520 118.490 189.580 ;
        RECT 119.190 189.520 119.510 189.580 ;
        RECT 118.170 189.380 119.510 189.520 ;
        RECT 118.170 189.320 118.490 189.380 ;
        RECT 119.190 189.320 119.510 189.380 ;
        RECT 125.310 189.520 125.630 189.580 ;
        RECT 130.750 189.520 131.070 189.580 ;
        RECT 133.130 189.520 133.450 189.580 ;
        RECT 134.150 189.520 134.470 189.580 ;
        RECT 125.310 189.380 126.050 189.520 ;
        RECT 125.310 189.320 125.630 189.380 ;
        RECT 114.235 189.310 114.605 189.320 ;
        RECT 124.435 188.600 124.805 188.670 ;
        RECT 125.310 188.600 125.630 188.660 ;
        RECT 124.435 188.460 125.630 188.600 ;
        RECT 125.910 188.600 126.050 189.380 ;
        RECT 130.750 189.380 134.470 189.520 ;
        RECT 130.750 189.320 131.070 189.380 ;
        RECT 133.130 189.320 133.450 189.380 ;
        RECT 134.150 189.320 134.470 189.380 ;
        RECT 139.250 189.320 139.765 189.580 ;
        RECT 139.395 189.310 139.765 189.320 ;
        RECT 137.210 189.060 137.530 189.120 ;
        RECT 138.570 189.060 138.890 189.120 ;
        RECT 141.630 189.060 141.950 189.120 ;
        RECT 137.210 188.920 141.950 189.060 ;
        RECT 137.210 188.860 137.530 188.920 ;
        RECT 138.570 188.860 138.890 188.920 ;
        RECT 141.630 188.860 141.950 188.920 ;
        RECT 131.430 188.600 131.750 188.660 ;
        RECT 125.910 188.460 131.750 188.600 ;
        RECT 124.435 188.390 124.805 188.460 ;
        RECT 125.310 188.400 125.630 188.460 ;
        RECT 131.430 188.400 131.750 188.460 ;
        RECT 109.330 188.140 109.650 188.200 ;
        RECT 111.710 188.140 112.030 188.200 ;
        RECT 113.750 188.140 114.070 188.200 ;
        RECT 109.330 188.000 114.070 188.140 ;
        RECT 109.330 187.940 109.650 188.000 ;
        RECT 111.710 187.940 112.030 188.000 ;
        RECT 113.750 187.940 114.070 188.000 ;
        RECT 120.210 188.140 120.530 188.200 ;
        RECT 123.270 188.140 123.590 188.200 ;
        RECT 124.970 188.140 125.290 188.200 ;
        RECT 127.350 188.140 127.670 188.200 ;
        RECT 120.210 188.000 127.670 188.140 ;
        RECT 120.210 187.940 120.530 188.000 ;
        RECT 123.270 187.940 123.590 188.000 ;
        RECT 124.970 187.940 125.290 188.000 ;
        RECT 127.350 187.940 127.670 188.000 ;
        RECT 107.435 187.680 107.805 187.750 ;
        RECT 108.990 187.680 109.310 187.740 ;
        RECT 107.435 187.540 109.310 187.680 ;
        RECT 107.435 187.470 107.805 187.540 ;
        RECT 108.990 187.480 109.310 187.540 ;
        RECT 112.050 187.680 112.370 187.740 ;
        RECT 113.750 187.680 114.070 187.740 ;
        RECT 112.050 187.540 114.070 187.680 ;
        RECT 112.050 187.480 112.370 187.540 ;
        RECT 113.750 187.480 114.070 187.540 ;
        RECT 115.450 187.680 115.770 187.740 ;
        RECT 117.150 187.680 117.470 187.740 ;
        RECT 119.870 187.680 120.190 187.740 ;
        RECT 115.450 187.540 120.190 187.680 ;
        RECT 115.450 187.480 115.770 187.540 ;
        RECT 117.150 187.480 117.470 187.540 ;
        RECT 119.870 187.480 120.190 187.540 ;
        RECT 120.890 187.680 121.210 187.740 ;
        RECT 131.090 187.680 131.410 187.740 ;
        RECT 120.890 187.540 131.410 187.680 ;
        RECT 120.890 187.480 121.210 187.540 ;
        RECT 131.090 187.480 131.410 187.540 ;
        RECT 117.635 187.280 118.005 187.290 ;
        RECT 109.670 187.220 109.990 187.280 ;
        RECT 115.110 187.220 115.430 187.280 ;
        RECT 109.670 187.080 115.430 187.220 ;
        RECT 109.670 187.020 109.990 187.080 ;
        RECT 115.110 187.020 115.430 187.080 ;
        RECT 117.490 187.020 118.005 187.280 ;
        RECT 136.190 187.220 136.510 187.280 ;
        RECT 138.230 187.220 138.550 187.280 ;
        RECT 136.190 187.080 138.550 187.220 ;
        RECT 136.190 187.020 136.510 187.080 ;
        RECT 138.230 187.020 138.550 187.080 ;
        RECT 117.635 187.010 118.005 187.020 ;
        RECT 110.010 186.760 110.330 186.820 ;
        RECT 114.430 186.760 114.750 186.820 ;
        RECT 116.470 186.760 116.790 186.820 ;
        RECT 122.930 186.760 123.250 186.820 ;
        RECT 110.010 186.620 123.250 186.760 ;
        RECT 110.010 186.560 110.330 186.620 ;
        RECT 114.430 186.560 114.750 186.620 ;
        RECT 116.470 186.560 116.790 186.620 ;
        RECT 122.930 186.560 123.250 186.620 ;
        RECT 130.750 186.760 131.070 186.820 ;
        RECT 133.810 186.760 134.130 186.820 ;
        RECT 134.490 186.760 134.810 186.820 ;
        RECT 140.950 186.760 141.270 186.820 ;
        RECT 130.750 186.620 141.270 186.760 ;
        RECT 130.750 186.560 131.070 186.620 ;
        RECT 133.810 186.560 134.130 186.620 ;
        RECT 134.490 186.560 134.810 186.620 ;
        RECT 140.950 186.560 141.270 186.620 ;
        RECT 115.450 186.300 115.770 186.360 ;
        RECT 122.930 186.300 123.250 186.360 ;
        RECT 115.450 186.160 123.250 186.300 ;
        RECT 115.450 186.100 115.770 186.160 ;
        RECT 122.930 186.100 123.250 186.160 ;
        RECT 123.610 186.300 123.930 186.360 ;
        RECT 125.310 186.300 125.630 186.360 ;
        RECT 123.610 186.160 125.630 186.300 ;
        RECT 123.610 186.100 123.930 186.160 ;
        RECT 125.310 186.100 125.630 186.160 ;
        RECT 125.990 186.300 126.310 186.360 ;
        RECT 130.750 186.300 131.070 186.360 ;
        RECT 137.210 186.300 137.530 186.360 ;
        RECT 139.250 186.300 139.570 186.360 ;
        RECT 125.990 186.160 136.930 186.300 ;
        RECT 125.990 186.100 126.310 186.160 ;
        RECT 130.750 186.100 131.070 186.160 ;
        RECT 114.430 185.840 114.750 185.900 ;
        RECT 117.490 185.840 117.810 185.900 ;
        RECT 114.430 185.700 117.810 185.840 ;
        RECT 114.430 185.640 114.750 185.700 ;
        RECT 117.490 185.640 117.810 185.700 ;
        RECT 118.170 185.840 118.490 185.900 ;
        RECT 122.590 185.840 122.910 185.900 ;
        RECT 118.170 185.700 122.910 185.840 ;
        RECT 118.170 185.640 118.490 185.700 ;
        RECT 122.590 185.640 122.910 185.700 ;
        RECT 125.310 185.840 125.630 185.900 ;
        RECT 128.370 185.840 128.690 185.900 ;
        RECT 125.310 185.700 128.690 185.840 ;
        RECT 125.310 185.640 125.630 185.700 ;
        RECT 128.370 185.640 128.690 185.700 ;
        RECT 131.235 185.840 131.605 185.910 ;
        RECT 136.190 185.840 136.510 185.900 ;
        RECT 131.235 185.700 136.510 185.840 ;
        RECT 136.790 185.840 136.930 186.160 ;
        RECT 137.210 186.160 139.570 186.300 ;
        RECT 137.210 186.100 137.530 186.160 ;
        RECT 139.250 186.100 139.570 186.160 ;
        RECT 141.630 186.300 141.950 186.360 ;
        RECT 144.835 186.300 145.205 186.370 ;
        RECT 141.630 186.160 145.205 186.300 ;
        RECT 141.630 186.100 141.950 186.160 ;
        RECT 144.835 186.090 145.205 186.160 ;
        RECT 138.570 185.840 138.890 185.900 ;
        RECT 136.790 185.700 138.890 185.840 ;
        RECT 131.235 185.630 131.605 185.700 ;
        RECT 136.190 185.640 136.510 185.700 ;
        RECT 138.570 185.640 138.890 185.700 ;
        RECT 117.830 185.380 118.150 185.440 ;
        RECT 119.870 185.380 120.190 185.440 ;
        RECT 124.970 185.380 125.290 185.440 ;
        RECT 117.830 185.240 125.290 185.380 ;
        RECT 117.830 185.180 118.150 185.240 ;
        RECT 119.870 185.180 120.190 185.240 ;
        RECT 124.970 185.180 125.290 185.240 ;
        RECT 131.770 185.380 132.090 185.440 ;
        RECT 133.810 185.380 134.130 185.440 ;
        RECT 131.770 185.240 134.130 185.380 ;
        RECT 131.770 185.180 132.090 185.240 ;
        RECT 133.810 185.180 134.130 185.240 ;
        RECT 141.435 184.980 141.805 184.990 ;
        RECT 112.730 184.920 113.050 184.980 ;
        RECT 119.870 184.920 120.190 184.980 ;
        RECT 112.730 184.780 120.190 184.920 ;
        RECT 112.730 184.720 113.050 184.780 ;
        RECT 119.870 184.720 120.190 184.780 ;
        RECT 126.330 184.920 126.650 184.980 ;
        RECT 130.750 184.920 131.070 184.980 ;
        RECT 135.510 184.920 135.830 184.980 ;
        RECT 126.330 184.780 131.070 184.920 ;
        RECT 126.330 184.720 126.650 184.780 ;
        RECT 130.750 184.720 131.070 184.780 ;
        RECT 131.350 184.780 135.830 184.920 ;
        RECT 110.010 184.460 110.330 184.520 ;
        RECT 114.430 184.460 114.750 184.520 ;
        RECT 110.010 184.320 114.750 184.460 ;
        RECT 110.010 184.260 110.330 184.320 ;
        RECT 114.430 184.260 114.750 184.320 ;
        RECT 117.150 184.460 117.470 184.520 ;
        RECT 122.930 184.460 123.250 184.520 ;
        RECT 117.150 184.320 123.250 184.460 ;
        RECT 117.150 184.260 117.470 184.320 ;
        RECT 122.930 184.260 123.250 184.320 ;
        RECT 128.370 184.460 128.690 184.520 ;
        RECT 130.750 184.460 131.070 184.520 ;
        RECT 131.350 184.460 131.490 184.780 ;
        RECT 135.510 184.720 135.830 184.780 ;
        RECT 141.435 184.720 141.950 184.980 ;
        RECT 141.435 184.710 141.805 184.720 ;
        RECT 128.370 184.320 131.490 184.460 ;
        RECT 134.490 184.460 134.810 184.520 ;
        RECT 135.510 184.460 135.830 184.520 ;
        RECT 134.490 184.320 135.830 184.460 ;
        RECT 128.370 184.260 128.690 184.320 ;
        RECT 130.750 184.260 131.070 184.320 ;
        RECT 134.490 184.260 134.810 184.320 ;
        RECT 135.510 184.260 135.830 184.320 ;
        RECT 104.035 184.025 104.405 184.070 ;
        RECT 98.665 184.000 104.965 184.025 ;
        RECT 114.770 184.000 115.090 184.060 ;
        RECT 98.665 183.860 115.090 184.000 ;
        RECT 98.665 183.835 104.965 183.860 ;
        RECT 97.860 169.020 98.360 170.590 ;
        RECT 98.665 101.925 98.855 183.835 ;
        RECT 104.035 183.790 104.405 183.835 ;
        RECT 114.770 183.800 115.090 183.860 ;
        RECT 131.430 184.000 131.750 184.060 ;
        RECT 133.810 184.000 134.130 184.060 ;
        RECT 140.950 184.000 141.270 184.060 ;
        RECT 131.430 183.860 141.270 184.000 ;
        RECT 131.430 183.800 131.750 183.860 ;
        RECT 133.810 183.800 134.130 183.860 ;
        RECT 140.950 183.800 141.270 183.860 ;
        RECT 111.710 183.540 112.030 183.600 ;
        RECT 114.430 183.540 114.750 183.600 ;
        RECT 116.810 183.540 117.130 183.600 ;
        RECT 111.710 183.400 117.130 183.540 ;
        RECT 111.710 183.340 112.030 183.400 ;
        RECT 114.430 183.340 114.750 183.400 ;
        RECT 116.810 183.340 117.130 183.400 ;
        RECT 127.835 183.540 128.205 183.610 ;
        RECT 128.370 183.540 128.690 183.600 ;
        RECT 127.835 183.400 128.690 183.540 ;
        RECT 127.835 183.330 128.205 183.400 ;
        RECT 128.370 183.340 128.690 183.400 ;
        RECT 134.635 183.540 135.005 183.610 ;
        RECT 136.190 183.540 136.510 183.600 ;
        RECT 134.635 183.400 136.510 183.540 ;
        RECT 134.635 183.330 135.005 183.400 ;
        RECT 136.190 183.340 136.510 183.400 ;
        RECT 138.035 183.540 138.405 183.610 ;
        RECT 139.250 183.540 139.570 183.600 ;
        RECT 138.035 183.400 139.570 183.540 ;
        RECT 138.035 183.330 138.405 183.400 ;
        RECT 139.250 183.340 139.570 183.400 ;
        RECT 141.630 183.540 141.950 183.600 ;
        RECT 148.235 183.540 148.605 183.610 ;
        RECT 141.630 183.400 148.605 183.540 ;
        RECT 141.630 183.340 141.950 183.400 ;
        RECT 114.230 181.455 114.670 181.590 ;
        RECT 99.115 181.280 114.670 181.455 ;
        RECT 143.820 181.430 143.960 183.400 ;
        RECT 148.235 183.330 148.605 183.400 ;
        RECT 99.115 117.000 99.290 181.280 ;
        RECT 114.230 181.150 114.670 181.280 ;
        RECT 138.630 181.290 143.960 181.430 ;
        RECT 117.600 180.905 118.040 181.060 ;
        RECT 99.525 180.730 118.040 180.905 ;
        RECT 99.525 132.040 99.700 180.730 ;
        RECT 117.600 180.620 118.040 180.730 ;
        RECT 120.990 180.510 121.430 180.950 ;
        RECT 110.830 180.390 111.270 180.490 ;
        RECT 100.030 180.185 111.270 180.390 ;
        RECT 121.140 180.370 121.300 180.510 ;
        RECT 100.030 147.055 100.235 180.185 ;
        RECT 110.830 180.050 111.270 180.185 ;
        RECT 116.920 180.210 121.300 180.370 ;
        RECT 124.380 180.350 124.800 180.810 ;
        RECT 127.810 180.430 128.230 180.890 ;
        RECT 131.220 180.580 131.670 181.020 ;
        RECT 138.010 180.590 138.460 181.030 ;
        RECT 107.435 179.765 107.805 179.810 ;
        RECT 100.535 179.575 107.805 179.765 ;
        RECT 100.535 162.060 100.725 179.575 ;
        RECT 107.435 179.530 107.805 179.575 ;
        RECT 115.310 173.470 116.450 174.140 ;
        RECT 104.640 173.010 105.340 173.020 ;
        RECT 104.300 172.270 105.650 173.010 ;
        RECT 104.640 162.840 105.340 172.270 ;
        RECT 114.320 168.875 114.640 168.920 ;
        RECT 114.320 168.705 116.715 168.875 ;
        RECT 114.320 168.660 114.640 168.705 ;
        RECT 106.690 167.320 114.680 167.710 ;
        RECT 106.650 165.435 106.970 165.490 ;
        RECT 105.850 165.285 106.970 165.435 ;
        RECT 100.500 161.740 100.760 162.060 ;
        RECT 104.550 162.050 105.410 162.840 ;
        RECT 104.640 158.020 105.340 158.030 ;
        RECT 104.300 157.280 105.650 158.020 ;
        RECT 104.640 147.850 105.340 157.280 ;
        RECT 105.850 150.415 106.000 165.285 ;
        RECT 106.650 165.230 106.970 165.285 ;
        RECT 109.230 164.260 111.890 167.320 ;
        RECT 115.430 164.570 116.370 166.200 ;
        RECT 106.730 163.810 114.670 164.260 ;
        RECT 114.300 153.850 114.620 153.910 ;
        RECT 114.300 153.710 116.400 153.850 ;
        RECT 114.300 153.650 114.620 153.710 ;
        RECT 106.690 152.330 114.680 152.720 ;
        RECT 106.720 150.415 107.040 150.470 ;
        RECT 105.850 150.265 107.040 150.415 ;
        RECT 100.600 147.055 100.920 147.080 ;
        RECT 104.550 147.060 105.410 147.850 ;
        RECT 100.030 146.850 100.920 147.055 ;
        RECT 100.600 146.820 100.920 146.850 ;
        RECT 104.640 143.040 105.340 143.050 ;
        RECT 104.300 142.300 105.650 143.040 ;
        RECT 104.640 132.870 105.340 142.300 ;
        RECT 105.850 135.425 106.000 150.265 ;
        RECT 106.720 150.210 107.040 150.265 ;
        RECT 109.230 149.270 111.890 152.330 ;
        RECT 106.730 148.820 114.670 149.270 ;
        RECT 114.375 138.925 114.695 138.955 ;
        RECT 114.375 138.730 115.945 138.925 ;
        RECT 114.375 138.695 114.695 138.730 ;
        RECT 106.690 137.350 114.680 137.740 ;
        RECT 106.750 135.425 107.070 135.480 ;
        RECT 105.850 135.275 107.070 135.425 ;
        RECT 104.550 132.080 105.410 132.870 ;
        RECT 100.650 132.040 100.970 132.080 ;
        RECT 99.525 131.865 100.970 132.040 ;
        RECT 100.650 131.820 100.970 131.865 ;
        RECT 104.640 128.010 105.340 128.020 ;
        RECT 104.300 127.270 105.650 128.010 ;
        RECT 104.640 117.840 105.340 127.270 ;
        RECT 105.850 124.775 106.000 135.275 ;
        RECT 106.750 135.220 107.070 135.275 ;
        RECT 109.230 134.290 111.890 137.350 ;
        RECT 106.730 133.840 114.670 134.290 ;
        RECT 105.850 124.625 107.775 124.775 ;
        RECT 106.510 123.970 106.830 124.000 ;
        RECT 105.790 123.770 106.830 123.970 ;
        RECT 104.550 117.050 105.410 117.840 ;
        RECT 100.570 117.000 100.890 117.040 ;
        RECT 99.115 116.825 100.890 117.000 ;
        RECT 100.570 116.780 100.890 116.825 ;
        RECT 104.640 113.020 105.340 113.030 ;
        RECT 104.300 112.280 105.650 113.020 ;
        RECT 104.640 102.850 105.340 112.280 ;
        RECT 105.790 109.350 105.990 123.770 ;
        RECT 106.510 123.740 106.830 123.770 ;
        RECT 107.625 123.375 107.775 124.625 ;
        RECT 106.285 123.225 107.775 123.375 ;
        RECT 106.285 120.455 106.435 123.225 ;
        RECT 106.690 122.320 114.680 122.710 ;
        RECT 106.680 120.455 107.000 120.510 ;
        RECT 106.285 120.305 107.000 120.455 ;
        RECT 106.310 120.250 107.000 120.305 ;
        RECT 106.310 120.170 106.900 120.250 ;
        RECT 106.310 114.000 106.570 120.170 ;
        RECT 109.230 119.260 111.890 122.320 ;
        RECT 106.730 118.810 114.670 119.260 ;
        RECT 106.335 113.850 106.545 114.000 ;
        RECT 114.790 113.850 115.070 113.885 ;
        RECT 106.335 113.550 115.080 113.850 ;
        RECT 106.335 110.525 106.545 113.550 ;
        RECT 114.790 113.515 115.070 113.550 ;
        RECT 106.335 110.315 108.075 110.525 ;
        RECT 105.790 109.150 107.580 109.350 ;
        RECT 106.810 108.980 107.130 109.005 ;
        RECT 105.575 108.775 107.130 108.980 ;
        RECT 100.290 101.925 100.750 102.360 ;
        RECT 104.550 102.060 105.410 102.850 ;
        RECT 98.665 101.735 100.750 101.925 ;
        RECT 100.290 101.300 100.750 101.735 ;
        RECT 105.575 101.230 105.780 108.775 ;
        RECT 106.810 108.745 107.130 108.775 ;
        RECT 107.380 108.510 107.580 109.150 ;
        RECT 103.700 101.025 105.780 101.230 ;
        RECT 105.970 108.310 107.580 108.510 ;
        RECT 103.700 96.850 103.905 101.025 ;
        RECT 105.970 100.740 106.170 108.310 ;
        RECT 107.865 108.130 108.075 110.315 ;
        RECT 106.400 108.015 108.075 108.130 ;
        RECT 106.400 107.990 108.040 108.015 ;
        RECT 106.400 105.340 106.540 107.990 ;
        RECT 106.690 107.330 114.680 107.720 ;
        RECT 106.790 105.340 107.110 105.400 ;
        RECT 106.400 105.200 107.110 105.340 ;
        RECT 106.790 105.140 107.110 105.200 ;
        RECT 109.230 104.270 111.890 107.330 ;
        RECT 106.730 103.820 114.670 104.270 ;
        RECT 115.750 101.055 115.945 138.730 ;
        RECT 105.080 100.540 106.170 100.740 ;
        RECT 108.385 100.860 115.945 101.055 ;
        RECT 105.080 97.530 105.280 100.540 ;
        RECT 104.960 96.970 105.410 97.530 ;
        RECT 108.385 97.520 108.580 100.860 ;
        RECT 116.260 100.460 116.400 153.710 ;
        RECT 111.270 100.320 116.400 100.460 ;
        RECT 108.260 96.960 108.710 97.520 ;
        RECT 111.270 97.470 111.410 100.320 ;
        RECT 116.545 100.015 116.715 168.705 ;
        RECT 116.920 102.160 117.080 180.210 ;
        RECT 124.545 180.000 124.700 180.350 ;
        RECT 117.345 179.845 124.700 180.000 ;
        RECT 117.345 117.030 117.500 179.845 ;
        RECT 127.915 179.590 128.100 180.430 ;
        RECT 117.690 179.405 128.100 179.590 ;
        RECT 117.690 132.205 117.875 179.405 ;
        RECT 131.345 179.160 131.500 180.580 ;
        RECT 118.115 179.005 131.500 179.160 ;
        RECT 118.115 147.100 118.270 179.005 ;
        RECT 138.130 178.750 138.310 180.590 ;
        RECT 118.450 178.570 138.310 178.750 ;
        RECT 118.450 162.120 118.630 178.570 ;
        RECT 138.630 178.340 138.770 181.290 ;
        RECT 141.400 180.835 141.850 180.960 ;
        RECT 144.790 180.875 145.240 181.020 ;
        RECT 136.520 178.200 138.770 178.340 ;
        RECT 138.985 180.640 141.850 180.835 ;
        RECT 123.680 173.040 124.380 173.050 ;
        RECT 123.340 172.300 124.690 173.040 ;
        RECT 123.680 162.870 124.380 172.300 ;
        RECT 135.590 169.180 136.250 170.640 ;
        RECT 133.285 168.925 133.605 168.955 ;
        RECT 133.285 168.730 136.275 168.925 ;
        RECT 133.285 168.695 133.605 168.730 ;
        RECT 125.730 167.350 133.720 167.740 ;
        RECT 125.700 165.485 126.020 165.540 ;
        RECT 124.760 165.335 126.020 165.485 ;
        RECT 119.630 162.120 119.950 162.160 ;
        RECT 118.450 161.940 119.950 162.120 ;
        RECT 123.590 162.080 124.450 162.870 ;
        RECT 119.630 161.900 119.950 161.940 ;
        RECT 124.760 159.685 124.910 165.335 ;
        RECT 125.700 165.280 126.020 165.335 ;
        RECT 128.270 164.290 130.930 167.350 ;
        RECT 134.600 166.100 135.380 166.120 ;
        RECT 134.550 166.020 135.380 166.100 ;
        RECT 134.510 164.600 135.380 166.020 ;
        RECT 134.510 164.540 135.290 164.600 ;
        RECT 125.770 163.840 133.710 164.290 ;
        RECT 124.760 159.370 125.015 159.685 ;
        RECT 123.680 158.020 124.380 158.030 ;
        RECT 123.340 157.280 124.690 158.020 ;
        RECT 123.680 147.850 124.380 157.280 ;
        RECT 124.865 150.395 125.015 159.370 ;
        RECT 133.460 153.905 133.780 153.960 ;
        RECT 133.460 153.755 135.875 153.905 ;
        RECT 133.460 153.700 133.780 153.755 ;
        RECT 125.730 152.330 133.720 152.720 ;
        RECT 125.690 150.395 126.010 150.450 ;
        RECT 124.865 150.245 126.010 150.395 ;
        RECT 119.580 147.100 119.900 147.150 ;
        RECT 118.115 146.945 119.900 147.100 ;
        RECT 123.590 147.060 124.450 147.850 ;
        RECT 119.580 146.890 119.900 146.945 ;
        RECT 123.630 143.000 124.330 143.010 ;
        RECT 123.290 142.260 124.640 143.000 ;
        RECT 123.630 132.830 124.330 142.260 ;
        RECT 124.865 135.405 125.015 150.245 ;
        RECT 125.690 150.190 126.010 150.245 ;
        RECT 128.270 149.270 130.930 152.330 ;
        RECT 125.770 148.820 133.710 149.270 ;
        RECT 133.340 138.875 133.660 138.930 ;
        RECT 133.340 138.725 135.515 138.875 ;
        RECT 133.340 138.670 133.660 138.725 ;
        RECT 125.680 137.310 133.670 137.700 ;
        RECT 125.620 135.405 125.940 135.460 ;
        RECT 124.865 135.255 125.940 135.405 ;
        RECT 117.690 132.190 119.740 132.205 ;
        RECT 117.690 132.020 119.820 132.190 ;
        RECT 123.540 132.040 124.400 132.830 ;
        RECT 117.710 131.990 119.820 132.020 ;
        RECT 119.500 131.930 119.820 131.990 ;
        RECT 123.630 127.980 124.330 127.990 ;
        RECT 123.290 127.240 124.640 127.980 ;
        RECT 123.630 117.810 124.330 127.240 ;
        RECT 124.865 120.395 125.015 135.255 ;
        RECT 125.620 135.200 125.940 135.255 ;
        RECT 128.220 134.250 130.880 137.310 ;
        RECT 125.720 133.800 133.660 134.250 ;
        RECT 133.225 123.930 133.545 123.965 ;
        RECT 133.225 123.745 135.180 123.930 ;
        RECT 133.225 123.705 133.545 123.745 ;
        RECT 125.680 122.290 133.670 122.680 ;
        RECT 125.710 120.395 126.030 120.450 ;
        RECT 124.865 120.245 126.030 120.395 ;
        RECT 119.490 117.030 119.810 117.080 ;
        RECT 117.345 116.875 119.810 117.030 ;
        RECT 123.540 117.020 124.400 117.810 ;
        RECT 119.490 116.820 119.810 116.875 ;
        RECT 124.865 113.850 125.015 120.245 ;
        RECT 125.710 120.190 126.030 120.245 ;
        RECT 128.220 119.230 130.880 122.290 ;
        RECT 125.720 118.780 133.660 119.230 ;
        RECT 133.510 113.850 133.790 113.885 ;
        RECT 117.525 113.550 133.800 113.850 ;
        RECT 123.630 113.000 124.330 113.010 ;
        RECT 123.290 112.260 124.640 113.000 ;
        RECT 123.630 102.830 124.330 112.260 ;
        RECT 124.865 105.395 125.015 113.550 ;
        RECT 133.510 113.515 133.790 113.550 ;
        RECT 133.425 108.850 133.745 108.895 ;
        RECT 133.425 108.685 134.750 108.850 ;
        RECT 133.425 108.635 133.745 108.685 ;
        RECT 125.680 107.310 133.670 107.700 ;
        RECT 125.670 105.395 125.990 105.450 ;
        RECT 124.865 105.245 125.990 105.395 ;
        RECT 125.670 105.190 125.990 105.245 ;
        RECT 128.220 104.250 130.880 107.310 ;
        RECT 125.720 103.800 133.660 104.250 ;
        RECT 119.580 102.160 119.900 102.210 ;
        RECT 116.920 102.000 119.900 102.160 ;
        RECT 123.540 102.040 124.400 102.830 ;
        RECT 119.580 101.950 119.900 102.000 ;
        RECT 134.585 101.060 134.750 108.685 ;
        RECT 114.415 99.845 116.715 100.015 ;
        RECT 117.300 100.895 134.750 101.060 ;
        RECT 114.415 97.520 114.585 99.845 ;
        RECT 111.090 96.910 111.540 97.470 ;
        RECT 114.280 96.960 114.730 97.520 ;
        RECT 117.300 97.430 117.465 100.895 ;
        RECT 134.995 100.590 135.180 123.745 ;
        RECT 120.140 100.405 135.180 100.590 ;
        RECT 120.140 97.450 120.325 100.405 ;
        RECT 135.365 100.155 135.515 138.725 ;
        RECT 123.015 100.005 135.515 100.155 ;
        RECT 123.015 97.450 123.165 100.005 ;
        RECT 135.725 99.745 135.875 153.755 ;
        RECT 126.435 99.595 135.875 99.745 ;
        RECT 126.435 97.500 126.585 99.595 ;
        RECT 136.080 99.385 136.275 168.730 ;
        RECT 136.520 102.020 136.660 178.200 ;
        RECT 138.985 177.980 139.180 180.640 ;
        RECT 141.400 180.520 141.850 180.640 ;
        RECT 142.235 180.700 145.240 180.875 ;
        RECT 142.235 180.210 142.410 180.700 ;
        RECT 144.790 180.580 145.240 180.700 ;
        RECT 136.820 177.820 139.180 177.980 ;
        RECT 136.820 117.030 136.980 177.820 ;
        RECT 138.985 177.805 139.180 177.820 ;
        RECT 139.425 180.035 142.410 180.210 ;
        RECT 139.425 177.590 139.600 180.035 ;
        RECT 143.785 179.960 144.155 180.240 ;
        RECT 143.870 179.765 144.075 179.960 ;
        RECT 137.220 177.215 137.500 177.585 ;
        RECT 137.725 177.415 139.600 177.590 ;
        RECT 139.850 179.560 144.075 179.765 ;
        RECT 137.270 132.080 137.450 177.215 ;
        RECT 137.725 147.010 137.900 177.415 ;
        RECT 139.850 177.215 140.055 179.560 ;
        RECT 138.050 177.010 140.055 177.215 ;
        RECT 138.050 162.185 138.255 177.010 ;
        RECT 142.630 173.080 143.330 173.090 ;
        RECT 142.290 172.340 143.640 173.080 ;
        RECT 142.630 162.910 143.330 172.340 ;
        RECT 152.310 168.945 152.630 168.980 ;
        RECT 152.310 168.755 154.195 168.945 ;
        RECT 152.310 168.720 152.630 168.755 ;
        RECT 144.680 167.390 152.670 167.780 ;
        RECT 144.660 165.485 144.980 165.540 ;
        RECT 143.770 165.335 144.980 165.485 ;
        RECT 138.510 162.185 138.830 162.210 ;
        RECT 138.050 161.980 138.830 162.185 ;
        RECT 142.540 162.120 143.400 162.910 ;
        RECT 138.510 161.950 138.830 161.980 ;
        RECT 143.770 159.345 143.920 165.335 ;
        RECT 144.660 165.280 144.980 165.335 ;
        RECT 147.220 164.330 149.880 167.390 ;
        RECT 144.720 163.880 152.660 164.330 ;
        RECT 143.770 159.090 144.025 159.345 ;
        RECT 142.680 158.020 143.380 158.030 ;
        RECT 142.340 157.280 143.690 158.020 ;
        RECT 142.680 147.850 143.380 157.280 ;
        RECT 143.875 150.275 144.025 159.090 ;
        RECT 152.180 158.420 153.540 159.710 ;
        RECT 152.345 153.840 152.665 153.865 ;
        RECT 152.345 153.635 153.695 153.840 ;
        RECT 152.345 153.605 152.665 153.635 ;
        RECT 144.730 152.330 152.720 152.720 ;
        RECT 144.690 150.275 145.010 150.330 ;
        RECT 143.875 150.125 145.010 150.275 ;
        RECT 142.590 147.060 143.450 147.850 ;
        RECT 138.640 147.010 138.960 147.050 ;
        RECT 137.725 146.835 138.960 147.010 ;
        RECT 138.640 146.790 138.960 146.835 ;
        RECT 142.630 143.000 143.330 143.010 ;
        RECT 142.290 142.260 143.640 143.000 ;
        RECT 142.630 132.830 143.330 142.260 ;
        RECT 143.875 135.335 144.025 150.125 ;
        RECT 144.690 150.070 145.010 150.125 ;
        RECT 147.270 149.270 149.930 152.330 ;
        RECT 144.770 148.820 152.710 149.270 ;
        RECT 153.490 139.590 153.695 153.635 ;
        RECT 154.005 140.155 154.195 168.755 ;
        RECT 154.005 139.965 154.715 140.155 ;
        RECT 153.490 139.385 154.380 139.590 ;
        RECT 152.340 138.865 152.660 138.920 ;
        RECT 152.340 138.715 153.935 138.865 ;
        RECT 152.340 138.660 152.660 138.715 ;
        RECT 144.680 137.310 152.670 137.700 ;
        RECT 144.660 135.335 144.980 135.390 ;
        RECT 143.875 135.185 144.980 135.335 ;
        RECT 138.630 132.080 138.950 132.120 ;
        RECT 137.270 131.900 138.950 132.080 ;
        RECT 142.540 132.040 143.400 132.830 ;
        RECT 138.630 131.860 138.950 131.900 ;
        RECT 142.630 127.980 143.330 127.990 ;
        RECT 142.290 127.240 143.640 127.980 ;
        RECT 142.630 117.810 143.330 127.240 ;
        RECT 143.875 120.335 144.025 135.185 ;
        RECT 144.660 135.130 144.980 135.185 ;
        RECT 147.220 134.250 149.880 137.310 ;
        RECT 144.720 133.800 152.660 134.250 ;
        RECT 152.355 123.840 152.675 123.865 ;
        RECT 152.355 123.635 153.560 123.840 ;
        RECT 152.355 123.605 152.675 123.635 ;
        RECT 144.680 122.290 152.670 122.680 ;
        RECT 144.620 120.335 144.940 120.390 ;
        RECT 143.875 120.185 144.940 120.335 ;
        RECT 138.620 117.030 138.940 117.080 ;
        RECT 136.820 116.870 138.940 117.030 ;
        RECT 142.540 117.020 143.400 117.810 ;
        RECT 138.620 116.820 138.940 116.870 ;
        RECT 143.875 114.410 144.025 120.185 ;
        RECT 144.620 120.130 144.940 120.185 ;
        RECT 147.220 119.230 149.880 122.290 ;
        RECT 144.720 118.780 152.660 119.230 ;
        RECT 143.070 114.360 144.380 114.410 ;
        RECT 143.060 113.915 144.380 114.360 ;
        RECT 136.965 113.775 137.355 113.850 ;
        RECT 143.070 113.775 144.380 113.915 ;
        RECT 136.965 113.625 144.380 113.775 ;
        RECT 136.965 113.550 137.355 113.625 ;
        RECT 143.070 113.550 144.380 113.625 ;
        RECT 142.680 113.000 143.380 113.010 ;
        RECT 142.340 112.260 143.690 113.000 ;
        RECT 142.680 102.830 143.380 112.260 ;
        RECT 143.875 110.035 144.025 113.550 ;
        RECT 143.875 109.885 145.475 110.035 ;
        RECT 144.790 108.930 145.110 108.990 ;
        RECT 143.760 108.790 145.110 108.930 ;
        RECT 138.660 102.020 138.980 102.080 ;
        RECT 142.590 102.040 143.450 102.830 ;
        RECT 136.520 101.880 138.980 102.020 ;
        RECT 138.660 101.820 138.980 101.880 ;
        RECT 143.760 100.630 143.900 108.790 ;
        RECT 144.790 108.730 145.110 108.790 ;
        RECT 145.325 108.315 145.475 109.885 ;
        RECT 144.215 108.165 145.475 108.315 ;
        RECT 144.215 105.405 144.365 108.165 ;
        RECT 144.730 107.310 152.720 107.700 ;
        RECT 144.710 105.405 145.030 105.460 ;
        RECT 144.215 105.255 145.030 105.405 ;
        RECT 144.710 105.200 145.030 105.255 ;
        RECT 147.270 104.250 149.930 107.310 ;
        RECT 144.770 103.800 152.710 104.250 ;
        RECT 129.205 99.190 136.275 99.385 ;
        RECT 136.700 100.490 143.900 100.630 ;
        RECT 117.130 96.960 117.630 97.430 ;
        RECT 120.140 97.300 120.650 97.450 ;
        RECT 120.150 96.980 120.650 97.300 ;
        RECT 122.840 96.980 123.340 97.450 ;
        RECT 126.280 97.030 126.780 97.500 ;
        RECT 129.205 97.480 129.400 99.190 ;
        RECT 136.700 98.970 136.840 100.490 ;
        RECT 153.355 100.040 153.560 123.635 ;
        RECT 132.390 98.830 136.840 98.970 ;
        RECT 137.175 99.835 153.560 100.040 ;
        RECT 129.090 97.010 129.590 97.480 ;
        RECT 132.390 97.440 132.530 98.830 ;
        RECT 137.175 98.500 137.380 99.835 ;
        RECT 153.785 99.545 153.935 138.715 ;
        RECT 134.960 98.295 137.380 98.500 ;
        RECT 138.445 99.395 153.935 99.545 ;
        RECT 132.200 96.970 132.700 97.440 ;
        RECT 134.960 97.430 135.165 98.295 ;
        RECT 134.820 96.960 135.320 97.430 ;
        RECT 138.445 97.400 138.595 99.395 ;
        RECT 154.175 99.160 154.380 139.385 ;
        RECT 141.775 98.955 154.380 99.160 ;
        RECT 141.775 97.810 141.980 98.955 ;
        RECT 154.525 98.755 154.715 139.965 ;
        RECT 148.025 98.565 154.715 98.755 ;
        RECT 148.025 97.820 148.215 98.565 ;
        RECT 141.775 97.475 142.290 97.810 ;
        RECT 117.300 96.940 117.465 96.960 ;
        RECT 138.300 96.930 138.800 97.400 ;
        RECT 141.790 97.340 142.290 97.475 ;
        RECT 147.910 97.350 148.410 97.820 ;
        RECT 103.580 96.380 104.000 96.850 ;
      LAYER met3 ;
        RECT 63.700 224.950 64.020 225.330 ;
        RECT 66.510 224.950 66.830 225.330 ;
        RECT 63.710 216.655 64.010 224.950 ;
        RECT 66.520 217.195 66.820 224.950 ;
        RECT 69.280 224.940 69.600 225.320 ;
        RECT 72.050 224.990 72.370 225.370 ;
        RECT 69.290 221.685 69.590 224.940 ;
        RECT 69.265 221.335 69.615 221.685 ;
        RECT 72.060 221.215 72.360 224.990 ;
        RECT 74.815 224.980 75.135 225.360 ;
        RECT 72.035 220.865 72.385 221.215 ;
        RECT 74.825 220.620 75.125 224.980 ;
        RECT 77.590 224.860 77.910 225.240 ;
        RECT 80.305 224.960 80.625 225.340 ;
        RECT 74.800 220.270 75.150 220.620 ;
        RECT 77.600 217.595 77.900 224.860 ;
        RECT 80.315 220.050 80.615 224.960 ;
        RECT 83.070 224.860 83.390 225.240 ;
        RECT 85.810 225.000 86.130 225.380 ;
        RECT 80.290 219.700 80.640 220.050 ;
        RECT 83.080 219.655 83.380 224.860 ;
        RECT 83.055 219.305 83.405 219.655 ;
        RECT 85.820 219.215 86.120 225.000 ;
        RECT 88.610 224.950 88.930 225.330 ;
        RECT 91.390 225.060 91.710 225.440 ;
        RECT 85.795 218.865 86.145 219.215 ;
        RECT 88.620 217.965 88.920 224.950 ;
        RECT 91.400 218.745 91.700 225.060 ;
        RECT 94.080 225.030 94.400 225.410 ;
        RECT 143.700 225.340 144.080 225.350 ;
        RECT 138.070 225.040 144.080 225.340 ;
        RECT 91.375 218.395 91.725 218.745 ;
        RECT 94.090 218.295 94.390 225.030 ;
        RECT 138.070 223.260 138.370 225.040 ;
        RECT 143.700 225.030 144.080 225.040 ;
        RECT 110.720 219.270 111.320 223.260 ;
        RECT 110.720 219.260 111.850 219.270 ;
        RECT 120.920 219.260 121.520 223.260 ;
        RECT 127.720 219.260 128.320 223.260 ;
        RECT 134.520 219.260 135.120 223.260 ;
        RECT 137.920 219.260 138.520 223.260 ;
        RECT 110.870 219.055 111.850 219.260 ;
        RECT 110.870 218.970 111.865 219.055 ;
        RECT 111.535 218.725 111.865 218.970 ;
        RECT 88.595 217.615 88.945 217.965 ;
        RECT 94.065 217.945 94.415 218.295 ;
        RECT 77.575 217.245 77.925 217.595 ;
        RECT 66.495 216.845 66.845 217.195 ;
        RECT 121.070 216.755 121.370 219.260 ;
        RECT 127.870 218.820 128.170 219.260 ;
        RECT 127.830 218.440 128.220 218.820 ;
        RECT 127.870 216.755 128.170 218.440 ;
        RECT 134.670 216.755 134.970 219.260 ;
        RECT 63.685 216.305 64.035 216.655 ;
        RECT 121.055 216.425 121.385 216.755 ;
        RECT 127.855 216.425 128.185 216.755 ;
        RECT 134.655 216.425 134.985 216.755 ;
        RECT 138.070 205.715 138.370 219.260 ;
        RECT 139.415 206.765 139.745 207.095 ;
        RECT 138.055 205.385 138.385 205.715 ;
        RECT 139.430 202.955 139.730 206.765 ;
        RECT 139.415 202.625 139.745 202.955 ;
        RECT 7.305 202.220 8.895 202.245 ;
        RECT 1.140 200.620 8.900 202.220 ;
        RECT 110.515 200.630 110.845 202.210 ;
        RECT 115.955 200.630 116.285 202.210 ;
        RECT 121.395 200.630 121.725 202.210 ;
        RECT 126.835 200.630 127.165 202.210 ;
        RECT 132.275 200.630 132.605 202.210 ;
        RECT 137.715 200.630 138.045 202.210 ;
        RECT 7.305 200.595 8.895 200.620 ;
        RECT 107.795 197.330 108.125 198.910 ;
        RECT 113.235 197.330 113.565 198.910 ;
        RECT 118.675 197.330 119.005 198.910 ;
        RECT 124.115 197.330 124.445 198.910 ;
        RECT 129.555 197.330 129.885 198.910 ;
        RECT 134.995 197.330 135.325 198.910 ;
        RECT 110.855 192.045 111.185 192.375 ;
        RECT 107.455 187.445 107.785 187.775 ;
        RECT 104.055 183.765 104.385 184.095 ;
        RECT 104.070 180.215 104.370 183.765 ;
        RECT 107.470 180.215 107.770 187.445 ;
        RECT 110.870 180.490 111.170 192.045 ;
        RECT 121.055 190.665 121.385 190.995 ;
        RECT 114.255 189.285 114.585 189.615 ;
        RECT 114.270 181.590 114.570 189.285 ;
        RECT 117.655 186.985 117.985 187.315 ;
        RECT 114.230 181.150 114.670 181.590 ;
        RECT 110.830 180.215 111.270 180.490 ;
        RECT 114.270 180.215 114.570 181.150 ;
        RECT 117.670 181.060 117.970 186.985 ;
        RECT 117.600 180.620 118.040 181.060 ;
        RECT 121.070 180.950 121.370 190.665 ;
        RECT 139.430 189.615 139.730 202.625 ;
        RECT 143.155 200.630 143.485 202.210 ;
        RECT 140.435 197.330 140.765 198.910 ;
        RECT 143.795 193.875 144.145 194.225 ;
        RECT 139.415 189.285 139.745 189.615 ;
        RECT 124.455 188.365 124.785 188.695 ;
        RECT 117.670 180.215 117.970 180.620 ;
        RECT 120.990 180.610 121.430 180.950 ;
        RECT 124.470 180.810 124.770 188.365 ;
        RECT 131.255 185.605 131.585 185.935 ;
        RECT 127.855 183.305 128.185 183.635 ;
        RECT 127.870 180.890 128.170 183.305 ;
        RECT 131.270 181.020 131.570 185.605 ;
        RECT 141.455 184.685 141.785 185.015 ;
        RECT 134.655 183.305 134.985 183.635 ;
        RECT 138.055 183.305 138.385 183.635 ;
        RECT 120.920 180.215 121.480 180.610 ;
        RECT 124.380 180.470 124.800 180.810 ;
        RECT 127.810 180.570 128.260 180.890 ;
        RECT 131.220 180.580 131.670 181.020 ;
        RECT 124.330 180.215 124.870 180.470 ;
        RECT 127.760 180.215 128.320 180.570 ;
        RECT 131.270 180.215 131.570 180.580 ;
        RECT 134.670 180.215 134.970 183.305 ;
        RECT 138.070 181.030 138.370 183.305 ;
        RECT 138.010 180.590 138.460 181.030 ;
        RECT 141.470 180.960 141.770 184.685 ;
        RECT 138.070 180.215 138.370 180.590 ;
        RECT 141.400 180.520 141.850 180.960 ;
        RECT 141.470 180.215 141.770 180.520 ;
        RECT 143.820 180.265 144.120 193.875 ;
        RECT 144.855 186.065 145.185 186.395 ;
        RECT 144.870 181.020 145.170 186.065 ;
        RECT 148.255 183.305 148.585 183.635 ;
        RECT 144.790 180.580 145.240 181.020 ;
        RECT 103.920 176.215 104.520 180.215 ;
        RECT 107.320 176.215 107.920 180.215 ;
        RECT 110.720 176.215 111.320 180.215 ;
        RECT 114.120 176.215 114.720 180.215 ;
        RECT 117.520 176.215 118.120 180.215 ;
        RECT 120.920 176.215 121.520 180.215 ;
        RECT 124.320 176.215 124.920 180.215 ;
        RECT 127.720 176.215 128.320 180.215 ;
        RECT 131.120 176.215 131.720 180.215 ;
        RECT 134.520 177.550 135.120 180.215 ;
        RECT 137.195 177.550 137.525 177.565 ;
        RECT 134.520 177.250 137.525 177.550 ;
        RECT 134.520 176.215 135.120 177.250 ;
        RECT 137.195 177.235 137.525 177.250 ;
        RECT 137.920 176.215 138.520 180.215 ;
        RECT 141.320 176.215 141.920 180.215 ;
        RECT 143.805 179.935 144.135 180.265 ;
        RECT 144.870 180.215 145.170 180.580 ;
        RECT 148.270 180.215 148.570 183.305 ;
        RECT 144.720 176.215 145.320 180.215 ;
        RECT 148.120 176.215 148.720 180.215 ;
        RECT 115.310 173.470 117.670 174.130 ;
        RECT 116.700 170.620 117.670 173.470 ;
        RECT 97.860 169.020 136.610 170.620 ;
        RECT 115.360 164.530 154.350 166.130 ;
        RECT 152.140 158.470 153.730 164.530 ;
        RECT 114.765 113.850 115.095 113.865 ;
        RECT 117.545 113.850 117.895 113.875 ;
        RECT 114.765 113.550 117.895 113.850 ;
        RECT 114.765 113.535 115.095 113.550 ;
        RECT 117.545 113.525 117.895 113.550 ;
        RECT 133.485 113.850 133.815 113.865 ;
        RECT 136.985 113.850 137.335 113.875 ;
        RECT 133.485 113.550 137.335 113.850 ;
        RECT 143.070 113.550 144.380 114.410 ;
        RECT 133.485 113.535 133.815 113.550 ;
        RECT 136.985 113.525 137.335 113.550 ;
      LAYER met4 ;
        RECT 42.010 224.930 44.470 225.470 ;
        RECT 44.770 224.930 47.230 225.470 ;
        RECT 47.530 224.930 49.990 225.470 ;
        RECT 63.695 224.975 63.790 225.305 ;
        RECT 66.505 224.975 66.550 225.305 ;
        RECT 69.275 224.965 69.310 225.295 ;
        RECT 72.045 225.015 72.070 225.345 ;
        RECT 72.370 225.015 72.375 225.345 ;
        RECT 74.810 225.005 74.830 225.335 ;
        RECT 75.130 225.005 75.140 225.335 ;
        RECT 42.945 224.145 43.395 224.930 ;
        RECT 77.585 224.885 77.590 225.215 ;
        RECT 77.890 224.885 77.915 225.215 ;
        RECT 80.300 224.985 80.350 225.315 ;
        RECT 83.065 224.885 83.110 225.215 ;
        RECT 85.805 225.025 85.870 225.355 ;
        RECT 88.605 224.975 88.630 225.305 ;
        RECT 88.930 224.975 88.935 225.305 ;
        RECT 91.385 225.085 91.390 225.415 ;
        RECT 91.690 225.085 91.715 225.415 ;
        RECT 94.075 225.055 94.150 225.385 ;
        RECT 143.725 225.025 143.830 225.355 ;
        RECT 1.945 223.695 43.395 224.145 ;
        RECT 1.945 220.760 2.395 223.695 ;
        RECT 7.300 200.620 146.450 202.220 ;
        RECT 6.000 198.920 134.860 198.930 ;
        RECT 6.000 197.330 143.560 198.920 ;
        RECT 107.720 197.320 143.560 197.330 ;
        RECT 133.260 168.930 134.860 197.320 ;
        RECT 144.850 164.530 146.450 200.620 ;
        RECT 143.750 113.915 152.485 114.360 ;
        RECT 152.040 1.000 152.485 113.915 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

