magic
tech sky130A
magscale 1 2
timestamp 1730796449
<< metal1 >>
rect 29076 44240 29082 44292
rect 29134 44240 29140 44292
rect 28996 44110 29048 44116
rect 28996 44052 29048 44058
rect 28872 43842 28924 43848
rect 28872 43784 28924 43790
rect 28770 43650 28822 43656
rect 28770 43592 28822 43598
rect 21092 41162 21144 41168
rect 21092 41104 21144 41110
rect 21104 38202 21132 41104
rect 21230 40984 21236 41036
rect 21288 41024 21294 41036
rect 21288 40984 21308 41024
rect 21280 39406 21308 40984
rect 21352 40868 21404 40874
rect 21352 40812 21404 40816
rect 21352 40810 21426 40812
rect 21364 40784 21426 40810
rect 21398 40216 21426 40784
rect 28781 40341 28811 43592
rect 21380 40164 21386 40216
rect 21438 40164 21444 40216
rect 28782 39952 28810 40341
rect 28762 39940 28832 39952
rect 28762 39888 28770 39940
rect 28822 39888 28832 39940
rect 28762 39874 28832 39888
rect 28884 39480 28912 43784
rect 28866 39428 28872 39480
rect 28924 39428 28930 39480
rect 21260 39388 21340 39406
rect 21260 39336 21268 39388
rect 21320 39336 21340 39388
rect 21260 39328 21340 39336
rect 21078 38192 21158 38202
rect 29008 38200 29036 44052
rect 29094 40774 29122 44240
rect 29076 40768 29140 40774
rect 29076 40716 29082 40768
rect 29134 40716 29140 40768
rect 29076 40710 29140 40716
rect 21078 38140 21092 38192
rect 21144 38140 21158 38192
rect 21078 38124 21158 38140
rect 28988 38192 29054 38200
rect 28988 38140 28996 38192
rect 29048 38140 29054 38192
rect 28988 38132 29054 38140
rect 23062 34814 23544 34828
rect 23062 34718 23078 34814
rect 23256 34718 23544 34814
rect 23062 34696 23544 34718
rect 23374 34470 23544 34696
rect 27118 34116 27250 34128
rect 19658 33834 19698 34098
rect 27118 33852 27140 34116
rect 27236 33852 27250 34116
rect 27118 33836 27250 33852
rect 30708 32924 30832 33186
rect 30436 31888 30708 31942
rect 30436 31722 30470 31888
rect 30640 31722 30708 31888
rect 30436 31684 30708 31722
rect 22349 21794 22444 21800
rect 22205 21699 22349 21794
rect 22349 21693 22444 21699
rect 19348 20166 19409 20167
rect 19330 20106 19630 20166
rect 19348 2249 19409 20106
rect 21234 20052 21426 20112
rect 21228 19860 21234 20052
rect 21321 19860 21426 20052
rect 7074 2188 19409 2249
rect 7074 598 7135 2188
rect 7042 571 7184 598
rect 7042 510 7074 571
rect 7135 510 7184 571
rect 7042 484 7184 510
<< via1 >>
rect 29082 44240 29134 44292
rect 28996 44058 29048 44110
rect 28872 43790 28924 43842
rect 28770 43598 28822 43650
rect 21092 41110 21144 41162
rect 21236 40984 21288 41036
rect 21352 40816 21404 40868
rect 21386 40164 21438 40216
rect 28770 39888 28822 39940
rect 28872 39428 28924 39480
rect 21268 39336 21320 39388
rect 29082 40716 29134 40768
rect 21092 38140 21144 38192
rect 28996 38140 29048 38192
rect 23078 34718 23256 34814
rect 19586 33820 19658 34104
rect 27140 33852 27236 34116
rect 23106 32924 23262 33226
rect 26926 32928 27048 33192
rect 30470 31722 30640 31888
rect 22349 21699 22444 21794
rect 22739 20992 22844 21097
rect 21234 19860 21321 20052
rect 7074 510 7135 571
<< metal2 >>
rect 13849 44272 13858 44332
rect 13918 44316 13927 44332
rect 13918 44288 14608 44316
rect 13918 44272 13927 44288
rect 14580 44280 14608 44288
rect 29082 44292 29134 44298
rect 14580 44252 29082 44280
rect 14403 44178 14412 44238
rect 14472 44222 14481 44238
rect 29082 44234 29134 44240
rect 14472 44194 24484 44222
rect 14472 44178 14481 44194
rect 14965 44119 15025 44128
rect 24207 44108 24216 44116
rect 15025 44069 24216 44108
rect 24207 44060 24216 44069
rect 24272 44060 24281 44116
rect 24456 44098 24484 44194
rect 28990 44098 28996 44110
rect 24456 44070 28996 44098
rect 14965 44050 15025 44059
rect 28990 44058 28996 44070
rect 29048 44058 29054 44110
rect 16063 44005 16123 44014
rect 26927 43995 26936 44002
rect 26256 43991 26936 43995
rect 16123 43958 26936 43991
rect 26256 43954 26936 43958
rect 26927 43946 26936 43954
rect 26992 43946 27001 44002
rect 16063 43936 16123 43945
rect 16607 43866 16616 43926
rect 16676 43910 16685 43926
rect 16676 43882 19248 43910
rect 16676 43866 16685 43882
rect 19220 43854 22528 43882
rect 17155 43778 17164 43838
rect 17224 43831 17233 43838
rect 17224 43800 19109 43831
rect 22500 43830 22528 43854
rect 28866 43830 28872 43842
rect 22220 43800 22334 43804
rect 22500 43802 28872 43830
rect 17224 43785 22334 43800
rect 28866 43790 28872 43802
rect 28924 43790 28930 43842
rect 17224 43778 17233 43785
rect 19063 43754 22334 43785
rect 22220 43750 22334 43754
rect 25566 43754 25644 43764
rect 18271 43684 18280 43744
rect 18340 43731 18349 43744
rect 18340 43709 18983 43731
rect 25566 43709 25576 43754
rect 18340 43698 25576 43709
rect 25632 43698 25644 43754
rect 18340 43697 25644 43698
rect 18340 43684 18349 43697
rect 18949 43688 25644 43697
rect 18949 43675 25621 43688
rect 18809 43594 18818 43654
rect 18878 43639 18887 43654
rect 28764 43639 28770 43650
rect 18878 43609 28770 43639
rect 18878 43594 18887 43609
rect 28764 43598 28770 43609
rect 28822 43598 28828 43650
rect 17715 43528 17724 43588
rect 17784 43572 17793 43588
rect 17784 43564 18780 43572
rect 18918 43564 21490 43572
rect 17784 43544 21490 43564
rect 17784 43528 17793 43544
rect 18748 43536 18944 43544
rect 15511 43454 15520 43514
rect 15580 43498 15589 43514
rect 15580 43470 21392 43498
rect 15580 43454 15589 43470
rect 13295 43374 13304 43434
rect 13364 43418 13373 43434
rect 13364 43390 21276 43418
rect 13364 43374 13373 43390
rect 12733 43266 12742 43326
rect 12802 43310 12811 43326
rect 12802 43282 21132 43310
rect 12802 43266 12811 43282
rect 21104 41162 21132 43282
rect 21086 41110 21092 41162
rect 21144 41110 21150 41162
rect 21248 41042 21276 43390
rect 21236 41036 21288 41042
rect 21236 40978 21288 40984
rect 21364 40868 21392 43470
rect 21346 40816 21352 40868
rect 21404 40816 21410 40868
rect 21462 40728 21490 43544
rect 29076 40768 29140 40774
rect 29076 40716 29082 40768
rect 29134 40716 29140 40768
rect 29076 40710 29140 40716
rect 21386 40216 21438 40222
rect 21386 40158 21438 40164
rect 28804 39952 28868 39954
rect 28762 39940 28868 39952
rect 28762 39888 28770 39940
rect 28822 39918 28868 39940
rect 28822 39888 28832 39918
rect 28762 39874 28832 39888
rect 28872 39480 28924 39486
rect 28872 39422 28924 39428
rect 21260 39388 21340 39406
rect 21260 39336 21268 39388
rect 21320 39336 21340 39388
rect 21260 39328 21340 39336
rect 21078 38192 21158 38202
rect 21078 38140 21092 38192
rect 21144 38140 21158 38192
rect 21078 38124 21158 38140
rect 28988 38192 29054 38200
rect 28988 38140 28996 38192
rect 29048 38140 29054 38192
rect 28988 38132 29054 38140
rect 23062 34814 23290 34828
rect 23062 34718 23078 34814
rect 23256 34718 23290 34814
rect 23062 34694 23290 34718
rect 19572 34104 19672 34118
rect 19572 33820 19586 34104
rect 19658 33820 19672 34104
rect 27118 34116 27250 34128
rect 27118 33852 27140 34116
rect 27236 33852 27250 34116
rect 27118 33836 27250 33852
rect 19572 33804 19672 33820
rect 23086 33226 23274 33240
rect 23086 32924 23106 33226
rect 23262 32924 23274 33226
rect 26920 33220 27076 33224
rect 26910 33204 27076 33220
rect 23086 32914 23274 32924
rect 26902 33192 27076 33204
rect 26902 32928 26926 33192
rect 27048 32928 27076 33192
rect 26902 32920 27076 32928
rect 26902 32908 27058 32920
rect 30436 31888 30708 31942
rect 30436 31722 30470 31888
rect 30640 31722 30708 31888
rect 30436 31684 30708 31722
rect 28614 22872 28876 22882
rect 28612 22867 28876 22872
rect 28612 22788 28755 22867
rect 28834 22788 28876 22867
rect 28612 22783 28876 22788
rect 28614 22710 28876 22783
rect 22376 21794 22556 21858
rect 22343 21699 22349 21794
rect 22444 21789 22556 21794
rect 22444 21704 22452 21789
rect 22537 21704 22556 21789
rect 22444 21699 22556 21704
rect 22376 21678 22556 21699
rect 22678 21097 22858 21140
rect 22678 20992 22739 21097
rect 22844 20992 22858 21097
rect 22678 20960 22858 20992
rect 18851 20347 20045 20385
rect 18851 2659 18889 20347
rect 21210 20052 21336 20080
rect 21210 19860 21234 20052
rect 21321 19860 21336 20052
rect 21210 19846 21336 19860
rect 3361 2621 18889 2659
rect 3361 258 3399 2621
rect 21164 2310 21390 2422
rect 11105 2305 21390 2310
rect 11105 2228 21239 2305
rect 21316 2228 21390 2305
rect 11105 2223 21390 2228
rect 11105 696 11192 2223
rect 21164 2172 21390 2223
rect 11105 600 11192 609
rect 7042 571 7184 598
rect 7042 510 7074 571
rect 7135 510 7184 571
rect 7042 484 7184 510
<< rmetal2 >>
rect 3316 188 3448 258
rect 3316 100 3340 188
rect 3424 100 3448 188
rect 3316 82 3448 100
<< via2 >>
rect 13858 44272 13918 44332
rect 14412 44178 14472 44238
rect 14965 44059 15025 44119
rect 24216 44060 24272 44116
rect 16063 43945 16123 44005
rect 26936 43946 26992 44002
rect 16616 43866 16676 43926
rect 17164 43778 17224 43838
rect 18280 43684 18340 43744
rect 25576 43698 25632 43754
rect 18818 43594 18878 43654
rect 17724 43528 17784 43588
rect 15520 43454 15580 43514
rect 13304 43374 13364 43434
rect 12742 43266 12802 43326
rect 23078 34718 23256 34814
rect 19586 33820 19658 34104
rect 27140 33852 27236 34116
rect 23124 32948 23246 33212
rect 26926 32928 27048 33192
rect 30470 31722 30640 31888
rect 28755 22788 28834 22867
rect 22452 21704 22537 21789
rect 22744 20997 22839 21092
rect 21234 19860 21321 20052
rect 21239 2228 21316 2305
rect 11105 609 11192 696
rect 7074 510 7135 571
rect 3340 100 3424 188
<< metal3 >>
rect 18278 45082 18342 45088
rect 14410 45068 14474 45074
rect 12740 45060 12804 45066
rect 12740 44990 12804 44996
rect 13302 45060 13366 45066
rect 13302 44990 13366 44996
rect 13856 45058 13920 45064
rect 14410 44998 14474 45004
rect 14963 45066 15027 45072
rect 17162 45070 17226 45076
rect 16061 45062 16125 45068
rect 12742 43331 12802 44990
rect 13304 43439 13364 44990
rect 13856 44988 13920 44994
rect 13858 44337 13918 44988
rect 13853 44332 13923 44337
rect 13853 44272 13858 44332
rect 13918 44272 13923 44332
rect 13853 44267 13923 44272
rect 14412 44243 14472 44998
rect 14963 44996 15027 45002
rect 15518 45042 15582 45048
rect 14407 44238 14477 44243
rect 14407 44178 14412 44238
rect 14472 44178 14477 44238
rect 14407 44173 14477 44178
rect 14965 44124 15025 44996
rect 16061 44992 16125 44998
rect 16614 45042 16678 45048
rect 15518 44972 15582 44978
rect 14960 44119 15030 44124
rect 14960 44059 14965 44119
rect 15025 44059 15030 44119
rect 14960 44054 15030 44059
rect 15520 43519 15580 44972
rect 16063 44010 16123 44992
rect 17162 45000 17226 45006
rect 17722 45060 17786 45066
rect 16614 44972 16678 44978
rect 16058 44005 16128 44010
rect 16058 43945 16063 44005
rect 16123 43945 16128 44005
rect 16058 43940 16128 43945
rect 16616 43931 16676 44972
rect 16611 43926 16681 43931
rect 16611 43866 16616 43926
rect 16676 43866 16681 43926
rect 16611 43861 16681 43866
rect 17164 43843 17224 45000
rect 18278 45012 18342 45018
rect 18816 45076 18880 45082
rect 28740 45068 28746 45070
rect 17722 44990 17786 44996
rect 17159 43838 17229 43843
rect 17159 43778 17164 43838
rect 17224 43778 17229 43838
rect 17159 43773 17229 43778
rect 17724 43593 17784 44990
rect 18280 43749 18340 45012
rect 18816 45006 18880 45012
rect 27614 45008 28746 45068
rect 18275 43744 18345 43749
rect 18275 43684 18280 43744
rect 18340 43684 18345 43744
rect 18275 43679 18345 43684
rect 18818 43659 18878 45006
rect 24211 44116 24277 44121
rect 24211 44060 24216 44116
rect 24272 44060 24277 44116
rect 24211 44055 24277 44060
rect 24214 43716 24274 44055
rect 26931 44002 26997 44007
rect 26931 43946 26936 44002
rect 26992 43946 26997 44002
rect 26931 43941 26997 43946
rect 25558 43754 25694 43772
rect 25558 43698 25576 43754
rect 25632 43698 25694 43754
rect 25558 43680 25694 43698
rect 26934 43684 26994 43941
rect 27614 43754 27674 45008
rect 28740 45006 28746 45008
rect 28810 45006 28816 45070
rect 18813 43654 18883 43659
rect 18813 43594 18818 43654
rect 18878 43594 18883 43654
rect 17719 43588 17789 43593
rect 18813 43589 18883 43594
rect 17719 43528 17724 43588
rect 17784 43528 17789 43588
rect 17719 43523 17789 43528
rect 15515 43514 15585 43519
rect 15515 43454 15520 43514
rect 15580 43454 15585 43514
rect 15515 43449 15585 43454
rect 13299 43434 13369 43439
rect 13299 43374 13304 43434
rect 13364 43374 13369 43434
rect 13299 43369 13369 43374
rect 12737 43326 12807 43331
rect 12737 43266 12742 43326
rect 12802 43266 12807 43326
rect 12737 43261 12807 43266
rect 1461 40444 1779 40449
rect 228 40124 234 40444
rect 554 40443 1780 40444
rect 554 40125 1461 40443
rect 1779 40125 1780 40443
rect 554 40124 1780 40125
rect 1461 40119 1779 40124
rect 23062 34814 23534 34826
rect 23062 34718 23078 34814
rect 23256 34718 23534 34814
rect 23062 34694 23534 34718
rect 23340 34124 23534 34694
rect 19572 34123 27322 34124
rect 19572 34104 26653 34123
rect 19572 33820 19586 34104
rect 19658 33820 26653 34104
rect 19572 33805 26653 33820
rect 26971 34116 27322 34123
rect 26971 33852 27140 34116
rect 27236 33852 27322 34116
rect 26971 33805 27322 33852
rect 19572 33804 27322 33805
rect 23072 33225 30870 33226
rect 23072 33212 28971 33225
rect 23072 32948 23124 33212
rect 23246 33192 28971 33212
rect 23246 32948 26926 33192
rect 23072 32928 26926 32948
rect 27048 32928 28971 33192
rect 23072 32907 28971 32928
rect 29289 32907 30870 33225
rect 23072 32906 30870 32907
rect 30428 31888 30746 32906
rect 30428 31722 30470 31888
rect 30640 31722 30746 31888
rect 30428 31694 30746 31722
rect 28614 22871 28876 22882
rect 28614 22784 28751 22871
rect 28838 22784 28876 22871
rect 28614 22710 28876 22784
rect 22376 21793 22556 21858
rect 22376 21700 22448 21793
rect 22541 21700 22556 21793
rect 22376 21678 22556 21700
rect 22678 21096 22858 21140
rect 22678 20993 22740 21096
rect 22843 20993 22858 21096
rect 22678 20960 22858 20993
rect 21210 20057 21336 20080
rect 21210 19855 21229 20057
rect 21326 19855 21336 20057
rect 21210 19846 21336 19855
rect 21164 2309 21390 2422
rect 21164 2224 21235 2309
rect 21320 2224 21390 2309
rect 21164 2172 21390 2224
rect 11100 696 11110 701
rect 11100 609 11105 696
rect 11100 604 11110 609
rect 11197 604 11203 701
rect 7042 576 7184 598
rect 7042 571 7076 576
rect 7042 510 7074 571
rect 7042 505 7076 510
rect 7140 505 7184 576
rect 7042 484 7184 505
rect 3304 188 3474 284
rect 3304 100 3340 188
rect 3424 100 3474 188
rect 3304 60 3474 100
<< via3 >>
rect 12740 44996 12804 45060
rect 13302 44996 13366 45060
rect 13856 44994 13920 45058
rect 14410 45004 14474 45068
rect 14963 45002 15027 45066
rect 15518 44978 15582 45042
rect 16061 44998 16125 45062
rect 16614 44978 16678 45042
rect 17162 45006 17226 45070
rect 17722 44996 17786 45060
rect 18278 45018 18342 45082
rect 18816 45012 18880 45076
rect 28746 45006 28810 45070
rect 234 40124 554 40444
rect 1461 40125 1779 40443
rect 26653 33805 26971 34123
rect 28971 32907 29289 33225
rect 28751 22867 28838 22871
rect 28751 22788 28755 22867
rect 28755 22788 28834 22867
rect 28834 22788 28838 22867
rect 28751 22784 28838 22788
rect 22448 21789 22541 21793
rect 22448 21704 22452 21789
rect 22452 21704 22537 21789
rect 22537 21704 22541 21789
rect 22448 21700 22541 21704
rect 22740 21092 22843 21096
rect 22740 20997 22744 21092
rect 22744 20997 22839 21092
rect 22839 20997 22843 21092
rect 22740 20993 22843 20997
rect 21229 20052 21326 20057
rect 21229 19860 21234 20052
rect 21234 19860 21321 20052
rect 21321 19860 21326 20052
rect 21229 19855 21326 19860
rect 21235 2305 21320 2309
rect 21235 2228 21239 2305
rect 21239 2228 21316 2305
rect 21316 2228 21320 2305
rect 21235 2224 21320 2228
rect 11110 696 11197 701
rect 11110 609 11192 696
rect 11192 609 11197 696
rect 11110 604 11197 609
rect 7076 571 7140 576
rect 7076 510 7135 571
rect 7135 510 7140 571
rect 7076 505 7140 510
rect 3340 100 3424 188
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 45094 8402 45152
rect 8894 45094 8954 45152
rect 9446 45094 9506 45152
rect 8342 44986 8404 45094
rect 8890 44986 8954 45094
rect 9444 44986 9506 45094
rect 8342 44952 8402 44986
rect 8894 44952 8954 44986
rect 9446 44952 9506 44986
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 45061 12818 45152
rect 13310 45061 13370 45152
rect 12739 45060 12818 45061
rect 12739 44996 12740 45060
rect 12804 44996 12818 45060
rect 12739 44995 12818 44996
rect 13301 45060 13370 45061
rect 13301 44996 13302 45060
rect 13366 44996 13370 45060
rect 13862 45059 13922 45152
rect 14414 45069 14474 45152
rect 13301 44995 13370 44996
rect 12758 44952 12818 44995
rect 13310 44952 13370 44995
rect 13855 45058 13922 45059
rect 13855 44994 13856 45058
rect 13920 44994 13922 45058
rect 14409 45068 14475 45069
rect 14409 45004 14410 45068
rect 14474 45004 14475 45068
rect 14966 45067 15026 45152
rect 14409 45003 14475 45004
rect 14962 45066 15028 45067
rect 13855 44993 13922 44994
rect 13862 44952 13922 44993
rect 14414 44952 14474 45003
rect 14962 45002 14963 45066
rect 15027 45002 15028 45066
rect 15518 45043 15578 45152
rect 16070 45063 16130 45152
rect 16060 45062 16130 45063
rect 14962 45001 15028 45002
rect 15517 45042 15583 45043
rect 14966 44952 15026 45001
rect 15517 44978 15518 45042
rect 15582 44978 15583 45042
rect 16060 44998 16061 45062
rect 16125 44998 16130 45062
rect 16622 45043 16682 45152
rect 17174 45071 17234 45152
rect 16060 44997 16130 44998
rect 15517 44977 15583 44978
rect 15518 44952 15578 44977
rect 16070 44952 16130 44997
rect 16613 45042 16682 45043
rect 16613 44978 16614 45042
rect 16678 44978 16682 45042
rect 17161 45070 17234 45071
rect 17161 45006 17162 45070
rect 17226 45006 17234 45070
rect 17726 45061 17786 45152
rect 18278 45083 18338 45152
rect 18277 45082 18343 45083
rect 17161 45005 17234 45006
rect 16613 44977 16682 44978
rect 16622 44952 16682 44977
rect 17174 44952 17234 45005
rect 17721 45060 17787 45061
rect 17721 44996 17722 45060
rect 17786 44996 17787 45060
rect 18277 45018 18278 45082
rect 18342 45018 18343 45082
rect 18830 45077 18890 45152
rect 18277 45017 18343 45018
rect 18815 45076 18890 45077
rect 17721 44995 17787 44996
rect 17726 44952 17786 44995
rect 18278 44952 18338 45017
rect 18815 45012 18816 45076
rect 18880 45012 18890 45076
rect 18815 45011 18890 45012
rect 18830 44952 18890 45011
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 45071 28826 45152
rect 28745 45070 28826 45071
rect 28745 45006 28746 45070
rect 28810 45006 28826 45070
rect 28745 45005 28826 45006
rect 28766 44952 28826 45005
rect 29318 44952 29378 45152
rect 200 40444 600 44152
rect 200 40124 234 40444
rect 554 40124 600 40444
rect 200 1000 600 40124
rect 800 39786 1200 44150
rect 1460 40443 29290 40444
rect 1460 40125 1461 40443
rect 1779 40125 29290 40443
rect 1460 40124 29290 40125
rect 800 39466 26972 39786
rect 800 1000 1200 39466
rect 26652 34123 26972 39466
rect 26652 33805 26653 34123
rect 26971 33805 26972 34123
rect 26652 33786 26972 33805
rect 28970 33225 29290 40124
rect 28970 32907 28971 33225
rect 29289 32907 29290 33225
rect 28970 32906 29290 32907
rect 28750 22871 30497 22872
rect 28750 22784 28751 22871
rect 28838 22784 30497 22871
rect 28750 22783 30497 22784
rect 21684 21793 22806 21836
rect 21684 21700 22448 21793
rect 22541 21700 22806 21793
rect 21684 21656 22806 21700
rect 21228 20057 21327 20058
rect 21228 19855 21229 20057
rect 21326 19855 21327 20057
rect 21228 19854 21327 19855
rect 21234 2309 21321 19854
rect 21234 2224 21235 2309
rect 21320 2224 21321 2309
rect 21234 2223 21321 2224
rect 21684 1496 21864 21656
rect 14906 1316 21864 1496
rect 22376 21097 22556 21134
rect 22376 21096 22844 21097
rect 22376 20993 22740 21096
rect 22843 20993 22844 21096
rect 22376 20992 22844 20993
rect 11109 701 11198 702
rect 11109 604 11110 701
rect 11197 604 11198 701
rect 11109 603 11198 604
rect 7075 576 7141 577
rect 7075 505 7076 576
rect 7140 571 7141 576
rect 7140 510 7342 571
rect 7140 505 7141 510
rect 7075 504 7141 505
rect 3304 200 3474 284
rect 7281 200 7342 510
rect 11110 200 11197 603
rect 3304 188 3494 200
rect 3304 100 3340 188
rect 3424 100 3494 188
rect 3304 60 3494 100
rect 3314 0 3494 60
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 1316
rect 22376 892 22556 20992
rect 18770 712 22556 892
rect 18770 0 18950 712
rect 30408 200 30497 22783
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 200
use flash_adc  flash_adc_0 ~/Documents/github_project/adc_dac2/mag
timestamp 1730795883
transform 0 1 17574 -1 0 22644
box -22008 1842 3604 13395
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 480 90 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 480 90 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 480 90 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 480 90 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 480 90 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 480 90 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 480 90 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 480 90 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
