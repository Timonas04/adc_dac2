magic
tech sky130A
magscale 1 2
timestamp 1730934983
<< pwell >>
rect 30680 18340 31040 18740
rect 28020 17760 28380 18160
<< locali >>
rect 25210 17291 25389 17652
<< metal1 >>
rect 28475 25361 29291 25461
rect 28475 23602 28575 25361
rect 30094 23840 30294 23846
rect 30728 23840 30928 23846
rect 29470 23834 29670 23840
rect 29170 23824 29370 23830
rect 29470 23776 29670 23782
rect 29772 23834 29972 23840
rect 30094 23782 30294 23788
rect 30404 23834 30604 23840
rect 30728 23782 30928 23788
rect 31042 23834 31242 23840
rect 29772 23776 29972 23782
rect 30404 23776 30604 23782
rect 31042 23776 31242 23782
rect 31374 23838 31574 23844
rect 31374 23780 31574 23786
rect 29170 23766 29370 23772
rect 24378 23502 28575 23602
rect 24378 23166 24478 23502
rect 26894 23208 26994 23502
rect 28768 22800 28774 22960
rect 28934 22800 29312 22960
rect 23718 22432 24539 22671
rect 23718 19825 23957 22432
rect 29036 21069 29114 21571
rect 26072 21056 26124 21062
rect 26072 20998 26124 21004
rect 28577 20991 29114 21069
rect 26864 20900 26916 20906
rect 24382 20894 24434 20900
rect 26864 20842 26916 20848
rect 24382 20836 24434 20842
rect 26032 20664 26038 20720
rect 26094 20664 26100 20720
rect 28552 20660 28558 20712
rect 28610 20660 28616 20712
rect 21304 19586 23957 19825
rect 28774 19910 28934 19916
rect 30084 19768 30154 19933
rect 13826 18057 14088 18068
rect 21304 18057 21543 19586
rect 24265 19316 24518 19634
rect 26822 19316 27062 19616
rect 24265 19286 27062 19316
rect 13826 17818 13837 18057
rect 14076 17818 21543 18057
rect 21781 19276 27062 19286
rect 28774 19276 28934 19750
rect 30015 19734 30154 19768
rect 30015 19712 30040 19734
rect 30006 19656 30040 19712
rect 30015 19641 30040 19656
rect 30109 19641 30154 19734
rect 30015 19612 30154 19641
rect 30084 19507 30154 19612
rect 30390 19510 30741 19933
rect 30980 19510 31331 19933
rect 31573 19738 31750 19929
rect 31573 19507 31772 19738
rect 21781 19116 28934 19276
rect 29952 19184 30008 19190
rect 21781 19076 27062 19116
rect 21781 19033 24518 19076
rect 25149 19045 26178 19076
rect 13826 17808 14088 17818
rect 15001 17587 18552 17645
rect 21781 17613 22034 19033
rect 19555 17587 22034 17613
rect 15001 17571 22034 17587
rect 24906 18934 26178 19045
rect 24906 18847 26156 18934
rect 24906 18190 25242 18847
rect 25360 18420 25720 18720
rect 25360 18360 25480 18420
rect 25560 18360 25720 18420
rect 25360 18320 25720 18360
rect 25940 18420 26300 18720
rect 25940 18360 26080 18420
rect 26140 18360 26300 18420
rect 25940 18320 26300 18360
rect 26540 18420 26900 18720
rect 26540 18360 26680 18420
rect 26740 18360 26900 18420
rect 26540 18320 26900 18360
rect 27140 18400 27500 18720
rect 27140 18340 27260 18400
rect 27320 18340 27500 18400
rect 27140 18320 27500 18340
rect 27720 18400 28080 18720
rect 27720 18340 27860 18400
rect 27920 18340 28080 18400
rect 27720 18320 28080 18340
rect 28320 18400 28680 18720
rect 28320 18340 28460 18400
rect 28520 18340 28680 18400
rect 28320 18320 28680 18340
rect 28900 18400 29260 18720
rect 28900 18340 29060 18400
rect 29120 18340 29260 18400
rect 28900 18320 29260 18340
rect 29500 18400 29860 18720
rect 29500 18340 29640 18400
rect 29700 18340 29860 18400
rect 29500 18320 29860 18340
rect 24906 17577 25402 18190
rect 25640 17880 26000 18160
rect 25640 17820 25780 17880
rect 25840 17820 26000 17880
rect 25640 17760 26000 17820
rect 26240 17840 26600 18160
rect 26240 17780 26380 17840
rect 26440 17780 26600 17840
rect 26840 17880 27200 18180
rect 26840 17820 26980 17880
rect 27040 17820 27200 17880
rect 26840 17780 27200 17820
rect 27420 17860 27780 18160
rect 27420 17800 27560 17860
rect 27620 17800 27780 17860
rect 26240 17760 26600 17780
rect 27420 17760 27780 17800
rect 28020 17840 28380 18160
rect 28020 17780 28160 17840
rect 28220 17780 28380 17840
rect 28600 17860 28960 18180
rect 28600 17800 28760 17860
rect 28820 17800 28960 17860
rect 28600 17780 28960 17800
rect 29200 17860 29560 18180
rect 29952 18160 30008 19128
rect 30087 18963 30438 19386
rect 30682 18966 31033 19389
rect 31276 18966 31627 19389
rect 30080 18320 30440 18720
rect 30680 18340 31040 18740
rect 31280 18320 31640 18720
rect 31704 18180 31772 19507
rect 29200 17800 29340 17860
rect 29400 17800 29560 17860
rect 29200 17780 29560 17800
rect 28020 17760 28380 17780
rect 29800 17760 30160 18160
rect 30380 17760 30740 18160
rect 30980 17760 31340 18160
rect 31580 17755 31772 18180
rect 31580 17745 31720 17755
rect 24906 17575 28975 17577
rect 22851 17571 28975 17575
rect 15001 17494 28975 17571
rect 15001 17391 16275 17494
rect 18401 17464 28975 17494
rect 18401 17462 24744 17464
rect 18401 17329 19706 17462
rect 21767 17458 24744 17462
rect 24948 17458 28140 17464
rect 21767 17424 24706 17458
rect 24958 17426 28094 17458
rect 28352 17426 28975 17464
rect 24958 17424 26521 17426
rect 21767 17384 23118 17424
rect 21767 17335 23002 17384
rect 25207 17372 26521 17424
rect 28690 17376 28975 17426
rect 25207 17341 26560 17372
rect 18401 17291 18552 17329
rect 21767 17327 22034 17335
rect 21767 17285 21918 17327
rect 25207 17285 25402 17341
rect 26442 17310 26560 17341
rect 28824 17280 28975 17376
rect 31580 17360 31720 17457
rect 31623 17344 31679 17350
rect 31623 17282 31679 17288
rect 16708 16242 16714 16294
rect 16766 16242 16772 16294
rect 20226 16246 20232 16298
rect 20284 16246 20290 16298
rect 23532 16234 23538 16286
rect 23590 16234 23596 16286
rect 26936 16234 26942 16286
rect 26994 16234 27000 16286
rect 30420 16244 30426 16296
rect 30478 16244 30484 16296
rect 17840 12819 18107 12914
rect 21112 12819 21497 12914
rect 24684 12819 24882 12914
rect 28010 12819 28292 12914
rect 31464 12819 31691 12914
rect 8411 12315 8463 12321
rect 8411 12257 8463 12263
rect 8423 12128 8451 12257
rect 15011 12224 15017 12323
rect 15116 12224 15122 12323
rect 18012 12284 18107 12819
rect 18439 12237 18445 12336
rect 18544 12237 18550 12336
rect 21402 12259 21497 12819
rect 18012 12183 18107 12189
rect 21816 12166 21822 12265
rect 21921 12166 21927 12265
rect 24787 12259 24882 12819
rect 21402 12158 21497 12164
rect 25240 12178 25246 12277
rect 25345 12178 25351 12277
rect 28197 12259 28292 12819
rect 31596 12279 31691 12819
rect 24787 12158 24882 12164
rect 28628 12179 28634 12278
rect 28733 12179 28739 12278
rect 31596 12178 31691 12184
rect 28197 12158 28292 12164
rect 9824 12140 9876 12146
rect 8423 12100 9824 12128
rect 9824 12082 9876 12088
rect 9216 11996 9222 12048
rect 9274 12047 9280 12048
rect 15958 12047 16008 12125
rect 9274 11997 16008 12047
rect 9274 11996 9280 11997
rect 12019 11888 12071 11894
rect 12143 11879 12149 11931
rect 12201 11925 12207 11931
rect 19363 11925 19404 12121
rect 12201 11884 19404 11925
rect 12201 11879 12207 11884
rect 22769 11847 22798 12115
rect 12071 11836 22798 11847
rect 12019 11830 22798 11836
rect 12030 11818 22798 11830
rect 11866 11734 11872 11786
rect 11924 11780 11930 11786
rect 26163 11780 26203 12120
rect 11924 11740 26203 11780
rect 11924 11734 11930 11740
rect 11733 11661 11739 11713
rect 11791 11706 11797 11713
rect 29564 11706 29603 12120
rect 11791 11667 29603 11706
rect 11791 11661 11797 11667
rect 15011 11506 15017 11605
rect 15116 11506 15505 11605
rect 18006 11425 18012 11520
rect 18107 11425 18113 11520
rect 18439 11506 18445 11605
rect 18544 11506 18803 11605
rect 21396 11455 21402 11550
rect 21497 11455 21503 11550
rect 21816 11506 21822 11605
rect 21921 11506 22237 11605
rect 24781 11480 24787 11575
rect 24882 11480 24888 11575
rect 25713 11506 25719 11605
rect 25818 11506 25914 11605
rect 28191 11465 28197 11560
rect 28292 11465 28298 11560
rect 28628 11506 28634 11605
rect 28733 11506 29039 11605
rect 31590 11484 31596 11579
rect 31691 11484 31697 11579
rect 16708 10436 16714 10488
rect 16766 10436 16772 10488
rect 20226 10442 20232 10494
rect 20284 10442 20290 10494
rect 23532 10440 23538 10492
rect 23590 10440 23596 10492
rect 26936 10440 26942 10492
rect 26994 10440 27000 10492
rect 30420 10428 30426 10480
rect 30478 10428 30484 10480
rect 17850 7019 18079 7114
rect 21157 7019 21500 7114
rect 24420 7019 24886 7114
rect 28069 7019 28287 7114
rect 31267 7019 31689 7114
rect 15050 6422 15056 6521
rect 15155 6422 15161 6521
rect 17984 6436 18079 7019
rect 21405 6436 21500 7019
rect 21392 6422 21516 6436
rect 17984 6335 18079 6341
rect 21392 6326 21402 6422
rect 21500 6326 21516 6422
rect 24791 6450 24886 7019
rect 25217 6871 25316 6877
rect 25217 6766 25316 6772
rect 24791 6349 24886 6355
rect 28192 6455 28287 7019
rect 31594 6480 31689 7019
rect 28192 6354 28287 6360
rect 28617 6388 28741 6398
rect 12521 6238 12573 6244
rect 12658 6224 12664 6276
rect 12716 6268 12722 6276
rect 15965 6268 16001 6318
rect 12716 6232 16001 6268
rect 12716 6224 12722 6232
rect 12573 6186 12576 6208
rect 12521 6180 12576 6186
rect 12530 6171 12576 6180
rect 19367 6171 19400 6317
rect 21392 6316 21516 6326
rect 12530 6138 19400 6171
rect 12390 6064 12396 6116
rect 12448 6113 12454 6116
rect 22760 6113 22806 6323
rect 12448 6110 12498 6113
rect 19618 6110 22806 6113
rect 12448 6067 22806 6110
rect 12448 6064 12454 6067
rect 12211 5967 12217 6019
rect 12269 6017 12275 6019
rect 26159 6017 26208 6325
rect 28617 6289 28627 6388
rect 28726 6289 28741 6388
rect 31594 6379 31689 6385
rect 28617 6279 28741 6289
rect 12269 5968 26208 6017
rect 12269 5967 12275 5968
rect 12054 5878 12060 5930
rect 12112 5927 12118 5930
rect 29560 5927 29606 6323
rect 12112 5881 29606 5927
rect 12112 5878 12118 5881
rect 15050 5706 15056 5805
rect 15155 5706 15370 5805
rect 18434 5706 18440 5805
rect 18539 5706 18808 5805
rect 21811 5706 21817 5805
rect 21916 5706 22141 5805
rect 24781 5751 24876 5757
rect 25712 5706 25718 5805
rect 25817 5706 25823 5805
rect 28621 5706 28627 5805
rect 28726 5706 28957 5805
rect 24781 5650 24876 5656
rect 31588 5646 31594 5741
rect 31689 5646 31695 5741
rect 28163 5235 28169 5330
rect 28264 5235 28270 5330
rect 7447 4633 7499 4639
rect 7139 4612 7447 4621
rect 7127 4606 7447 4612
rect 7179 4593 7447 4606
rect 16708 4630 16714 4682
rect 16766 4630 16772 4682
rect 20226 4630 20232 4682
rect 20284 4630 20290 4682
rect 23532 4634 23538 4686
rect 23590 4634 23596 4686
rect 26934 4640 26940 4692
rect 26992 4640 26998 4692
rect 30420 4644 30426 4696
rect 30478 4644 30484 4696
rect 7447 4575 7499 4581
rect 7127 4548 7179 4554
rect 8192 4514 8244 4520
rect 6938 4462 6944 4514
rect 6996 4502 7002 4514
rect 6996 4474 8192 4502
rect 6996 4462 7002 4474
rect 8192 4456 8244 4462
rect 8834 4435 8886 4441
rect 6377 4383 6383 4435
rect 6435 4423 6441 4435
rect 6435 4395 8834 4423
rect 6435 4383 6441 4395
rect 8834 4377 8886 4383
rect 29968 3983 29985 3989
rect 29925 3917 29985 3923
rect 17959 2492 18132 2507
rect 17959 2355 17974 2492
rect 18111 2355 18132 2492
rect 17959 2340 18132 2355
rect 21364 2492 21519 2500
rect 21364 2355 21372 2492
rect 21509 2355 21519 2492
rect 21364 2345 21519 2355
rect 24743 2492 24908 2506
rect 24743 2355 24757 2492
rect 24894 2355 24908 2492
rect 24743 2342 24908 2355
rect 28136 2492 28301 2507
rect 28136 2355 28152 2492
rect 28289 2355 28301 2492
rect 28136 2343 28301 2355
rect 31484 2492 31649 2502
rect 31484 2355 31501 2492
rect 31638 2355 31724 2492
rect 31484 2338 31649 2355
rect 12170 390 12176 442
rect 12228 438 12234 442
rect 15961 438 16005 522
rect 12228 394 16005 438
rect 12228 390 12234 394
rect 11791 379 11843 385
rect 11217 360 11269 366
rect 12049 354 12125 387
rect 11791 321 11843 327
rect 12045 348 12125 354
rect 11217 302 11269 308
rect 11224 102 11262 302
rect 11800 175 11834 321
rect 12097 327 12125 348
rect 19363 327 19404 521
rect 12097 296 19404 327
rect 11915 289 11967 295
rect 12045 290 19404 296
rect 12049 286 19404 290
rect 22765 243 22802 519
rect 11967 237 22802 243
rect 11915 231 22802 237
rect 11922 206 22802 231
rect 26166 175 26200 517
rect 11800 141 26200 175
rect 29564 102 29602 519
rect 11224 64 29602 102
<< via1 >>
rect 29170 23772 29370 23824
rect 29470 23782 29670 23834
rect 29772 23782 29972 23834
rect 30094 23788 30294 23840
rect 30404 23782 30604 23834
rect 30728 23788 30928 23840
rect 31042 23782 31242 23834
rect 31374 23786 31574 23838
rect 28774 22800 28934 22960
rect 26072 21004 26124 21056
rect 24382 20842 24434 20894
rect 26864 20848 26916 20900
rect 26038 20664 26094 20720
rect 28558 20660 28610 20712
rect 28774 19750 28934 19910
rect 13837 17818 14076 18057
rect 30040 19641 30109 19734
rect 29952 19128 30008 19184
rect 25480 18360 25560 18420
rect 26080 18360 26140 18420
rect 26680 18360 26740 18420
rect 27260 18340 27320 18400
rect 27860 18340 27920 18400
rect 28460 18340 28520 18400
rect 29060 18340 29120 18400
rect 29640 18340 29700 18400
rect 25780 17820 25840 17880
rect 26380 17780 26440 17840
rect 26980 17820 27040 17880
rect 27560 17800 27620 17860
rect 28160 17780 28220 17840
rect 28760 17800 28820 17860
rect 29340 17800 29400 17860
rect 31623 17288 31679 17344
rect 16714 16242 16766 16294
rect 20232 16246 20284 16298
rect 23538 16234 23590 16286
rect 26942 16234 26994 16286
rect 30426 16244 30478 16296
rect 17636 15554 17696 15614
rect 21003 15498 21072 15567
rect 23854 15516 23914 15576
rect 27974 15528 28034 15588
rect 29938 15517 29998 15577
rect 8411 12263 8463 12315
rect 15017 12224 15116 12323
rect 18012 12189 18107 12284
rect 18445 12237 18544 12336
rect 21402 12164 21497 12259
rect 21822 12166 21921 12265
rect 24787 12164 24882 12259
rect 25246 12178 25345 12277
rect 28197 12164 28292 12259
rect 28634 12179 28733 12278
rect 31596 12184 31691 12279
rect 9824 12088 9876 12140
rect 9222 11996 9274 12048
rect 12019 11836 12071 11888
rect 12149 11879 12201 11931
rect 11872 11734 11924 11786
rect 11739 11661 11791 11713
rect 15017 11506 15116 11605
rect 18012 11425 18107 11520
rect 18445 11506 18544 11605
rect 21402 11455 21497 11550
rect 21822 11506 21921 11605
rect 24787 11480 24882 11575
rect 25719 11506 25818 11605
rect 28197 11465 28292 11560
rect 28634 11506 28733 11605
rect 31596 11484 31691 11579
rect 16714 10436 16766 10488
rect 20232 10442 20284 10494
rect 23538 10440 23590 10492
rect 26942 10440 26994 10492
rect 30426 10428 30478 10480
rect 21063 9803 21123 9807
rect 17107 9781 17167 9796
rect 17092 9736 17167 9781
rect 21060 9747 21123 9803
rect 24395 9796 24460 9800
rect 21060 9743 21120 9747
rect 24395 9736 24484 9796
rect 27600 9743 27660 9803
rect 17092 9721 17152 9736
rect 24395 9735 24460 9736
rect 30169 9734 30229 9794
rect 15056 6422 15155 6521
rect 17984 6426 18079 6436
rect 17984 6346 18080 6426
rect 18440 6400 18539 6499
rect 17984 6341 18079 6346
rect 21402 6326 21500 6422
rect 21817 6415 21916 6514
rect 25217 6772 25316 6871
rect 24791 6355 24886 6450
rect 28192 6360 28287 6455
rect 12521 6186 12573 6238
rect 12664 6224 12716 6276
rect 12396 6064 12448 6116
rect 12217 5967 12269 6019
rect 28627 6289 28726 6388
rect 31594 6385 31689 6480
rect 12060 5878 12112 5930
rect 15056 5706 15155 5805
rect 17984 5676 18079 5771
rect 18440 5706 18539 5805
rect 21405 5656 21500 5751
rect 21817 5706 21916 5805
rect 24781 5656 24876 5751
rect 25718 5706 25817 5805
rect 28627 5706 28726 5805
rect 31594 5646 31689 5741
rect 28169 5235 28264 5330
rect 7127 4554 7179 4606
rect 7447 4581 7499 4633
rect 16714 4630 16766 4682
rect 20232 4630 20284 4682
rect 23538 4634 23590 4686
rect 26940 4640 26992 4692
rect 30426 4644 30478 4696
rect 6944 4462 6996 4514
rect 8192 4462 8244 4514
rect 6383 4383 6435 4435
rect 8834 4383 8886 4435
rect 17631 3946 17691 4006
rect 20992 3946 21052 4006
rect 24487 3906 24552 3971
rect 26529 3941 26589 4001
rect 29908 3983 29968 3991
rect 29908 3931 29985 3983
rect 29925 3923 29985 3931
rect 17974 2355 18111 2492
rect 21372 2355 21509 2492
rect 24757 2355 24894 2492
rect 28152 2355 28289 2492
rect 31501 2355 31638 2492
rect 12176 390 12228 442
rect 11217 308 11269 360
rect 11791 327 11843 379
rect 12045 296 12097 348
rect 11915 237 11967 289
<< metal2 >>
rect 4320 44858 28769 44860
rect 4313 44802 4322 44858
rect 4378 44802 28769 44858
rect 4320 44800 28769 44802
rect 28829 44800 28838 44860
rect 4451 44684 18816 44686
rect 4444 44628 4453 44684
rect 4509 44628 18816 44684
rect 4451 44626 18816 44628
rect 18876 44626 18885 44686
rect 27641 44643 27650 44703
rect 27710 44692 27719 44703
rect 27710 44654 31493 44692
rect 27710 44643 27719 44654
rect 27100 44559 27109 44619
rect 27169 44610 27178 44619
rect 27169 44567 31404 44610
rect 27169 44559 27178 44567
rect 4625 44525 18270 44527
rect 4618 44469 4627 44525
rect 4683 44469 18270 44525
rect 4625 44467 18270 44469
rect 18330 44467 18339 44527
rect 26546 44469 26555 44529
rect 26615 44519 26624 44529
rect 26615 44479 31313 44519
rect 26615 44469 26624 44479
rect 4151 44390 17720 44392
rect 4144 44334 4153 44390
rect 4209 44334 17720 44390
rect 4151 44332 17720 44334
rect 17780 44332 17789 44392
rect 25983 44379 25992 44439
rect 26052 44433 26061 44439
rect 26052 44385 31219 44433
rect 26052 44379 26061 44385
rect 25447 44278 25456 44338
rect 25516 44329 25525 44338
rect 25516 44287 31126 44329
rect 25516 44278 25525 44287
rect 3999 44239 17162 44241
rect 3992 44183 4001 44239
rect 4057 44183 17162 44239
rect 3999 44181 17162 44183
rect 17222 44181 17231 44241
rect 24897 44186 24906 44246
rect 24966 44236 24975 44246
rect 24966 44196 31041 44236
rect 24966 44186 24975 44196
rect 24344 44159 24404 44168
rect 4799 44128 16611 44130
rect 4792 44072 4801 44128
rect 4857 44072 16611 44128
rect 4799 44070 16611 44072
rect 16671 44070 16680 44130
rect 24404 44105 30962 44152
rect 24344 44090 24404 44099
rect 3843 44003 4121 44008
rect 3838 43947 3847 44003
rect 3903 43998 4121 44003
rect 16047 43998 16056 44005
rect 3903 43952 16056 43998
rect 3903 43947 4121 43952
rect 3843 43943 4121 43947
rect 16047 43945 16056 43952
rect 16116 43945 16125 44005
rect 23792 44004 23801 44064
rect 23861 44058 23870 44064
rect 23861 44010 30868 44058
rect 23861 44004 23870 44010
rect 21019 43893 21028 43953
rect 21088 43940 21097 43953
rect 21088 43906 30763 43940
rect 21088 43893 21097 43906
rect 3714 43879 3984 43881
rect 3707 43823 3716 43879
rect 3772 43874 3984 43879
rect 15499 43874 15508 43881
rect 3772 43828 15508 43874
rect 3772 43823 3984 43828
rect 3714 43821 3984 43823
rect 15499 43821 15508 43828
rect 15568 43821 15577 43881
rect 20473 43801 20482 43861
rect 20542 43848 20551 43861
rect 20542 43814 30669 43848
rect 20542 43801 20551 43814
rect 3557 43782 3685 43785
rect 3551 43726 3560 43782
rect 3616 43779 3685 43782
rect 14953 43779 14962 43785
rect 3616 43730 14962 43779
rect 3616 43726 3685 43730
rect 3557 43723 3685 43726
rect 14953 43725 14962 43730
rect 15022 43725 15031 43785
rect 4946 43665 5136 43667
rect 4939 43609 4948 43665
rect 5004 43660 5136 43665
rect 14406 43660 14415 43668
rect 5004 43615 14415 43660
rect 5004 43609 5136 43615
rect 4946 43607 5136 43609
rect 14406 43608 14415 43615
rect 14475 43608 14484 43668
rect 5077 43545 13859 43547
rect 5070 43489 5079 43545
rect 5135 43489 13859 43545
rect 5077 43487 13859 43489
rect 13919 43487 13928 43547
rect 3423 43464 3479 43471
rect 3421 43462 3711 43464
rect 3421 43406 3423 43462
rect 3479 43457 3711 43462
rect 3479 43411 13362 43457
rect 3479 43406 3711 43411
rect 3421 43404 3711 43406
rect 3423 43397 3479 43404
rect 13270 43399 13362 43411
rect 13270 43390 13369 43399
rect 13270 43375 13309 43390
rect 3285 43343 12762 43345
rect 3278 43287 3287 43343
rect 3343 43287 12762 43343
rect 3285 43285 12762 43287
rect 12822 43285 12831 43345
rect 13309 43321 13369 43330
rect 30635 26230 30669 43814
rect 26036 26196 30669 26230
rect 26036 23615 26070 26196
rect 30729 26141 30763 43906
rect 27331 26107 30763 26141
rect 27331 23621 27365 26107
rect 30820 26068 30868 44010
rect 29246 26020 30868 26068
rect 29246 23824 29294 26020
rect 30915 25958 30962 44105
rect 29547 25911 30962 25958
rect 29547 23834 29594 25911
rect 31001 25863 31041 44196
rect 29852 25823 31041 25863
rect 29852 23834 29892 25823
rect 31084 25779 31126 44287
rect 30173 25737 31126 25779
rect 30173 23840 30215 25737
rect 31171 25698 31219 44385
rect 30480 25650 31219 25698
rect 29164 23772 29170 23824
rect 29370 23772 29376 23824
rect 29464 23782 29470 23834
rect 29670 23782 29676 23834
rect 29766 23782 29772 23834
rect 29972 23782 29978 23834
rect 30088 23788 30094 23840
rect 30294 23788 30300 23840
rect 30480 23834 30528 25650
rect 31273 25620 31313 44479
rect 30808 25580 31313 25620
rect 30808 23840 30848 25580
rect 31361 25544 31404 44567
rect 31121 25501 31404 25544
rect 30398 23782 30404 23834
rect 30604 23782 30610 23834
rect 30722 23788 30728 23840
rect 30928 23788 30934 23840
rect 31121 23834 31164 25501
rect 31455 23838 31493 44654
rect 31036 23782 31042 23834
rect 31242 23782 31248 23834
rect 31368 23786 31374 23838
rect 31574 23786 31580 23838
rect 24075 23581 26070 23615
rect 24075 20885 24109 23581
rect 26036 23568 26070 23581
rect 26549 23587 27365 23621
rect 26066 21004 26072 21056
rect 26124 21053 26130 21056
rect 26124 21007 26439 21053
rect 26124 21004 26130 21007
rect 24376 20885 24382 20894
rect 24075 20851 24382 20885
rect 24376 20842 24382 20851
rect 24434 20842 24440 20894
rect 26038 20720 26094 20726
rect 26038 19184 26094 20664
rect 26393 19334 26439 21007
rect 26549 20891 26583 23587
rect 27331 23568 27365 23587
rect 28774 22960 28934 22966
rect 26858 20891 26864 20900
rect 26549 20857 26864 20891
rect 26858 20848 26864 20857
rect 26916 20848 26922 20900
rect 28558 20712 28610 20718
rect 28558 20654 28610 20660
rect 28561 19334 28607 20654
rect 28774 19910 28934 22800
rect 28768 19750 28774 19910
rect 28934 19750 28940 19910
rect 30015 19734 30129 19768
rect 30015 19641 30040 19734
rect 30109 19712 30129 19734
rect 30109 19656 31760 19712
rect 30109 19641 30129 19656
rect 30015 19612 30129 19641
rect 26393 19288 30475 19334
rect 26038 19128 29952 19184
rect 30008 19128 30014 19184
rect 23465 19018 23474 19078
rect 23534 19070 23543 19078
rect 23534 19026 29691 19070
rect 23534 19018 23543 19026
rect 23660 18911 23669 18980
rect 23738 18911 29408 18980
rect 23845 18789 23854 18849
rect 23914 18843 23923 18849
rect 23914 18794 29110 18843
rect 23914 18789 23923 18794
rect 24066 18702 24075 18762
rect 24135 18753 24144 18762
rect 24135 18711 28208 18753
rect 24135 18702 24144 18711
rect 24247 18599 24256 18659
rect 24316 18654 24325 18659
rect 24316 18604 27921 18654
rect 24316 18599 24325 18604
rect 24415 18506 24424 18566
rect 24484 18565 24493 18566
rect 24484 18507 27626 18565
rect 24484 18506 24493 18507
rect 25460 18420 25580 18440
rect 25460 18415 25480 18420
rect 25440 18406 25480 18415
rect 25560 18360 25580 18420
rect 26060 18420 26160 18440
rect 26060 18401 26080 18420
rect 25500 18346 25580 18360
rect 25440 18340 25580 18346
rect 26038 18360 26080 18401
rect 26140 18360 26160 18420
rect 26660 18420 26760 18440
rect 26660 18397 26680 18420
rect 26740 18398 26760 18420
rect 26038 18340 26160 18360
rect 26641 18360 26680 18397
rect 25440 18337 25500 18340
rect 13826 18057 14088 18068
rect 13826 17818 13837 18057
rect 14076 17818 14088 18057
rect 26038 18054 26103 18340
rect 26641 18339 26681 18360
rect 26672 18338 26681 18339
rect 26741 18340 26760 18398
rect 27240 18400 27340 18420
rect 27240 18381 27260 18400
rect 27227 18340 27260 18381
rect 27320 18340 27340 18400
rect 26741 18338 26750 18340
rect 27227 18334 27340 18340
rect 27240 18320 27340 18334
rect 27272 18120 27319 18320
rect 25024 17989 25033 18054
rect 25098 17989 26103 18054
rect 26804 18073 27319 18120
rect 25760 17880 25860 17900
rect 25760 17874 25780 17880
rect 13826 17808 14088 17818
rect 25243 17814 25252 17874
rect 25312 17820 25780 17874
rect 25840 17820 25860 17880
rect 25312 17814 25860 17820
rect 26360 17840 26460 17860
rect 26360 17815 26380 17840
rect 25760 17800 25860 17814
rect 26342 17780 26380 17815
rect 26440 17780 26460 17840
rect 26342 17760 26460 17780
rect 24805 17643 24814 17703
rect 24874 17701 24883 17703
rect 26342 17701 26398 17760
rect 24874 17645 26398 17701
rect 24874 17643 24883 17645
rect 26804 17460 26851 18073
rect 26960 17880 27060 17900
rect 27568 17880 27626 18507
rect 27871 18420 27921 18604
rect 27840 18400 27940 18420
rect 27840 18340 27860 18400
rect 27920 18340 27940 18400
rect 27840 18320 27940 18340
rect 26960 17820 26980 17880
rect 27040 17820 27060 17880
rect 26960 17800 27060 17820
rect 27540 17860 27640 17880
rect 28166 17860 28208 18711
rect 29061 18420 29110 18794
rect 28440 18400 28540 18420
rect 28440 18340 28460 18400
rect 28520 18340 28540 18400
rect 28440 18320 28540 18340
rect 29040 18400 29140 18420
rect 29040 18340 29060 18400
rect 29120 18340 29140 18400
rect 29040 18320 29140 18340
rect 27540 17800 27560 17860
rect 27620 17800 27640 17860
rect 26980 17623 27030 17800
rect 27540 17780 27640 17800
rect 28140 17840 28240 17860
rect 28140 17780 28160 17840
rect 28220 17780 28240 17840
rect 27568 17779 27626 17780
rect 28140 17760 28240 17780
rect 26975 17614 27035 17623
rect 26975 17545 27035 17554
rect 26798 17451 26858 17460
rect 26798 17382 26858 17391
rect 16714 16294 16766 16300
rect 16714 16236 16766 16242
rect 20232 16298 20284 16304
rect 20232 16240 20284 16246
rect 23538 16286 23590 16292
rect 7140 12494 7200 12503
rect 7200 12434 7324 12454
rect 7140 12426 7324 12434
rect 7140 12425 7200 12426
rect 8407 12362 8467 12371
rect 15017 12323 15116 12329
rect 8405 12302 8407 12315
rect 8467 12302 8469 12315
rect 4625 12266 4685 12275
rect 8405 12263 8411 12302
rect 8463 12263 8469 12302
rect 4625 12205 4685 12206
rect 4349 12145 4685 12205
rect 12146 12220 12206 12229
rect 4142 11736 4151 11796
rect 4211 11780 4220 11796
rect 4211 11752 4302 11780
rect 4211 11736 4220 11752
rect 3990 11605 3999 11665
rect 4059 11605 4223 11665
rect 3549 11492 3558 11552
rect 3618 11539 3627 11552
rect 3618 11504 3711 11539
rect 3618 11492 3627 11504
rect 3412 11182 3421 11242
rect 3481 11226 3490 11242
rect 3481 11198 3597 11226
rect 3481 11182 3490 11198
rect 3276 11033 3285 11093
rect 3345 11077 3354 11093
rect 3345 11049 3523 11077
rect 3345 11033 3354 11049
rect 3495 6415 3523 11049
rect 3569 6547 3597 11198
rect 3676 7617 3711 11504
rect 3844 11492 3904 11501
rect 3904 11432 4068 11492
rect 3844 11423 3904 11432
rect 3743 11293 3803 11302
rect 3743 11224 3803 11233
rect 3759 10010 3787 11224
rect 4008 10176 4068 11432
rect 4008 10120 4010 10176
rect 4066 10120 4068 10176
rect 4008 10118 4068 10120
rect 4010 10111 4066 10118
rect 3759 9982 4090 10010
rect 3663 7456 3723 7617
rect 3663 7400 3665 7456
rect 3721 7400 3723 7456
rect 3663 7398 3723 7400
rect 3665 7391 3721 7398
rect 3569 6519 4004 6547
rect 3495 6387 3835 6415
rect 3807 4423 3835 6387
rect 3976 4502 4004 6519
rect 4062 5312 4090 9982
rect 4163 5573 4223 11605
rect 4274 8694 4302 11752
rect 4349 8816 4409 12145
rect 8212 12110 8221 12170
rect 8281 12154 8290 12170
rect 15017 12219 15116 12224
rect 8281 12126 8612 12154
rect 12146 12151 12206 12160
rect 8281 12110 8290 12126
rect 9818 12088 9824 12140
rect 9876 12128 9882 12140
rect 9876 12100 9900 12128
rect 9876 12088 9882 12100
rect 7924 12067 7984 12076
rect 7924 11998 7984 12007
rect 9222 12048 9274 12054
rect 9222 11990 9274 11996
rect 11345 11918 11785 11957
rect 12155 11937 12196 12151
rect 14852 12028 14861 12219
rect 15052 12028 15162 12219
rect 11746 11719 11785 11918
rect 12149 11931 12201 11937
rect 12013 11836 12019 11888
rect 12071 11836 12077 11888
rect 12149 11873 12201 11879
rect 11872 11786 11924 11792
rect 11872 11728 11924 11734
rect 11739 11713 11791 11719
rect 11739 11655 11791 11661
rect 11878 11543 11918 11728
rect 11868 11534 11928 11543
rect 11868 11465 11928 11474
rect 12031 10182 12060 11836
rect 15017 11605 15116 12028
rect 15017 11500 15116 11506
rect 12660 10858 12720 10867
rect 12660 10789 12720 10798
rect 12016 10173 12076 10182
rect 12016 10104 12076 10113
rect 12518 9494 12578 9503
rect 12518 9425 12578 9434
rect 12392 8820 12452 8829
rect 4342 8760 4351 8816
rect 4407 8760 4416 8816
rect 4349 8758 4409 8760
rect 12392 8751 12452 8760
rect 4274 8666 4450 8694
rect 4163 5453 4291 5573
rect 4062 5284 4379 5312
rect 4351 4594 4379 5284
rect 4422 4680 4450 8666
rect 12214 8138 12274 8147
rect 12214 8069 12274 8078
rect 12056 7462 12116 7471
rect 12056 7393 12116 7402
rect 11912 6777 11972 6786
rect 11912 6708 11972 6717
rect 11787 6098 11847 6107
rect 11787 6029 11847 6038
rect 4422 4652 7324 4680
rect 7121 4594 7127 4606
rect 4351 4566 7127 4594
rect 7121 4554 7127 4566
rect 7179 4554 7185 4606
rect 7441 4581 7447 4633
rect 7499 4621 7505 4633
rect 7499 4593 7876 4621
rect 7499 4581 7505 4593
rect 6944 4514 6996 4520
rect 3976 4474 6944 4502
rect 8186 4462 8192 4514
rect 8244 4502 8250 4514
rect 8244 4474 8704 4502
rect 8244 4462 8250 4474
rect 6944 4456 6996 4462
rect 6383 4435 6435 4441
rect 3807 4395 6383 4423
rect 8828 4383 8834 4435
rect 8886 4423 8892 4435
rect 8886 4395 9900 4423
rect 8886 4383 8892 4395
rect 6383 4377 6435 4383
rect 11224 360 11262 4201
rect 11800 379 11834 6029
rect 11211 308 11217 360
rect 11269 308 11275 360
rect 11785 327 11791 379
rect 11843 327 11849 379
rect 11923 289 11960 6708
rect 12063 5936 12109 7393
rect 12219 6025 12268 8069
rect 12399 6122 12445 8751
rect 12531 6238 12564 9425
rect 12672 6282 12708 10789
rect 16717 10494 16763 16236
rect 17614 15614 17711 15630
rect 17614 15554 17636 15614
rect 17696 15554 17711 15614
rect 17614 15537 17711 15554
rect 18445 12336 18544 12342
rect 18006 12189 18012 12284
rect 18107 12189 18113 12284
rect 18012 11520 18107 12189
rect 18445 11605 18544 12237
rect 18445 11500 18544 11506
rect 18012 11419 18107 11425
rect 20235 10500 20281 16240
rect 23538 16228 23590 16234
rect 26942 16286 26994 16292
rect 26942 16228 26994 16234
rect 20987 15567 21084 15579
rect 20987 15498 21003 15567
rect 21072 15498 21084 15567
rect 20987 15486 21084 15498
rect 21822 12265 21921 12271
rect 21396 12164 21402 12259
rect 21497 12164 21503 12259
rect 21402 11550 21497 12164
rect 21822 11605 21921 12166
rect 21822 11500 21921 11506
rect 21402 11449 21497 11455
rect 20232 10494 20284 10500
rect 23541 10498 23587 16228
rect 23837 15576 23934 15591
rect 23837 15516 23854 15576
rect 23914 15516 23934 15576
rect 23837 15498 23934 15516
rect 25246 12277 25345 12283
rect 24781 12164 24787 12259
rect 24882 12164 24888 12259
rect 24787 11575 24882 12164
rect 25246 11605 25345 12178
rect 25719 11605 25818 11611
rect 25246 11506 25719 11605
rect 25719 11500 25818 11506
rect 24787 11474 24882 11480
rect 26945 10498 26991 16228
rect 27950 15588 28085 15608
rect 27950 15528 27974 15588
rect 28034 15528 28085 15588
rect 28460 15586 28515 18320
rect 29061 18306 29110 18320
rect 29339 17880 29408 18911
rect 29647 18420 29691 19026
rect 29620 18400 29720 18420
rect 29620 18340 29640 18400
rect 29700 18340 29720 18400
rect 29620 18320 29720 18340
rect 29647 18314 29691 18320
rect 28740 17860 28840 17880
rect 28740 17800 28760 17860
rect 28820 17800 28840 17860
rect 28740 17780 28840 17800
rect 29320 17860 29420 17880
rect 29320 17800 29340 17860
rect 29400 17800 29420 17860
rect 29320 17780 29420 17800
rect 28759 17570 28816 17780
rect 29339 17756 29408 17780
rect 28749 17510 28758 17570
rect 28818 17510 28827 17570
rect 30429 16302 30475 19288
rect 31704 17344 31760 19656
rect 31617 17288 31623 17344
rect 31679 17288 31760 17344
rect 30426 16296 30478 16302
rect 30426 16238 30478 16244
rect 27950 15514 28085 15528
rect 28458 15577 28518 15586
rect 28458 15508 28518 15517
rect 29926 15577 30013 15591
rect 29926 15517 29938 15577
rect 29998 15517 30013 15577
rect 29926 15504 30013 15517
rect 28634 12278 28733 12284
rect 28191 12164 28197 12259
rect 28292 12164 28298 12259
rect 28197 11560 28292 12164
rect 28634 11605 28733 12179
rect 28634 11500 28733 11506
rect 28197 11459 28292 11465
rect 16714 10488 16766 10494
rect 20232 10436 20284 10442
rect 23538 10492 23590 10498
rect 16714 10430 16766 10436
rect 15056 6521 15155 6527
rect 12664 6276 12716 6282
rect 12515 6186 12521 6238
rect 12573 6186 12579 6238
rect 12664 6218 12716 6224
rect 12396 6116 12448 6122
rect 12396 6058 12448 6064
rect 12217 6019 12269 6025
rect 12217 5961 12269 5967
rect 12060 5930 12112 5936
rect 12060 5872 12112 5878
rect 15056 5805 15155 6422
rect 15056 5700 15155 5706
rect 16717 6057 16763 10430
rect 17080 9796 17188 9810
rect 17080 9781 17107 9796
rect 17080 9721 17092 9781
rect 17167 9736 17188 9796
rect 17152 9721 17188 9736
rect 17080 9708 17188 9721
rect 18429 6499 18557 6515
rect 17970 6436 18098 6452
rect 17970 6341 17984 6436
rect 18079 6426 18098 6436
rect 18080 6346 18098 6426
rect 18429 6400 18440 6499
rect 18539 6400 18557 6499
rect 18429 6391 18557 6400
rect 18079 6341 18098 6346
rect 17970 6328 18098 6341
rect 20235 6057 20281 10436
rect 23538 10434 23590 10440
rect 26942 10492 26994 10498
rect 30429 10486 30475 16238
rect 31590 12184 31596 12279
rect 31691 12184 31697 12279
rect 31596 11579 31691 12184
rect 31596 11478 31691 11484
rect 26942 10434 26994 10440
rect 30426 10480 30478 10486
rect 21045 9807 21141 9820
rect 21045 9803 21063 9807
rect 21045 9743 21060 9803
rect 21123 9747 21141 9807
rect 21120 9743 21141 9747
rect 21045 9730 21141 9743
rect 21803 6514 21931 6524
rect 21803 6415 21817 6514
rect 21916 6415 21931 6514
rect 21803 6400 21931 6415
rect 23541 6057 23587 10434
rect 24367 9800 24503 9810
rect 24367 9735 24395 9800
rect 24460 9796 24503 9800
rect 24484 9736 24503 9796
rect 24460 9735 24503 9736
rect 24367 9716 24503 9735
rect 25211 6772 25217 6871
rect 25316 6772 25760 6871
rect 24321 6355 24791 6450
rect 24886 6355 24892 6450
rect 24321 6317 24416 6355
rect 25661 6326 25760 6772
rect 25661 6321 25962 6326
rect 25661 6232 25868 6321
rect 25957 6232 25966 6321
rect 25661 6227 25962 6232
rect 24321 6213 24416 6222
rect 26945 6057 26991 10434
rect 30426 10422 30478 10428
rect 27590 9803 27677 9823
rect 27590 9743 27600 9803
rect 27660 9743 27677 9803
rect 27590 9736 27677 9743
rect 30157 9794 30244 9807
rect 30157 9734 30169 9794
rect 30229 9734 30244 9794
rect 30157 9720 30244 9734
rect 28186 6360 28192 6455
rect 28287 6360 28331 6455
rect 28426 6360 28435 6455
rect 28612 6388 28736 6397
rect 28612 6289 28627 6388
rect 28726 6289 28736 6388
rect 28612 6278 28736 6289
rect 30429 6057 30475 10422
rect 31588 6385 31594 6480
rect 31689 6385 31695 6480
rect 16717 6011 30475 6057
rect 12042 5419 12102 5428
rect 12042 5350 12102 5359
rect 12051 348 12092 5350
rect 12172 4737 12232 4746
rect 16717 4688 16763 6011
rect 18440 5805 18539 5811
rect 17967 5771 18091 5780
rect 17967 5676 17984 5771
rect 18079 5676 18091 5771
rect 18431 5706 18440 5805
rect 18539 5706 18548 5805
rect 18440 5700 18539 5706
rect 17967 5666 18091 5676
rect 20235 4688 20281 6011
rect 21805 5805 21929 5819
rect 21397 5751 21509 5759
rect 21397 5656 21405 5751
rect 21500 5656 21509 5751
rect 21805 5706 21817 5805
rect 21916 5706 21929 5805
rect 21805 5692 21929 5706
rect 21397 5647 21509 5656
rect 23541 4692 23587 6011
rect 25863 5877 25962 5886
rect 25718 5805 25817 5811
rect 24321 5746 24781 5751
rect 24317 5661 24326 5746
rect 24411 5661 24781 5746
rect 24321 5656 24781 5661
rect 24876 5656 24882 5751
rect 25817 5778 25863 5805
rect 25817 5706 25962 5778
rect 25718 5700 25817 5706
rect 26943 4698 26989 6011
rect 28174 5895 28259 5899
rect 28169 5890 28264 5895
rect 28169 5805 28174 5890
rect 28259 5805 28264 5890
rect 28169 5330 28264 5805
rect 28627 5887 28726 5896
rect 28627 5700 28726 5706
rect 28169 5229 28264 5235
rect 30429 4702 30475 6011
rect 31594 5741 31689 6385
rect 31594 5640 31689 5646
rect 26940 4692 26992 4698
rect 12172 4668 12232 4677
rect 16714 4682 16766 4688
rect 12180 448 12224 4668
rect 16714 4624 16766 4630
rect 20232 4682 20284 4688
rect 20232 4624 20284 4630
rect 23538 4686 23590 4692
rect 26940 4634 26992 4640
rect 30426 4696 30478 4702
rect 30426 4638 30478 4644
rect 23538 4628 23590 4634
rect 17614 4006 17722 4033
rect 17614 3946 17631 4006
rect 17691 3946 17722 4006
rect 17614 3931 17722 3946
rect 20973 4006 21081 4032
rect 20973 3946 20992 4006
rect 21052 3946 21081 4006
rect 26515 4001 26623 4022
rect 20973 3930 21081 3946
rect 24472 3971 24580 3992
rect 24472 3906 24487 3971
rect 24552 3906 24580 3971
rect 26515 3941 26529 4001
rect 26589 3941 26623 4001
rect 26515 3920 26623 3941
rect 29889 3991 29997 4010
rect 29889 3931 29908 3991
rect 29968 3983 29997 3991
rect 29889 3923 29925 3931
rect 29985 3923 29997 3983
rect 29889 3908 29997 3923
rect 24472 3890 24580 3906
rect 17959 2492 18132 2507
rect 17959 2355 17974 2492
rect 18111 2355 18132 2492
rect 17959 2340 18132 2355
rect 21364 2492 21519 2500
rect 21364 2355 21372 2492
rect 21509 2355 21519 2492
rect 21364 2345 21519 2355
rect 24743 2492 24908 2506
rect 24743 2355 24757 2492
rect 24894 2355 24908 2492
rect 24743 2342 24908 2355
rect 28136 2492 28301 2507
rect 28136 2355 28152 2492
rect 28289 2355 28301 2492
rect 28136 2343 28301 2355
rect 12176 442 12228 448
rect 12176 384 12228 390
rect 12039 296 12045 348
rect 12097 296 12103 348
rect 11909 237 11915 289
rect 11967 237 11973 289
rect 30429 195 30475 4638
rect 31484 2492 31649 2502
rect 31484 2355 31501 2492
rect 31638 2355 31649 2492
rect 31484 2338 31649 2355
rect 30359 130 30368 195
rect 30536 130 30545 195
<< rmetal2 >>
rect 21391 6422 21519 6439
rect 21391 6326 21402 6422
rect 21500 6326 21519 6422
rect 21391 6315 21519 6326
<< via2 >>
rect 4322 44802 4378 44858
rect 28769 44800 28829 44860
rect 4453 44628 4509 44684
rect 18816 44626 18876 44686
rect 27650 44643 27710 44703
rect 27109 44559 27169 44619
rect 4627 44469 4683 44525
rect 18270 44467 18330 44527
rect 26555 44469 26615 44529
rect 4153 44334 4209 44390
rect 17720 44332 17780 44392
rect 25992 44379 26052 44439
rect 25456 44278 25516 44338
rect 4001 44183 4057 44239
rect 17162 44181 17222 44241
rect 24906 44186 24966 44246
rect 4801 44072 4857 44128
rect 16611 44070 16671 44130
rect 24344 44099 24404 44159
rect 3847 43947 3903 44003
rect 16056 43945 16116 44005
rect 23801 44004 23861 44064
rect 21028 43893 21088 43953
rect 3716 43823 3772 43879
rect 15508 43821 15568 43881
rect 20482 43801 20542 43861
rect 3560 43726 3616 43782
rect 14962 43725 15022 43785
rect 4948 43609 5004 43665
rect 14415 43608 14475 43668
rect 5079 43489 5135 43545
rect 13859 43487 13919 43547
rect 3423 43406 3479 43462
rect 3287 43287 3343 43343
rect 12762 43285 12822 43345
rect 13309 43330 13369 43390
rect 23474 19018 23534 19078
rect 23669 18911 23738 18980
rect 23854 18789 23914 18849
rect 24075 18702 24135 18762
rect 24256 18599 24316 18659
rect 24424 18506 24484 18566
rect 25440 18360 25480 18406
rect 25480 18360 25500 18406
rect 25440 18346 25500 18360
rect 26681 18360 26740 18398
rect 26740 18360 26741 18398
rect 13842 17823 14071 18052
rect 26681 18338 26741 18360
rect 25033 17989 25098 18054
rect 25252 17814 25312 17874
rect 24814 17643 24874 17703
rect 26975 17554 27035 17614
rect 26798 17391 26858 17451
rect 7140 12434 7200 12494
rect 8407 12315 8467 12362
rect 8407 12302 8411 12315
rect 8411 12302 8463 12315
rect 8463 12302 8467 12315
rect 4625 12206 4685 12266
rect 4151 11736 4211 11796
rect 3999 11605 4059 11665
rect 3558 11492 3618 11552
rect 3421 11182 3481 11242
rect 3285 11033 3345 11093
rect 3844 11432 3904 11492
rect 3743 11233 3803 11293
rect 4010 10120 4066 10176
rect 3665 7400 3721 7456
rect 8221 12110 8281 12170
rect 12146 12160 12206 12220
rect 7924 12007 7984 12067
rect 14861 12028 15052 12219
rect 11868 11474 11928 11534
rect 12660 10798 12720 10858
rect 12016 10113 12076 10173
rect 12518 9434 12578 9494
rect 4351 8760 4407 8816
rect 12392 8760 12452 8820
rect 12214 8078 12274 8138
rect 12056 7402 12116 7462
rect 11912 6717 11972 6777
rect 11787 6038 11847 6098
rect 17638 15556 17694 15612
rect 21008 15503 21067 15562
rect 23856 15518 23912 15574
rect 27976 15530 28032 15586
rect 28758 17510 28818 17570
rect 28458 15517 28518 15577
rect 29940 15519 29996 15575
rect 17094 9723 17150 9779
rect 17984 6341 18079 6436
rect 18445 6405 18534 6494
rect 21062 9745 21118 9801
rect 21405 6326 21500 6421
rect 21822 6420 21911 6509
rect 24426 9738 24482 9794
rect 24321 6222 24416 6317
rect 25868 6232 25957 6321
rect 27602 9745 27658 9801
rect 30171 9736 30227 9792
rect 28331 6360 28426 6455
rect 28632 6294 28721 6383
rect 12042 5359 12102 5419
rect 12172 4677 12232 4737
rect 17989 5681 18074 5766
rect 18440 5706 18539 5805
rect 21410 5661 21495 5746
rect 21817 5706 21916 5805
rect 24326 5661 24411 5746
rect 25863 5778 25962 5877
rect 28174 5805 28259 5890
rect 28627 5805 28726 5887
rect 28627 5788 28726 5805
rect 17633 3948 17689 4004
rect 20994 3948 21050 4004
rect 24491 3910 24547 3966
rect 26531 3943 26587 3999
rect 29927 3925 29983 3981
rect 17979 2360 18106 2487
rect 21377 2360 21504 2487
rect 24762 2360 24889 2487
rect 28157 2360 28284 2487
rect 31506 2360 31633 2487
rect 30368 130 30536 195
<< metal3 >>
rect 20480 45087 20544 45093
rect 17718 45067 17782 45073
rect 13307 45053 13371 45059
rect 12760 45042 12824 45048
rect 13307 44983 13371 44989
rect 13857 45054 13921 45060
rect 13857 44984 13921 44990
rect 14413 45055 14477 45061
rect 15506 45056 15570 45062
rect 14413 44985 14477 44991
rect 14960 45041 15024 45047
rect 12760 44972 12824 44978
rect 4317 44858 4383 44863
rect 4317 44802 4322 44858
rect 4378 44802 4383 44858
rect 4317 44797 4383 44802
rect 4148 44390 4214 44395
rect 4148 44334 4153 44390
rect 4209 44334 4214 44390
rect 4148 44329 4214 44334
rect 3996 44239 4062 44244
rect 3996 44183 4001 44239
rect 4057 44183 4062 44239
rect 3996 44178 4062 44183
rect 3842 44003 3908 44008
rect 3842 43947 3847 44003
rect 3903 43947 3908 44003
rect 3842 43942 3908 43947
rect 3711 43879 3777 43884
rect 3711 43823 3716 43879
rect 3772 43823 3777 43879
rect 3711 43818 3777 43823
rect 3555 43782 3621 43787
rect 3555 43726 3560 43782
rect 3616 43726 3621 43782
rect 3555 43721 3621 43726
rect 3418 43462 3484 43467
rect 3418 43406 3423 43462
rect 3479 43406 3484 43462
rect 3418 43401 3484 43406
rect 3282 43343 3348 43348
rect 3282 43287 3287 43343
rect 3343 43287 3348 43343
rect 3282 43282 3348 43287
rect 3285 11098 3345 43282
rect 3421 11247 3481 43401
rect 3557 11676 3619 43721
rect 3558 11557 3618 11676
rect 3553 11552 3623 11557
rect 3553 11492 3558 11552
rect 3618 11492 3623 11552
rect 3553 11487 3623 11492
rect 3714 11455 3774 43818
rect 3842 11649 3907 43942
rect 3999 11670 4059 44178
rect 4151 11801 4211 44329
rect 4146 11796 4216 11801
rect 4146 11736 4151 11796
rect 4211 11736 4216 11796
rect 4146 11731 4216 11736
rect 3994 11665 4064 11670
rect 3844 11497 3904 11649
rect 3994 11605 3999 11665
rect 4059 11605 4064 11665
rect 3994 11600 4064 11605
rect 3681 11395 3774 11455
rect 3839 11492 3909 11497
rect 3839 11432 3844 11492
rect 3904 11432 3909 11492
rect 3839 11427 3909 11432
rect 3681 11298 3741 11395
rect 3681 11293 3808 11298
rect 3416 11242 3486 11247
rect 3416 11182 3421 11242
rect 3481 11182 3486 11242
rect 3681 11233 3743 11293
rect 3803 11233 3808 11293
rect 3738 11228 3808 11233
rect 3416 11177 3486 11182
rect 3280 11093 3350 11098
rect 3280 11033 3285 11093
rect 3345 11033 3350 11093
rect 3280 11028 3350 11033
rect 4320 10798 4380 44797
rect 4448 44684 4514 44689
rect 4448 44628 4453 44684
rect 4509 44628 4514 44684
rect 4448 44623 4514 44628
rect 4451 12067 4511 44623
rect 4622 44525 4688 44530
rect 4622 44469 4627 44525
rect 4683 44469 4688 44525
rect 4622 44464 4688 44469
rect 4625 12271 4685 44464
rect 4796 44128 4862 44133
rect 4796 44072 4801 44128
rect 4857 44072 4862 44128
rect 4796 44067 4862 44072
rect 4620 12266 4690 12271
rect 4620 12206 4625 12266
rect 4685 12206 4690 12266
rect 4620 12201 4690 12206
rect 4799 12214 4859 44067
rect 4943 43665 5009 43670
rect 4943 43609 4948 43665
rect 5004 43609 5009 43665
rect 4943 43604 5009 43609
rect 4946 12362 5006 43604
rect 5074 43545 5140 43550
rect 5074 43489 5079 43545
rect 5135 43489 5140 43545
rect 5074 43484 5140 43489
rect 5077 12494 5137 43484
rect 12762 43350 12822 44972
rect 13309 43395 13369 44983
rect 13859 43552 13919 44984
rect 14415 43673 14475 44985
rect 15506 44986 15570 44992
rect 16054 45049 16118 45055
rect 14960 44971 15024 44977
rect 14962 43790 15022 44971
rect 15508 43886 15568 44986
rect 16054 44979 16118 44985
rect 16609 45046 16673 45052
rect 16056 44010 16116 44979
rect 16609 44976 16673 44982
rect 17160 45041 17224 45047
rect 18814 45061 18878 45067
rect 17718 44997 17782 45003
rect 18268 45041 18332 45047
rect 16611 44135 16671 44976
rect 17160 44971 17224 44977
rect 17162 44246 17222 44971
rect 17720 44397 17780 44997
rect 20480 45017 20544 45023
rect 21026 45087 21090 45093
rect 21026 45017 21090 45023
rect 23799 45083 23863 45089
rect 25990 45086 26054 45092
rect 18814 44991 18878 44997
rect 18268 44971 18332 44977
rect 18270 44532 18330 44971
rect 18816 44691 18876 44991
rect 18811 44686 18881 44691
rect 18811 44626 18816 44686
rect 18876 44626 18881 44686
rect 18811 44621 18881 44626
rect 18265 44527 18335 44532
rect 18265 44467 18270 44527
rect 18330 44467 18335 44527
rect 18265 44462 18335 44467
rect 17715 44392 17785 44397
rect 17715 44332 17720 44392
rect 17780 44332 17785 44392
rect 17715 44327 17785 44332
rect 17157 44241 17227 44246
rect 17157 44181 17162 44241
rect 17222 44181 17227 44241
rect 17157 44176 17227 44181
rect 16606 44130 16676 44135
rect 16606 44070 16611 44130
rect 16671 44070 16676 44130
rect 16606 44065 16676 44070
rect 16051 44005 16121 44010
rect 16051 43945 16056 44005
rect 16116 43945 16121 44005
rect 16051 43940 16121 43945
rect 15503 43881 15573 43886
rect 15503 43821 15508 43881
rect 15568 43821 15573 43881
rect 20482 43866 20542 45017
rect 21028 43958 21088 45017
rect 23799 45013 23863 45019
rect 24342 45070 24406 45076
rect 23801 44069 23861 45013
rect 24342 45000 24406 45006
rect 24904 45073 24968 45079
rect 24904 45003 24968 45009
rect 25454 45075 25518 45081
rect 27107 45065 27171 45071
rect 25990 45016 26054 45022
rect 26553 45059 26617 45065
rect 25454 45005 25518 45011
rect 24344 44164 24404 45000
rect 24906 44251 24966 45003
rect 25456 44343 25516 45005
rect 25992 44444 26052 45016
rect 27107 44995 27171 45001
rect 27648 45067 27712 45073
rect 27648 44997 27712 45003
rect 28767 45023 28831 45029
rect 26553 44989 26617 44995
rect 26555 44534 26615 44989
rect 27109 44624 27169 44995
rect 27650 44708 27710 44997
rect 28767 44953 28831 44959
rect 28769 44865 28829 44953
rect 28764 44860 28834 44865
rect 28764 44800 28769 44860
rect 28829 44800 28834 44860
rect 28764 44795 28834 44800
rect 27645 44703 27715 44708
rect 27645 44643 27650 44703
rect 27710 44643 27715 44703
rect 27645 44638 27715 44643
rect 27104 44619 27174 44624
rect 27104 44559 27109 44619
rect 27169 44559 27174 44619
rect 27104 44554 27174 44559
rect 26550 44529 26620 44534
rect 26550 44469 26555 44529
rect 26615 44469 26620 44529
rect 26550 44464 26620 44469
rect 25987 44439 26057 44444
rect 25987 44379 25992 44439
rect 26052 44379 26057 44439
rect 25987 44374 26057 44379
rect 25451 44338 25521 44343
rect 25451 44278 25456 44338
rect 25516 44278 25521 44338
rect 25451 44273 25521 44278
rect 24901 44246 24971 44251
rect 24901 44186 24906 44246
rect 24966 44186 24971 44246
rect 24901 44181 24971 44186
rect 24339 44159 24409 44164
rect 24339 44099 24344 44159
rect 24404 44099 24409 44159
rect 24339 44094 24409 44099
rect 23796 44064 23866 44069
rect 23796 44004 23801 44064
rect 23861 44004 23866 44064
rect 23796 43999 23866 44004
rect 21023 43953 21093 43958
rect 21023 43893 21028 43953
rect 21088 43893 21093 43953
rect 21023 43888 21093 43893
rect 15503 43816 15573 43821
rect 20477 43861 20547 43866
rect 20477 43801 20482 43861
rect 20542 43801 20547 43861
rect 20477 43796 20547 43801
rect 14957 43785 15027 43790
rect 14957 43725 14962 43785
rect 15022 43725 15027 43785
rect 14957 43720 15027 43725
rect 14410 43668 14480 43673
rect 14410 43608 14415 43668
rect 14475 43608 14480 43668
rect 14410 43603 14480 43608
rect 13854 43547 13924 43552
rect 13854 43487 13859 43547
rect 13919 43487 13924 43547
rect 13854 43482 13924 43487
rect 13304 43390 13374 43395
rect 12757 43345 12827 43350
rect 12757 43285 12762 43345
rect 12822 43285 12827 43345
rect 13304 43330 13309 43390
rect 13369 43330 13374 43390
rect 13304 43325 13374 43330
rect 12757 43280 12827 43285
rect 23469 19078 23539 19083
rect 23469 19018 23474 19078
rect 23534 19018 23539 19078
rect 23469 19013 23539 19018
rect 13837 18052 14076 18057
rect 13837 17823 13842 18052
rect 14071 17823 14076 18052
rect 7135 12494 7205 12499
rect 5077 12434 7140 12494
rect 7200 12434 7205 12494
rect 7135 12429 7205 12434
rect 8402 12362 8472 12367
rect 4946 12302 8407 12362
rect 8467 12302 8472 12362
rect 8402 12297 8472 12302
rect 12141 12220 12211 12225
rect 4799 12175 8281 12214
rect 4799 12170 8286 12175
rect 4799 12154 8221 12170
rect 8216 12110 8221 12154
rect 8281 12110 8286 12170
rect 12141 12160 12146 12220
rect 12206 12160 12211 12220
rect 12141 12155 12211 12160
rect 8216 12105 8286 12110
rect 7919 12067 7989 12072
rect 4451 12007 7924 12067
rect 7984 12007 7989 12067
rect 7919 12002 7989 12007
rect 11863 11534 11933 11539
rect 11863 11474 11868 11534
rect 11928 11474 11933 11534
rect 11863 11469 11933 11474
rect 12655 10858 12725 10863
rect 12655 10798 12660 10858
rect 12720 10798 12725 10858
rect 12655 10793 12725 10798
rect 4005 10178 4071 10181
rect 4005 10176 4494 10178
rect 4005 10120 4010 10176
rect 4066 10120 4494 10176
rect 4005 10118 4494 10120
rect 12011 10173 12081 10178
rect 4005 10115 4071 10118
rect 12011 10113 12016 10173
rect 12076 10113 12081 10173
rect 12011 10108 12081 10113
rect 12513 9494 12583 9499
rect 12513 9434 12518 9494
rect 12578 9434 12583 9494
rect 12513 9429 12583 9434
rect 4346 8816 4412 8821
rect 4346 8760 4351 8816
rect 4407 8760 4412 8816
rect 4346 8755 4412 8760
rect 12387 8820 12457 8825
rect 12387 8760 12392 8820
rect 12452 8760 12457 8820
rect 12387 8755 12457 8760
rect 12209 8138 12279 8143
rect 12209 8078 12214 8138
rect 12274 8078 12279 8138
rect 12209 8073 12279 8078
rect 12051 7462 12121 7467
rect 3660 7458 3726 7461
rect 4160 7458 4226 7461
rect 3660 7456 4411 7458
rect 3660 7400 3665 7456
rect 3721 7400 4411 7456
rect 3660 7398 4411 7400
rect 12051 7402 12056 7462
rect 12116 7402 12121 7462
rect 3660 7395 3726 7398
rect 4160 7395 4226 7398
rect 12051 7397 12121 7402
rect 11879 6777 12054 6811
rect 11879 6717 11912 6777
rect 11972 6717 12054 6777
rect 11879 6683 12039 6717
rect 11782 6098 11852 6103
rect 11782 6038 11787 6098
rect 11847 6038 11852 6098
rect 11782 6033 11852 6038
rect 12037 5419 12107 5424
rect 12037 5359 12042 5419
rect 12102 5359 12107 5419
rect 12037 5354 12107 5359
rect 12167 4737 12237 4742
rect 12167 4677 12172 4737
rect 12232 4677 12237 4737
rect 12167 4672 12237 4677
rect 13837 4340 14076 17823
rect 23474 15771 23534 19013
rect 23664 18980 23743 18985
rect 23664 18911 23669 18980
rect 23738 18911 23743 18980
rect 23664 18906 23743 18911
rect 17636 15711 23534 15771
rect 17636 15630 17696 15711
rect 17614 15612 17711 15630
rect 17614 15556 17638 15612
rect 17694 15556 17711 15612
rect 17614 15537 17711 15556
rect 20987 15567 21084 15579
rect 23669 15567 23738 18906
rect 23849 18849 23919 18854
rect 23849 18789 23854 18849
rect 23914 18789 23919 18849
rect 23849 18784 23919 18789
rect 23854 15591 23914 18784
rect 24070 18762 24140 18767
rect 24070 18702 24075 18762
rect 24135 18702 24140 18762
rect 24070 18697 24140 18702
rect 20987 15562 23738 15567
rect 20987 15503 21008 15562
rect 21067 15503 23738 15562
rect 20987 15498 23738 15503
rect 23837 15574 23934 15591
rect 23837 15518 23856 15574
rect 23912 15518 23934 15574
rect 23837 15498 23934 15518
rect 20987 15486 21084 15498
rect 14823 12224 15085 12245
rect 14823 12023 14856 12224
rect 15057 12023 15085 12224
rect 14823 11999 15085 12023
rect 24075 10308 24135 18697
rect 24251 18659 24321 18664
rect 24251 18599 24256 18659
rect 24316 18599 24321 18659
rect 24251 18594 24321 18599
rect 17092 10248 24135 10308
rect 17092 9784 17152 10248
rect 24256 10022 24316 18594
rect 24624 18577 26741 18637
rect 24419 18566 24489 18571
rect 24419 18506 24424 18566
rect 24484 18506 24489 18566
rect 24419 18501 24489 18506
rect 21060 9962 24316 10022
rect 21060 9806 21120 9962
rect 21057 9801 21123 9806
rect 17089 9779 17155 9784
rect 17089 9723 17094 9779
rect 17150 9723 17155 9779
rect 21057 9745 21062 9801
rect 21118 9745 21123 9801
rect 24424 9799 24484 18501
rect 21057 9740 21123 9745
rect 24421 9794 24487 9799
rect 24421 9738 24426 9794
rect 24482 9738 24487 9794
rect 24421 9733 24487 9738
rect 17089 9718 17155 9723
rect 21817 6509 21916 6514
rect 18440 6494 18539 6499
rect 17979 6436 18084 6441
rect 17979 6341 17984 6436
rect 18079 6341 18084 6436
rect 17979 6336 18084 6341
rect 18440 6405 18445 6494
rect 18534 6405 18539 6494
rect 17984 5766 18079 6336
rect 18440 5810 18539 6405
rect 21400 6421 21505 6426
rect 21400 6326 21405 6421
rect 21500 6326 21505 6421
rect 21400 6321 21505 6326
rect 21817 6420 21822 6509
rect 21911 6420 21916 6509
rect 17984 5681 17989 5766
rect 18074 5681 18079 5766
rect 18435 5805 18544 5810
rect 18435 5706 18440 5805
rect 18539 5706 18544 5805
rect 18435 5701 18544 5706
rect 21405 5746 21500 6321
rect 21817 5810 21916 6420
rect 24316 6317 24421 6322
rect 24316 6222 24321 6317
rect 24416 6222 24421 6317
rect 24316 6217 24421 6222
rect 17984 5676 18079 5681
rect 21405 5661 21410 5746
rect 21495 5661 21500 5746
rect 21812 5805 21921 5810
rect 21812 5706 21817 5805
rect 21916 5706 21921 5805
rect 21812 5701 21921 5706
rect 24321 5746 24416 6217
rect 21405 5656 21500 5661
rect 24321 5661 24326 5746
rect 24411 5661 24416 5746
rect 24321 5656 24416 5661
rect 24624 4597 24684 18577
rect 25435 18406 25505 18411
rect 25435 18346 25440 18406
rect 25500 18346 25505 18406
rect 26681 18403 26741 18577
rect 25435 18341 25505 18346
rect 26676 18398 26746 18403
rect 25028 18054 25103 18059
rect 25028 17989 25033 18054
rect 25098 17989 25103 18054
rect 25028 17984 25103 17989
rect 24809 17703 24879 17708
rect 24809 17643 24814 17703
rect 24874 17643 24879 17703
rect 24809 17638 24879 17643
rect 17631 4537 24684 4597
rect 13824 4330 14084 4340
rect 201 4320 599 4325
rect 7547 4320 7947 4326
rect 200 4319 7547 4320
rect 200 3921 201 4319
rect 599 4081 7547 4319
rect 13824 4093 13833 4330
rect 14080 4093 14084 4330
rect 13824 4086 14084 4093
rect 599 3921 7947 4081
rect 17631 4009 17691 4537
rect 24814 4248 24874 17638
rect 20992 4188 24874 4248
rect 20992 4009 21052 4188
rect 17628 4004 17694 4009
rect 17628 3948 17633 4004
rect 17689 3948 17694 4004
rect 17628 3943 17694 3948
rect 20989 4004 21055 4009
rect 20989 3948 20994 4004
rect 21050 3948 21055 4004
rect 20989 3943 21055 3948
rect 24486 3970 24552 3971
rect 25033 3970 25098 17984
rect 25247 17874 25317 17879
rect 25247 17814 25252 17874
rect 25312 17814 25317 17874
rect 25247 17809 25317 17814
rect 24486 3966 25098 3970
rect 200 3920 7947 3921
rect 201 3915 599 3920
rect 24486 3910 24491 3966
rect 24547 3910 25098 3966
rect 25252 4001 25312 17809
rect 25440 5661 25500 18341
rect 26676 18338 26681 18398
rect 26741 18338 26746 18398
rect 26676 18333 26746 18338
rect 26970 17614 27040 17619
rect 26970 17554 26975 17614
rect 27035 17554 27854 17614
rect 28753 17570 28823 17575
rect 26970 17549 27040 17554
rect 26793 17451 26863 17456
rect 26793 17391 26798 17451
rect 26858 17391 27660 17451
rect 26793 17386 26863 17391
rect 27600 9823 27660 17391
rect 27590 9801 27677 9823
rect 27590 9745 27602 9801
rect 27658 9745 27677 9801
rect 27590 9736 27677 9745
rect 27794 9794 27854 17554
rect 28062 17510 28758 17570
rect 28818 17510 28823 17570
rect 28062 15608 28122 17510
rect 28753 17505 28823 17510
rect 27950 15586 28122 15608
rect 27950 15530 27976 15586
rect 28032 15530 28122 15586
rect 27950 15528 28122 15530
rect 28453 15577 28523 15582
rect 29926 15577 30013 15591
rect 27950 15514 28085 15528
rect 28453 15517 28458 15577
rect 28518 15575 30013 15577
rect 28518 15519 29940 15575
rect 29996 15519 30013 15575
rect 28518 15517 30013 15519
rect 28453 15512 28523 15517
rect 29926 15504 30013 15517
rect 30157 9794 30244 9807
rect 27794 9792 30244 9794
rect 27794 9736 30171 9792
rect 30227 9736 30244 9792
rect 27794 9734 30244 9736
rect 30157 9720 30244 9734
rect 28326 6455 28431 6460
rect 28326 6360 28331 6455
rect 28426 6360 28431 6455
rect 28326 6355 28431 6360
rect 28612 6383 28736 6397
rect 25863 6321 25962 6326
rect 25863 6232 25868 6321
rect 25957 6232 25962 6321
rect 25863 5882 25962 6232
rect 28331 5895 28426 6355
rect 28612 6294 28632 6383
rect 28721 6294 28736 6383
rect 28612 6278 28736 6294
rect 28169 5890 28426 5895
rect 28627 5892 28726 6278
rect 25858 5877 25967 5882
rect 25858 5778 25863 5877
rect 25962 5778 25967 5877
rect 28169 5805 28174 5890
rect 28259 5805 28426 5890
rect 28169 5800 28426 5805
rect 28622 5887 28731 5892
rect 28622 5788 28627 5887
rect 28726 5788 28731 5887
rect 28622 5783 28731 5788
rect 25858 5773 25967 5778
rect 25440 5601 29985 5661
rect 26526 4001 26592 4004
rect 25252 3999 26592 4001
rect 25252 3943 26531 3999
rect 26587 3943 26592 3999
rect 29925 3986 29985 5601
rect 25252 3941 26592 3943
rect 26526 3938 26592 3941
rect 29922 3981 29988 3986
rect 29922 3925 29927 3981
rect 29983 3925 29988 3981
rect 29922 3920 29988 3925
rect 24486 3905 25098 3910
rect 17959 2492 18132 2507
rect 21364 2492 21519 2500
rect 17959 2491 31638 2492
rect 17957 2356 17963 2491
rect 18098 2487 31638 2491
rect 18106 2360 21377 2487
rect 21504 2360 24762 2487
rect 24889 2360 28157 2487
rect 28284 2360 31506 2487
rect 31633 2360 31638 2487
rect 18098 2356 31638 2360
rect 17959 2355 31638 2356
rect 17959 2340 18132 2355
rect 21364 2345 21519 2355
rect 30363 199 30541 200
rect 30357 126 30363 199
rect 30541 126 30547 199
rect 30363 125 30541 126
<< via3 >>
rect 12760 44978 12824 45042
rect 13307 44989 13371 45053
rect 13857 44990 13921 45054
rect 14413 44991 14477 45055
rect 14960 44977 15024 45041
rect 15506 44992 15570 45056
rect 16054 44985 16118 45049
rect 16609 44982 16673 45046
rect 17160 44977 17224 45041
rect 17718 45003 17782 45067
rect 18268 44977 18332 45041
rect 18814 44997 18878 45061
rect 20480 45023 20544 45087
rect 21026 45023 21090 45087
rect 23799 45019 23863 45083
rect 24342 45006 24406 45070
rect 24904 45009 24968 45073
rect 25454 45011 25518 45075
rect 25990 45022 26054 45086
rect 26553 44995 26617 45059
rect 27107 45001 27171 45065
rect 27648 45003 27712 45067
rect 28767 44959 28831 45023
rect 14856 12219 15057 12224
rect 14856 12028 14861 12219
rect 14861 12028 15052 12219
rect 15052 12028 15057 12219
rect 14856 12023 15057 12028
rect 201 3921 599 4319
rect 7547 4081 7947 4320
rect 13833 4093 14080 4330
rect 17963 2487 18098 2491
rect 17963 2360 17979 2487
rect 17979 2360 18098 2487
rect 17963 2356 18098 2360
rect 30363 195 30541 199
rect 30363 130 30368 195
rect 30368 130 30536 195
rect 30536 130 30541 195
rect 30363 126 30541 130
<< metal4 >>
rect 6134 44952 6194 45152
rect 6686 44952 6746 45152
rect 7238 44952 7298 45152
rect 7790 44952 7850 45152
rect 8342 44952 8402 45152
rect 8894 44952 8954 45152
rect 9446 44952 9506 45152
rect 9998 44952 10058 45152
rect 10550 44952 10610 45152
rect 11102 44952 11162 45152
rect 11654 44952 11714 45152
rect 12206 44952 12266 45152
rect 12758 45077 12818 45152
rect 12758 45042 12829 45077
rect 13310 45059 13370 45152
rect 13862 45093 13922 45152
rect 12758 44978 12760 45042
rect 12824 45011 12829 45042
rect 13291 45054 13370 45059
rect 13861 45055 13927 45093
rect 14414 45056 14474 45152
rect 13856 45054 13927 45055
rect 13291 45053 13372 45054
rect 12824 44978 12825 45011
rect 13291 44993 13307 45053
rect 13306 44989 13307 44993
rect 13371 44989 13372 45053
rect 13856 44990 13857 45054
rect 13921 45027 13927 45054
rect 14412 45055 14478 45056
rect 14966 45055 15026 45152
rect 15518 45057 15578 45152
rect 14412 45045 14413 45055
rect 13921 44990 13922 45027
rect 13856 44989 13922 44990
rect 13306 44988 13372 44989
rect 12758 44977 12825 44978
rect 12758 44952 12818 44977
rect 13310 44952 13370 44988
rect 13862 44952 13922 44989
rect 14399 44991 14413 45045
rect 14477 44991 14478 45055
rect 14399 44990 14478 44991
rect 14957 45041 15026 45055
rect 14399 44979 14474 44990
rect 14957 44989 14960 45041
rect 14414 44952 14474 44979
rect 14959 44977 14960 44989
rect 15024 44977 15026 45041
rect 15505 45056 15578 45057
rect 15505 45017 15506 45056
rect 14959 44976 15026 44977
rect 14966 44952 15026 44976
rect 15503 44992 15506 45017
rect 15570 44992 15578 45056
rect 16070 45051 16130 45152
rect 16059 45050 16130 45051
rect 15503 44952 15578 44992
rect 16053 45049 16130 45050
rect 16053 44985 16054 45049
rect 16118 44985 16130 45049
rect 16622 45047 16682 45152
rect 17174 45049 17234 45152
rect 17726 45068 17786 45152
rect 17717 45067 17786 45068
rect 17717 45049 17718 45067
rect 16608 45046 16682 45047
rect 16608 45017 16609 45046
rect 16053 44984 16130 44985
rect 16070 44952 16130 44984
rect 16605 44982 16609 45017
rect 16673 44982 16682 45046
rect 16605 44952 16682 44982
rect 17159 45041 17234 45049
rect 17159 44977 17160 45041
rect 17224 44977 17234 45041
rect 17707 45003 17718 45049
rect 17782 45003 17786 45067
rect 18278 45042 18338 45152
rect 18830 45062 18890 45152
rect 17707 44983 17786 45003
rect 17159 44976 17234 44977
rect 17174 44952 17234 44976
rect 17726 44952 17786 44983
rect 18267 45041 18338 45042
rect 18267 44977 18268 45041
rect 18332 44977 18338 45041
rect 18813 45061 18890 45062
rect 18813 44997 18814 45061
rect 18878 45029 18890 45061
rect 18878 44997 18891 45029
rect 18813 44996 18891 44997
rect 18267 44976 18338 44977
rect 18270 44967 18338 44976
rect 18278 44952 18338 44967
rect 18825 44963 18891 44996
rect 18830 44952 18890 44963
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 45088 20546 45152
rect 21038 45088 21098 45152
rect 20479 45087 20546 45088
rect 20479 45023 20480 45087
rect 20544 45023 20546 45087
rect 20479 45022 20546 45023
rect 21025 45087 21098 45088
rect 21025 45023 21026 45087
rect 21090 45023 21098 45087
rect 21025 45022 21098 45023
rect 20486 44952 20546 45022
rect 21038 44952 21098 45022
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 45084 23858 45152
rect 23798 45083 23864 45084
rect 23798 45019 23799 45083
rect 23863 45019 23864 45083
rect 24350 45071 24410 45152
rect 23798 45018 23864 45019
rect 24341 45070 24410 45071
rect 23798 44952 23858 45018
rect 24341 45006 24342 45070
rect 24406 45006 24410 45070
rect 24341 45005 24410 45006
rect 24350 44952 24410 45005
rect 24902 45074 24962 45152
rect 25454 45076 25514 45152
rect 26006 45087 26066 45152
rect 25989 45086 26066 45087
rect 25453 45075 25519 45076
rect 24902 45073 24969 45074
rect 24902 45009 24904 45073
rect 24968 45009 24969 45073
rect 25453 45011 25454 45075
rect 25518 45011 25519 45075
rect 25989 45022 25990 45086
rect 26054 45022 26066 45086
rect 26558 45060 26618 45152
rect 27110 45066 27170 45152
rect 27662 45068 27722 45152
rect 27647 45067 27722 45068
rect 25989 45021 26066 45022
rect 25453 45010 25519 45011
rect 24902 45008 24969 45009
rect 24902 44952 24962 45008
rect 25454 44952 25514 45010
rect 26006 44952 26066 45021
rect 26552 45059 26618 45060
rect 26552 44995 26553 45059
rect 26617 44995 26618 45059
rect 27106 45065 27172 45066
rect 27106 45001 27107 45065
rect 27171 45001 27172 45065
rect 27647 45003 27648 45067
rect 27712 45003 27722 45067
rect 27647 45002 27722 45003
rect 27106 45000 27172 45001
rect 26552 44994 26618 44995
rect 26558 44952 26618 44994
rect 27110 44952 27170 45000
rect 27662 44952 27722 45002
rect 28214 44952 28274 45152
rect 28766 45024 28826 45152
rect 28766 45023 28832 45024
rect 28766 44959 28767 45023
rect 28831 44959 28832 45023
rect 28766 44958 28832 44959
rect 28766 44952 28826 44958
rect 29318 44952 29378 45152
rect 15503 44951 15569 44952
rect 16605 44951 16671 44952
rect 200 4319 600 44152
rect 200 3921 201 4319
rect 599 3921 600 4319
rect 200 1000 600 3921
rect 800 12289 1200 44152
rect 1776 12289 2844 12290
rect 800 12224 15207 12289
rect 800 12023 14856 12224
rect 15057 12023 15207 12224
rect 800 11968 15207 12023
rect 800 1000 1200 11968
rect 1776 11954 2844 11968
rect 8268 11735 8589 11968
rect 7628 4572 7867 5027
rect 7628 4356 7866 4572
rect 7628 4331 7867 4356
rect 13824 4331 14084 4340
rect 7628 4330 18150 4331
rect 7628 4321 13833 4330
rect 7546 4320 13833 4321
rect 7546 4081 7547 4320
rect 7947 4093 13833 4320
rect 14080 4093 18150 4330
rect 7947 4092 18150 4093
rect 7947 4081 7948 4092
rect 13824 4086 14084 4092
rect 7546 4080 7948 4081
rect 17962 2491 18099 4092
rect 17962 2356 17963 2491
rect 18098 2356 18099 2491
rect 17962 2355 18099 2356
rect 3314 0 3494 204
rect 7178 0 7358 204
rect 11042 0 11222 204
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 199 30542 200
rect 30362 126 30363 199
rect 30541 126 30542 199
rect 30362 0 30542 126
use bit4_encoder  bit4_encoder_0 ~/Documents/github_project/adc_dac2/mag
timestamp 1730889744
transform 1 0 3400 0 1 2600
box 0 0 9409 11553
use compr2  compr2_0
timestamp 1730933686
transform 0 1 30003 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_1
timestamp 1730933686
transform 0 1 26603 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_2
timestamp 1730933686
transform 0 1 23203 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_3
timestamp 1730933686
transform 0 1 19803 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_4
timestamp 1730933686
transform 0 1 16403 -1 0 6375
box 510 -1403 5975 1713
use compr2  compr2_5
timestamp 1730933686
transform 0 1 30003 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_6
timestamp 1730933686
transform 0 1 26603 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_7
timestamp 1730933686
transform 0 1 23203 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_8
timestamp 1730933686
transform 0 1 19803 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_9
timestamp 1730933686
transform 0 1 16403 -1 0 12175
box 510 -1403 5975 1713
use compr2  compr2_10
timestamp 1730933686
transform 0 1 30003 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_11
timestamp 1730933686
transform 0 1 26603 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_12
timestamp 1730933686
transform 0 1 23203 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_13
timestamp 1730933686
transform 0 1 19803 -1 0 17975
box 510 -1403 5975 1713
use compr2  compr2_14
timestamp 1730933686
transform 0 1 16403 -1 0 17975
box 510 -1403 5975 1713
use pass_gate2  pass_gate2_0 ~/Documents/github_project/adc_dac2/mag
timestamp 1730933686
transform 1 0 21997 0 1 23096
box 2195 -3712 4186 290
use pass_gate2  pass_gate2_1
timestamp 1730933686
transform 1 0 24483 0 1 23096
box 2195 -3712 4186 290
use r2r_dac  r2r_dac_0 ~/Documents/github_project/adc_dac2/mag
timestamp 1730882523
transform 1 0 28000 0 1 25658
box 1000 -5458 3772 -192
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR1
timestamp 1730882523
transform 1 0 28049 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR2
timestamp 1730882523
transform 1 0 26273 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR3
timestamp 1730882523
transform 1 0 26865 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR4
timestamp 1730882523
transform 1 0 27753 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR5
timestamp 1730882523
transform 1 0 27457 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR6
timestamp 1730882523
transform 1 0 30417 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR7
timestamp 1730882523
transform 1 0 27161 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR8
timestamp 1730882523
transform 1 0 29529 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR9
timestamp 1730882523
transform 1 0 28345 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR10
timestamp 1730882523
transform 1 0 29233 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR11
timestamp 1730882523
transform 1 0 28641 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR12
timestamp 1730882523
transform 1 0 28937 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR13
timestamp 1730882523
transform 1 0 29825 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR14
timestamp 1730882523
transform 1 0 26569 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR15
timestamp 1730882523
transform 1 0 25977 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR16
timestamp 1730882523
transform 1 0 30121 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR17
timestamp 1730882523
transform 1 0 30713 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR18
timestamp 1730882523
transform 1 0 31305 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR19
timestamp 1730882523
transform 1 0 31009 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR20
timestamp 1730882523
transform 1 0 31601 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR21
timestamp 1730882523
transform 1 0 25681 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR22
timestamp 1730882523
transform 1 0 25385 0 1 18252
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR23
timestamp 1730882523
transform 1 0 31305 0 1 19450
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR24
timestamp 1730882523
transform 1 0 30121 0 1 19450
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR25
timestamp 1730882523
transform 1 0 30713 0 1 19450
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR26
timestamp 1730882523
transform 1 0 31009 0 1 19450
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR27
timestamp 1730882523
transform 1 0 30417 0 1 19450
box -201 -652 201 652
use sky130_fd_pr__res_xhigh_po_0p35_MGD972  XR28
timestamp 1730882523
transform 1 0 31601 0 1 19450
box -201 -652 201 652
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
