VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_tim2305_adc_dac
  CLASS BLOCK ;
  FOREIGN tt_um_tim2305_adc_dac ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 17.575 204.525 17.745 204.715 ;
        RECT 18.955 204.525 19.125 204.715 ;
        RECT 24.475 204.525 24.645 204.715 ;
        RECT 29.990 204.575 30.110 204.685 ;
        RECT 30.915 204.525 31.085 204.715 ;
        RECT 36.435 204.525 36.605 204.715 ;
        RECT 41.955 204.525 42.125 204.715 ;
        RECT 43.795 204.525 43.965 204.715 ;
        RECT 49.315 204.525 49.485 204.715 ;
        RECT 54.835 204.525 55.005 204.715 ;
        RECT 56.675 204.525 56.845 204.715 ;
        RECT 62.195 204.525 62.365 204.715 ;
        RECT 67.715 204.525 67.885 204.715 ;
        RECT 69.555 204.525 69.725 204.715 ;
        RECT 75.075 204.525 75.245 204.715 ;
        RECT 78.295 204.525 78.465 204.715 ;
        RECT 78.755 204.525 78.925 204.715 ;
        RECT 81.510 204.575 81.630 204.685 ;
        RECT 82.435 204.525 82.605 204.715 ;
        RECT 87.955 204.525 88.125 204.715 ;
        RECT 93.475 204.525 93.645 204.715 ;
        RECT 95.315 204.525 95.485 204.715 ;
        RECT 100.835 204.525 101.005 204.715 ;
        RECT 106.355 204.525 106.525 204.715 ;
        RECT 108.195 204.525 108.365 204.715 ;
        RECT 113.715 204.525 113.885 204.715 ;
        RECT 119.235 204.525 119.405 204.715 ;
        RECT 121.075 204.525 121.245 204.715 ;
        RECT 126.595 204.525 126.765 204.715 ;
        RECT 132.115 204.525 132.285 204.715 ;
        RECT 133.955 204.525 134.125 204.715 ;
        RECT 139.475 204.525 139.645 204.715 ;
        RECT 141.310 204.575 141.430 204.685 ;
        RECT 142.695 204.525 142.865 204.715 ;
        RECT 17.435 203.715 18.805 204.525 ;
        RECT 18.815 203.715 24.325 204.525 ;
        RECT 24.335 203.715 29.845 204.525 ;
        RECT 30.325 203.655 30.755 204.440 ;
        RECT 30.775 203.715 36.285 204.525 ;
        RECT 36.295 203.715 41.805 204.525 ;
        RECT 41.815 203.715 43.185 204.525 ;
        RECT 43.205 203.655 43.635 204.440 ;
        RECT 43.655 203.715 49.165 204.525 ;
        RECT 49.175 203.715 54.685 204.525 ;
        RECT 54.695 203.715 56.065 204.525 ;
        RECT 56.085 203.655 56.515 204.440 ;
        RECT 56.535 203.715 62.045 204.525 ;
        RECT 62.055 203.715 67.565 204.525 ;
        RECT 67.575 203.715 68.945 204.525 ;
        RECT 68.965 203.655 69.395 204.440 ;
        RECT 69.415 203.715 74.925 204.525 ;
        RECT 74.935 203.715 76.765 204.525 ;
        RECT 76.775 203.845 78.605 204.525 ;
        RECT 76.775 203.615 78.120 203.845 ;
        RECT 78.615 203.715 81.365 204.525 ;
        RECT 81.845 203.655 82.275 204.440 ;
        RECT 82.295 203.715 87.805 204.525 ;
        RECT 87.815 203.715 93.325 204.525 ;
        RECT 93.335 203.715 94.705 204.525 ;
        RECT 94.725 203.655 95.155 204.440 ;
        RECT 95.175 203.715 100.685 204.525 ;
        RECT 100.695 203.715 106.205 204.525 ;
        RECT 106.215 203.715 107.585 204.525 ;
        RECT 107.605 203.655 108.035 204.440 ;
        RECT 108.055 203.715 113.565 204.525 ;
        RECT 113.575 203.715 119.085 204.525 ;
        RECT 119.095 203.715 120.465 204.525 ;
        RECT 120.485 203.655 120.915 204.440 ;
        RECT 120.935 203.715 126.445 204.525 ;
        RECT 126.455 203.715 131.965 204.525 ;
        RECT 131.975 203.715 133.345 204.525 ;
        RECT 133.365 203.655 133.795 204.440 ;
        RECT 133.815 203.715 139.325 204.525 ;
        RECT 139.335 203.715 141.165 204.525 ;
        RECT 141.635 203.715 143.005 204.525 ;
      LAYER nwell ;
        RECT 17.240 200.495 143.200 203.325 ;
      LAYER pwell ;
        RECT 17.435 199.295 18.805 200.105 ;
        RECT 18.815 199.295 24.325 200.105 ;
        RECT 24.335 199.295 29.845 200.105 ;
        RECT 30.325 199.380 30.755 200.165 ;
        RECT 30.775 199.295 36.285 200.105 ;
        RECT 36.295 199.295 41.805 200.105 ;
        RECT 41.815 199.295 47.325 200.105 ;
        RECT 47.335 199.295 52.845 200.105 ;
        RECT 52.855 199.295 55.605 200.105 ;
        RECT 56.085 199.380 56.515 200.165 ;
        RECT 56.535 199.295 62.045 200.105 ;
        RECT 62.055 199.295 67.565 200.105 ;
        RECT 67.575 199.295 73.085 200.105 ;
        RECT 73.095 199.295 78.605 200.105 ;
        RECT 78.615 199.295 81.365 200.105 ;
        RECT 81.845 199.380 82.275 200.165 ;
        RECT 82.295 199.295 87.805 200.105 ;
        RECT 87.815 199.295 93.325 200.105 ;
        RECT 93.335 199.295 98.845 200.105 ;
        RECT 98.855 199.295 104.365 200.105 ;
        RECT 104.375 199.295 107.125 200.105 ;
        RECT 107.605 199.380 108.035 200.165 ;
        RECT 108.055 199.295 113.565 200.105 ;
        RECT 113.575 199.295 119.085 200.105 ;
        RECT 119.095 199.295 124.605 200.105 ;
        RECT 124.615 199.295 130.125 200.105 ;
        RECT 130.135 199.295 132.885 200.105 ;
        RECT 133.365 199.380 133.795 200.165 ;
        RECT 133.815 199.295 139.325 200.105 ;
        RECT 139.335 199.295 141.165 200.105 ;
        RECT 141.635 199.295 143.005 200.105 ;
        RECT 17.575 199.085 17.745 199.295 ;
        RECT 18.955 199.085 19.125 199.295 ;
        RECT 24.475 199.085 24.645 199.295 ;
        RECT 29.995 199.245 30.165 199.275 ;
        RECT 29.990 199.135 30.165 199.245 ;
        RECT 29.995 199.085 30.165 199.135 ;
        RECT 30.915 199.105 31.085 199.295 ;
        RECT 35.515 199.085 35.685 199.275 ;
        RECT 36.435 199.105 36.605 199.295 ;
        RECT 41.035 199.085 41.205 199.275 ;
        RECT 41.955 199.105 42.125 199.295 ;
        RECT 42.870 199.135 42.990 199.245 ;
        RECT 43.795 199.085 43.965 199.275 ;
        RECT 47.475 199.105 47.645 199.295 ;
        RECT 49.315 199.085 49.485 199.275 ;
        RECT 52.995 199.105 53.165 199.295 ;
        RECT 54.835 199.085 55.005 199.275 ;
        RECT 55.750 199.135 55.870 199.245 ;
        RECT 56.675 199.105 56.845 199.295 ;
        RECT 60.355 199.085 60.525 199.275 ;
        RECT 62.195 199.105 62.365 199.295 ;
        RECT 65.875 199.085 66.045 199.275 ;
        RECT 67.715 199.105 67.885 199.295 ;
        RECT 68.630 199.135 68.750 199.245 ;
        RECT 69.555 199.085 69.725 199.275 ;
        RECT 73.235 199.105 73.405 199.295 ;
        RECT 75.075 199.085 75.245 199.275 ;
        RECT 78.755 199.105 78.925 199.295 ;
        RECT 80.595 199.085 80.765 199.275 ;
        RECT 81.510 199.135 81.630 199.245 ;
        RECT 82.435 199.105 82.605 199.295 ;
        RECT 86.115 199.085 86.285 199.275 ;
        RECT 87.955 199.105 88.125 199.295 ;
        RECT 91.635 199.085 91.805 199.275 ;
        RECT 93.475 199.105 93.645 199.295 ;
        RECT 94.390 199.135 94.510 199.245 ;
        RECT 95.315 199.085 95.485 199.275 ;
        RECT 98.995 199.105 99.165 199.295 ;
        RECT 100.835 199.085 101.005 199.275 ;
        RECT 104.515 199.105 104.685 199.295 ;
        RECT 106.355 199.085 106.525 199.275 ;
        RECT 107.270 199.135 107.390 199.245 ;
        RECT 108.195 199.105 108.365 199.295 ;
        RECT 111.875 199.085 112.045 199.275 ;
        RECT 113.715 199.105 113.885 199.295 ;
        RECT 117.395 199.085 117.565 199.275 ;
        RECT 119.235 199.105 119.405 199.295 ;
        RECT 120.150 199.135 120.270 199.245 ;
        RECT 121.075 199.085 121.245 199.275 ;
        RECT 124.755 199.105 124.925 199.295 ;
        RECT 126.595 199.085 126.765 199.275 ;
        RECT 130.275 199.105 130.445 199.295 ;
        RECT 132.115 199.085 132.285 199.275 ;
        RECT 133.030 199.135 133.150 199.245 ;
        RECT 133.955 199.105 134.125 199.295 ;
        RECT 137.635 199.085 137.805 199.275 ;
        RECT 139.475 199.105 139.645 199.295 ;
        RECT 141.310 199.135 141.430 199.245 ;
        RECT 142.695 199.085 142.865 199.295 ;
        RECT 17.435 198.275 18.805 199.085 ;
        RECT 18.815 198.275 24.325 199.085 ;
        RECT 24.335 198.275 29.845 199.085 ;
        RECT 29.855 198.275 35.365 199.085 ;
        RECT 35.375 198.275 40.885 199.085 ;
        RECT 40.895 198.275 42.725 199.085 ;
        RECT 43.205 198.215 43.635 199.000 ;
        RECT 43.655 198.275 49.165 199.085 ;
        RECT 49.175 198.275 54.685 199.085 ;
        RECT 54.695 198.275 60.205 199.085 ;
        RECT 60.215 198.275 65.725 199.085 ;
        RECT 65.735 198.275 68.485 199.085 ;
        RECT 68.965 198.215 69.395 199.000 ;
        RECT 69.415 198.275 74.925 199.085 ;
        RECT 74.935 198.275 80.445 199.085 ;
        RECT 80.455 198.275 85.965 199.085 ;
        RECT 85.975 198.275 91.485 199.085 ;
        RECT 91.495 198.275 94.245 199.085 ;
        RECT 94.725 198.215 95.155 199.000 ;
        RECT 95.175 198.275 100.685 199.085 ;
        RECT 100.695 198.275 106.205 199.085 ;
        RECT 106.215 198.275 111.725 199.085 ;
        RECT 111.735 198.275 117.245 199.085 ;
        RECT 117.255 198.275 120.005 199.085 ;
        RECT 120.485 198.215 120.915 199.000 ;
        RECT 120.935 198.275 126.445 199.085 ;
        RECT 126.455 198.275 131.965 199.085 ;
        RECT 131.975 198.275 137.485 199.085 ;
        RECT 137.495 198.275 141.165 199.085 ;
        RECT 141.635 198.275 143.005 199.085 ;
      LAYER nwell ;
        RECT 17.240 195.055 143.200 197.885 ;
      LAYER pwell ;
        RECT 17.435 193.855 18.805 194.665 ;
        RECT 18.815 193.855 24.325 194.665 ;
        RECT 24.335 193.855 29.845 194.665 ;
        RECT 30.325 193.940 30.755 194.725 ;
        RECT 30.775 193.855 36.285 194.665 ;
        RECT 36.295 193.855 41.805 194.665 ;
        RECT 41.815 193.855 47.325 194.665 ;
        RECT 47.335 193.855 52.845 194.665 ;
        RECT 52.855 193.855 55.605 194.665 ;
        RECT 56.085 193.940 56.515 194.725 ;
        RECT 56.535 193.855 62.045 194.665 ;
        RECT 62.055 193.855 67.565 194.665 ;
        RECT 67.575 193.855 73.085 194.665 ;
        RECT 73.095 193.855 78.605 194.665 ;
        RECT 78.615 193.855 81.365 194.665 ;
        RECT 81.845 193.940 82.275 194.725 ;
        RECT 82.295 193.855 87.805 194.665 ;
        RECT 87.815 193.855 93.325 194.665 ;
        RECT 93.335 193.855 98.845 194.665 ;
        RECT 98.855 193.855 104.365 194.665 ;
        RECT 104.375 193.855 107.125 194.665 ;
        RECT 107.605 193.940 108.035 194.725 ;
        RECT 108.055 193.855 113.565 194.665 ;
        RECT 113.575 193.855 119.085 194.665 ;
        RECT 119.095 193.855 124.605 194.665 ;
        RECT 124.615 193.855 130.125 194.665 ;
        RECT 130.135 193.855 132.885 194.665 ;
        RECT 133.365 193.940 133.795 194.725 ;
        RECT 133.815 193.855 139.325 194.665 ;
        RECT 139.335 193.855 141.165 194.665 ;
        RECT 141.635 193.855 143.005 194.665 ;
        RECT 17.575 193.645 17.745 193.855 ;
        RECT 18.955 193.645 19.125 193.855 ;
        RECT 24.475 193.645 24.645 193.855 ;
        RECT 29.995 193.805 30.165 193.835 ;
        RECT 29.990 193.695 30.165 193.805 ;
        RECT 29.995 193.645 30.165 193.695 ;
        RECT 30.915 193.665 31.085 193.855 ;
        RECT 35.515 193.645 35.685 193.835 ;
        RECT 36.435 193.665 36.605 193.855 ;
        RECT 41.035 193.645 41.205 193.835 ;
        RECT 41.955 193.665 42.125 193.855 ;
        RECT 42.870 193.695 42.990 193.805 ;
        RECT 43.795 193.645 43.965 193.835 ;
        RECT 47.475 193.665 47.645 193.855 ;
        RECT 49.315 193.645 49.485 193.835 ;
        RECT 52.995 193.665 53.165 193.855 ;
        RECT 54.835 193.645 55.005 193.835 ;
        RECT 55.750 193.695 55.870 193.805 ;
        RECT 56.675 193.665 56.845 193.855 ;
        RECT 60.355 193.645 60.525 193.835 ;
        RECT 62.195 193.665 62.365 193.855 ;
        RECT 65.875 193.645 66.045 193.835 ;
        RECT 67.715 193.665 67.885 193.855 ;
        RECT 68.175 193.645 68.345 193.835 ;
        RECT 68.630 193.695 68.750 193.805 ;
        RECT 70.475 193.645 70.645 193.835 ;
        RECT 70.935 193.645 71.105 193.835 ;
        RECT 73.235 193.665 73.405 193.855 ;
        RECT 78.755 193.665 78.925 193.855 ;
        RECT 81.515 193.805 81.685 193.835 ;
        RECT 81.510 193.695 81.685 193.805 ;
        RECT 81.515 193.645 81.685 193.695 ;
        RECT 82.435 193.665 82.605 193.855 ;
        RECT 84.275 193.645 84.445 193.835 ;
        RECT 84.735 193.645 84.905 193.835 ;
        RECT 87.955 193.665 88.125 193.855 ;
        RECT 90.255 193.645 90.425 193.835 ;
        RECT 93.475 193.665 93.645 193.855 ;
        RECT 93.945 193.690 94.105 193.800 ;
        RECT 95.315 193.645 95.485 193.835 ;
        RECT 98.995 193.665 99.165 193.855 ;
        RECT 100.835 193.645 101.005 193.835 ;
        RECT 104.515 193.665 104.685 193.855 ;
        RECT 106.355 193.645 106.525 193.835 ;
        RECT 107.270 193.695 107.390 193.805 ;
        RECT 108.195 193.665 108.365 193.855 ;
        RECT 111.875 193.645 112.045 193.835 ;
        RECT 113.715 193.665 113.885 193.855 ;
        RECT 118.775 193.645 118.945 193.835 ;
        RECT 119.235 193.645 119.405 193.855 ;
        RECT 121.075 193.645 121.245 193.835 ;
        RECT 124.755 193.665 124.925 193.855 ;
        RECT 126.595 193.645 126.765 193.835 ;
        RECT 130.275 193.665 130.445 193.855 ;
        RECT 132.115 193.645 132.285 193.835 ;
        RECT 133.030 193.695 133.150 193.805 ;
        RECT 133.955 193.665 134.125 193.855 ;
        RECT 137.635 193.645 137.805 193.835 ;
        RECT 139.475 193.665 139.645 193.855 ;
        RECT 141.310 193.695 141.430 193.805 ;
        RECT 142.695 193.645 142.865 193.855 ;
        RECT 17.435 192.835 18.805 193.645 ;
        RECT 18.815 192.835 24.325 193.645 ;
        RECT 24.335 192.835 29.845 193.645 ;
        RECT 29.855 192.835 35.365 193.645 ;
        RECT 35.375 192.835 40.885 193.645 ;
        RECT 40.895 192.835 42.725 193.645 ;
        RECT 43.205 192.775 43.635 193.560 ;
        RECT 43.655 192.835 49.165 193.645 ;
        RECT 49.175 192.835 54.685 193.645 ;
        RECT 54.695 192.835 60.205 193.645 ;
        RECT 60.215 192.835 65.725 193.645 ;
        RECT 65.735 192.835 67.105 193.645 ;
        RECT 67.115 192.865 68.485 193.645 ;
        RECT 68.965 192.775 69.395 193.560 ;
        RECT 69.425 192.735 70.775 193.645 ;
        RECT 70.795 192.965 78.105 193.645 ;
        RECT 74.310 192.745 75.220 192.965 ;
        RECT 76.755 192.735 78.105 192.965 ;
        RECT 78.250 192.965 81.715 193.645 ;
        RECT 81.845 192.965 84.585 193.645 ;
        RECT 78.250 192.735 79.170 192.965 ;
        RECT 84.595 192.835 90.105 193.645 ;
        RECT 90.115 192.835 93.785 193.645 ;
        RECT 94.725 192.775 95.155 193.560 ;
        RECT 95.175 192.835 100.685 193.645 ;
        RECT 100.695 192.835 106.205 193.645 ;
        RECT 106.215 192.835 111.725 193.645 ;
        RECT 111.735 192.835 117.245 193.645 ;
        RECT 117.255 192.965 119.085 193.645 ;
        RECT 117.255 192.735 118.600 192.965 ;
        RECT 119.095 192.835 120.465 193.645 ;
        RECT 120.485 192.775 120.915 193.560 ;
        RECT 120.935 192.835 126.445 193.645 ;
        RECT 126.455 192.835 131.965 193.645 ;
        RECT 131.975 192.835 137.485 193.645 ;
        RECT 137.495 192.835 141.165 193.645 ;
        RECT 141.635 192.835 143.005 193.645 ;
      LAYER nwell ;
        RECT 17.240 189.615 143.200 192.445 ;
      LAYER pwell ;
        RECT 17.435 188.415 18.805 189.225 ;
        RECT 18.815 188.415 24.325 189.225 ;
        RECT 24.335 188.415 29.845 189.225 ;
        RECT 30.325 188.500 30.755 189.285 ;
        RECT 30.775 188.415 36.285 189.225 ;
        RECT 36.295 188.415 41.805 189.225 ;
        RECT 41.815 188.415 47.325 189.225 ;
        RECT 47.335 188.415 52.845 189.225 ;
        RECT 52.855 188.415 55.605 189.225 ;
        RECT 56.085 188.500 56.515 189.285 ;
        RECT 56.535 188.415 62.045 189.225 ;
        RECT 62.055 188.415 64.805 189.225 ;
        RECT 65.370 189.095 66.290 189.325 ;
        RECT 65.370 188.415 68.835 189.095 ;
        RECT 69.895 188.415 71.245 189.325 ;
        RECT 71.355 188.415 74.465 189.325 ;
        RECT 77.990 189.095 78.900 189.315 ;
        RECT 80.435 189.095 81.785 189.325 ;
        RECT 74.475 188.415 81.785 189.095 ;
        RECT 81.845 188.500 82.275 189.285 ;
        RECT 83.345 189.095 84.275 189.325 ;
        RECT 82.440 188.415 84.275 189.095 ;
        RECT 84.595 188.415 90.105 189.225 ;
        RECT 90.115 188.415 92.865 189.225 ;
        RECT 93.355 188.415 94.705 189.325 ;
        RECT 95.675 189.095 97.025 189.325 ;
        RECT 98.560 189.095 99.470 189.315 ;
        RECT 95.675 188.415 102.985 189.095 ;
        RECT 102.995 188.415 105.285 189.325 ;
        RECT 105.295 188.415 107.125 189.325 ;
        RECT 107.605 188.500 108.035 189.285 ;
        RECT 108.055 188.415 111.725 189.225 ;
        RECT 112.695 189.095 114.045 189.325 ;
        RECT 115.580 189.095 116.490 189.315 ;
        RECT 120.055 189.095 121.405 189.325 ;
        RECT 122.940 189.095 123.850 189.315 ;
        RECT 112.695 188.415 120.005 189.095 ;
        RECT 120.055 188.415 127.365 189.095 ;
        RECT 127.375 188.415 132.885 189.225 ;
        RECT 133.365 188.500 133.795 189.285 ;
        RECT 133.815 188.415 139.325 189.225 ;
        RECT 139.335 188.415 141.165 189.225 ;
        RECT 141.635 188.415 143.005 189.225 ;
        RECT 17.575 188.205 17.745 188.415 ;
        RECT 18.955 188.205 19.125 188.415 ;
        RECT 24.475 188.205 24.645 188.415 ;
        RECT 29.995 188.365 30.165 188.395 ;
        RECT 29.990 188.255 30.165 188.365 ;
        RECT 29.995 188.205 30.165 188.255 ;
        RECT 30.915 188.225 31.085 188.415 ;
        RECT 35.525 188.250 35.685 188.360 ;
        RECT 36.435 188.205 36.605 188.415 ;
        RECT 40.115 188.205 40.285 188.395 ;
        RECT 41.955 188.225 42.125 188.415 ;
        RECT 42.870 188.255 42.990 188.365 ;
        RECT 43.795 188.205 43.965 188.395 ;
        RECT 47.475 188.225 47.645 188.415 ;
        RECT 49.315 188.205 49.485 188.395 ;
        RECT 52.995 188.225 53.165 188.415 ;
        RECT 55.750 188.255 55.870 188.365 ;
        RECT 56.215 188.205 56.385 188.395 ;
        RECT 56.675 188.205 56.845 188.415 ;
        RECT 58.510 188.255 58.630 188.365 ;
        RECT 62.195 188.225 62.365 188.415 ;
        RECT 64.950 188.255 65.070 188.365 ;
        RECT 65.875 188.205 66.045 188.395 ;
        RECT 66.335 188.205 66.505 188.395 ;
        RECT 68.635 188.225 68.805 188.415 ;
        RECT 69.105 188.260 69.265 188.370 ;
        RECT 69.555 188.205 69.725 188.395 ;
        RECT 70.930 188.225 71.100 188.415 ;
        RECT 71.395 188.225 71.565 188.415 ;
        RECT 74.615 188.225 74.785 188.415 ;
        RECT 82.440 188.395 82.605 188.415 ;
        RECT 76.920 188.205 77.090 188.395 ;
        RECT 82.435 188.225 82.605 188.395 ;
        RECT 83.815 188.205 83.985 188.395 ;
        RECT 84.270 188.255 84.390 188.365 ;
        RECT 84.735 188.225 84.905 188.415 ;
        RECT 85.650 188.205 85.820 188.395 ;
        RECT 86.115 188.205 86.285 188.395 ;
        RECT 89.790 188.255 89.910 188.365 ;
        RECT 90.255 188.225 90.425 188.415 ;
        RECT 93.010 188.255 93.130 188.365 ;
        RECT 93.475 188.205 93.645 188.395 ;
        RECT 93.945 188.250 94.105 188.360 ;
        RECT 94.390 188.225 94.560 188.415 ;
        RECT 94.865 188.260 95.025 188.370 ;
        RECT 102.215 188.205 102.385 188.395 ;
        RECT 102.675 188.205 102.845 188.415 ;
        RECT 103.135 188.225 103.305 188.415 ;
        RECT 105.440 188.225 105.610 188.415 ;
        RECT 107.275 188.365 107.445 188.395 ;
        RECT 106.365 188.250 106.525 188.360 ;
        RECT 107.270 188.255 107.445 188.365 ;
        RECT 107.275 188.205 107.445 188.255 ;
        RECT 108.195 188.225 108.365 188.415 ;
        RECT 111.885 188.260 112.045 188.370 ;
        RECT 114.630 188.255 114.750 188.365 ;
        RECT 118.500 188.205 118.670 188.395 ;
        RECT 119.235 188.205 119.405 188.395 ;
        RECT 119.695 188.225 119.865 188.415 ;
        RECT 121.075 188.205 121.245 188.395 ;
        RECT 126.595 188.205 126.765 188.395 ;
        RECT 127.055 188.225 127.225 188.415 ;
        RECT 127.515 188.225 127.685 188.415 ;
        RECT 132.115 188.205 132.285 188.395 ;
        RECT 133.030 188.255 133.150 188.365 ;
        RECT 133.955 188.225 134.125 188.415 ;
        RECT 137.635 188.205 137.805 188.395 ;
        RECT 139.475 188.225 139.645 188.415 ;
        RECT 141.310 188.255 141.430 188.365 ;
        RECT 142.695 188.205 142.865 188.415 ;
        RECT 17.435 187.395 18.805 188.205 ;
        RECT 18.815 187.395 24.325 188.205 ;
        RECT 24.335 187.395 29.845 188.205 ;
        RECT 29.855 187.395 35.365 188.205 ;
        RECT 36.295 187.525 39.965 188.205 ;
        RECT 39.035 187.295 39.965 187.525 ;
        RECT 39.975 187.395 42.725 188.205 ;
        RECT 43.205 187.335 43.635 188.120 ;
        RECT 43.655 187.395 49.165 188.205 ;
        RECT 49.175 187.395 54.685 188.205 ;
        RECT 54.695 187.525 56.525 188.205 ;
        RECT 56.535 187.395 58.365 188.205 ;
        RECT 58.875 187.525 66.185 188.205 ;
        RECT 58.875 187.295 60.225 187.525 ;
        RECT 61.760 187.305 62.670 187.525 ;
        RECT 66.195 187.295 68.915 188.205 ;
        RECT 68.965 187.335 69.395 188.120 ;
        RECT 69.415 187.525 76.725 188.205 ;
        RECT 72.930 187.305 73.840 187.525 ;
        RECT 75.375 187.295 76.725 187.525 ;
        RECT 76.775 187.525 80.360 188.205 ;
        RECT 80.550 187.525 84.015 188.205 ;
        RECT 76.775 187.295 77.695 187.525 ;
        RECT 80.550 187.295 81.470 187.525 ;
        RECT 84.615 187.295 85.965 188.205 ;
        RECT 85.975 187.395 89.645 188.205 ;
        RECT 90.210 187.525 93.675 188.205 ;
        RECT 90.210 187.295 91.130 187.525 ;
        RECT 94.725 187.335 95.155 188.120 ;
        RECT 95.215 187.525 102.525 188.205 ;
        RECT 102.645 187.525 106.110 188.205 ;
        RECT 107.135 187.525 114.445 188.205 ;
        RECT 115.185 187.525 119.085 188.205 ;
        RECT 95.215 187.295 96.565 187.525 ;
        RECT 98.100 187.305 99.010 187.525 ;
        RECT 105.190 187.295 106.110 187.525 ;
        RECT 110.650 187.305 111.560 187.525 ;
        RECT 113.095 187.295 114.445 187.525 ;
        RECT 118.155 187.295 119.085 187.525 ;
        RECT 119.095 187.395 120.465 188.205 ;
        RECT 120.485 187.335 120.915 188.120 ;
        RECT 120.935 187.395 126.445 188.205 ;
        RECT 126.455 187.395 131.965 188.205 ;
        RECT 131.975 187.395 137.485 188.205 ;
        RECT 137.495 187.395 141.165 188.205 ;
        RECT 141.635 187.395 143.005 188.205 ;
      LAYER nwell ;
        RECT 17.240 184.175 143.200 187.005 ;
      LAYER pwell ;
        RECT 17.435 182.975 18.805 183.785 ;
        RECT 18.815 182.975 22.485 183.785 ;
        RECT 26.470 183.655 27.380 183.875 ;
        RECT 28.915 183.655 30.265 183.885 ;
        RECT 22.955 182.975 30.265 183.655 ;
        RECT 30.325 183.060 30.755 183.845 ;
        RECT 30.775 182.975 32.605 183.785 ;
        RECT 35.815 183.655 36.745 183.885 ;
        RECT 40.270 183.655 41.180 183.875 ;
        RECT 42.715 183.655 44.065 183.885 ;
        RECT 33.075 182.975 36.745 183.655 ;
        RECT 36.755 182.975 44.065 183.655 ;
        RECT 44.115 182.975 47.785 183.785 ;
        RECT 51.310 183.655 52.220 183.875 ;
        RECT 53.755 183.655 55.105 183.885 ;
        RECT 47.795 182.975 55.105 183.655 ;
        RECT 56.085 183.060 56.515 183.845 ;
        RECT 60.050 183.655 60.960 183.875 ;
        RECT 62.495 183.655 63.845 183.885 ;
        RECT 56.535 182.975 63.845 183.655 ;
        RECT 64.355 183.655 65.275 183.885 ;
        RECT 64.355 182.975 67.940 183.655 ;
        RECT 68.055 182.975 69.405 183.885 ;
        RECT 72.070 183.655 72.990 183.885 ;
        RECT 69.525 182.975 72.990 183.655 ;
        RECT 73.105 182.975 76.765 183.885 ;
        RECT 76.775 182.975 78.145 183.785 ;
        RECT 79.490 183.685 80.445 183.885 ;
        RECT 78.165 183.005 80.445 183.685 ;
        RECT 17.575 182.765 17.745 182.975 ;
        RECT 18.955 182.765 19.125 182.975 ;
        RECT 22.630 182.815 22.750 182.925 ;
        RECT 23.095 182.785 23.265 182.975 ;
        RECT 27.695 182.765 27.865 182.955 ;
        RECT 30.915 182.765 31.085 182.975 ;
        RECT 31.375 182.765 31.545 182.955 ;
        RECT 32.755 182.925 32.925 182.955 ;
        RECT 32.750 182.815 32.925 182.925 ;
        RECT 32.755 182.765 32.925 182.815 ;
        RECT 33.215 182.785 33.385 182.975 ;
        RECT 35.055 182.765 35.225 182.955 ;
        RECT 36.895 182.785 37.065 182.975 ;
        RECT 42.425 182.810 42.585 182.920 ;
        RECT 43.795 182.765 43.965 182.955 ;
        RECT 44.255 182.785 44.425 182.975 ;
        RECT 47.935 182.785 48.105 182.975 ;
        RECT 50.235 182.765 50.405 182.955 ;
        RECT 50.695 182.765 50.865 182.955 ;
        RECT 55.305 182.820 55.465 182.930 ;
        RECT 55.755 182.765 55.925 182.955 ;
        RECT 56.215 182.765 56.385 182.955 ;
        RECT 56.675 182.785 56.845 182.975 ;
        RECT 61.735 182.765 61.905 182.955 ;
        RECT 64.030 182.815 64.150 182.925 ;
        RECT 64.500 182.785 64.670 182.975 ;
        RECT 67.250 182.815 67.370 182.925 ;
        RECT 68.170 182.785 68.340 182.975 ;
        RECT 68.635 182.765 68.805 182.955 ;
        RECT 69.555 182.785 69.725 182.975 ;
        RECT 17.435 181.955 18.805 182.765 ;
        RECT 18.815 181.955 24.325 182.765 ;
        RECT 24.335 182.085 28.005 182.765 ;
        RECT 24.335 181.855 25.265 182.085 ;
        RECT 28.015 181.855 31.185 182.765 ;
        RECT 31.235 181.955 32.605 182.765 ;
        RECT 32.615 182.085 34.905 182.765 ;
        RECT 34.915 182.085 42.225 182.765 ;
        RECT 33.985 181.855 34.905 182.085 ;
        RECT 38.430 181.865 39.340 182.085 ;
        RECT 40.875 181.855 42.225 182.085 ;
        RECT 43.205 181.895 43.635 182.680 ;
        RECT 43.695 181.855 46.865 182.765 ;
        RECT 46.875 182.085 50.545 182.765 ;
        RECT 46.875 181.855 47.805 182.085 ;
        RECT 50.555 181.955 54.225 182.765 ;
        RECT 54.235 181.855 56.050 182.765 ;
        RECT 56.075 181.955 61.585 182.765 ;
        RECT 61.595 181.955 67.105 182.765 ;
        RECT 67.585 181.855 68.935 182.765 ;
        RECT 69.415 182.735 70.370 182.765 ;
        RECT 71.400 182.735 71.570 182.955 ;
        RECT 71.855 182.785 72.025 182.955 ;
        RECT 73.230 182.785 73.400 182.975 ;
        RECT 71.860 182.765 72.025 182.785 ;
        RECT 74.155 182.765 74.325 182.955 ;
        RECT 76.915 182.785 77.085 182.975 ;
        RECT 78.290 182.785 78.460 183.005 ;
        RECT 79.490 182.975 80.445 183.005 ;
        RECT 80.455 182.975 81.805 183.885 ;
        RECT 81.845 183.060 82.275 183.845 ;
        RECT 83.255 183.655 84.605 183.885 ;
        RECT 86.140 183.655 87.050 183.875 ;
        RECT 93.230 183.655 94.150 183.885 ;
        RECT 97.770 183.655 98.680 183.875 ;
        RECT 100.215 183.655 101.565 183.885 ;
        RECT 83.255 182.975 90.565 183.655 ;
        RECT 90.685 182.975 94.150 183.655 ;
        RECT 94.255 182.975 101.565 183.655 ;
        RECT 101.710 183.655 102.630 183.885 ;
        RECT 106.630 183.685 107.585 183.885 ;
        RECT 101.710 182.975 105.175 183.655 ;
        RECT 105.305 183.005 107.585 183.685 ;
        RECT 107.605 183.060 108.035 183.845 ;
        RECT 79.675 182.765 79.845 182.955 ;
        RECT 81.520 182.785 81.690 182.975 ;
        RECT 82.445 182.820 82.605 182.930 ;
        RECT 87.035 182.765 87.205 182.955 ;
        RECT 90.255 182.785 90.425 182.975 ;
        RECT 90.715 182.955 90.885 182.975 ;
        RECT 90.715 182.785 90.890 182.955 ;
        RECT 94.395 182.925 94.565 182.975 ;
        RECT 94.390 182.815 94.565 182.925 ;
        RECT 95.310 182.815 95.430 182.925 ;
        RECT 94.395 182.785 94.565 182.815 ;
        RECT 90.720 182.765 90.890 182.785 ;
        RECT 95.775 182.765 95.945 182.955 ;
        RECT 68.965 181.895 69.395 182.680 ;
        RECT 69.415 182.055 71.695 182.735 ;
        RECT 71.860 182.085 73.695 182.765 ;
        RECT 69.415 181.855 70.370 182.055 ;
        RECT 72.765 181.855 73.695 182.085 ;
        RECT 74.015 181.955 79.525 182.765 ;
        RECT 79.535 182.085 86.845 182.765 ;
        RECT 83.050 181.865 83.960 182.085 ;
        RECT 85.495 181.855 86.845 182.085 ;
        RECT 86.895 181.955 90.565 182.765 ;
        RECT 90.575 181.855 94.050 182.765 ;
        RECT 94.725 181.895 95.155 182.680 ;
        RECT 95.635 182.085 99.305 182.765 ;
        RECT 99.460 182.735 99.630 182.955 ;
        RECT 104.975 182.785 105.145 182.975 ;
        RECT 105.430 182.955 105.600 183.005 ;
        RECT 106.630 182.975 107.585 183.005 ;
        RECT 108.055 182.975 111.265 183.885 ;
        RECT 111.275 182.975 113.465 183.885 ;
        RECT 114.035 182.975 117.705 183.885 ;
        RECT 118.025 183.655 118.955 183.885 ;
        RECT 118.025 182.975 119.860 183.655 ;
        RECT 120.015 182.975 121.365 183.885 ;
        RECT 121.395 182.975 122.745 183.885 ;
        RECT 122.775 182.975 128.285 183.785 ;
        RECT 128.295 182.975 131.965 183.785 ;
        RECT 131.975 182.975 133.345 183.785 ;
        RECT 133.365 183.060 133.795 183.845 ;
        RECT 133.815 182.975 137.485 183.785 ;
        RECT 137.955 182.975 139.325 183.755 ;
        RECT 140.255 182.975 141.625 183.755 ;
        RECT 141.635 182.975 143.005 183.785 ;
        RECT 105.430 182.785 105.605 182.955 ;
        RECT 105.435 182.765 105.605 182.785 ;
        RECT 105.895 182.765 106.065 182.955 ;
        RECT 108.185 182.785 108.355 182.975 ;
        RECT 108.660 182.765 108.830 182.955 ;
        RECT 111.420 182.785 111.590 182.975 ;
        RECT 112.795 182.765 112.965 182.955 ;
        RECT 113.265 182.810 113.425 182.920 ;
        RECT 113.710 182.815 113.830 182.925 ;
        RECT 114.175 182.765 114.345 182.955 ;
        RECT 101.590 182.735 102.525 182.765 ;
        RECT 99.460 182.535 102.525 182.735 ;
        RECT 98.375 181.855 99.305 182.085 ;
        RECT 99.315 182.055 102.525 182.535 ;
        RECT 99.315 181.855 100.245 182.055 ;
        RECT 101.575 181.855 102.525 182.055 ;
        RECT 102.535 181.855 105.745 182.765 ;
        RECT 105.755 181.855 108.505 182.765 ;
        RECT 108.515 181.855 110.705 182.765 ;
        RECT 110.815 182.085 113.105 182.765 ;
        RECT 114.035 182.085 116.325 182.765 ;
        RECT 116.480 182.735 116.650 182.955 ;
        RECT 117.390 182.785 117.560 182.975 ;
        RECT 119.695 182.955 119.860 182.975 ;
        RECT 119.695 182.785 119.865 182.955 ;
        RECT 120.160 182.785 120.330 182.975 ;
        RECT 121.075 182.765 121.245 182.955 ;
        RECT 122.460 182.785 122.630 182.975 ;
        RECT 122.915 182.785 123.085 182.975 ;
        RECT 126.595 182.765 126.765 182.955 ;
        RECT 128.435 182.925 128.605 182.975 ;
        RECT 128.430 182.815 128.605 182.925 ;
        RECT 128.435 182.785 128.605 182.815 ;
        RECT 128.895 182.765 129.065 182.955 ;
        RECT 132.115 182.785 132.285 182.975 ;
        RECT 133.955 182.785 134.125 182.975 ;
        RECT 137.630 182.815 137.750 182.925 ;
        RECT 138.095 182.785 138.265 182.975 ;
        RECT 139.475 182.765 139.645 182.955 ;
        RECT 139.935 182.765 140.105 182.955 ;
        RECT 141.305 182.785 141.475 182.975 ;
        RECT 142.695 182.765 142.865 182.975 ;
        RECT 118.610 182.735 119.545 182.765 ;
        RECT 116.480 182.535 119.545 182.735 ;
        RECT 110.815 181.855 111.735 182.085 ;
        RECT 115.405 181.855 116.325 182.085 ;
        RECT 116.335 182.055 119.545 182.535 ;
        RECT 116.335 181.855 117.265 182.055 ;
        RECT 118.595 181.855 119.545 182.055 ;
        RECT 120.485 181.895 120.915 182.680 ;
        RECT 120.935 181.955 126.445 182.765 ;
        RECT 126.455 181.955 128.285 182.765 ;
        RECT 128.755 182.085 136.065 182.765 ;
        RECT 132.270 181.865 133.180 182.085 ;
        RECT 134.715 181.855 136.065 182.085 ;
        RECT 136.210 182.085 139.675 182.765 ;
        RECT 139.795 182.085 141.625 182.765 ;
        RECT 136.210 181.855 137.130 182.085 ;
        RECT 140.280 181.855 141.625 182.085 ;
        RECT 141.635 181.955 143.005 182.765 ;
      LAYER nwell ;
        RECT 17.240 178.735 143.200 181.565 ;
      LAYER pwell ;
        RECT 17.435 177.535 18.805 178.345 ;
        RECT 18.815 177.535 22.485 178.345 ;
        RECT 22.495 178.215 23.425 178.445 ;
        RECT 22.495 177.535 26.165 178.215 ;
        RECT 26.175 177.535 29.845 178.345 ;
        RECT 30.325 177.620 30.755 178.405 ;
        RECT 30.775 177.535 34.445 178.345 ;
        RECT 34.935 177.535 36.285 178.445 ;
        RECT 36.310 177.535 38.125 178.445 ;
        RECT 40.210 178.215 41.345 178.445 ;
        RECT 38.135 177.535 41.345 178.215 ;
        RECT 41.375 177.535 42.725 178.445 ;
        RECT 42.735 177.535 44.085 178.445 ;
        RECT 44.115 177.535 49.625 178.345 ;
        RECT 52.375 178.215 53.305 178.445 ;
        RECT 49.635 177.535 53.305 178.215 ;
        RECT 53.315 177.535 54.665 178.445 ;
        RECT 54.695 177.535 56.065 178.345 ;
        RECT 56.085 177.620 56.515 178.405 ;
        RECT 56.535 177.535 62.045 178.345 ;
        RECT 62.975 177.535 65.895 178.445 ;
        RECT 66.290 178.215 67.210 178.445 ;
        RECT 69.970 178.215 70.890 178.445 ;
        RECT 66.290 177.535 69.755 178.215 ;
        RECT 69.970 177.535 73.435 178.215 ;
        RECT 73.575 177.535 74.925 178.445 ;
        RECT 74.935 177.535 76.285 178.445 ;
        RECT 76.315 177.535 81.825 178.345 ;
        RECT 81.845 177.620 82.275 178.405 ;
        RECT 84.950 178.215 85.870 178.445 ;
        RECT 82.405 177.535 85.870 178.215 ;
        RECT 85.975 177.535 91.485 178.345 ;
        RECT 91.955 177.535 93.305 178.445 ;
        RECT 93.355 177.535 94.705 178.445 ;
        RECT 94.715 177.535 96.545 178.345 ;
        RECT 98.375 178.215 99.305 178.445 ;
        RECT 96.555 177.535 99.305 178.215 ;
        RECT 99.325 177.535 100.675 178.445 ;
        RECT 101.165 177.535 102.515 178.445 ;
        RECT 102.535 177.535 103.905 178.345 ;
        RECT 104.370 177.765 106.205 178.445 ;
        RECT 104.370 177.535 106.060 177.765 ;
        RECT 106.215 177.535 107.585 178.345 ;
        RECT 107.605 177.620 108.035 178.405 ;
        RECT 108.055 177.535 110.805 178.345 ;
        RECT 111.275 178.215 112.195 178.445 ;
        RECT 115.395 178.215 116.325 178.445 ;
        RECT 111.275 177.535 113.565 178.215 ;
        RECT 113.575 177.535 116.325 178.215 ;
        RECT 116.335 178.215 117.265 178.445 ;
        RECT 120.430 178.245 121.385 178.445 ;
        RECT 116.335 177.535 119.085 178.215 ;
        RECT 119.105 177.565 121.385 178.245 ;
        RECT 17.575 177.325 17.745 177.535 ;
        RECT 18.955 177.325 19.125 177.535 ;
        RECT 20.335 177.325 20.505 177.515 ;
        RECT 22.175 177.325 22.345 177.515 ;
        RECT 25.855 177.345 26.025 177.535 ;
        RECT 26.315 177.345 26.485 177.535 ;
        RECT 29.540 177.325 29.710 177.515 ;
        RECT 29.990 177.375 30.110 177.485 ;
        RECT 30.915 177.325 31.085 177.535 ;
        RECT 34.590 177.375 34.710 177.485 ;
        RECT 35.970 177.345 36.140 177.535 ;
        RECT 36.435 177.325 36.605 177.535 ;
        RECT 38.275 177.345 38.445 177.535 ;
        RECT 41.955 177.325 42.125 177.515 ;
        RECT 42.410 177.345 42.580 177.535 ;
        RECT 42.880 177.345 43.050 177.535 ;
        RECT 43.795 177.325 43.965 177.515 ;
        RECT 44.255 177.345 44.425 177.535 ;
        RECT 45.630 177.375 45.750 177.485 ;
        RECT 47.475 177.325 47.645 177.515 ;
        RECT 47.935 177.325 48.105 177.515 ;
        RECT 49.775 177.345 49.945 177.535 ;
        RECT 50.235 177.325 50.405 177.515 ;
        RECT 53.460 177.345 53.630 177.535 ;
        RECT 54.835 177.345 55.005 177.535 ;
        RECT 56.675 177.345 56.845 177.535 ;
        RECT 57.595 177.325 57.765 177.515 ;
        RECT 61.270 177.375 61.390 177.485 ;
        RECT 61.735 177.325 61.905 177.515 ;
        RECT 62.205 177.380 62.365 177.490 ;
        RECT 63.120 177.345 63.290 177.535 ;
        RECT 69.555 177.325 69.725 177.535 ;
        RECT 72.315 177.325 72.485 177.515 ;
        RECT 73.235 177.345 73.405 177.535 ;
        RECT 73.690 177.345 73.860 177.535 ;
        RECT 76.000 177.345 76.170 177.535 ;
        RECT 76.455 177.345 76.625 177.535 ;
        RECT 82.435 177.345 82.605 177.535 ;
        RECT 86.115 177.345 86.285 177.535 ;
        RECT 86.575 177.325 86.745 177.515 ;
        RECT 90.255 177.325 90.425 177.515 ;
        RECT 90.715 177.325 90.885 177.515 ;
        RECT 91.630 177.375 91.750 177.485 ;
        RECT 93.020 177.345 93.190 177.535 ;
        RECT 94.390 177.345 94.560 177.535 ;
        RECT 94.855 177.345 95.025 177.535 ;
        RECT 95.315 177.325 95.485 177.515 ;
        RECT 96.695 177.345 96.865 177.535 ;
        RECT 100.375 177.345 100.545 177.535 ;
        RECT 100.835 177.485 101.005 177.515 ;
        RECT 100.830 177.375 101.005 177.485 ;
        RECT 100.835 177.325 101.005 177.375 ;
        RECT 101.295 177.345 101.465 177.535 ;
        RECT 102.675 177.345 102.845 177.535 ;
        RECT 105.890 177.345 106.060 177.535 ;
        RECT 106.355 177.325 106.525 177.535 ;
        RECT 108.195 177.345 108.365 177.535 ;
        RECT 110.030 177.375 110.150 177.485 ;
        RECT 110.950 177.375 111.070 177.485 ;
        RECT 113.255 177.325 113.425 177.535 ;
        RECT 113.715 177.515 113.885 177.535 ;
        RECT 113.715 177.345 113.890 177.515 ;
        RECT 113.720 177.325 113.890 177.345 ;
        RECT 116.020 177.325 116.190 177.515 ;
        RECT 118.775 177.345 118.945 177.535 ;
        RECT 119.230 177.345 119.400 177.565 ;
        RECT 120.430 177.535 121.385 177.565 ;
        RECT 121.395 177.535 123.225 178.445 ;
        RECT 123.720 178.215 125.065 178.445 ;
        RECT 123.235 177.535 125.065 178.215 ;
        RECT 125.075 177.535 130.585 178.345 ;
        RECT 130.595 177.535 133.345 178.345 ;
        RECT 133.365 177.620 133.795 178.405 ;
        RECT 133.815 178.215 134.745 178.445 ;
        RECT 138.440 178.215 139.785 178.445 ;
        RECT 140.280 178.215 141.625 178.445 ;
        RECT 133.815 177.535 137.715 178.215 ;
        RECT 137.955 177.535 139.785 178.215 ;
        RECT 139.795 177.535 141.625 178.215 ;
        RECT 141.635 177.535 143.005 178.345 ;
        RECT 119.690 177.325 119.860 177.515 ;
        RECT 120.150 177.375 120.270 177.485 ;
        RECT 121.540 177.345 121.710 177.535 ;
        RECT 123.375 177.345 123.545 177.535 ;
        RECT 124.290 177.325 124.460 177.515 ;
        RECT 124.760 177.325 124.930 177.515 ;
        RECT 125.215 177.345 125.385 177.535 ;
        RECT 127.055 177.325 127.225 177.515 ;
        RECT 128.890 177.375 129.010 177.485 ;
        RECT 129.355 177.325 129.525 177.515 ;
        RECT 130.735 177.325 130.905 177.535 ;
        RECT 134.230 177.345 134.400 177.535 ;
        RECT 138.095 177.345 138.265 177.535 ;
        RECT 139.935 177.345 140.105 177.535 ;
        RECT 141.315 177.325 141.485 177.515 ;
        RECT 142.695 177.325 142.865 177.535 ;
        RECT 17.435 176.515 18.805 177.325 ;
        RECT 18.815 176.545 20.185 177.325 ;
        RECT 20.195 176.515 22.025 177.325 ;
        RECT 22.035 176.645 29.345 177.325 ;
        RECT 25.550 176.425 26.460 176.645 ;
        RECT 27.995 176.415 29.345 176.645 ;
        RECT 29.395 176.415 30.745 177.325 ;
        RECT 30.775 176.515 36.285 177.325 ;
        RECT 36.295 176.515 41.805 177.325 ;
        RECT 41.815 176.515 43.185 177.325 ;
        RECT 43.205 176.455 43.635 177.240 ;
        RECT 43.655 176.515 45.485 177.325 ;
        RECT 45.955 176.415 47.770 177.325 ;
        RECT 47.795 176.645 50.085 177.325 ;
        RECT 50.095 176.645 57.405 177.325 ;
        RECT 49.165 176.415 50.085 176.645 ;
        RECT 53.610 176.425 54.520 176.645 ;
        RECT 56.055 176.415 57.405 176.645 ;
        RECT 57.455 176.515 61.125 177.325 ;
        RECT 61.595 176.645 68.905 177.325 ;
        RECT 65.110 176.425 66.020 176.645 ;
        RECT 67.555 176.415 68.905 176.645 ;
        RECT 68.965 176.455 69.395 177.240 ;
        RECT 69.425 176.415 72.155 177.325 ;
        RECT 72.175 176.645 79.485 177.325 ;
        RECT 75.690 176.425 76.600 176.645 ;
        RECT 78.135 176.415 79.485 176.645 ;
        RECT 79.575 176.645 86.885 177.325 ;
        RECT 86.990 176.645 90.455 177.325 ;
        RECT 79.575 176.415 80.925 176.645 ;
        RECT 82.460 176.425 83.370 176.645 ;
        RECT 86.990 176.415 87.910 176.645 ;
        RECT 90.575 176.515 94.245 177.325 ;
        RECT 94.725 176.455 95.155 177.240 ;
        RECT 95.175 176.515 100.685 177.325 ;
        RECT 100.695 176.515 106.205 177.325 ;
        RECT 106.215 176.515 109.885 177.325 ;
        RECT 110.485 176.415 113.485 177.325 ;
        RECT 113.575 176.645 115.850 177.325 ;
        RECT 114.480 176.415 115.850 176.645 ;
        RECT 115.875 176.415 117.705 177.325 ;
        RECT 117.730 176.645 120.005 177.325 ;
        RECT 117.730 176.415 119.100 176.645 ;
        RECT 120.485 176.455 120.915 177.240 ;
        RECT 121.130 176.415 124.605 177.325 ;
        RECT 124.615 176.415 126.825 177.325 ;
        RECT 126.915 176.515 128.745 177.325 ;
        RECT 129.215 176.545 130.585 177.325 ;
        RECT 130.595 176.645 137.905 177.325 ;
        RECT 134.110 176.425 135.020 176.645 ;
        RECT 136.555 176.415 137.905 176.645 ;
        RECT 138.050 176.645 141.515 177.325 ;
        RECT 138.050 176.415 138.970 176.645 ;
        RECT 141.635 176.515 143.005 177.325 ;
      LAYER nwell ;
        RECT 17.240 173.295 143.200 176.125 ;
      LAYER pwell ;
        RECT 17.435 172.095 18.805 172.905 ;
        RECT 18.815 172.095 20.645 172.905 ;
        RECT 24.630 172.775 25.540 172.995 ;
        RECT 27.075 172.775 28.425 173.005 ;
        RECT 21.115 172.095 28.425 172.775 ;
        RECT 28.475 172.095 29.825 173.005 ;
        RECT 30.325 172.180 30.755 172.965 ;
        RECT 30.775 172.095 32.605 172.905 ;
        RECT 33.560 172.775 34.905 173.005 ;
        RECT 33.075 172.095 34.905 172.775 ;
        RECT 35.370 172.325 37.205 173.005 ;
        RECT 35.370 172.095 37.060 172.325 ;
        RECT 37.215 172.095 39.965 173.005 ;
        RECT 39.975 172.095 43.185 173.005 ;
        RECT 46.155 172.915 47.105 173.005 ;
        RECT 43.205 172.095 45.945 172.775 ;
        RECT 46.155 172.095 48.085 172.915 ;
        RECT 48.755 172.775 50.105 173.005 ;
        RECT 51.640 172.775 52.550 172.995 ;
        RECT 48.755 172.095 56.065 172.775 ;
        RECT 56.085 172.180 56.515 172.965 ;
        RECT 56.535 172.775 57.670 173.005 ;
        RECT 56.535 172.095 59.745 172.775 ;
        RECT 59.755 172.095 61.125 172.905 ;
        RECT 64.650 172.775 65.560 172.995 ;
        RECT 67.095 172.775 68.445 173.005 ;
        RECT 61.135 172.095 68.445 172.775 ;
        RECT 68.515 172.095 69.865 173.005 ;
        RECT 69.875 172.095 71.245 172.905 ;
        RECT 71.350 172.775 72.270 173.005 ;
        RECT 71.350 172.095 74.815 172.775 ;
        RECT 75.105 172.095 78.605 173.005 ;
        RECT 78.615 172.805 79.560 173.005 ;
        RECT 80.895 172.805 81.825 173.005 ;
        RECT 78.615 172.325 81.825 172.805 ;
        RECT 78.615 172.125 81.685 172.325 ;
        RECT 81.845 172.180 82.275 172.965 ;
        RECT 85.955 172.775 86.885 173.005 ;
        RECT 78.615 172.095 79.560 172.125 ;
        RECT 17.575 171.885 17.745 172.095 ;
        RECT 18.955 171.885 19.125 172.095 ;
        RECT 20.790 171.935 20.910 172.045 ;
        RECT 21.255 171.905 21.425 172.095 ;
        RECT 21.710 171.885 21.880 172.075 ;
        RECT 25.395 171.885 25.565 172.075 ;
        RECT 27.695 171.885 27.865 172.075 ;
        RECT 28.155 171.885 28.325 172.075 ;
        RECT 28.620 171.905 28.790 172.095 ;
        RECT 29.990 171.935 30.110 172.045 ;
        RECT 30.915 171.905 31.085 172.095 ;
        RECT 31.375 171.885 31.545 172.075 ;
        RECT 32.750 171.935 32.870 172.045 ;
        RECT 33.215 171.905 33.385 172.095 ;
        RECT 36.890 171.905 37.060 172.095 ;
        RECT 37.350 171.885 37.520 172.075 ;
        RECT 37.810 171.935 37.930 172.045 ;
        RECT 39.655 171.905 39.825 172.095 ;
        RECT 40.115 171.905 40.285 172.095 ;
        RECT 42.875 171.885 43.045 172.075 ;
        RECT 43.800 171.885 43.970 172.075 ;
        RECT 45.635 171.905 45.805 172.095 ;
        RECT 47.935 172.075 48.085 172.095 ;
        RECT 47.935 171.905 48.105 172.075 ;
        RECT 48.390 171.935 48.510 172.045 ;
        RECT 55.755 171.905 55.925 172.095 ;
        RECT 59.435 171.885 59.605 172.095 ;
        RECT 59.895 172.075 60.065 172.095 ;
        RECT 59.895 171.905 60.070 172.075 ;
        RECT 59.900 171.885 60.070 171.905 ;
        RECT 61.275 171.885 61.445 172.095 ;
        RECT 66.795 171.885 66.965 172.075 ;
        RECT 68.630 171.905 68.800 172.095 ;
        RECT 70.015 171.905 70.185 172.095 ;
        RECT 74.615 171.905 74.785 172.095 ;
        RECT 75.105 172.075 75.240 172.095 ;
        RECT 75.070 171.905 75.240 172.075 ;
        RECT 76.455 171.885 76.625 172.075 ;
        RECT 76.915 171.885 77.085 172.075 ;
        RECT 81.515 171.905 81.685 172.125 ;
        RECT 82.985 172.095 86.885 172.775 ;
        RECT 86.895 172.095 88.245 173.005 ;
        RECT 88.275 172.095 93.785 172.905 ;
        RECT 93.795 172.095 95.165 172.905 ;
        RECT 95.175 172.775 96.105 173.005 ;
        RECT 99.410 172.775 100.330 173.005 ;
        RECT 105.650 172.775 106.570 173.005 ;
        RECT 95.175 172.095 99.075 172.775 ;
        RECT 99.410 172.095 102.875 172.775 ;
        RECT 103.105 172.095 106.570 172.775 ;
        RECT 107.605 172.180 108.035 172.965 ;
        RECT 108.135 172.095 110.345 173.005 ;
        RECT 110.355 172.095 111.705 173.005 ;
        RECT 111.735 172.095 113.085 173.005 ;
        RECT 114.910 172.805 115.865 173.005 ;
        RECT 113.585 172.125 115.865 172.805 ;
        RECT 82.430 171.935 82.550 172.045 ;
        RECT 83.815 171.905 83.985 172.075 ;
        RECT 81.515 171.885 81.680 171.905 ;
        RECT 83.815 171.885 83.965 171.905 ;
        RECT 84.275 171.885 84.445 172.075 ;
        RECT 86.300 171.905 86.470 172.095 ;
        RECT 87.040 171.905 87.210 172.095 ;
        RECT 88.230 171.885 88.400 172.075 ;
        RECT 88.415 171.905 88.585 172.095 ;
        RECT 92.095 171.885 92.265 172.075 ;
        RECT 93.935 171.905 94.105 172.095 ;
        RECT 95.590 171.905 95.760 172.095 ;
        RECT 102.215 171.885 102.385 172.075 ;
        RECT 102.675 171.905 102.845 172.095 ;
        RECT 103.135 171.905 103.305 172.095 ;
        RECT 105.435 171.885 105.605 172.075 ;
        RECT 105.885 171.885 106.055 172.075 ;
        RECT 106.825 171.940 106.985 172.050 ;
        RECT 109.115 171.885 109.285 172.075 ;
        RECT 110.030 171.905 110.200 172.095 ;
        RECT 110.500 171.905 110.670 172.095 ;
        RECT 112.800 171.905 112.970 172.095 ;
        RECT 113.710 172.075 113.880 172.125 ;
        RECT 114.910 172.095 115.865 172.125 ;
        RECT 116.025 172.095 119.680 173.005 ;
        RECT 121.350 172.805 122.305 173.005 ;
        RECT 120.025 172.125 122.305 172.805 ;
        RECT 123.365 172.775 124.295 173.005 ;
        RECT 116.025 172.075 116.185 172.095 ;
        RECT 113.250 171.935 113.370 172.045 ;
        RECT 113.710 171.905 113.885 172.075 ;
        RECT 116.015 171.905 116.185 172.075 ;
        RECT 113.715 171.885 113.885 171.905 ;
        RECT 116.935 171.885 117.105 172.075 ;
        RECT 119.705 171.930 119.865 172.040 ;
        RECT 120.150 171.905 120.320 172.125 ;
        RECT 121.350 172.095 122.305 172.125 ;
        RECT 122.460 172.095 124.295 172.775 ;
        RECT 124.615 172.095 125.985 172.905 ;
        RECT 125.995 172.095 129.205 173.005 ;
        RECT 132.415 172.775 133.345 173.005 ;
        RECT 129.445 172.095 133.345 172.775 ;
        RECT 133.365 172.180 133.795 172.965 ;
        RECT 137.330 172.775 138.240 172.995 ;
        RECT 139.775 172.775 141.125 173.005 ;
        RECT 133.815 172.095 141.125 172.775 ;
        RECT 141.635 172.095 143.005 172.905 ;
        RECT 122.460 172.075 122.625 172.095 ;
        RECT 121.075 171.905 121.245 172.075 ;
        RECT 122.455 171.905 122.625 172.075 ;
        RECT 124.755 171.905 124.925 172.095 ;
        RECT 121.085 171.885 121.245 171.905 ;
        RECT 125.215 171.885 125.385 172.075 ;
        RECT 126.135 171.905 126.305 172.095 ;
        RECT 128.435 171.885 128.605 172.075 ;
        RECT 132.760 171.905 132.930 172.095 ;
        RECT 133.955 171.905 134.125 172.095 ;
        RECT 135.060 171.885 135.230 172.075 ;
        RECT 135.795 171.885 135.965 172.075 ;
        RECT 140.395 171.885 140.565 172.075 ;
        RECT 140.865 171.930 141.025 172.040 ;
        RECT 141.310 171.935 141.430 172.045 ;
        RECT 142.695 171.885 142.865 172.095 ;
        RECT 17.435 171.075 18.805 171.885 ;
        RECT 18.815 171.075 20.645 171.885 ;
        RECT 20.675 170.975 22.025 171.885 ;
        RECT 22.035 171.205 25.705 171.885 ;
        RECT 25.715 171.205 28.005 171.885 ;
        RECT 28.015 171.205 31.225 171.885 ;
        RECT 22.035 170.975 22.965 171.205 ;
        RECT 25.715 170.975 26.635 171.205 ;
        RECT 30.090 170.975 31.225 171.205 ;
        RECT 31.235 171.075 33.985 171.885 ;
        RECT 34.190 170.975 37.665 171.885 ;
        RECT 38.370 171.205 43.185 171.885 ;
        RECT 43.205 171.015 43.635 171.800 ;
        RECT 43.655 170.975 54.665 171.885 ;
        RECT 54.930 171.205 59.745 171.885 ;
        RECT 59.755 170.975 61.105 171.885 ;
        RECT 61.135 171.075 66.645 171.885 ;
        RECT 66.655 171.075 68.485 171.885 ;
        RECT 68.965 171.015 69.395 171.800 ;
        RECT 69.455 171.205 76.765 171.885 ;
        RECT 69.455 170.975 70.805 171.205 ;
        RECT 72.340 170.985 73.250 171.205 ;
        RECT 76.785 170.975 79.515 171.885 ;
        RECT 79.845 171.205 81.680 171.885 ;
        RECT 79.845 170.975 80.775 171.205 ;
        RECT 82.035 171.065 83.965 171.885 ;
        RECT 84.245 171.205 87.710 171.885 ;
        RECT 82.035 170.975 82.985 171.065 ;
        RECT 86.790 170.975 87.710 171.205 ;
        RECT 87.815 171.205 91.715 171.885 ;
        RECT 87.815 170.975 88.745 171.205 ;
        RECT 91.955 171.075 94.705 171.885 ;
        RECT 94.725 171.015 95.155 171.800 ;
        RECT 95.215 171.205 102.525 171.885 ;
        RECT 95.215 170.975 96.565 171.205 ;
        RECT 98.100 170.985 99.010 171.205 ;
        RECT 102.535 170.975 105.745 171.885 ;
        RECT 105.755 170.975 108.965 171.885 ;
        RECT 108.975 171.075 112.645 171.885 ;
        RECT 113.575 170.975 116.785 171.885 ;
        RECT 116.805 170.975 119.535 171.885 ;
        RECT 120.485 171.015 120.915 171.800 ;
        RECT 121.085 170.975 124.740 171.885 ;
        RECT 125.075 170.975 128.285 171.885 ;
        RECT 128.295 170.975 131.505 171.885 ;
        RECT 131.745 171.205 135.645 171.885 ;
        RECT 134.715 170.975 135.645 171.205 ;
        RECT 135.655 171.105 137.025 171.885 ;
        RECT 137.130 171.205 140.595 171.885 ;
        RECT 137.130 170.975 138.050 171.205 ;
        RECT 141.635 171.075 143.005 171.885 ;
      LAYER nwell ;
        RECT 17.240 167.855 143.200 170.685 ;
      LAYER pwell ;
        RECT 17.435 166.655 18.805 167.465 ;
        RECT 18.815 166.655 24.325 167.465 ;
        RECT 25.255 166.655 27.070 167.565 ;
        RECT 27.095 166.655 29.845 167.465 ;
        RECT 30.325 166.740 30.755 167.525 ;
        RECT 30.775 166.655 32.605 167.465 ;
        RECT 34.410 167.365 35.365 167.565 ;
        RECT 33.085 166.685 35.365 167.365 ;
        RECT 17.575 166.445 17.745 166.655 ;
        RECT 18.955 166.445 19.125 166.655 ;
        RECT 21.710 166.495 21.830 166.605 ;
        RECT 22.175 166.445 22.345 166.635 ;
        RECT 24.485 166.500 24.645 166.610 ;
        RECT 26.775 166.445 26.945 166.655 ;
        RECT 27.235 166.445 27.405 166.655 ;
        RECT 29.995 166.605 30.165 166.635 ;
        RECT 29.990 166.495 30.165 166.605 ;
        RECT 29.995 166.445 30.165 166.495 ;
        RECT 30.915 166.465 31.085 166.655 ;
        RECT 33.210 166.635 33.380 166.685 ;
        RECT 34.410 166.655 35.365 166.685 ;
        RECT 36.315 166.655 37.665 167.565 ;
        RECT 37.870 166.655 41.345 167.565 ;
        RECT 41.355 167.365 42.300 167.565 ;
        RECT 43.635 167.365 44.565 167.565 ;
        RECT 41.355 166.885 44.565 167.365 ;
        RECT 45.625 167.335 46.555 167.565 ;
        RECT 41.355 166.685 44.425 166.885 ;
        RECT 41.355 166.655 42.300 166.685 ;
        RECT 36.430 166.635 36.600 166.655 ;
        RECT 32.750 166.495 32.870 166.605 ;
        RECT 33.210 166.465 33.385 166.635 ;
        RECT 35.525 166.500 35.685 166.610 ;
        RECT 36.430 166.465 36.605 166.635 ;
        RECT 39.190 166.495 39.310 166.605 ;
        RECT 33.215 166.445 33.385 166.465 ;
        RECT 36.435 166.445 36.605 166.465 ;
        RECT 17.435 165.635 18.805 166.445 ;
        RECT 18.815 165.635 21.565 166.445 ;
        RECT 22.075 165.535 25.245 166.445 ;
        RECT 25.255 165.765 27.085 166.445 ;
        RECT 27.095 165.635 29.845 166.445 ;
        RECT 29.955 165.535 33.065 166.445 ;
        RECT 33.175 165.535 36.285 166.445 ;
        RECT 36.295 165.635 39.045 166.445 ;
        RECT 39.650 166.415 39.820 166.635 ;
        RECT 41.030 166.465 41.200 166.655 ;
        RECT 41.955 166.445 42.125 166.635 ;
        RECT 43.800 166.445 43.970 166.635 ;
        RECT 44.255 166.465 44.425 166.685 ;
        RECT 44.720 166.655 46.555 167.335 ;
        RECT 46.875 166.655 50.545 167.465 ;
        RECT 53.295 167.335 54.225 167.565 ;
        RECT 50.555 166.655 54.225 167.335 ;
        RECT 54.255 166.655 55.605 167.565 ;
        RECT 56.085 166.740 56.515 167.525 ;
        RECT 56.915 166.655 59.340 167.335 ;
        RECT 59.755 166.655 63.425 167.465 ;
        RECT 64.355 166.655 69.170 167.335 ;
        RECT 69.415 166.655 80.425 167.565 ;
        RECT 80.455 166.655 81.805 167.565 ;
        RECT 81.845 166.740 82.275 167.525 ;
        RECT 82.795 167.335 84.145 167.565 ;
        RECT 85.680 167.335 86.590 167.555 ;
        RECT 93.630 167.335 94.540 167.555 ;
        RECT 96.075 167.335 97.425 167.565 ;
        RECT 82.795 166.655 90.105 167.335 ;
        RECT 90.115 166.655 97.425 167.335 ;
        RECT 97.475 166.655 99.305 167.465 ;
        RECT 99.355 167.335 100.705 167.565 ;
        RECT 102.240 167.335 103.150 167.555 ;
        RECT 99.355 166.655 106.665 167.335 ;
        RECT 107.605 166.740 108.035 167.525 ;
        RECT 110.710 167.335 111.630 167.565 ;
        RECT 108.165 166.655 111.630 167.335 ;
        RECT 111.815 166.655 114.815 167.565 ;
        RECT 114.955 166.655 117.875 167.565 ;
        RECT 118.175 166.655 120.005 167.465 ;
        RECT 120.025 166.655 122.755 167.565 ;
        RECT 123.085 167.335 124.015 167.565 ;
        RECT 123.085 166.655 124.920 167.335 ;
        RECT 125.075 166.655 130.585 167.465 ;
        RECT 132.000 167.335 133.345 167.565 ;
        RECT 131.515 166.655 133.345 167.335 ;
        RECT 133.365 166.740 133.795 167.525 ;
        RECT 133.815 167.335 134.745 167.565 ;
        RECT 138.050 167.335 138.970 167.565 ;
        RECT 133.815 166.655 137.715 167.335 ;
        RECT 138.050 166.655 141.515 167.335 ;
        RECT 141.635 166.655 143.005 167.465 ;
        RECT 44.720 166.635 44.885 166.655 ;
        RECT 44.715 166.465 44.885 166.635 ;
        RECT 47.015 166.465 47.185 166.655 ;
        RECT 47.475 166.445 47.645 166.635 ;
        RECT 50.695 166.465 50.865 166.655 ;
        RECT 52.995 166.445 53.165 166.635 ;
        RECT 55.290 166.465 55.460 166.655 ;
        RECT 55.750 166.495 55.870 166.605 ;
        RECT 57.595 166.445 57.765 166.635 ;
        RECT 58.055 166.445 58.225 166.635 ;
        RECT 59.435 166.465 59.605 166.635 ;
        RECT 59.895 166.465 60.065 166.655 ;
        RECT 63.575 166.445 63.745 166.635 ;
        RECT 64.495 166.465 64.665 166.655 ;
        RECT 69.560 166.635 69.730 166.655 ;
        RECT 65.420 166.445 65.590 166.635 ;
        RECT 67.255 166.445 67.425 166.635 ;
        RECT 69.555 166.465 69.730 166.635 ;
        RECT 69.555 166.445 69.725 166.465 ;
        RECT 76.915 166.445 77.085 166.635 ;
        RECT 78.295 166.445 78.465 166.635 ;
        RECT 81.520 166.465 81.690 166.655 ;
        RECT 82.250 166.445 82.420 166.635 ;
        RECT 82.430 166.495 82.550 166.605 ;
        RECT 86.390 166.445 86.560 166.635 ;
        RECT 89.795 166.465 89.965 166.655 ;
        RECT 90.255 166.445 90.425 166.655 ;
        RECT 93.945 166.490 94.105 166.600 ;
        RECT 95.315 166.445 95.485 166.635 ;
        RECT 97.615 166.465 97.785 166.655 ;
        RECT 106.355 166.635 106.525 166.655 ;
        RECT 98.075 166.445 98.245 166.635 ;
        RECT 103.135 166.445 103.305 166.635 ;
        RECT 105.890 166.495 106.010 166.605 ;
        RECT 106.350 166.465 106.525 166.635 ;
        RECT 106.825 166.500 106.985 166.610 ;
        RECT 106.350 166.445 106.520 166.465 ;
        RECT 107.735 166.445 107.905 166.635 ;
        RECT 108.195 166.465 108.365 166.655 ;
        RECT 111.875 166.465 112.045 166.655 ;
        RECT 113.255 166.445 113.425 166.635 ;
        RECT 115.100 166.465 115.270 166.655 ;
        RECT 116.930 166.495 117.050 166.605 ;
        RECT 118.315 166.465 118.485 166.655 ;
        RECT 119.235 166.445 119.405 166.635 ;
        RECT 119.705 166.490 119.865 166.600 ;
        RECT 122.455 166.465 122.625 166.655 ;
        RECT 124.755 166.635 124.920 166.655 ;
        RECT 124.290 166.445 124.460 166.635 ;
        RECT 124.755 166.445 124.925 166.635 ;
        RECT 125.215 166.465 125.385 166.655 ;
        RECT 128.435 166.445 128.605 166.635 ;
        RECT 129.815 166.445 129.985 166.635 ;
        RECT 130.745 166.500 130.905 166.610 ;
        RECT 131.195 166.445 131.365 166.635 ;
        RECT 131.655 166.465 131.825 166.655 ;
        RECT 134.230 166.465 134.400 166.655 ;
        RECT 139.475 166.445 139.645 166.635 ;
        RECT 139.935 166.445 140.105 166.635 ;
        RECT 141.315 166.465 141.485 166.655 ;
        RECT 142.695 166.445 142.865 166.655 ;
        RECT 40.850 166.415 41.805 166.445 ;
        RECT 39.525 165.735 41.805 166.415 ;
        RECT 40.850 165.535 41.805 165.735 ;
        RECT 41.815 165.635 43.185 166.445 ;
        RECT 43.205 165.575 43.635 166.360 ;
        RECT 43.655 165.535 47.310 166.445 ;
        RECT 47.335 165.635 52.845 166.445 ;
        RECT 52.895 165.535 56.065 166.445 ;
        RECT 56.075 165.765 57.905 166.445 ;
        RECT 57.915 165.635 63.425 166.445 ;
        RECT 63.435 165.635 65.265 166.445 ;
        RECT 65.275 165.535 67.105 166.445 ;
        RECT 67.115 165.635 68.945 166.445 ;
        RECT 68.965 165.575 69.395 166.360 ;
        RECT 69.415 165.765 76.725 166.445 ;
        RECT 72.930 165.545 73.840 165.765 ;
        RECT 75.375 165.535 76.725 165.765 ;
        RECT 76.775 165.635 78.145 166.445 ;
        RECT 78.265 165.765 81.730 166.445 ;
        RECT 80.810 165.535 81.730 165.765 ;
        RECT 81.835 165.765 85.735 166.445 ;
        RECT 85.975 165.765 89.875 166.445 ;
        RECT 81.835 165.535 82.765 165.765 ;
        RECT 85.975 165.535 86.905 165.765 ;
        RECT 90.115 165.635 93.785 166.445 ;
        RECT 94.725 165.575 95.155 166.360 ;
        RECT 95.175 165.635 97.925 166.445 ;
        RECT 97.935 165.765 102.750 166.445 ;
        RECT 102.995 165.635 105.745 166.445 ;
        RECT 106.235 165.535 107.585 166.445 ;
        RECT 107.595 165.635 113.105 166.445 ;
        RECT 113.115 165.635 116.785 166.445 ;
        RECT 117.255 165.765 119.545 166.445 ;
        RECT 117.255 165.535 118.175 165.765 ;
        RECT 120.485 165.575 120.915 166.360 ;
        RECT 121.130 165.535 124.605 166.445 ;
        RECT 124.615 165.635 128.285 166.445 ;
        RECT 128.295 165.635 129.665 166.445 ;
        RECT 129.675 165.665 131.045 166.445 ;
        RECT 131.055 165.765 138.365 166.445 ;
        RECT 134.570 165.545 135.480 165.765 ;
        RECT 137.015 165.535 138.365 165.765 ;
        RECT 138.415 165.665 139.785 166.445 ;
        RECT 139.795 165.765 141.625 166.445 ;
        RECT 140.280 165.535 141.625 165.765 ;
        RECT 141.635 165.635 143.005 166.445 ;
      LAYER nwell ;
        RECT 17.240 162.415 143.200 165.245 ;
      LAYER pwell ;
        RECT 17.435 161.215 18.805 162.025 ;
        RECT 18.815 161.215 20.185 161.995 ;
        RECT 20.195 161.215 21.565 162.025 ;
        RECT 21.585 161.895 24.585 162.125 ;
        RECT 26.175 161.895 27.105 162.125 ;
        RECT 21.585 161.805 26.165 161.895 ;
        RECT 21.575 161.445 26.165 161.805 ;
        RECT 21.575 161.255 22.505 161.445 ;
        RECT 21.585 161.215 22.505 161.255 ;
        RECT 24.595 161.215 26.165 161.445 ;
        RECT 26.175 161.215 29.845 161.895 ;
        RECT 30.325 161.300 30.755 162.085 ;
        RECT 31.255 161.215 32.605 162.125 ;
        RECT 32.615 161.215 35.365 162.025 ;
        RECT 35.375 161.215 38.585 162.125 ;
        RECT 41.315 161.925 42.265 162.125 ;
        RECT 38.595 161.245 42.265 161.925 ;
        RECT 17.575 161.005 17.745 161.215 ;
        RECT 18.965 161.195 19.135 161.215 ;
        RECT 18.955 161.025 19.135 161.195 ;
        RECT 20.335 161.025 20.505 161.215 ;
        RECT 20.790 161.055 20.910 161.165 ;
        RECT 25.855 161.025 26.025 161.215 ;
        RECT 18.955 161.005 19.125 161.025 ;
        RECT 28.155 161.005 28.325 161.195 ;
        RECT 28.615 161.005 28.785 161.195 ;
        RECT 29.535 161.025 29.705 161.215 ;
        RECT 29.990 161.055 30.110 161.165 ;
        RECT 30.910 161.055 31.030 161.165 ;
        RECT 31.370 161.055 31.490 161.165 ;
        RECT 31.840 161.005 32.010 161.195 ;
        RECT 32.290 161.025 32.460 161.215 ;
        RECT 32.755 161.025 32.925 161.215 ;
        RECT 34.135 161.005 34.305 161.195 ;
        RECT 37.355 161.005 37.525 161.195 ;
        RECT 38.285 161.025 38.455 161.215 ;
        RECT 38.740 161.005 38.910 161.245 ;
        RECT 41.315 161.215 42.265 161.245 ;
        RECT 43.505 161.895 44.435 162.125 ;
        RECT 43.505 161.215 45.340 161.895 ;
        RECT 45.495 161.215 49.165 162.025 ;
        RECT 49.645 161.215 52.375 162.125 ;
        RECT 53.145 161.215 56.065 162.125 ;
        RECT 56.085 161.300 56.515 162.085 ;
        RECT 56.575 161.895 57.925 162.125 ;
        RECT 59.460 161.895 60.370 162.115 ;
        RECT 56.575 161.215 63.885 161.895 ;
        RECT 63.895 161.215 69.405 162.025 ;
        RECT 70.785 161.895 71.705 162.125 ;
        RECT 73.545 161.895 74.465 162.125 ;
        RECT 69.415 161.215 71.705 161.895 ;
        RECT 72.175 161.215 74.465 161.895 ;
        RECT 74.475 161.215 77.950 162.125 ;
        RECT 78.155 161.925 79.105 162.125 ;
        RECT 78.155 161.245 81.825 161.925 ;
        RECT 81.845 161.300 82.275 162.085 ;
        RECT 85.870 161.895 86.790 162.125 ;
        RECT 90.095 161.895 91.025 162.125 ;
        RECT 93.690 161.895 94.610 162.125 ;
        RECT 78.155 161.215 79.105 161.245 ;
        RECT 45.175 161.195 45.340 161.215 ;
        RECT 42.425 161.050 42.585 161.170 ;
        RECT 43.795 161.005 43.965 161.195 ;
        RECT 45.175 161.025 45.345 161.195 ;
        RECT 45.635 161.005 45.805 161.215 ;
        RECT 49.310 161.055 49.430 161.165 ;
        RECT 49.775 161.025 49.945 161.215 ;
        RECT 51.160 161.005 51.330 161.195 ;
        RECT 51.615 161.005 51.785 161.195 ;
        RECT 52.530 161.055 52.650 161.165 ;
        RECT 55.750 161.025 55.920 161.215 ;
        RECT 62.195 161.005 62.365 161.195 ;
        RECT 63.575 161.025 63.745 161.215 ;
        RECT 64.035 161.025 64.205 161.215 ;
        RECT 65.875 161.005 66.045 161.195 ;
        RECT 66.335 161.005 66.505 161.195 ;
        RECT 69.555 161.005 69.725 161.215 ;
        RECT 71.395 161.005 71.565 161.195 ;
        RECT 71.850 161.055 71.970 161.165 ;
        RECT 72.315 161.025 72.485 161.215 ;
        RECT 17.435 160.195 18.805 161.005 ;
        RECT 18.815 160.195 20.645 161.005 ;
        RECT 21.155 160.325 28.465 161.005 ;
        RECT 21.155 160.095 22.505 160.325 ;
        RECT 24.040 160.105 24.950 160.325 ;
        RECT 28.475 160.195 31.225 161.005 ;
        RECT 31.840 160.775 33.530 161.005 ;
        RECT 31.695 160.095 33.530 160.775 ;
        RECT 33.995 160.095 37.205 161.005 ;
        RECT 37.215 160.195 38.585 161.005 ;
        RECT 38.595 160.325 42.265 161.005 ;
        RECT 38.595 160.095 39.520 160.325 ;
        RECT 43.205 160.135 43.635 160.920 ;
        RECT 43.655 160.195 45.485 161.005 ;
        RECT 45.495 160.095 50.045 161.005 ;
        RECT 50.095 160.095 51.445 161.005 ;
        RECT 51.475 160.325 55.145 161.005 ;
        RECT 54.215 160.095 55.145 160.325 ;
        RECT 55.195 160.325 62.505 161.005 ;
        RECT 62.515 160.325 66.185 161.005 ;
        RECT 55.195 160.095 56.545 160.325 ;
        RECT 58.080 160.105 58.990 160.325 ;
        RECT 62.515 160.095 63.445 160.325 ;
        RECT 66.195 160.195 68.945 161.005 ;
        RECT 68.965 160.135 69.395 160.920 ;
        RECT 69.415 160.195 71.245 161.005 ;
        RECT 71.255 160.325 74.005 161.005 ;
        RECT 74.160 160.975 74.330 161.195 ;
        RECT 74.620 161.025 74.790 161.215 ;
        RECT 79.685 161.005 79.855 161.195 ;
        RECT 80.145 161.050 80.305 161.160 ;
        RECT 81.510 161.025 81.680 161.245 ;
        RECT 83.325 161.215 86.790 161.895 ;
        RECT 87.125 161.215 91.025 161.895 ;
        RECT 91.145 161.215 94.610 161.895 ;
        RECT 95.175 161.895 96.105 162.125 ;
        RECT 95.175 161.215 99.075 161.895 ;
        RECT 99.315 161.215 100.685 162.025 ;
        RECT 103.350 161.895 104.270 162.125 ;
        RECT 100.805 161.215 104.270 161.895 ;
        RECT 104.375 161.215 107.125 162.025 ;
        RECT 107.605 161.300 108.035 162.085 ;
        RECT 118.855 162.035 119.805 162.125 ;
        RECT 108.055 161.215 113.565 162.025 ;
        RECT 113.575 161.215 117.245 162.025 ;
        RECT 117.875 161.215 119.805 162.035 ;
        RECT 120.015 161.895 120.935 162.125 ;
        RECT 120.015 161.215 123.600 161.895 ;
        RECT 123.890 161.215 127.365 162.125 ;
        RECT 127.375 161.215 130.585 162.125 ;
        RECT 130.595 161.215 133.345 162.025 ;
        RECT 133.365 161.300 133.795 162.085 ;
        RECT 133.815 161.895 134.745 162.125 ;
        RECT 138.050 161.895 138.970 162.125 ;
        RECT 133.815 161.215 137.715 161.895 ;
        RECT 138.050 161.215 141.515 161.895 ;
        RECT 141.635 161.215 143.005 162.025 ;
        RECT 82.445 161.060 82.605 161.170 ;
        RECT 83.355 161.025 83.525 161.215 ;
        RECT 75.820 160.975 76.765 161.005 ;
        RECT 73.075 160.095 74.005 160.325 ;
        RECT 74.015 160.295 76.765 160.975 ;
        RECT 75.820 160.095 76.765 160.295 ;
        RECT 76.775 160.095 79.985 161.005 ;
        RECT 80.915 160.975 81.850 161.005 ;
        RECT 83.810 160.975 83.980 161.195 ;
        RECT 90.440 161.025 90.610 161.215 ;
        RECT 91.175 161.005 91.345 161.215 ;
        RECT 91.635 161.005 91.805 161.195 ;
        RECT 94.390 161.055 94.510 161.165 ;
        RECT 94.850 161.055 94.970 161.165 ;
        RECT 95.325 161.050 95.485 161.160 ;
        RECT 95.590 161.025 95.760 161.215 ;
        RECT 99.455 161.025 99.625 161.215 ;
        RECT 100.835 161.025 101.005 161.215 ;
        RECT 103.135 161.005 103.305 161.195 ;
        RECT 103.595 161.005 103.765 161.195 ;
        RECT 104.515 161.025 104.685 161.215 ;
        RECT 106.815 161.005 106.985 161.195 ;
        RECT 107.270 161.055 107.390 161.165 ;
        RECT 108.195 161.025 108.365 161.215 ;
        RECT 113.715 161.195 113.885 161.215 ;
        RECT 117.875 161.195 118.025 161.215 ;
        RECT 108.650 161.055 108.770 161.165 ;
        RECT 109.115 161.025 109.285 161.195 ;
        RECT 109.135 161.005 109.285 161.025 ;
        RECT 112.335 161.005 112.505 161.195 ;
        RECT 113.715 161.025 113.890 161.195 ;
        RECT 113.720 161.005 113.890 161.025 ;
        RECT 115.090 161.005 115.260 161.195 ;
        RECT 116.480 161.005 116.650 161.195 ;
        RECT 116.945 161.050 117.105 161.160 ;
        RECT 117.390 161.055 117.510 161.165 ;
        RECT 117.855 161.025 118.025 161.195 ;
        RECT 120.160 161.025 120.330 161.215 ;
        RECT 118.005 161.005 118.025 161.025 ;
        RECT 80.915 160.775 83.980 160.975 ;
        RECT 80.915 160.295 84.125 160.775 ;
        RECT 80.915 160.095 81.865 160.295 ;
        RECT 83.195 160.095 84.125 160.295 ;
        RECT 84.175 160.325 91.485 161.005 ;
        RECT 84.175 160.095 85.525 160.325 ;
        RECT 87.060 160.105 87.970 160.325 ;
        RECT 91.495 160.195 94.245 161.005 ;
        RECT 94.725 160.135 95.155 160.920 ;
        RECT 96.135 160.325 103.445 161.005 ;
        RECT 96.135 160.095 97.485 160.325 ;
        RECT 99.020 160.105 99.930 160.325 ;
        RECT 103.455 160.095 106.665 161.005 ;
        RECT 106.675 160.195 108.505 161.005 ;
        RECT 109.135 160.185 111.065 161.005 ;
        RECT 110.115 160.095 111.065 160.185 ;
        RECT 111.285 160.095 112.635 161.005 ;
        RECT 112.655 160.095 114.005 161.005 ;
        RECT 114.055 160.095 115.405 161.005 ;
        RECT 115.415 160.095 116.765 161.005 ;
        RECT 118.005 160.325 120.455 161.005 ;
        RECT 121.070 160.975 121.240 161.195 ;
        RECT 123.375 161.005 123.545 161.195 ;
        RECT 127.050 161.025 127.220 161.215 ;
        RECT 127.515 161.025 127.685 161.215 ;
        RECT 129.360 161.005 129.530 161.195 ;
        RECT 129.825 161.050 129.985 161.160 ;
        RECT 130.735 161.005 130.905 161.215 ;
        RECT 134.230 161.025 134.400 161.215 ;
        RECT 138.095 161.005 138.265 161.195 ;
        RECT 139.935 161.005 140.105 161.195 ;
        RECT 141.315 161.025 141.485 161.215 ;
        RECT 142.695 161.005 142.865 161.215 ;
        RECT 122.270 160.975 123.225 161.005 ;
        RECT 118.495 160.095 120.455 160.325 ;
        RECT 120.485 160.135 120.915 160.920 ;
        RECT 120.945 160.295 123.225 160.975 ;
        RECT 123.235 160.325 128.050 161.005 ;
        RECT 122.270 160.095 123.225 160.295 ;
        RECT 128.295 160.095 129.645 161.005 ;
        RECT 130.595 160.325 137.905 161.005 ;
        RECT 137.955 160.325 139.785 161.005 ;
        RECT 139.795 160.325 141.625 161.005 ;
        RECT 134.110 160.105 135.020 160.325 ;
        RECT 136.555 160.095 137.905 160.325 ;
        RECT 138.440 160.095 139.785 160.325 ;
        RECT 140.280 160.095 141.625 160.325 ;
        RECT 141.635 160.195 143.005 161.005 ;
      LAYER nwell ;
        RECT 17.240 156.975 143.200 159.805 ;
      LAYER pwell ;
        RECT 17.435 155.775 18.805 156.585 ;
        RECT 23.250 156.455 24.160 156.675 ;
        RECT 25.695 156.455 27.045 156.685 ;
        RECT 19.735 155.775 27.045 156.455 ;
        RECT 27.095 155.775 29.845 156.585 ;
        RECT 30.325 155.860 30.755 156.645 ;
        RECT 30.785 155.775 33.525 156.455 ;
        RECT 33.535 155.775 39.045 156.585 ;
        RECT 39.055 155.775 41.805 156.685 ;
        RECT 41.815 155.775 43.645 156.585 ;
        RECT 43.655 156.485 44.600 156.685 ;
        RECT 43.655 155.805 46.405 156.485 ;
        RECT 43.655 155.775 44.600 155.805 ;
        RECT 17.575 155.565 17.745 155.775 ;
        RECT 18.955 155.565 19.125 155.755 ;
        RECT 19.875 155.585 20.045 155.775 ;
        RECT 24.475 155.565 24.645 155.755 ;
        RECT 26.310 155.615 26.430 155.725 ;
        RECT 26.775 155.565 26.945 155.755 ;
        RECT 27.235 155.585 27.405 155.775 ;
        RECT 33.215 155.755 33.385 155.775 ;
        RECT 29.995 155.725 30.165 155.755 ;
        RECT 29.990 155.615 30.165 155.725 ;
        RECT 32.750 155.615 32.870 155.725 ;
        RECT 29.995 155.565 30.165 155.615 ;
        RECT 33.215 155.585 33.390 155.755 ;
        RECT 33.675 155.585 33.845 155.775 ;
        RECT 33.220 155.565 33.390 155.585 ;
        RECT 35.515 155.565 35.685 155.755 ;
        RECT 39.195 155.585 39.365 155.775 ;
        RECT 41.035 155.565 41.205 155.755 ;
        RECT 41.955 155.585 42.125 155.775 ;
        RECT 42.870 155.615 42.990 155.725 ;
        RECT 43.795 155.565 43.965 155.755 ;
        RECT 45.170 155.615 45.290 155.725 ;
        RECT 45.635 155.565 45.805 155.755 ;
        RECT 46.090 155.585 46.260 155.805 ;
        RECT 46.545 155.775 49.545 156.685 ;
        RECT 49.635 155.775 50.985 156.685 ;
        RECT 54.675 156.455 55.605 156.685 ;
        RECT 51.935 155.775 55.605 156.455 ;
        RECT 56.085 155.860 56.515 156.645 ;
        RECT 56.575 156.455 57.925 156.685 ;
        RECT 59.460 156.455 60.370 156.675 ;
        RECT 72.175 156.485 73.105 156.685 ;
        RECT 74.435 156.485 75.385 156.685 ;
        RECT 56.575 155.775 63.885 156.455 ;
        RECT 64.355 155.775 67.095 156.455 ;
        RECT 67.115 155.775 71.930 156.455 ;
        RECT 72.175 156.005 75.385 156.485 ;
        RECT 77.215 156.455 78.145 156.685 ;
        RECT 80.810 156.455 81.730 156.685 ;
        RECT 72.320 155.805 75.385 156.005 ;
        RECT 17.435 154.755 18.805 155.565 ;
        RECT 18.815 154.755 24.325 155.565 ;
        RECT 24.335 154.755 26.165 155.565 ;
        RECT 26.675 154.655 29.845 155.565 ;
        RECT 29.855 154.755 32.605 155.565 ;
        RECT 33.220 155.335 34.910 155.565 ;
        RECT 33.075 154.655 34.910 155.335 ;
        RECT 35.375 154.755 40.885 155.565 ;
        RECT 40.895 154.755 42.725 155.565 ;
        RECT 43.205 154.695 43.635 155.480 ;
        RECT 43.665 154.655 45.015 155.565 ;
        RECT 45.595 154.655 48.705 155.565 ;
        RECT 48.860 155.535 49.030 155.755 ;
        RECT 49.315 155.585 49.485 155.775 ;
        RECT 49.780 155.585 49.950 155.775 ;
        RECT 51.165 155.620 51.325 155.730 ;
        RECT 51.615 155.565 51.785 155.755 ;
        RECT 52.075 155.585 52.245 155.775 ;
        RECT 55.750 155.615 55.870 155.725 ;
        RECT 56.215 155.565 56.385 155.755 ;
        RECT 56.675 155.565 56.845 155.755 ;
        RECT 62.195 155.565 62.365 155.755 ;
        RECT 63.575 155.585 63.745 155.775 ;
        RECT 64.030 155.615 64.150 155.725 ;
        RECT 64.495 155.585 64.665 155.775 ;
        RECT 67.255 155.585 67.425 155.775 ;
        RECT 67.715 155.565 67.885 155.755 ;
        RECT 69.555 155.565 69.725 155.755 ;
        RECT 72.320 155.585 72.490 155.805 ;
        RECT 74.450 155.775 75.385 155.805 ;
        RECT 75.395 155.775 78.145 156.455 ;
        RECT 78.265 155.775 81.730 156.455 ;
        RECT 81.845 155.860 82.275 156.645 ;
        RECT 82.335 156.455 83.685 156.685 ;
        RECT 85.220 156.455 86.130 156.675 ;
        RECT 89.655 156.455 90.585 156.685 ;
        RECT 82.335 155.775 89.645 156.455 ;
        RECT 89.655 155.775 93.555 156.455 ;
        RECT 93.795 155.775 95.625 156.585 ;
        RECT 101.155 156.455 102.085 156.685 ;
        RECT 96.095 155.775 100.910 156.455 ;
        RECT 101.155 155.775 105.055 156.455 ;
        RECT 105.295 155.775 107.125 156.585 ;
        RECT 107.605 155.860 108.035 156.645 ;
        RECT 108.055 155.775 109.885 156.685 ;
        RECT 110.365 155.775 111.715 156.685 ;
        RECT 111.735 155.775 115.405 156.585 ;
        RECT 116.025 155.775 119.680 156.685 ;
        RECT 120.015 155.775 121.845 156.685 ;
        RECT 122.315 155.775 133.325 156.685 ;
        RECT 133.365 155.860 133.795 156.645 ;
        RECT 133.815 156.455 134.745 156.685 ;
        RECT 138.050 156.455 138.970 156.685 ;
        RECT 133.815 155.775 137.715 156.455 ;
        RECT 138.050 155.775 141.515 156.455 ;
        RECT 141.635 155.775 143.005 156.585 ;
        RECT 75.535 155.585 75.705 155.775 ;
        RECT 78.295 155.585 78.465 155.775 ;
        RECT 80.135 155.565 80.305 155.755 ;
        RECT 80.595 155.565 80.765 155.755 ;
        RECT 89.335 155.565 89.505 155.775 ;
        RECT 90.070 155.565 90.240 155.775 ;
        RECT 93.935 155.585 94.105 155.775 ;
        RECT 95.325 155.610 95.485 155.720 ;
        RECT 95.770 155.615 95.890 155.725 ;
        RECT 96.235 155.565 96.405 155.775 ;
        RECT 101.570 155.565 101.740 155.775 ;
        RECT 105.435 155.585 105.605 155.775 ;
        RECT 105.710 155.565 105.880 155.755 ;
        RECT 107.270 155.615 107.390 155.725 ;
        RECT 108.200 155.585 108.370 155.775 ;
        RECT 110.030 155.615 110.150 155.725 ;
        RECT 110.495 155.585 110.665 155.775 ;
        RECT 111.875 155.585 112.045 155.775 ;
        RECT 116.025 155.755 116.185 155.775 ;
        RECT 112.795 155.565 112.965 155.755 ;
        RECT 113.255 155.565 113.425 155.755 ;
        RECT 115.550 155.615 115.670 155.725 ;
        RECT 116.015 155.585 116.185 155.755 ;
        RECT 116.480 155.565 116.650 155.755 ;
        RECT 119.705 155.610 119.865 155.720 ;
        RECT 120.160 155.585 120.330 155.775 ;
        RECT 50.520 155.535 51.465 155.565 ;
        RECT 48.715 154.855 51.465 155.535 ;
        RECT 50.520 154.655 51.465 154.855 ;
        RECT 51.475 154.755 53.305 155.565 ;
        RECT 53.315 154.655 56.425 155.565 ;
        RECT 56.535 154.755 62.045 155.565 ;
        RECT 62.055 154.755 67.565 155.565 ;
        RECT 67.575 154.755 68.945 155.565 ;
        RECT 68.965 154.695 69.395 155.480 ;
        RECT 69.415 154.885 76.725 155.565 ;
        RECT 72.930 154.665 73.840 154.885 ;
        RECT 75.375 154.655 76.725 154.885 ;
        RECT 76.870 154.885 80.335 155.565 ;
        RECT 76.870 154.655 77.790 154.885 ;
        RECT 80.455 154.755 82.285 155.565 ;
        RECT 82.335 154.885 89.645 155.565 ;
        RECT 89.655 154.885 93.555 155.565 ;
        RECT 82.335 154.655 83.685 154.885 ;
        RECT 85.220 154.665 86.130 154.885 ;
        RECT 89.655 154.655 90.585 154.885 ;
        RECT 94.725 154.695 95.155 155.480 ;
        RECT 96.095 154.885 100.910 155.565 ;
        RECT 101.155 154.885 105.055 155.565 ;
        RECT 105.295 154.885 109.195 155.565 ;
        RECT 109.530 154.885 112.995 155.565 ;
        RECT 101.155 154.655 102.085 154.885 ;
        RECT 105.295 154.655 106.225 154.885 ;
        RECT 109.530 154.655 110.450 154.885 ;
        RECT 113.115 154.655 116.325 155.565 ;
        RECT 116.335 154.655 119.255 155.565 ;
        RECT 121.070 155.535 121.240 155.755 ;
        RECT 121.990 155.615 122.110 155.725 ;
        RECT 122.460 155.585 122.630 155.775 ;
        RECT 123.375 155.565 123.545 155.755 ;
        RECT 128.435 155.585 128.605 155.755 ;
        RECT 128.440 155.565 128.605 155.585 ;
        RECT 130.735 155.565 130.905 155.755 ;
        RECT 134.230 155.585 134.400 155.775 ;
        RECT 138.095 155.565 138.265 155.755 ;
        RECT 139.470 155.615 139.590 155.725 ;
        RECT 139.935 155.565 140.105 155.755 ;
        RECT 141.315 155.585 141.485 155.775 ;
        RECT 142.695 155.565 142.865 155.775 ;
        RECT 122.270 155.535 123.225 155.565 ;
        RECT 120.485 154.695 120.915 155.480 ;
        RECT 120.945 154.855 123.225 155.535 ;
        RECT 123.235 154.885 128.050 155.565 ;
        RECT 128.440 154.885 130.275 155.565 ;
        RECT 130.595 154.885 137.905 155.565 ;
        RECT 122.270 154.655 123.225 154.855 ;
        RECT 129.345 154.655 130.275 154.885 ;
        RECT 134.110 154.665 135.020 154.885 ;
        RECT 136.555 154.655 137.905 154.885 ;
        RECT 137.955 154.785 139.325 155.565 ;
        RECT 139.795 154.885 141.625 155.565 ;
        RECT 140.280 154.655 141.625 154.885 ;
        RECT 141.635 154.755 143.005 155.565 ;
      LAYER nwell ;
        RECT 17.240 151.535 143.200 154.365 ;
      LAYER pwell ;
        RECT 17.435 150.335 18.805 151.145 ;
        RECT 18.815 150.335 24.325 151.145 ;
        RECT 24.335 150.335 29.845 151.145 ;
        RECT 30.325 150.420 30.755 151.205 ;
        RECT 30.775 150.335 36.285 151.145 ;
        RECT 36.295 150.335 38.125 151.145 ;
        RECT 38.190 150.335 48.210 151.245 ;
        RECT 48.255 150.335 53.765 151.145 ;
        RECT 53.775 150.335 55.605 151.145 ;
        RECT 56.085 150.420 56.515 151.205 ;
        RECT 56.535 150.335 62.045 151.145 ;
        RECT 62.055 150.335 67.565 151.145 ;
        RECT 67.575 150.335 70.325 151.145 ;
        RECT 70.795 151.015 71.725 151.245 ;
        RECT 70.795 150.335 74.695 151.015 ;
        RECT 74.935 150.335 76.305 151.145 ;
        RECT 76.410 151.015 77.330 151.245 ;
        RECT 76.410 150.335 79.875 151.015 ;
        RECT 79.995 150.335 81.825 151.145 ;
        RECT 81.845 150.420 82.275 151.205 ;
        RECT 82.295 150.335 87.805 151.145 ;
        RECT 87.815 150.335 89.185 151.145 ;
        RECT 92.395 151.015 93.325 151.245 ;
        RECT 89.425 150.335 93.325 151.015 ;
        RECT 93.335 150.335 96.085 151.145 ;
        RECT 100.070 151.015 100.980 151.235 ;
        RECT 102.515 151.015 103.865 151.245 ;
        RECT 96.555 150.335 103.865 151.015 ;
        RECT 103.915 150.335 107.585 151.145 ;
        RECT 107.605 150.420 108.035 151.205 ;
        RECT 110.710 151.015 111.630 151.245 ;
        RECT 108.165 150.335 111.630 151.015 ;
        RECT 111.735 150.335 113.565 151.245 ;
        RECT 113.595 150.335 114.945 151.245 ;
        RECT 118.530 151.015 119.450 151.245 ;
        RECT 115.985 150.335 119.450 151.015 ;
        RECT 119.555 150.335 122.765 151.245 ;
        RECT 132.415 151.015 133.345 151.245 ;
        RECT 123.235 150.335 128.050 151.015 ;
        RECT 129.445 150.335 133.345 151.015 ;
        RECT 133.365 150.420 133.795 151.205 ;
        RECT 137.330 151.015 138.240 151.235 ;
        RECT 139.775 151.015 141.125 151.245 ;
        RECT 133.815 150.335 141.125 151.015 ;
        RECT 141.635 150.335 143.005 151.145 ;
        RECT 17.575 150.125 17.745 150.335 ;
        RECT 18.955 150.125 19.125 150.335 ;
        RECT 20.795 150.125 20.965 150.315 ;
        RECT 23.555 150.125 23.725 150.315 ;
        RECT 24.475 150.145 24.645 150.335 ;
        RECT 29.990 150.175 30.110 150.285 ;
        RECT 30.915 150.145 31.085 150.335 ;
        RECT 35.050 150.125 35.220 150.315 ;
        RECT 35.515 150.125 35.685 150.315 ;
        RECT 36.435 150.145 36.605 150.335 ;
        RECT 38.275 150.145 38.445 150.335 ;
        RECT 39.205 150.170 39.365 150.280 ;
        RECT 40.115 150.125 40.285 150.315 ;
        RECT 42.870 150.175 42.990 150.285 ;
        RECT 43.795 150.145 43.965 150.315 ;
        RECT 43.800 150.125 43.965 150.145 ;
        RECT 46.095 150.125 46.265 150.315 ;
        RECT 48.395 150.145 48.565 150.335 ;
        RECT 51.615 150.125 51.785 150.315 ;
        RECT 53.915 150.145 54.085 150.335 ;
        RECT 55.750 150.175 55.870 150.285 ;
        RECT 56.675 150.145 56.845 150.335 ;
        RECT 57.135 150.125 57.305 150.315 ;
        RECT 62.195 150.145 62.365 150.335 ;
        RECT 62.655 150.125 62.825 150.315 ;
        RECT 67.715 150.145 67.885 150.335 ;
        RECT 68.185 150.170 68.345 150.280 ;
        RECT 69.555 150.125 69.725 150.315 ;
        RECT 70.470 150.175 70.590 150.285 ;
        RECT 71.210 150.145 71.380 150.335 ;
        RECT 75.075 150.145 75.245 150.335 ;
        RECT 77.190 150.125 77.360 150.315 ;
        RECT 79.675 150.145 79.845 150.335 ;
        RECT 80.135 150.145 80.305 150.335 ;
        RECT 82.435 150.145 82.605 150.335 ;
        RECT 84.275 150.125 84.445 150.315 ;
        RECT 84.735 150.125 84.905 150.315 ;
        RECT 87.955 150.145 88.125 150.335 ;
        RECT 90.255 150.125 90.425 150.315 ;
        RECT 92.740 150.145 92.910 150.335 ;
        RECT 93.475 150.145 93.645 150.335 ;
        RECT 93.945 150.170 94.105 150.280 ;
        RECT 95.315 150.125 95.485 150.315 ;
        RECT 96.230 150.175 96.350 150.285 ;
        RECT 96.695 150.125 96.865 150.335 ;
        RECT 104.055 150.145 104.225 150.335 ;
        RECT 108.195 150.145 108.365 150.335 ;
        RECT 111.880 150.315 112.050 150.335 ;
        RECT 111.875 150.145 112.050 150.315 ;
        RECT 112.345 150.170 112.505 150.280 ;
        RECT 113.710 150.145 113.880 150.335 ;
        RECT 115.105 150.180 115.265 150.290 ;
        RECT 116.015 150.145 116.185 150.335 ;
        RECT 111.875 150.125 112.045 150.145 ;
        RECT 120.155 150.125 120.325 150.315 ;
        RECT 121.070 150.125 121.240 150.315 ;
        RECT 122.455 150.145 122.625 150.335 ;
        RECT 122.910 150.175 123.030 150.285 ;
        RECT 123.375 150.125 123.545 150.335 ;
        RECT 126.595 150.125 126.765 150.315 ;
        RECT 128.445 150.180 128.605 150.290 ;
        RECT 129.815 150.125 129.985 150.315 ;
        RECT 132.760 150.145 132.930 150.335 ;
        RECT 133.035 150.125 133.205 150.315 ;
        RECT 133.955 150.145 134.125 150.335 ;
        RECT 134.875 150.125 135.045 150.315 ;
        RECT 139.475 150.125 139.645 150.315 ;
        RECT 139.935 150.125 140.105 150.315 ;
        RECT 141.310 150.175 141.430 150.285 ;
        RECT 142.695 150.125 142.865 150.335 ;
        RECT 17.435 149.315 18.805 150.125 ;
        RECT 18.815 149.445 20.645 150.125 ;
        RECT 19.300 149.215 20.645 149.445 ;
        RECT 20.655 149.315 23.405 150.125 ;
        RECT 23.415 149.445 30.725 150.125 ;
        RECT 31.695 149.445 35.365 150.125 ;
        RECT 26.930 149.225 27.840 149.445 ;
        RECT 29.375 149.215 30.725 149.445 ;
        RECT 34.440 149.215 35.365 149.445 ;
        RECT 35.375 149.315 39.045 150.125 ;
        RECT 39.975 149.445 42.725 150.125 ;
        RECT 41.795 149.215 42.725 149.445 ;
        RECT 43.205 149.255 43.635 150.040 ;
        RECT 43.800 149.445 45.635 150.125 ;
        RECT 44.705 149.215 45.635 149.445 ;
        RECT 45.955 149.315 51.465 150.125 ;
        RECT 51.475 149.315 56.985 150.125 ;
        RECT 56.995 149.315 62.505 150.125 ;
        RECT 62.515 149.315 68.025 150.125 ;
        RECT 68.965 149.255 69.395 150.040 ;
        RECT 69.415 149.445 76.725 150.125 ;
        RECT 72.930 149.225 73.840 149.445 ;
        RECT 75.375 149.215 76.725 149.445 ;
        RECT 76.775 149.445 80.675 150.125 ;
        RECT 81.010 149.445 84.475 150.125 ;
        RECT 76.775 149.215 77.705 149.445 ;
        RECT 81.010 149.215 81.930 149.445 ;
        RECT 84.595 149.315 90.105 150.125 ;
        RECT 90.115 149.315 93.785 150.125 ;
        RECT 94.725 149.255 95.155 150.040 ;
        RECT 95.175 149.315 96.545 150.125 ;
        RECT 96.555 149.445 103.865 150.125 ;
        RECT 100.070 149.225 100.980 149.445 ;
        RECT 102.515 149.215 103.865 149.445 ;
        RECT 104.875 149.445 112.185 150.125 ;
        RECT 113.155 149.445 120.465 150.125 ;
        RECT 104.875 149.215 106.225 149.445 ;
        RECT 107.760 149.225 108.670 149.445 ;
        RECT 113.155 149.215 114.505 149.445 ;
        RECT 116.040 149.225 116.950 149.445 ;
        RECT 120.485 149.255 120.915 150.040 ;
        RECT 120.955 149.215 122.305 150.125 ;
        RECT 123.235 149.215 126.445 150.125 ;
        RECT 126.455 149.215 129.665 150.125 ;
        RECT 129.675 149.215 132.885 150.125 ;
        RECT 132.895 149.315 134.725 150.125 ;
        RECT 134.735 149.345 136.105 150.125 ;
        RECT 136.210 149.445 139.675 150.125 ;
        RECT 139.795 149.445 141.625 150.125 ;
        RECT 136.210 149.215 137.130 149.445 ;
        RECT 140.280 149.215 141.625 149.445 ;
        RECT 141.635 149.315 143.005 150.125 ;
      LAYER nwell ;
        RECT 17.240 146.095 143.200 148.925 ;
      LAYER pwell ;
        RECT 17.435 144.895 18.805 145.705 ;
        RECT 18.815 144.895 20.645 145.575 ;
        RECT 20.655 144.895 22.485 145.705 ;
        RECT 22.515 144.895 23.865 145.805 ;
        RECT 23.875 145.575 24.795 145.805 ;
        RECT 23.875 144.895 26.165 145.575 ;
        RECT 26.175 144.895 27.525 145.805 ;
        RECT 27.865 145.575 28.795 145.805 ;
        RECT 27.865 144.895 29.700 145.575 ;
        RECT 30.325 144.980 30.755 145.765 ;
        RECT 30.775 145.575 31.910 145.805 ;
        RECT 30.775 144.895 33.985 145.575 ;
        RECT 33.995 144.895 37.665 145.705 ;
        RECT 39.050 145.125 40.885 145.805 ;
        RECT 39.050 144.895 40.740 145.125 ;
        RECT 40.895 144.895 43.645 145.705 ;
        RECT 45.980 145.575 47.325 145.805 ;
        RECT 43.655 144.895 45.485 145.575 ;
        RECT 45.495 144.895 47.325 145.575 ;
        RECT 47.335 144.895 52.845 145.705 ;
        RECT 52.855 144.895 55.605 145.705 ;
        RECT 56.085 144.980 56.515 145.765 ;
        RECT 56.535 144.895 58.365 145.705 ;
        RECT 58.375 144.895 60.205 145.575 ;
        RECT 60.215 144.895 62.045 145.575 ;
        RECT 62.075 144.895 63.425 145.805 ;
        RECT 63.435 144.895 66.185 145.705 ;
        RECT 66.695 145.575 68.045 145.805 ;
        RECT 69.580 145.575 70.490 145.795 ;
        RECT 74.015 145.575 74.945 145.805 ;
        RECT 66.695 144.895 74.005 145.575 ;
        RECT 74.015 144.895 77.915 145.575 ;
        RECT 78.165 144.895 80.905 145.575 ;
        RECT 81.845 144.980 82.275 145.765 ;
        RECT 82.295 144.895 84.125 145.705 ;
        RECT 84.135 145.575 85.065 145.805 ;
        RECT 90.930 145.575 91.850 145.805 ;
        RECT 84.135 144.895 88.035 145.575 ;
        RECT 88.385 144.895 91.850 145.575 ;
        RECT 91.955 144.895 97.465 145.705 ;
        RECT 97.475 144.895 98.845 145.705 ;
        RECT 98.855 145.575 99.785 145.805 ;
        RECT 102.995 145.575 103.925 145.805 ;
        RECT 98.855 144.895 102.755 145.575 ;
        RECT 102.995 144.895 106.895 145.575 ;
        RECT 107.605 144.980 108.035 145.765 ;
        RECT 111.170 145.575 112.090 145.805 ;
        RECT 108.625 144.895 112.090 145.575 ;
        RECT 112.205 144.895 113.555 145.805 ;
        RECT 114.495 144.895 115.845 145.805 ;
        RECT 115.875 144.895 119.545 145.705 ;
        RECT 122.755 145.575 123.685 145.805 ;
        RECT 119.785 144.895 123.685 145.575 ;
        RECT 123.695 145.575 125.040 145.805 ;
        RECT 129.510 145.575 130.420 145.795 ;
        RECT 131.955 145.575 133.305 145.805 ;
        RECT 123.695 144.895 125.525 145.575 ;
        RECT 125.995 144.895 133.305 145.575 ;
        RECT 133.365 144.980 133.795 145.765 ;
        RECT 133.910 145.575 134.830 145.805 ;
        RECT 138.440 145.575 139.785 145.805 ;
        RECT 140.280 145.575 141.625 145.805 ;
        RECT 133.910 144.895 137.375 145.575 ;
        RECT 137.955 144.895 139.785 145.575 ;
        RECT 139.795 144.895 141.625 145.575 ;
        RECT 141.635 144.895 143.005 145.705 ;
        RECT 17.575 144.685 17.745 144.895 ;
        RECT 18.955 144.685 19.125 144.895 ;
        RECT 20.795 144.705 20.965 144.895 ;
        RECT 17.435 143.875 18.805 144.685 ;
        RECT 18.815 143.875 20.645 144.685 ;
        RECT 20.655 144.655 21.590 144.685 ;
        RECT 23.550 144.655 23.720 144.895 ;
        RECT 24.015 144.685 24.185 144.875 ;
        RECT 25.855 144.705 26.025 144.895 ;
        RECT 26.320 144.705 26.490 144.895 ;
        RECT 29.535 144.875 29.700 144.895 ;
        RECT 27.235 144.685 27.405 144.875 ;
        RECT 29.535 144.705 29.705 144.875 ;
        RECT 29.990 144.735 30.110 144.845 ;
        RECT 33.675 144.705 33.845 144.895 ;
        RECT 34.135 144.705 34.305 144.895 ;
        RECT 34.595 144.685 34.765 144.875 ;
        RECT 37.810 144.850 37.980 144.875 ;
        RECT 35.985 144.730 36.145 144.840 ;
        RECT 37.810 144.740 37.985 144.850 ;
        RECT 37.810 144.685 37.980 144.740 ;
        RECT 38.275 144.685 38.445 144.875 ;
        RECT 40.570 144.705 40.740 144.895 ;
        RECT 41.035 144.705 41.205 144.895 ;
        RECT 41.495 144.685 41.665 144.875 ;
        RECT 43.795 144.685 43.965 144.875 ;
        RECT 45.175 144.705 45.345 144.895 ;
        RECT 45.635 144.705 45.805 144.895 ;
        RECT 46.095 144.685 46.265 144.875 ;
        RECT 47.475 144.705 47.645 144.895 ;
        RECT 51.615 144.685 51.785 144.875 ;
        RECT 52.995 144.705 53.165 144.895 ;
        RECT 55.750 144.735 55.870 144.845 ;
        RECT 56.675 144.705 56.845 144.895 ;
        RECT 59.895 144.705 60.065 144.895 ;
        RECT 61.275 144.685 61.445 144.875 ;
        RECT 61.735 144.685 61.905 144.895 ;
        RECT 62.190 144.705 62.360 144.895 ;
        RECT 63.575 144.705 63.745 144.895 ;
        RECT 66.330 144.735 66.450 144.845 ;
        RECT 69.550 144.735 69.670 144.845 ;
        RECT 70.020 144.685 70.190 144.875 ;
        RECT 73.695 144.705 73.865 144.895 ;
        RECT 74.430 144.705 74.600 144.895 ;
        RECT 80.135 144.685 80.305 144.875 ;
        RECT 80.595 144.685 80.765 144.895 ;
        RECT 81.065 144.740 81.225 144.850 ;
        RECT 82.435 144.705 82.605 144.895 ;
        RECT 84.550 144.705 84.720 144.895 ;
        RECT 88.230 144.685 88.400 144.875 ;
        RECT 88.415 144.705 88.585 144.895 ;
        RECT 92.095 144.685 92.265 144.895 ;
        RECT 95.590 144.685 95.760 144.875 ;
        RECT 97.615 144.705 97.785 144.895 ;
        RECT 99.270 144.705 99.440 144.895 ;
        RECT 102.675 144.685 102.845 144.875 ;
        RECT 103.135 144.685 103.305 144.875 ;
        RECT 103.410 144.705 103.580 144.895 ;
        RECT 107.270 144.735 107.390 144.845 ;
        RECT 108.190 144.735 108.310 144.845 ;
        RECT 108.655 144.685 108.825 144.895 ;
        RECT 112.335 144.705 112.505 144.895 ;
        RECT 113.725 144.740 113.885 144.850 ;
        RECT 114.175 144.685 114.345 144.875 ;
        RECT 115.560 144.705 115.730 144.895 ;
        RECT 116.015 144.705 116.185 144.895 ;
        RECT 119.705 144.730 119.865 144.840 ;
        RECT 121.085 144.730 121.245 144.840 ;
        RECT 121.990 144.685 122.160 144.875 ;
        RECT 123.100 144.705 123.270 144.895 ;
        RECT 123.375 144.685 123.545 144.875 ;
        RECT 125.215 144.705 125.385 144.895 ;
        RECT 125.670 144.735 125.790 144.845 ;
        RECT 126.135 144.705 126.305 144.895 ;
        RECT 127.055 144.685 127.225 144.875 ;
        RECT 128.710 144.685 128.880 144.875 ;
        RECT 132.575 144.685 132.745 144.875 ;
        RECT 136.250 144.735 136.370 144.845 ;
        RECT 136.715 144.685 136.885 144.875 ;
        RECT 137.175 144.705 137.345 144.895 ;
        RECT 137.630 144.735 137.750 144.845 ;
        RECT 138.095 144.685 138.265 144.895 ;
        RECT 139.935 144.705 140.105 144.895 ;
        RECT 142.695 144.685 142.865 144.895 ;
        RECT 20.655 144.455 23.720 144.655 ;
        RECT 20.655 143.975 23.865 144.455 ;
        RECT 23.875 144.005 27.085 144.685 ;
        RECT 27.095 144.005 34.405 144.685 ;
        RECT 20.655 143.775 21.605 143.975 ;
        RECT 22.935 143.775 23.865 143.975 ;
        RECT 25.950 143.775 27.085 144.005 ;
        RECT 30.610 143.785 31.520 144.005 ;
        RECT 33.055 143.775 34.405 144.005 ;
        RECT 34.465 143.775 35.815 144.685 ;
        RECT 36.775 143.775 38.125 144.685 ;
        RECT 38.135 143.775 41.345 144.685 ;
        RECT 41.355 143.875 43.185 144.685 ;
        RECT 43.205 143.815 43.635 144.600 ;
        RECT 43.655 143.775 45.945 144.685 ;
        RECT 45.955 143.875 51.465 144.685 ;
        RECT 51.475 143.875 54.225 144.685 ;
        RECT 54.275 144.005 61.585 144.685 ;
        RECT 61.595 144.005 68.905 144.685 ;
        RECT 54.275 143.775 55.625 144.005 ;
        RECT 57.160 143.785 58.070 144.005 ;
        RECT 65.110 143.785 66.020 144.005 ;
        RECT 67.555 143.775 68.905 144.005 ;
        RECT 68.965 143.815 69.395 144.600 ;
        RECT 69.875 143.775 72.990 144.685 ;
        RECT 73.135 144.005 80.445 144.685 ;
        RECT 80.455 144.005 87.765 144.685 ;
        RECT 73.135 143.775 74.485 144.005 ;
        RECT 76.020 143.785 76.930 144.005 ;
        RECT 83.970 143.785 84.880 144.005 ;
        RECT 86.415 143.775 87.765 144.005 ;
        RECT 87.815 144.005 91.715 144.685 ;
        RECT 87.815 143.775 88.745 144.005 ;
        RECT 91.955 143.875 94.705 144.685 ;
        RECT 94.725 143.815 95.155 144.600 ;
        RECT 95.175 144.005 99.075 144.685 ;
        RECT 99.410 144.005 102.875 144.685 ;
        RECT 95.175 143.775 96.105 144.005 ;
        RECT 99.410 143.775 100.330 144.005 ;
        RECT 102.995 143.875 108.505 144.685 ;
        RECT 108.515 143.875 114.025 144.685 ;
        RECT 114.035 143.875 119.545 144.685 ;
        RECT 120.485 143.815 120.915 144.600 ;
        RECT 121.875 143.775 123.225 144.685 ;
        RECT 123.235 143.875 126.905 144.685 ;
        RECT 126.915 143.875 128.285 144.685 ;
        RECT 128.295 144.005 132.195 144.685 ;
        RECT 128.295 143.775 129.225 144.005 ;
        RECT 132.435 143.875 136.105 144.685 ;
        RECT 136.575 143.905 137.945 144.685 ;
        RECT 137.955 143.875 141.625 144.685 ;
        RECT 141.635 143.875 143.005 144.685 ;
      LAYER nwell ;
        RECT 17.240 140.655 143.200 143.485 ;
      LAYER pwell ;
        RECT 17.435 139.455 18.805 140.265 ;
        RECT 18.815 139.455 20.645 140.265 ;
        RECT 24.170 140.135 25.080 140.355 ;
        RECT 26.615 140.135 27.965 140.365 ;
        RECT 20.655 139.455 27.965 140.135 ;
        RECT 28.215 140.275 29.165 140.365 ;
        RECT 28.215 139.455 30.145 140.275 ;
        RECT 30.325 139.540 30.755 140.325 ;
        RECT 30.775 139.455 32.125 140.365 ;
        RECT 32.155 140.165 33.085 140.365 ;
        RECT 34.420 140.165 35.365 140.365 ;
        RECT 32.155 139.685 35.365 140.165 ;
        RECT 32.295 139.485 35.365 139.685 ;
        RECT 17.575 139.245 17.745 139.455 ;
        RECT 18.955 139.265 19.125 139.455 ;
        RECT 19.875 139.245 20.045 139.435 ;
        RECT 20.795 139.265 20.965 139.455 ;
        RECT 29.995 139.435 30.145 139.455 ;
        RECT 27.240 139.245 27.410 139.435 ;
        RECT 28.620 139.245 28.790 139.435 ;
        RECT 29.995 139.245 30.165 139.435 ;
        RECT 31.840 139.265 32.010 139.455 ;
        RECT 32.295 139.265 32.465 139.485 ;
        RECT 34.420 139.455 35.365 139.485 ;
        RECT 35.570 139.455 39.045 140.365 ;
        RECT 39.055 140.165 40.005 140.365 ;
        RECT 41.335 140.165 42.265 140.365 ;
        RECT 39.055 139.685 42.265 140.165 ;
        RECT 39.055 139.485 42.120 139.685 ;
        RECT 39.055 139.455 39.990 139.485 ;
        RECT 38.730 139.435 38.900 139.455 ;
        RECT 35.525 139.290 35.685 139.400 ;
        RECT 36.435 139.245 36.605 139.435 ;
        RECT 38.730 139.265 38.910 139.435 ;
        RECT 41.950 139.265 42.120 139.485 ;
        RECT 42.335 139.455 44.105 140.365 ;
        RECT 44.115 139.455 46.865 140.265 ;
        RECT 47.345 139.455 50.075 140.365 ;
        RECT 50.095 139.455 53.765 140.265 ;
        RECT 55.145 140.135 56.065 140.365 ;
        RECT 53.775 139.455 56.065 140.135 ;
        RECT 56.085 139.540 56.515 140.325 ;
        RECT 60.050 140.135 60.960 140.355 ;
        RECT 62.495 140.135 63.845 140.365 ;
        RECT 56.535 139.455 63.845 140.135 ;
        RECT 63.895 139.455 67.565 140.265 ;
        RECT 69.865 140.135 70.785 140.365 ;
        RECT 68.495 139.455 70.785 140.135 ;
        RECT 70.795 139.455 77.905 140.365 ;
        RECT 78.250 140.135 79.170 140.365 ;
        RECT 78.250 139.455 81.715 140.135 ;
        RECT 81.845 139.540 82.275 140.325 ;
        RECT 83.255 140.135 84.605 140.365 ;
        RECT 86.140 140.135 87.050 140.355 ;
        RECT 94.090 140.135 95.000 140.355 ;
        RECT 96.535 140.135 97.885 140.365 ;
        RECT 102.370 140.135 103.280 140.355 ;
        RECT 104.815 140.135 106.165 140.365 ;
        RECT 83.255 139.455 90.565 140.135 ;
        RECT 90.575 139.455 97.885 140.135 ;
        RECT 98.855 139.455 106.165 140.135 ;
        RECT 106.215 139.455 107.585 140.265 ;
        RECT 107.605 139.540 108.035 140.325 ;
        RECT 108.150 140.135 109.070 140.365 ;
        RECT 111.830 140.135 112.750 140.365 ;
        RECT 108.150 139.455 111.615 140.135 ;
        RECT 111.830 139.455 115.295 140.135 ;
        RECT 115.610 139.455 119.085 140.365 ;
        RECT 119.405 140.135 120.335 140.365 ;
        RECT 119.405 139.455 121.240 140.135 ;
        RECT 121.395 139.455 126.905 140.265 ;
        RECT 126.915 139.455 132.425 140.265 ;
        RECT 133.365 139.540 133.795 140.325 ;
        RECT 137.330 140.135 138.240 140.355 ;
        RECT 139.775 140.135 141.125 140.365 ;
        RECT 133.815 139.455 141.125 140.135 ;
        RECT 141.635 139.455 143.005 140.265 ;
        RECT 43.790 139.435 43.960 139.455 ;
        RECT 38.740 139.245 38.910 139.265 ;
        RECT 42.415 139.245 42.585 139.435 ;
        RECT 42.870 139.295 42.990 139.405 ;
        RECT 43.790 139.265 43.965 139.435 ;
        RECT 44.255 139.265 44.425 139.455 ;
        RECT 43.795 139.245 43.965 139.265 ;
        RECT 46.095 139.245 46.265 139.435 ;
        RECT 47.010 139.295 47.130 139.405 ;
        RECT 47.480 139.245 47.650 139.435 ;
        RECT 49.775 139.265 49.945 139.455 ;
        RECT 50.235 139.265 50.405 139.455 ;
        RECT 53.450 139.245 53.620 139.435 ;
        RECT 53.915 139.265 54.085 139.455 ;
        RECT 54.840 139.245 55.010 139.435 ;
        RECT 56.675 139.265 56.845 139.455 ;
        RECT 58.510 139.245 58.680 139.435 ;
        RECT 58.975 139.245 59.145 139.435 ;
        RECT 61.280 139.245 61.450 139.435 ;
        RECT 62.655 139.245 62.825 139.435 ;
        RECT 64.035 139.265 64.205 139.455 ;
        RECT 67.725 139.300 67.885 139.410 ;
        RECT 68.185 139.290 68.345 139.400 ;
        RECT 68.635 139.265 68.805 139.455 ;
        RECT 69.555 139.245 69.725 139.435 ;
        RECT 17.435 138.435 18.805 139.245 ;
        RECT 19.735 138.565 27.045 139.245 ;
        RECT 23.250 138.345 24.160 138.565 ;
        RECT 25.695 138.335 27.045 138.565 ;
        RECT 27.095 138.335 28.445 139.245 ;
        RECT 28.475 138.335 29.825 139.245 ;
        RECT 29.855 138.435 35.365 139.245 ;
        RECT 36.305 138.335 37.655 139.245 ;
        RECT 37.675 138.335 39.025 139.245 ;
        RECT 39.055 138.335 42.725 139.245 ;
        RECT 43.205 138.375 43.635 139.160 ;
        RECT 43.655 138.565 45.945 139.245 ;
        RECT 45.025 138.335 45.945 138.565 ;
        RECT 45.955 138.435 47.325 139.245 ;
        RECT 47.335 138.335 51.725 139.245 ;
        RECT 51.935 138.335 53.765 139.245 ;
        RECT 53.775 138.335 55.125 139.245 ;
        RECT 55.350 138.335 58.825 139.245 ;
        RECT 58.835 138.565 61.125 139.245 ;
        RECT 60.205 138.335 61.125 138.565 ;
        RECT 61.135 138.335 62.485 139.245 ;
        RECT 62.515 138.435 68.025 139.245 ;
        RECT 68.965 138.375 69.395 139.160 ;
        RECT 69.415 138.435 70.785 139.245 ;
        RECT 70.940 139.215 71.110 139.455 ;
        RECT 74.155 139.245 74.325 139.435 ;
        RECT 77.375 139.245 77.545 139.435 ;
        RECT 77.830 139.295 77.950 139.405 ;
        RECT 78.295 139.245 78.465 139.435 ;
        RECT 81.515 139.265 81.685 139.455 ;
        RECT 82.445 139.300 82.605 139.410 ;
        RECT 87.495 139.245 87.665 139.435 ;
        RECT 90.255 139.265 90.425 139.455 ;
        RECT 90.715 139.265 90.885 139.455 ;
        RECT 95.315 139.245 95.485 139.435 ;
        RECT 97.150 139.295 97.270 139.405 ;
        RECT 97.615 139.245 97.785 139.435 ;
        RECT 98.085 139.300 98.245 139.410 ;
        RECT 98.995 139.265 99.165 139.455 ;
        RECT 105.250 139.245 105.420 139.435 ;
        RECT 106.355 139.265 106.525 139.455 ;
        RECT 109.390 139.245 109.560 139.435 ;
        RECT 111.415 139.265 111.585 139.455 ;
        RECT 113.255 139.245 113.425 139.435 ;
        RECT 115.095 139.265 115.265 139.455 ;
        RECT 118.770 139.265 118.940 139.455 ;
        RECT 121.075 139.435 121.240 139.455 ;
        RECT 121.075 139.245 121.245 139.435 ;
        RECT 121.535 139.265 121.705 139.455 ;
        RECT 127.055 139.265 127.225 139.455 ;
        RECT 128.435 139.245 128.605 139.435 ;
        RECT 132.585 139.300 132.745 139.410 ;
        RECT 133.490 139.245 133.660 139.435 ;
        RECT 133.955 139.265 134.125 139.455 ;
        RECT 133.960 139.245 134.125 139.265 ;
        RECT 136.255 139.245 136.425 139.435 ;
        RECT 138.095 139.245 138.265 139.435 ;
        RECT 139.935 139.245 140.105 139.435 ;
        RECT 141.310 139.295 141.430 139.405 ;
        RECT 142.695 139.245 142.865 139.455 ;
        RECT 73.070 139.215 74.005 139.245 ;
        RECT 70.940 139.015 74.005 139.215 ;
        RECT 70.795 138.535 74.005 139.015 ;
        RECT 74.015 138.565 76.305 139.245 ;
        RECT 70.795 138.335 71.725 138.535 ;
        RECT 73.055 138.335 74.005 138.535 ;
        RECT 75.385 138.335 76.305 138.565 ;
        RECT 76.325 138.335 77.675 139.245 ;
        RECT 78.155 138.565 87.260 139.245 ;
        RECT 87.355 138.565 94.665 139.245 ;
        RECT 90.870 138.345 91.780 138.565 ;
        RECT 93.315 138.335 94.665 138.565 ;
        RECT 94.725 138.375 95.155 139.160 ;
        RECT 95.175 138.435 97.005 139.245 ;
        RECT 97.475 138.565 104.785 139.245 ;
        RECT 100.990 138.345 101.900 138.565 ;
        RECT 103.435 138.335 104.785 138.565 ;
        RECT 104.835 138.565 108.735 139.245 ;
        RECT 108.975 138.565 112.875 139.245 ;
        RECT 113.115 138.565 120.425 139.245 ;
        RECT 104.835 138.335 105.765 138.565 ;
        RECT 108.975 138.335 109.905 138.565 ;
        RECT 116.630 138.345 117.540 138.565 ;
        RECT 119.075 138.335 120.425 138.565 ;
        RECT 120.485 138.375 120.915 139.160 ;
        RECT 120.935 138.565 128.245 139.245 ;
        RECT 124.450 138.345 125.360 138.565 ;
        RECT 126.895 138.335 128.245 138.565 ;
        RECT 128.295 138.435 130.125 139.245 ;
        RECT 130.330 138.335 133.805 139.245 ;
        RECT 133.960 138.565 135.795 139.245 ;
        RECT 134.865 138.335 135.795 138.565 ;
        RECT 136.115 138.435 137.945 139.245 ;
        RECT 137.955 138.565 139.785 139.245 ;
        RECT 139.795 138.565 141.625 139.245 ;
        RECT 138.440 138.335 139.785 138.565 ;
        RECT 140.280 138.335 141.625 138.565 ;
        RECT 141.635 138.435 143.005 139.245 ;
      LAYER nwell ;
        RECT 17.240 135.215 143.200 138.045 ;
      LAYER pwell ;
        RECT 17.435 134.015 18.805 134.825 ;
        RECT 18.815 134.015 22.485 134.825 ;
        RECT 22.495 134.695 23.415 134.925 ;
        RECT 22.495 134.015 24.785 134.695 ;
        RECT 24.795 134.015 30.305 134.825 ;
        RECT 30.325 134.100 30.755 134.885 ;
        RECT 30.775 134.015 36.285 134.825 ;
        RECT 36.295 134.015 37.665 134.825 ;
        RECT 37.685 134.015 41.345 134.925 ;
        RECT 42.495 134.835 43.445 134.925 ;
        RECT 41.515 134.015 43.445 134.835 ;
        RECT 43.655 134.015 46.405 134.825 ;
        RECT 46.415 134.725 47.360 134.925 ;
        RECT 46.415 134.045 49.165 134.725 ;
        RECT 49.175 134.695 50.105 134.925 ;
        RECT 46.415 134.015 47.360 134.045 ;
        RECT 17.575 133.805 17.745 134.015 ;
        RECT 18.955 133.805 19.125 134.015 ;
        RECT 24.475 133.805 24.645 134.015 ;
        RECT 24.935 133.825 25.105 134.015 ;
        RECT 27.230 133.805 27.400 133.995 ;
        RECT 27.695 133.805 27.865 133.995 ;
        RECT 30.915 133.825 31.085 134.015 ;
        RECT 33.215 133.805 33.385 133.995 ;
        RECT 36.435 133.825 36.605 134.015 ;
        RECT 36.890 133.855 37.010 133.965 ;
        RECT 37.810 133.825 37.980 134.015 ;
        RECT 41.515 133.995 41.665 134.015 ;
        RECT 38.730 133.805 38.900 133.995 ;
        RECT 40.575 133.805 40.745 133.995 ;
        RECT 41.035 133.805 41.205 133.995 ;
        RECT 41.495 133.825 41.665 133.995 ;
        RECT 42.870 133.855 42.990 133.965 ;
        RECT 43.795 133.805 43.965 134.015 ;
        RECT 48.850 133.825 49.020 134.045 ;
        RECT 49.175 134.015 52.845 134.695 ;
        RECT 52.855 134.015 56.065 134.925 ;
        RECT 56.085 134.100 56.515 134.885 ;
        RECT 56.535 134.015 58.350 134.925 ;
        RECT 72.375 134.835 73.325 134.925 ;
        RECT 58.375 134.015 63.885 134.825 ;
        RECT 63.895 134.015 69.405 134.825 ;
        RECT 69.415 134.015 72.165 134.825 ;
        RECT 72.375 134.015 74.305 134.835 ;
        RECT 74.475 134.015 77.225 134.825 ;
        RECT 80.895 134.695 81.825 134.925 ;
        RECT 77.925 134.015 81.825 134.695 ;
        RECT 81.845 134.100 82.275 134.885 ;
        RECT 82.295 134.015 85.965 134.825 ;
        RECT 89.175 134.695 90.105 134.925 ;
        RECT 86.205 134.015 90.105 134.695 ;
        RECT 90.210 134.695 91.130 134.925 ;
        RECT 90.210 134.015 93.675 134.695 ;
        RECT 93.795 134.015 97.465 134.825 ;
        RECT 100.990 134.695 101.900 134.915 ;
        RECT 103.435 134.695 104.785 134.925 ;
        RECT 97.475 134.015 104.785 134.695 ;
        RECT 104.835 134.015 107.585 134.825 ;
        RECT 107.605 134.100 108.035 134.885 ;
        RECT 108.150 134.695 109.070 134.925 ;
        RECT 108.150 134.015 111.615 134.695 ;
        RECT 112.655 134.015 116.130 134.925 ;
        RECT 119.850 134.695 120.760 134.915 ;
        RECT 122.295 134.695 123.645 134.925 ;
        RECT 124.745 134.695 125.675 134.925 ;
        RECT 116.335 134.015 123.645 134.695 ;
        RECT 123.840 134.015 125.675 134.695 ;
        RECT 125.995 134.015 127.365 134.825 ;
        RECT 128.425 134.695 129.355 134.925 ;
        RECT 127.520 134.015 129.355 134.695 ;
        RECT 129.870 134.015 133.345 134.925 ;
        RECT 133.365 134.100 133.795 134.885 ;
        RECT 137.330 134.695 138.240 134.915 ;
        RECT 139.775 134.695 141.125 134.925 ;
        RECT 133.815 134.015 141.125 134.695 ;
        RECT 141.635 134.015 143.005 134.825 ;
        RECT 49.325 133.850 49.485 133.960 ;
        RECT 50.235 133.825 50.405 133.995 ;
        RECT 52.535 133.825 52.705 134.015 ;
        RECT 52.995 133.825 53.165 134.015 ;
        RECT 54.375 133.825 54.545 133.995 ;
        RECT 54.845 133.850 55.005 133.960 ;
        RECT 50.240 133.805 50.405 133.825 ;
        RECT 54.375 133.805 54.540 133.825 ;
        RECT 55.755 133.805 55.925 133.995 ;
        RECT 58.055 133.825 58.225 134.015 ;
        RECT 58.515 133.825 58.685 134.015 ;
        RECT 64.035 133.825 64.205 134.015 ;
        RECT 64.955 133.805 65.125 133.995 ;
        RECT 65.415 133.805 65.585 133.995 ;
        RECT 69.555 133.825 69.725 134.015 ;
        RECT 74.155 133.995 74.305 134.015 ;
        RECT 70.475 133.805 70.645 133.995 ;
        RECT 74.155 133.825 74.325 133.995 ;
        RECT 74.615 133.825 74.785 134.015 ;
        RECT 77.370 133.855 77.490 133.965 ;
        RECT 77.835 133.805 78.005 133.995 ;
        RECT 81.240 133.825 81.410 134.015 ;
        RECT 82.435 133.825 82.605 134.015 ;
        RECT 83.355 133.805 83.525 133.995 ;
        RECT 88.875 133.805 89.045 133.995 ;
        RECT 89.520 133.825 89.690 134.015 ;
        RECT 93.475 133.825 93.645 134.015 ;
        RECT 93.935 133.825 94.105 134.015 ;
        RECT 94.390 133.855 94.510 133.965 ;
        RECT 95.315 133.805 95.485 133.995 ;
        RECT 97.615 133.825 97.785 134.015 ;
        RECT 100.830 133.855 100.950 133.965 ;
        RECT 101.570 133.805 101.740 133.995 ;
        RECT 104.975 133.825 105.145 134.015 ;
        RECT 105.435 133.805 105.605 133.995 ;
        RECT 109.110 133.855 109.230 133.965 ;
        RECT 109.565 133.805 109.735 133.995 ;
        RECT 111.415 133.825 111.585 134.015 ;
        RECT 112.800 133.995 112.970 134.015 ;
        RECT 111.885 133.860 112.045 133.970 ;
        RECT 112.795 133.825 112.970 133.995 ;
        RECT 116.475 133.825 116.645 134.015 ;
        RECT 123.840 133.995 124.005 134.015 ;
        RECT 112.795 133.805 112.965 133.825 ;
        RECT 117.850 133.805 118.020 133.995 ;
        RECT 120.155 133.825 120.325 133.995 ;
        RECT 120.155 133.805 120.320 133.825 ;
        RECT 121.075 133.805 121.245 133.995 ;
        RECT 123.835 133.825 124.005 133.995 ;
        RECT 126.135 133.825 126.305 134.015 ;
        RECT 127.520 133.995 127.685 134.015 ;
        RECT 126.595 133.805 126.765 133.995 ;
        RECT 127.515 133.825 127.685 133.995 ;
        RECT 128.430 133.855 128.550 133.965 ;
        RECT 131.655 133.805 131.825 133.995 ;
        RECT 132.115 133.805 132.285 133.995 ;
        RECT 133.030 133.825 133.200 134.015 ;
        RECT 133.955 133.825 134.125 134.015 ;
        RECT 139.470 133.855 139.590 133.965 ;
        RECT 139.935 133.805 140.105 133.995 ;
        RECT 141.310 133.855 141.430 133.965 ;
        RECT 142.695 133.805 142.865 134.015 ;
        RECT 17.435 132.995 18.805 133.805 ;
        RECT 18.815 132.995 24.325 133.805 ;
        RECT 24.335 132.995 26.165 133.805 ;
        RECT 26.195 132.895 27.545 133.805 ;
        RECT 27.555 132.995 33.065 133.805 ;
        RECT 33.075 132.995 36.745 133.805 ;
        RECT 37.215 132.895 39.045 133.805 ;
        RECT 39.055 132.895 40.870 133.805 ;
        RECT 40.895 132.995 42.725 133.805 ;
        RECT 43.205 132.935 43.635 133.720 ;
        RECT 43.655 132.995 49.165 133.805 ;
        RECT 50.240 133.125 52.075 133.805 ;
        RECT 51.145 132.895 52.075 133.125 ;
        RECT 52.705 133.125 54.540 133.805 ;
        RECT 55.615 133.125 57.905 133.805 ;
        RECT 52.705 132.895 53.635 133.125 ;
        RECT 56.985 132.895 57.905 133.125 ;
        RECT 57.955 133.125 65.265 133.805 ;
        RECT 57.955 132.895 59.305 133.125 ;
        RECT 60.840 132.905 61.750 133.125 ;
        RECT 65.275 132.995 68.945 133.805 ;
        RECT 68.965 132.935 69.395 133.720 ;
        RECT 70.335 133.125 77.645 133.805 ;
        RECT 73.850 132.905 74.760 133.125 ;
        RECT 76.295 132.895 77.645 133.125 ;
        RECT 77.695 132.995 83.205 133.805 ;
        RECT 83.215 132.995 88.725 133.805 ;
        RECT 88.735 132.995 94.245 133.805 ;
        RECT 94.725 132.935 95.155 133.720 ;
        RECT 95.175 132.995 100.685 133.805 ;
        RECT 101.155 133.125 105.055 133.805 ;
        RECT 101.155 132.895 102.085 133.125 ;
        RECT 105.295 132.995 108.965 133.805 ;
        RECT 109.435 132.895 112.645 133.805 ;
        RECT 112.655 132.995 114.485 133.805 ;
        RECT 114.690 132.895 118.165 133.805 ;
        RECT 118.485 133.125 120.320 133.805 ;
        RECT 118.485 132.895 119.415 133.125 ;
        RECT 120.485 132.935 120.915 133.720 ;
        RECT 120.935 132.995 126.445 133.805 ;
        RECT 126.455 132.995 128.285 133.805 ;
        RECT 128.755 132.895 131.965 133.805 ;
        RECT 131.975 133.125 139.285 133.805 ;
        RECT 139.795 133.125 141.625 133.805 ;
        RECT 135.490 132.905 136.400 133.125 ;
        RECT 137.935 132.895 139.285 133.125 ;
        RECT 140.280 132.895 141.625 133.125 ;
        RECT 141.635 132.995 143.005 133.805 ;
      LAYER nwell ;
        RECT 17.240 129.775 143.200 132.605 ;
      LAYER pwell ;
        RECT 17.435 128.575 18.805 129.385 ;
        RECT 18.815 128.575 22.485 129.385 ;
        RECT 22.495 129.255 23.630 129.485 ;
        RECT 26.025 129.255 26.955 129.485 ;
        RECT 28.015 129.255 28.935 129.485 ;
        RECT 22.495 128.575 25.705 129.255 ;
        RECT 26.025 128.575 27.860 129.255 ;
        RECT 28.015 128.575 30.305 129.255 ;
        RECT 30.325 128.660 30.755 129.445 ;
        RECT 30.775 128.575 32.125 129.485 ;
        RECT 32.155 128.575 37.665 129.385 ;
        RECT 37.690 128.575 39.505 129.485 ;
        RECT 39.515 128.575 45.025 129.385 ;
        RECT 45.035 128.575 50.545 129.385 ;
        RECT 50.555 128.575 53.305 129.385 ;
        RECT 53.315 128.575 54.665 129.485 ;
        RECT 54.695 128.575 56.045 129.485 ;
        RECT 56.085 128.660 56.515 129.445 ;
        RECT 56.535 128.575 59.705 129.485 ;
        RECT 59.755 128.575 65.265 129.385 ;
        RECT 65.275 128.575 68.025 129.385 ;
        RECT 72.010 129.255 72.920 129.475 ;
        RECT 74.455 129.255 76.225 129.485 ;
        RECT 68.495 128.575 76.225 129.255 ;
        RECT 76.315 129.255 77.245 129.485 ;
        RECT 76.315 128.575 80.215 129.255 ;
        RECT 80.455 128.575 81.825 129.385 ;
        RECT 81.845 128.660 82.275 129.445 ;
        RECT 85.810 129.255 86.720 129.475 ;
        RECT 88.255 129.255 90.025 129.485 ;
        RECT 82.295 128.575 90.025 129.255 ;
        RECT 90.115 129.255 91.045 129.485 ;
        RECT 90.115 128.575 94.015 129.255 ;
        RECT 94.255 128.575 97.925 129.385 ;
        RECT 98.395 129.255 99.325 129.485 ;
        RECT 102.630 129.255 103.550 129.485 ;
        RECT 98.395 128.575 102.295 129.255 ;
        RECT 102.630 128.575 106.095 129.255 ;
        RECT 106.215 128.575 107.585 129.385 ;
        RECT 107.605 128.660 108.035 129.445 ;
        RECT 108.055 128.575 110.805 129.385 ;
        RECT 111.275 128.575 114.485 129.485 ;
        RECT 114.495 128.575 117.705 129.485 ;
        RECT 118.025 129.255 118.955 129.485 ;
        RECT 118.025 128.575 119.860 129.255 ;
        RECT 120.015 128.575 121.845 129.385 ;
        RECT 121.855 128.575 125.065 129.485 ;
        RECT 125.075 128.575 130.585 129.385 ;
        RECT 132.105 129.255 133.035 129.485 ;
        RECT 131.200 128.575 133.035 129.255 ;
        RECT 133.365 128.660 133.795 129.445 ;
        RECT 134.010 128.575 137.485 129.485 ;
        RECT 137.495 128.575 140.705 129.485 ;
        RECT 141.635 128.575 143.005 129.385 ;
        RECT 17.575 128.365 17.745 128.575 ;
        RECT 18.955 128.555 19.125 128.575 ;
        RECT 18.950 128.385 19.125 128.555 ;
        RECT 18.950 128.365 19.120 128.385 ;
        RECT 20.335 128.365 20.505 128.555 ;
        RECT 25.395 128.385 25.565 128.575 ;
        RECT 27.695 128.555 27.860 128.575 ;
        RECT 27.695 128.385 27.865 128.555 ;
        RECT 29.535 128.365 29.705 128.555 ;
        RECT 29.995 128.365 30.165 128.575 ;
        RECT 30.920 128.385 31.090 128.575 ;
        RECT 32.295 128.385 32.465 128.575 ;
        RECT 34.595 128.365 34.765 128.555 ;
        RECT 37.355 128.365 37.525 128.555 ;
        RECT 37.815 128.385 37.985 128.575 ;
        RECT 39.655 128.385 39.825 128.575 ;
        RECT 40.575 128.365 40.745 128.555 ;
        RECT 41.035 128.365 41.205 128.555 ;
        RECT 42.870 128.415 42.990 128.525 ;
        RECT 43.795 128.365 43.965 128.555 ;
        RECT 45.175 128.385 45.345 128.575 ;
        RECT 49.325 128.410 49.485 128.520 ;
        RECT 50.235 128.365 50.405 128.555 ;
        RECT 50.695 128.385 50.865 128.575 ;
        RECT 53.460 128.385 53.630 128.575 ;
        RECT 54.840 128.385 55.010 128.575 ;
        RECT 59.435 128.385 59.605 128.575 ;
        RECT 59.895 128.385 60.065 128.575 ;
        RECT 60.355 128.365 60.525 128.555 ;
        RECT 60.815 128.365 60.985 128.555 ;
        RECT 65.415 128.385 65.585 128.575 ;
        RECT 66.335 128.365 66.505 128.555 ;
        RECT 68.170 128.415 68.290 128.525 ;
        RECT 68.635 128.385 68.805 128.575 ;
        RECT 69.555 128.365 69.725 128.555 ;
        RECT 76.730 128.385 76.900 128.575 ;
        RECT 76.920 128.365 77.090 128.555 ;
        RECT 17.435 127.555 18.805 128.365 ;
        RECT 18.835 127.455 20.185 128.365 ;
        RECT 20.195 127.685 27.505 128.365 ;
        RECT 23.710 127.465 24.620 127.685 ;
        RECT 26.155 127.455 27.505 127.685 ;
        RECT 27.555 127.685 29.845 128.365 ;
        RECT 29.855 127.685 33.065 128.365 ;
        RECT 27.555 127.455 28.475 127.685 ;
        RECT 31.930 127.455 33.065 127.685 ;
        RECT 33.075 127.455 34.890 128.365 ;
        RECT 34.915 127.455 37.665 128.365 ;
        RECT 37.675 127.455 40.885 128.365 ;
        RECT 40.895 127.555 42.725 128.365 ;
        RECT 43.205 127.495 43.635 128.280 ;
        RECT 43.655 127.555 49.165 128.365 ;
        RECT 50.095 127.685 53.305 128.365 ;
        RECT 52.170 127.455 53.305 127.685 ;
        RECT 53.355 127.685 60.665 128.365 ;
        RECT 53.355 127.455 54.705 127.685 ;
        RECT 56.240 127.465 57.150 127.685 ;
        RECT 60.675 127.555 66.185 128.365 ;
        RECT 66.195 127.555 68.945 128.365 ;
        RECT 68.965 127.495 69.395 128.280 ;
        RECT 69.415 127.685 76.725 128.365 ;
        RECT 72.930 127.465 73.840 127.685 ;
        RECT 75.375 127.455 76.725 127.685 ;
        RECT 76.775 127.455 78.125 128.365 ;
        RECT 78.300 128.335 78.470 128.555 ;
        RECT 80.595 128.385 80.765 128.575 ;
        RECT 82.435 128.385 82.605 128.575 ;
        RECT 84.920 128.365 85.090 128.555 ;
        RECT 85.655 128.365 85.825 128.555 ;
        RECT 90.530 128.385 90.700 128.575 ;
        RECT 93.475 128.365 93.645 128.555 ;
        RECT 94.395 128.385 94.565 128.575 ;
        RECT 95.315 128.365 95.485 128.555 ;
        RECT 97.155 128.365 97.325 128.555 ;
        RECT 98.070 128.415 98.190 128.525 ;
        RECT 98.810 128.385 98.980 128.575 ;
        RECT 104.790 128.365 104.960 128.555 ;
        RECT 105.895 128.385 106.065 128.575 ;
        RECT 106.355 128.385 106.525 128.575 ;
        RECT 108.195 128.385 108.365 128.575 ;
        RECT 108.655 128.365 108.825 128.555 ;
        RECT 110.035 128.365 110.205 128.555 ;
        RECT 110.950 128.415 111.070 128.525 ;
        RECT 111.405 128.385 111.575 128.575 ;
        RECT 114.625 128.385 114.795 128.575 ;
        RECT 119.695 128.555 119.860 128.575 ;
        RECT 117.395 128.365 117.565 128.555 ;
        RECT 119.695 128.385 119.865 128.555 ;
        RECT 120.155 128.525 120.325 128.575 ;
        RECT 120.150 128.415 120.325 128.525 ;
        RECT 120.155 128.385 120.325 128.415 ;
        RECT 121.075 128.365 121.245 128.555 ;
        RECT 124.755 128.385 124.925 128.575 ;
        RECT 125.215 128.385 125.385 128.575 ;
        RECT 131.200 128.555 131.365 128.575 ;
        RECT 128.435 128.365 128.605 128.555 ;
        RECT 130.730 128.415 130.850 128.525 ;
        RECT 131.195 128.365 131.365 128.555 ;
        RECT 137.170 128.385 137.340 128.575 ;
        RECT 138.555 128.365 138.725 128.555 ;
        RECT 139.935 128.365 140.105 128.555 ;
        RECT 140.395 128.385 140.565 128.575 ;
        RECT 140.865 128.420 141.025 128.530 ;
        RECT 142.695 128.365 142.865 128.575 ;
        RECT 80.430 128.335 81.365 128.365 ;
        RECT 78.300 128.135 81.365 128.335 ;
        RECT 78.155 127.655 81.365 128.135 ;
        RECT 81.605 127.685 85.505 128.365 ;
        RECT 85.515 127.685 93.245 128.365 ;
        RECT 78.155 127.455 79.085 127.655 ;
        RECT 80.415 127.455 81.365 127.655 ;
        RECT 84.575 127.455 85.505 127.685 ;
        RECT 89.030 127.465 89.940 127.685 ;
        RECT 91.475 127.455 93.245 127.685 ;
        RECT 93.335 127.555 94.705 128.365 ;
        RECT 94.725 127.495 95.155 128.280 ;
        RECT 95.175 127.555 97.005 128.365 ;
        RECT 97.015 127.685 104.325 128.365 ;
        RECT 100.530 127.465 101.440 127.685 ;
        RECT 102.975 127.455 104.325 127.685 ;
        RECT 104.375 127.685 108.275 128.365 ;
        RECT 104.375 127.455 105.305 127.685 ;
        RECT 108.515 127.555 109.885 128.365 ;
        RECT 109.895 127.685 117.205 128.365 ;
        RECT 117.255 127.685 119.995 128.365 ;
        RECT 113.410 127.465 114.320 127.685 ;
        RECT 115.855 127.455 117.205 127.685 ;
        RECT 120.485 127.495 120.915 128.280 ;
        RECT 120.935 127.685 128.245 128.365 ;
        RECT 124.450 127.465 125.360 127.685 ;
        RECT 126.895 127.455 128.245 127.685 ;
        RECT 128.295 127.555 131.045 128.365 ;
        RECT 131.055 127.685 138.365 128.365 ;
        RECT 134.570 127.465 135.480 127.685 ;
        RECT 137.015 127.455 138.365 127.685 ;
        RECT 138.415 127.555 139.785 128.365 ;
        RECT 139.795 127.685 141.625 128.365 ;
        RECT 140.280 127.455 141.625 127.685 ;
        RECT 141.635 127.555 143.005 128.365 ;
      LAYER nwell ;
        RECT 17.240 124.335 143.200 127.165 ;
      LAYER pwell ;
        RECT 17.435 123.135 18.805 123.945 ;
        RECT 18.815 123.135 21.565 123.945 ;
        RECT 25.550 123.815 26.460 124.035 ;
        RECT 27.995 123.815 29.345 124.045 ;
        RECT 22.035 123.135 29.345 123.815 ;
        RECT 30.325 123.220 30.755 124.005 ;
        RECT 32.145 123.815 33.065 124.045 ;
        RECT 30.775 123.135 33.065 123.815 ;
        RECT 33.075 123.135 34.425 124.045 ;
        RECT 35.415 123.135 38.585 124.045 ;
        RECT 42.110 123.815 43.020 124.035 ;
        RECT 44.555 123.815 45.905 124.045 ;
        RECT 38.595 123.135 45.905 123.815 ;
        RECT 45.955 123.135 47.770 124.045 ;
        RECT 49.165 123.815 50.085 124.045 ;
        RECT 51.465 123.815 52.385 124.045 ;
        RECT 47.795 123.135 50.085 123.815 ;
        RECT 50.095 123.135 52.385 123.815 ;
        RECT 52.395 123.135 53.745 124.045 ;
        RECT 55.145 123.815 56.065 124.045 ;
        RECT 53.775 123.135 56.065 123.815 ;
        RECT 56.085 123.220 56.515 124.005 ;
        RECT 56.535 123.135 62.045 123.945 ;
        RECT 62.055 123.135 67.565 123.945 ;
        RECT 67.575 123.135 71.245 123.945 ;
        RECT 72.025 123.815 72.955 124.045 ;
        RECT 75.065 123.815 75.995 124.045 ;
        RECT 72.025 123.135 73.860 123.815 ;
        RECT 17.575 122.925 17.745 123.135 ;
        RECT 18.955 122.925 19.125 123.135 ;
        RECT 21.710 122.975 21.830 123.085 ;
        RECT 22.175 122.945 22.345 123.135 ;
        RECT 24.475 122.925 24.645 123.115 ;
        RECT 29.545 122.980 29.705 123.090 ;
        RECT 30.915 122.945 31.085 123.135 ;
        RECT 33.220 123.115 33.390 123.135 ;
        RECT 33.215 122.945 33.390 123.115 ;
        RECT 33.215 122.925 33.385 122.945 ;
        RECT 33.675 122.925 33.845 123.115 ;
        RECT 34.605 122.980 34.765 123.090 ;
        RECT 35.515 122.945 35.685 123.135 ;
        RECT 38.735 122.945 38.905 123.135 ;
        RECT 41.035 122.925 41.205 123.115 ;
        RECT 41.495 122.925 41.665 123.115 ;
        RECT 43.795 122.925 43.965 123.115 ;
        RECT 45.175 122.925 45.345 123.115 ;
        RECT 47.475 122.945 47.645 123.135 ;
        RECT 47.935 122.945 48.105 123.135 ;
        RECT 48.395 122.925 48.565 123.115 ;
        RECT 50.235 122.945 50.405 123.135 ;
        RECT 52.540 122.945 52.710 123.135 ;
        RECT 53.915 122.945 54.085 123.135 ;
        RECT 56.675 122.925 56.845 123.135 ;
        RECT 57.135 122.925 57.305 123.115 ;
        RECT 62.195 122.945 62.365 123.135 ;
        RECT 62.650 122.975 62.770 123.085 ;
        RECT 63.115 122.925 63.285 123.115 ;
        RECT 67.715 122.945 67.885 123.135 ;
        RECT 73.695 123.115 73.860 123.135 ;
        RECT 74.160 123.135 75.995 123.815 ;
        RECT 76.515 123.955 77.465 124.045 ;
        RECT 76.515 123.135 78.445 123.955 ;
        RECT 78.615 123.135 81.365 123.945 ;
        RECT 81.845 123.220 82.275 124.005 ;
        RECT 82.755 123.845 83.685 124.045 ;
        RECT 85.020 123.845 85.965 124.045 ;
        RECT 82.755 123.365 85.965 123.845 ;
        RECT 87.345 123.815 88.265 124.045 ;
        RECT 91.790 123.815 92.700 124.035 ;
        RECT 94.235 123.815 96.005 124.045 ;
        RECT 82.895 123.165 85.965 123.365 ;
        RECT 74.160 123.115 74.325 123.135 ;
        RECT 78.295 123.115 78.445 123.135 ;
        RECT 68.185 122.970 68.345 123.080 ;
        RECT 70.470 122.925 70.640 123.115 ;
        RECT 70.935 122.925 71.105 123.115 ;
        RECT 71.390 122.975 71.510 123.085 ;
        RECT 73.240 122.925 73.410 123.115 ;
        RECT 73.695 123.085 73.865 123.115 ;
        RECT 73.690 122.975 73.865 123.085 ;
        RECT 73.695 122.945 73.865 122.975 ;
        RECT 74.150 122.945 74.325 123.115 ;
        RECT 74.150 122.925 74.320 122.945 ;
        RECT 75.535 122.925 75.705 123.115 ;
        RECT 78.295 122.945 78.465 123.115 ;
        RECT 78.755 122.945 78.925 123.135 ;
        RECT 81.055 122.925 81.225 123.115 ;
        RECT 82.895 123.085 83.065 123.165 ;
        RECT 85.020 123.135 85.965 123.165 ;
        RECT 85.975 123.135 88.265 123.815 ;
        RECT 88.275 123.135 96.005 123.815 ;
        RECT 96.095 123.135 97.925 123.945 ;
        RECT 101.910 123.815 102.820 124.035 ;
        RECT 104.355 123.815 105.705 124.045 ;
        RECT 98.395 123.135 105.705 123.815 ;
        RECT 105.755 123.135 107.585 123.945 ;
        RECT 107.605 123.220 108.035 124.005 ;
        RECT 108.150 123.815 109.070 124.045 ;
        RECT 108.150 123.135 111.615 123.815 ;
        RECT 111.735 123.135 115.210 124.045 ;
        RECT 115.415 123.135 118.625 124.045 ;
        RECT 118.635 123.135 120.465 123.945 ;
        RECT 120.475 123.135 123.950 124.045 ;
        RECT 124.465 123.815 125.395 124.045 ;
        RECT 124.465 123.135 126.300 123.815 ;
        RECT 126.455 123.135 129.205 123.945 ;
        RECT 129.870 123.135 133.345 124.045 ;
        RECT 133.365 123.220 133.795 124.005 ;
        RECT 134.125 123.815 135.055 124.045 ;
        RECT 136.425 123.815 137.355 124.045 ;
        RECT 134.125 123.135 135.960 123.815 ;
        RECT 136.425 123.135 138.260 123.815 ;
        RECT 138.415 123.135 139.785 123.945 ;
        RECT 140.280 123.815 141.625 124.045 ;
        RECT 139.795 123.135 141.625 123.815 ;
        RECT 141.635 123.135 143.005 123.945 ;
        RECT 81.510 122.975 81.630 123.085 ;
        RECT 82.430 122.975 82.550 123.085 ;
        RECT 82.890 122.975 83.065 123.085 ;
        RECT 82.895 122.945 83.065 122.975 ;
        RECT 83.355 122.925 83.525 123.115 ;
        RECT 17.435 122.115 18.805 122.925 ;
        RECT 18.815 122.115 24.325 122.925 ;
        RECT 24.335 122.115 26.165 122.925 ;
        RECT 26.215 122.245 33.525 122.925 ;
        RECT 26.215 122.015 27.565 122.245 ;
        RECT 29.100 122.025 30.010 122.245 ;
        RECT 33.535 122.115 39.045 122.925 ;
        RECT 39.055 122.245 41.345 122.925 ;
        RECT 39.055 122.015 39.975 122.245 ;
        RECT 41.355 122.115 43.185 122.925 ;
        RECT 43.205 122.055 43.635 122.840 ;
        RECT 43.655 122.115 45.025 122.925 ;
        RECT 45.135 122.015 48.245 122.925 ;
        RECT 48.255 122.115 49.625 122.925 ;
        RECT 49.675 122.245 56.985 122.925 ;
        RECT 49.675 122.015 51.025 122.245 ;
        RECT 52.560 122.025 53.470 122.245 ;
        RECT 56.995 122.115 62.505 122.925 ;
        RECT 62.975 122.245 67.790 122.925 ;
        RECT 68.965 122.055 69.395 122.840 ;
        RECT 69.435 122.015 70.785 122.925 ;
        RECT 70.795 122.115 72.165 122.925 ;
        RECT 72.175 122.015 73.525 122.925 ;
        RECT 74.035 122.015 75.385 122.925 ;
        RECT 75.395 122.115 80.905 122.925 ;
        RECT 80.915 122.115 82.745 122.925 ;
        RECT 83.225 122.015 84.575 122.925 ;
        RECT 84.735 122.895 84.905 123.115 ;
        RECT 86.115 122.945 86.285 123.135 ;
        RECT 87.965 122.970 88.125 123.080 ;
        RECT 88.415 122.945 88.585 123.135 ;
        RECT 89.150 122.925 89.320 123.115 ;
        RECT 93.015 122.925 93.185 123.115 ;
        RECT 95.315 122.925 95.485 123.115 ;
        RECT 96.235 122.945 96.405 123.135 ;
        RECT 98.070 122.975 98.190 123.085 ;
        RECT 98.535 122.945 98.705 123.135 ;
        RECT 100.845 122.970 101.005 123.080 ;
        RECT 102.030 122.925 102.200 123.115 ;
        RECT 105.895 122.925 106.065 123.135 ;
        RECT 111.415 122.925 111.585 123.135 ;
        RECT 111.880 122.945 112.050 123.135 ;
        RECT 115.545 122.945 115.715 123.135 ;
        RECT 116.940 122.925 117.110 123.115 ;
        RECT 118.775 122.945 118.945 123.135 ;
        RECT 120.620 122.945 120.790 123.135 ;
        RECT 126.135 123.115 126.300 123.135 ;
        RECT 122.915 122.945 123.085 123.115 ;
        RECT 122.915 122.925 123.080 122.945 ;
        RECT 123.375 122.925 123.545 123.115 ;
        RECT 126.135 122.945 126.305 123.115 ;
        RECT 126.595 122.945 126.765 123.135 ;
        RECT 129.350 122.975 129.470 123.085 ;
        RECT 132.110 122.925 132.280 123.115 ;
        RECT 132.575 122.925 132.745 123.115 ;
        RECT 133.030 122.945 133.200 123.135 ;
        RECT 135.795 123.115 135.960 123.135 ;
        RECT 138.095 123.115 138.260 123.135 ;
        RECT 135.795 122.945 135.965 123.115 ;
        RECT 138.095 122.945 138.265 123.115 ;
        RECT 138.555 122.945 138.725 123.135 ;
        RECT 139.935 122.925 140.105 123.135 ;
        RECT 142.695 122.925 142.865 123.135 ;
        RECT 86.860 122.895 87.805 122.925 ;
        RECT 84.735 122.695 87.805 122.895 ;
        RECT 84.595 122.215 87.805 122.695 ;
        RECT 84.595 122.015 85.525 122.215 ;
        RECT 86.860 122.015 87.805 122.215 ;
        RECT 88.735 122.245 92.635 122.925 ;
        RECT 88.735 122.015 89.665 122.245 ;
        RECT 92.875 122.115 94.705 122.925 ;
        RECT 94.725 122.055 95.155 122.840 ;
        RECT 95.175 122.115 100.685 122.925 ;
        RECT 101.615 122.245 105.515 122.925 ;
        RECT 101.615 122.015 102.545 122.245 ;
        RECT 105.755 122.115 111.265 122.925 ;
        RECT 111.275 122.115 116.785 122.925 ;
        RECT 116.795 122.015 120.270 122.925 ;
        RECT 120.485 122.055 120.915 122.840 ;
        RECT 121.245 122.245 123.080 122.925 ;
        RECT 121.245 122.015 122.175 122.245 ;
        RECT 123.235 122.115 128.745 122.925 ;
        RECT 128.950 122.015 132.425 122.925 ;
        RECT 132.435 122.245 139.745 122.925 ;
        RECT 139.795 122.245 141.625 122.925 ;
        RECT 135.950 122.025 136.860 122.245 ;
        RECT 138.395 122.015 139.745 122.245 ;
        RECT 140.280 122.015 141.625 122.245 ;
        RECT 141.635 122.115 143.005 122.925 ;
      LAYER nwell ;
        RECT 17.240 118.895 143.200 121.725 ;
      LAYER pwell ;
        RECT 17.435 117.695 18.805 118.505 ;
        RECT 18.815 117.695 24.325 118.505 ;
        RECT 24.335 117.695 27.085 118.505 ;
        RECT 28.215 117.695 30.305 118.505 ;
        RECT 30.325 117.780 30.755 118.565 ;
        RECT 31.010 117.695 35.825 118.375 ;
        RECT 35.835 117.695 41.345 118.505 ;
        RECT 41.355 117.695 46.865 118.505 ;
        RECT 46.875 117.695 52.385 118.505 ;
        RECT 52.395 117.695 56.065 118.505 ;
        RECT 56.085 117.780 56.515 118.565 ;
        RECT 56.535 117.695 60.205 118.505 ;
        RECT 60.215 117.695 61.565 118.605 ;
        RECT 61.595 117.695 62.965 118.505 ;
        RECT 62.975 117.695 73.985 118.605 ;
        RECT 74.015 117.695 75.385 118.505 ;
        RECT 75.490 118.375 76.410 118.605 ;
        RECT 79.075 118.375 79.995 118.605 ;
        RECT 75.490 117.695 78.955 118.375 ;
        RECT 79.075 117.695 81.365 118.375 ;
        RECT 81.845 117.780 82.275 118.565 ;
        RECT 83.630 118.405 84.585 118.605 ;
        RECT 82.305 117.725 84.585 118.405 ;
        RECT 85.055 118.405 85.985 118.605 ;
        RECT 87.320 118.405 88.265 118.605 ;
        RECT 85.055 117.925 88.265 118.405 ;
        RECT 17.575 117.485 17.745 117.695 ;
        RECT 18.955 117.485 19.125 117.695 ;
        RECT 24.475 117.485 24.645 117.695 ;
        RECT 27.230 117.535 27.350 117.645 ;
        RECT 29.535 117.485 29.705 117.675 ;
        RECT 29.995 117.485 30.165 117.695 ;
        RECT 31.830 117.535 31.950 117.645 ;
        RECT 32.300 117.485 32.470 117.675 ;
        RECT 35.515 117.505 35.685 117.695 ;
        RECT 35.975 117.505 36.145 117.695 ;
        RECT 41.495 117.505 41.665 117.695 ;
        RECT 43.795 117.485 43.965 117.675 ;
        RECT 47.015 117.505 47.185 117.695 ;
        RECT 49.315 117.485 49.485 117.675 ;
        RECT 52.535 117.505 52.705 117.695 ;
        RECT 54.835 117.485 55.005 117.675 ;
        RECT 56.675 117.505 56.845 117.695 ;
        RECT 57.590 117.535 57.710 117.645 ;
        RECT 58.055 117.485 58.225 117.675 ;
        RECT 60.360 117.505 60.530 117.695 ;
        RECT 61.735 117.485 61.905 117.695 ;
        RECT 63.120 117.505 63.290 117.695 ;
        RECT 69.555 117.485 69.725 117.675 ;
        RECT 74.155 117.505 74.325 117.695 ;
        RECT 76.915 117.485 77.085 117.675 ;
        RECT 78.755 117.505 78.925 117.695 ;
        RECT 80.595 117.485 80.765 117.675 ;
        RECT 81.055 117.505 81.225 117.695 ;
        RECT 81.510 117.535 81.630 117.645 ;
        RECT 82.430 117.505 82.600 117.725 ;
        RECT 83.630 117.695 84.585 117.725 ;
        RECT 85.195 117.725 88.265 117.925 ;
        RECT 82.710 117.485 82.880 117.675 ;
        RECT 84.730 117.535 84.850 117.645 ;
        RECT 85.195 117.505 85.365 117.725 ;
        RECT 87.320 117.695 88.265 117.725 ;
        RECT 88.735 118.375 89.665 118.605 ;
        RECT 88.735 117.695 92.635 118.375 ;
        RECT 92.875 117.695 98.385 118.505 ;
        RECT 98.395 117.695 99.765 118.505 ;
        RECT 103.290 118.375 104.200 118.595 ;
        RECT 105.735 118.375 107.085 118.605 ;
        RECT 99.775 117.695 107.085 118.375 ;
        RECT 107.605 117.780 108.035 118.565 ;
        RECT 108.055 118.375 108.985 118.605 ;
        RECT 112.290 118.375 113.210 118.605 ;
        RECT 119.850 118.375 120.760 118.595 ;
        RECT 122.295 118.375 123.645 118.605 ;
        RECT 108.055 117.695 111.955 118.375 ;
        RECT 112.290 117.695 115.755 118.375 ;
        RECT 116.335 117.695 123.645 118.375 ;
        RECT 123.695 117.695 129.205 118.505 ;
        RECT 129.215 117.695 132.885 118.505 ;
        RECT 133.365 117.780 133.795 118.565 ;
        RECT 133.815 117.695 137.025 118.605 ;
        RECT 138.440 118.375 139.785 118.605 ;
        RECT 140.280 118.375 141.625 118.605 ;
        RECT 137.955 117.695 139.785 118.375 ;
        RECT 139.795 117.695 141.625 118.375 ;
        RECT 141.635 117.695 143.005 118.505 ;
        RECT 86.570 117.535 86.690 117.645 ;
        RECT 87.035 117.485 87.205 117.675 ;
        RECT 88.410 117.535 88.530 117.645 ;
        RECT 89.150 117.505 89.320 117.695 ;
        RECT 93.015 117.505 93.185 117.695 ;
        RECT 95.590 117.485 95.760 117.675 ;
        RECT 98.535 117.505 98.705 117.695 ;
        RECT 99.450 117.535 99.570 117.645 ;
        RECT 99.915 117.485 100.085 117.695 ;
        RECT 107.270 117.535 107.390 117.645 ;
        RECT 108.470 117.505 108.640 117.695 ;
        RECT 110.490 117.485 110.660 117.675 ;
        RECT 110.955 117.485 111.125 117.675 ;
        RECT 115.555 117.505 115.725 117.695 ;
        RECT 116.010 117.535 116.130 117.645 ;
        RECT 116.475 117.485 116.645 117.695 ;
        RECT 120.150 117.535 120.270 117.645 ;
        RECT 121.070 117.535 121.190 117.645 ;
        RECT 121.535 117.485 121.705 117.675 ;
        RECT 123.375 117.485 123.545 117.675 ;
        RECT 123.835 117.505 124.005 117.695 ;
        RECT 127.050 117.535 127.170 117.645 ;
        RECT 129.355 117.505 129.525 117.695 ;
        RECT 130.730 117.485 130.900 117.675 ;
        RECT 131.195 117.485 131.365 117.675 ;
        RECT 133.030 117.535 133.150 117.645 ;
        RECT 136.715 117.505 136.885 117.695 ;
        RECT 137.185 117.540 137.345 117.650 ;
        RECT 138.095 117.505 138.265 117.695 ;
        RECT 138.555 117.485 138.725 117.675 ;
        RECT 139.935 117.505 140.105 117.695 ;
        RECT 141.310 117.535 141.430 117.645 ;
        RECT 142.695 117.485 142.865 117.695 ;
        RECT 17.435 116.675 18.805 117.485 ;
        RECT 18.815 116.675 24.325 117.485 ;
        RECT 24.335 116.675 27.085 117.485 ;
        RECT 27.555 116.805 29.845 117.485 ;
        RECT 27.555 116.575 28.475 116.805 ;
        RECT 29.855 116.675 31.685 117.485 ;
        RECT 32.155 116.575 43.165 117.485 ;
        RECT 43.205 116.615 43.635 117.400 ;
        RECT 43.655 116.675 49.165 117.485 ;
        RECT 49.175 116.675 54.685 117.485 ;
        RECT 54.695 116.675 57.445 117.485 ;
        RECT 58.025 116.805 61.490 117.485 ;
        RECT 61.595 116.805 68.905 117.485 ;
        RECT 60.570 116.575 61.490 116.805 ;
        RECT 65.110 116.585 66.020 116.805 ;
        RECT 67.555 116.575 68.905 116.805 ;
        RECT 68.965 116.615 69.395 117.400 ;
        RECT 69.415 116.805 76.725 117.485 ;
        RECT 76.885 116.805 80.350 117.485 ;
        RECT 72.930 116.585 73.840 116.805 ;
        RECT 75.375 116.575 76.725 116.805 ;
        RECT 79.430 116.575 80.350 116.805 ;
        RECT 80.455 116.675 82.285 117.485 ;
        RECT 82.295 116.805 86.195 117.485 ;
        RECT 86.895 116.805 94.625 117.485 ;
        RECT 82.295 116.575 83.225 116.805 ;
        RECT 90.410 116.585 91.320 116.805 ;
        RECT 92.855 116.575 94.625 116.805 ;
        RECT 94.725 116.615 95.155 117.400 ;
        RECT 95.175 116.805 99.075 117.485 ;
        RECT 99.775 116.805 107.085 117.485 ;
        RECT 95.175 116.575 96.105 116.805 ;
        RECT 103.290 116.585 104.200 116.805 ;
        RECT 105.735 116.575 107.085 116.805 ;
        RECT 107.215 116.575 110.800 117.485 ;
        RECT 110.815 116.675 116.325 117.485 ;
        RECT 116.335 116.675 120.005 117.485 ;
        RECT 120.485 116.615 120.915 117.400 ;
        RECT 121.395 116.805 123.225 117.485 ;
        RECT 121.880 116.575 123.225 116.805 ;
        RECT 123.235 116.675 126.905 117.485 ;
        RECT 127.570 116.575 131.045 117.485 ;
        RECT 131.055 116.805 138.365 117.485 ;
        RECT 134.570 116.585 135.480 116.805 ;
        RECT 137.015 116.575 138.365 116.805 ;
        RECT 138.415 116.675 141.165 117.485 ;
        RECT 141.635 116.675 143.005 117.485 ;
      LAYER nwell ;
        RECT 17.240 113.455 143.200 116.285 ;
      LAYER pwell ;
        RECT 17.435 112.255 18.805 113.065 ;
        RECT 18.815 112.255 20.185 113.065 ;
        RECT 20.235 112.935 21.585 113.165 ;
        RECT 23.120 112.935 24.030 113.155 ;
        RECT 20.235 112.255 27.545 112.935 ;
        RECT 27.565 112.255 30.295 113.165 ;
        RECT 30.325 112.340 30.755 113.125 ;
        RECT 30.775 112.255 32.145 113.065 ;
        RECT 37.215 112.935 38.350 113.165 ;
        RECT 42.255 112.935 43.185 113.165 ;
        RECT 32.155 112.255 36.970 112.935 ;
        RECT 37.215 112.255 40.425 112.935 ;
        RECT 40.435 112.255 43.185 112.935 ;
        RECT 43.195 112.255 45.945 113.165 ;
        RECT 45.955 112.485 47.790 113.165 ;
        RECT 46.100 112.255 47.790 112.485 ;
        RECT 48.255 112.255 53.765 113.065 ;
        RECT 53.775 112.255 55.605 113.065 ;
        RECT 56.085 112.340 56.515 113.125 ;
        RECT 56.535 112.255 58.350 113.165 ;
        RECT 61.890 112.935 62.800 113.155 ;
        RECT 64.335 112.935 65.685 113.165 ;
        RECT 73.535 112.935 74.465 113.165 ;
        RECT 58.375 112.255 65.685 112.935 ;
        RECT 65.735 112.255 70.550 112.935 ;
        RECT 70.795 112.255 74.465 112.935 ;
        RECT 74.570 112.935 75.490 113.165 ;
        RECT 79.495 112.965 80.875 113.165 ;
        RECT 74.570 112.255 78.035 112.935 ;
        RECT 78.170 112.285 80.875 112.965 ;
        RECT 81.845 112.340 82.275 113.125 ;
        RECT 17.575 112.045 17.745 112.255 ;
        RECT 18.955 112.045 19.125 112.255 ;
        RECT 22.635 112.065 22.805 112.235 ;
        RECT 22.635 112.045 22.800 112.065 ;
        RECT 17.435 111.235 18.805 112.045 ;
        RECT 18.815 111.235 20.645 112.045 ;
        RECT 20.965 111.365 22.800 112.045 ;
        RECT 23.100 112.015 23.270 112.235 ;
        RECT 26.315 112.045 26.485 112.235 ;
        RECT 27.235 112.065 27.405 112.255 ;
        RECT 29.995 112.065 30.165 112.255 ;
        RECT 30.915 112.065 31.085 112.255 ;
        RECT 32.295 112.065 32.465 112.255 ;
        RECT 33.675 112.065 33.845 112.235 ;
        RECT 33.680 112.045 33.845 112.065 ;
        RECT 35.975 112.045 36.145 112.235 ;
        RECT 40.115 112.065 40.285 112.255 ;
        RECT 40.575 112.065 40.745 112.255 ;
        RECT 43.335 112.065 43.505 112.255 ;
        RECT 43.795 112.045 43.965 112.235 ;
        RECT 46.100 112.065 46.270 112.255 ;
        RECT 46.555 112.065 46.725 112.235 ;
        RECT 48.395 112.065 48.565 112.255 ;
        RECT 46.575 112.045 46.725 112.065 ;
        RECT 48.855 112.045 49.025 112.235 ;
        RECT 50.690 112.095 50.810 112.205 ;
        RECT 52.535 112.045 52.705 112.235 ;
        RECT 52.995 112.045 53.165 112.235 ;
        RECT 53.915 112.065 54.085 112.255 ;
        RECT 55.750 112.095 55.870 112.205 ;
        RECT 58.055 112.065 58.225 112.255 ;
        RECT 58.515 112.065 58.685 112.255 ;
        RECT 60.355 112.045 60.525 112.235 ;
        RECT 65.415 112.045 65.585 112.235 ;
        RECT 65.875 112.065 66.045 112.255 ;
        RECT 69.555 112.045 69.725 112.235 ;
        RECT 70.935 112.065 71.105 112.255 ;
        RECT 77.835 112.065 78.005 112.255 ;
        RECT 78.295 112.065 78.465 112.285 ;
        RECT 79.495 112.255 80.875 112.285 ;
        RECT 82.295 112.255 83.645 113.165 ;
        RECT 83.675 112.255 87.345 113.065 ;
        RECT 91.330 112.935 92.240 113.155 ;
        RECT 93.775 112.935 95.545 113.165 ;
        RECT 87.815 112.255 95.545 112.935 ;
        RECT 95.635 112.255 101.145 113.065 ;
        RECT 101.155 112.255 104.825 113.065 ;
        RECT 105.765 112.255 107.115 113.165 ;
        RECT 107.605 112.340 108.035 113.125 ;
        RECT 109.395 112.965 110.805 113.165 ;
        RECT 108.070 112.285 110.805 112.965 ;
        RECT 78.755 112.065 78.925 112.235 ;
        RECT 78.755 112.045 78.920 112.065 ;
        RECT 79.220 112.045 79.390 112.235 ;
        RECT 81.055 112.045 81.225 112.235 ;
        RECT 83.360 112.065 83.530 112.255 ;
        RECT 83.815 112.065 83.985 112.255 ;
        RECT 87.490 112.095 87.610 112.205 ;
        RECT 87.955 112.065 88.125 112.255 ;
        RECT 88.875 112.045 89.045 112.235 ;
        RECT 91.635 112.045 91.805 112.235 ;
        RECT 94.390 112.095 94.510 112.205 ;
        RECT 95.315 112.045 95.485 112.235 ;
        RECT 95.775 112.065 95.945 112.255 ;
        RECT 100.375 112.045 100.545 112.235 ;
        RECT 101.295 112.065 101.465 112.255 ;
        RECT 101.755 112.045 101.925 112.235 ;
        RECT 104.985 112.100 105.145 112.210 ;
        RECT 25.230 112.015 26.165 112.045 ;
        RECT 23.100 111.815 26.165 112.015 ;
        RECT 20.965 111.135 21.895 111.365 ;
        RECT 22.955 111.335 26.165 111.815 ;
        RECT 26.175 111.365 33.485 112.045 ;
        RECT 33.680 111.365 35.515 112.045 ;
        RECT 35.835 111.365 43.145 112.045 ;
        RECT 22.955 111.135 23.885 111.335 ;
        RECT 25.215 111.135 26.165 111.335 ;
        RECT 29.690 111.145 30.600 111.365 ;
        RECT 32.135 111.135 33.485 111.365 ;
        RECT 34.585 111.135 35.515 111.365 ;
        RECT 39.350 111.145 40.260 111.365 ;
        RECT 41.795 111.135 43.145 111.365 ;
        RECT 43.205 111.175 43.635 111.960 ;
        RECT 43.655 111.135 46.405 112.045 ;
        RECT 46.575 111.225 48.505 112.045 ;
        RECT 48.715 111.235 50.545 112.045 ;
        RECT 47.555 111.135 48.505 111.225 ;
        RECT 51.015 111.135 52.830 112.045 ;
        RECT 52.855 111.365 60.165 112.045 ;
        RECT 60.215 111.365 65.030 112.045 ;
        RECT 65.385 111.365 68.850 112.045 ;
        RECT 56.370 111.145 57.280 111.365 ;
        RECT 58.815 111.135 60.165 111.365 ;
        RECT 67.930 111.135 68.850 111.365 ;
        RECT 68.965 111.175 69.395 111.960 ;
        RECT 69.415 111.365 76.725 112.045 ;
        RECT 72.930 111.145 73.840 111.365 ;
        RECT 75.375 111.135 76.725 111.365 ;
        RECT 77.085 111.365 78.920 112.045 ;
        RECT 77.085 111.135 78.015 111.365 ;
        RECT 79.075 111.135 80.905 112.045 ;
        RECT 80.915 111.365 88.645 112.045 ;
        RECT 84.430 111.145 85.340 111.365 ;
        RECT 86.875 111.135 88.645 111.365 ;
        RECT 88.735 111.235 91.485 112.045 ;
        RECT 91.495 111.365 94.235 112.045 ;
        RECT 94.725 111.175 95.155 111.960 ;
        RECT 95.175 111.365 99.990 112.045 ;
        RECT 100.245 111.135 101.595 112.045 ;
        RECT 101.615 111.235 102.985 112.045 ;
        RECT 102.995 112.015 104.390 112.045 ;
        RECT 105.435 112.015 105.605 112.235 ;
        RECT 106.815 112.065 106.985 112.255 ;
        RECT 107.270 112.095 107.390 112.205 ;
        RECT 108.195 112.065 108.365 112.285 ;
        RECT 109.410 112.255 110.805 112.285 ;
        RECT 110.815 112.255 113.565 113.065 ;
        RECT 113.575 112.255 117.050 113.165 ;
        RECT 120.770 112.935 121.680 113.155 ;
        RECT 123.215 112.935 124.565 113.165 ;
        RECT 117.255 112.255 124.565 112.935 ;
        RECT 124.925 112.935 125.855 113.165 ;
        RECT 124.925 112.255 126.760 112.935 ;
        RECT 126.915 112.255 132.425 113.065 ;
        RECT 133.365 112.340 133.795 113.125 ;
        RECT 134.865 112.935 135.795 113.165 ;
        RECT 133.960 112.255 135.795 112.935 ;
        RECT 136.425 112.935 137.355 113.165 ;
        RECT 136.425 112.255 138.260 112.935 ;
        RECT 138.415 112.255 139.785 113.065 ;
        RECT 140.280 112.935 141.625 113.165 ;
        RECT 139.795 112.255 141.625 112.935 ;
        RECT 141.635 112.255 143.005 113.065 ;
        RECT 110.955 112.065 111.125 112.255 ;
        RECT 113.720 112.235 113.890 112.255 ;
        RECT 111.410 112.045 111.580 112.235 ;
        RECT 111.875 112.045 112.045 112.235 ;
        RECT 113.715 112.065 113.890 112.235 ;
        RECT 117.395 112.065 117.565 112.255 ;
        RECT 126.595 112.235 126.760 112.255 ;
        RECT 113.715 112.045 113.885 112.065 ;
        RECT 120.150 112.045 120.320 112.235 ;
        RECT 123.835 112.045 124.005 112.235 ;
        RECT 124.295 112.045 124.465 112.235 ;
        RECT 126.595 112.065 126.765 112.235 ;
        RECT 127.055 112.205 127.225 112.255 ;
        RECT 133.960 112.235 134.125 112.255 ;
        RECT 127.050 112.095 127.225 112.205 ;
        RECT 127.055 112.065 127.225 112.095 ;
        RECT 130.730 112.045 130.900 112.235 ;
        RECT 131.195 112.045 131.365 112.235 ;
        RECT 132.585 112.100 132.745 112.210 ;
        RECT 133.955 112.065 134.125 112.235 ;
        RECT 138.095 112.235 138.260 112.255 ;
        RECT 138.095 112.065 138.265 112.235 ;
        RECT 138.555 112.065 138.725 112.255 ;
        RECT 139.935 112.065 140.105 112.255 ;
        RECT 140.865 112.090 141.025 112.200 ;
        RECT 138.560 112.045 138.725 112.065 ;
        RECT 142.695 112.045 142.865 112.255 ;
        RECT 102.995 111.335 105.730 112.015 ;
        RECT 102.995 111.135 104.405 111.335 ;
        RECT 106.155 111.135 111.725 112.045 ;
        RECT 111.735 111.365 113.565 112.045 ;
        RECT 113.575 111.235 117.245 112.045 ;
        RECT 118.275 111.135 120.465 112.045 ;
        RECT 120.485 111.175 120.915 111.960 ;
        RECT 120.935 111.135 124.145 112.045 ;
        RECT 124.155 111.365 126.895 112.045 ;
        RECT 127.570 111.135 131.045 112.045 ;
        RECT 131.055 111.365 138.365 112.045 ;
        RECT 138.560 111.365 140.395 112.045 ;
        RECT 134.570 111.145 135.480 111.365 ;
        RECT 137.015 111.135 138.365 111.365 ;
        RECT 139.465 111.135 140.395 111.365 ;
        RECT 141.635 111.235 143.005 112.045 ;
      LAYER nwell ;
        RECT 17.240 108.015 143.200 110.845 ;
      LAYER pwell ;
        RECT 17.435 106.815 18.805 107.625 ;
        RECT 18.815 106.815 22.485 107.625 ;
        RECT 22.955 107.525 23.905 107.725 ;
        RECT 25.235 107.525 26.165 107.725 ;
        RECT 22.955 107.045 26.165 107.525 ;
        RECT 22.955 106.845 26.020 107.045 ;
        RECT 22.955 106.815 23.890 106.845 ;
        RECT 17.575 106.605 17.745 106.815 ;
        RECT 18.955 106.605 19.125 106.815 ;
        RECT 21.710 106.655 21.830 106.765 ;
        RECT 22.175 106.605 22.345 106.795 ;
        RECT 22.630 106.655 22.750 106.765 ;
        RECT 25.850 106.625 26.020 106.845 ;
        RECT 26.195 106.815 27.545 107.725 ;
        RECT 27.565 106.815 30.295 107.725 ;
        RECT 30.325 106.900 30.755 107.685 ;
        RECT 30.905 106.815 33.905 107.725 ;
        RECT 33.995 106.815 35.825 107.625 ;
        RECT 35.985 106.815 39.640 107.725 ;
        RECT 39.975 107.525 40.925 107.725 ;
        RECT 42.255 107.525 43.185 107.725 ;
        RECT 39.975 107.045 43.185 107.525 ;
        RECT 39.975 106.845 43.040 107.045 ;
        RECT 39.975 106.815 40.910 106.845 ;
        RECT 26.310 106.625 26.480 106.815 ;
        RECT 27.695 106.625 27.865 106.815 ;
        RECT 29.535 106.605 29.705 106.795 ;
        RECT 33.215 106.605 33.385 106.795 ;
        RECT 33.675 106.625 33.845 106.815 ;
        RECT 34.135 106.625 34.305 106.815 ;
        RECT 35.985 106.795 36.145 106.815 ;
        RECT 35.515 106.625 35.685 106.795 ;
        RECT 35.515 106.605 35.665 106.625 ;
        RECT 35.975 106.605 36.145 106.795 ;
        RECT 41.495 106.605 41.665 106.795 ;
        RECT 42.870 106.625 43.040 106.845 ;
        RECT 43.195 106.815 44.565 107.625 ;
        RECT 44.575 106.815 48.230 107.725 ;
        RECT 49.175 107.525 50.125 107.725 ;
        RECT 51.455 107.525 52.385 107.725 ;
        RECT 49.175 107.045 52.385 107.525 ;
        RECT 55.050 107.495 55.970 107.725 ;
        RECT 49.175 106.845 52.240 107.045 ;
        RECT 49.175 106.815 50.110 106.845 ;
        RECT 43.335 106.625 43.505 106.815 ;
        RECT 43.795 106.605 43.965 106.795 ;
        RECT 44.720 106.625 44.890 106.815 ;
        RECT 45.630 106.655 45.750 106.765 ;
        RECT 48.405 106.660 48.565 106.770 ;
        RECT 48.850 106.605 49.020 106.795 ;
        RECT 49.315 106.605 49.485 106.795 ;
        RECT 52.070 106.625 52.240 106.845 ;
        RECT 52.505 106.815 55.970 107.495 ;
        RECT 56.085 106.900 56.515 107.685 ;
        RECT 56.575 107.495 57.925 107.725 ;
        RECT 59.460 107.495 60.370 107.715 ;
        RECT 56.575 106.815 63.885 107.495 ;
        RECT 63.895 106.815 65.265 107.625 ;
        RECT 65.275 106.815 68.025 107.725 ;
        RECT 68.035 106.815 69.405 107.625 ;
        RECT 69.415 107.525 70.370 107.725 ;
        RECT 69.415 106.845 71.695 107.525 ;
        RECT 71.715 107.495 72.635 107.725 ;
        RECT 74.110 107.495 75.030 107.725 ;
        RECT 80.895 107.495 81.825 107.725 ;
        RECT 69.415 106.815 70.370 106.845 ;
        RECT 52.535 106.625 52.705 106.815 ;
        RECT 17.435 105.795 18.805 106.605 ;
        RECT 18.815 105.795 21.565 106.605 ;
        RECT 22.035 105.925 29.345 106.605 ;
        RECT 25.550 105.705 26.460 105.925 ;
        RECT 27.995 105.695 29.345 105.925 ;
        RECT 29.395 105.795 31.225 106.605 ;
        RECT 31.235 105.925 33.525 106.605 ;
        RECT 31.235 105.695 32.155 105.925 ;
        RECT 33.735 105.785 35.665 106.605 ;
        RECT 35.835 105.795 41.345 106.605 ;
        RECT 41.355 105.795 43.185 106.605 ;
        RECT 33.735 105.695 34.685 105.785 ;
        RECT 43.205 105.735 43.635 106.520 ;
        RECT 43.655 105.795 45.485 106.605 ;
        RECT 46.100 105.695 49.165 106.605 ;
        RECT 49.185 105.695 51.915 106.605 ;
        RECT 51.935 106.575 52.885 106.605 ;
        RECT 55.290 106.575 55.460 106.795 ;
        RECT 55.755 106.625 55.925 106.795 ;
        RECT 55.760 106.605 55.925 106.625 ;
        RECT 58.055 106.605 58.225 106.795 ;
        RECT 63.575 106.765 63.745 106.815 ;
        RECT 63.570 106.655 63.745 106.765 ;
        RECT 63.575 106.625 63.745 106.655 ;
        RECT 64.035 106.795 64.205 106.815 ;
        RECT 64.035 106.625 64.210 106.795 ;
        RECT 65.415 106.625 65.585 106.815 ;
        RECT 64.040 106.605 64.210 106.625 ;
        RECT 65.875 106.605 66.045 106.795 ;
        RECT 68.175 106.625 68.345 106.815 ;
        RECT 70.480 106.605 70.650 106.795 ;
        RECT 71.400 106.625 71.570 106.845 ;
        RECT 71.715 106.815 74.005 107.495 ;
        RECT 74.110 106.815 77.575 107.495 ;
        RECT 77.925 106.815 81.825 107.495 ;
        RECT 81.845 106.900 82.275 107.685 ;
        RECT 85.810 107.495 86.720 107.715 ;
        RECT 88.255 107.495 90.025 107.725 ;
        RECT 82.295 106.815 90.025 107.495 ;
        RECT 90.585 106.815 93.325 107.495 ;
        RECT 93.335 106.815 97.005 107.625 ;
        RECT 97.015 106.815 98.385 107.625 ;
        RECT 98.410 107.495 99.780 107.725 ;
        RECT 98.410 106.815 100.685 107.495 ;
        RECT 100.695 106.815 102.905 107.725 ;
        RECT 103.005 106.815 104.355 107.725 ;
        RECT 106.435 107.635 107.385 107.725 ;
        RECT 105.455 106.815 107.385 107.635 ;
        RECT 107.605 106.900 108.035 107.685 ;
        RECT 108.055 106.815 110.245 107.725 ;
        RECT 110.355 106.815 114.025 107.625 ;
        RECT 114.035 106.815 115.405 107.625 ;
        RECT 118.930 107.495 119.840 107.715 ;
        RECT 121.375 107.495 122.725 107.725 ;
        RECT 115.415 106.815 122.725 107.495 ;
        RECT 122.775 106.815 127.590 107.495 ;
        RECT 128.030 106.815 131.505 107.725 ;
        RECT 131.515 106.815 133.345 107.625 ;
        RECT 133.365 106.900 133.795 107.685 ;
        RECT 137.330 107.495 138.240 107.715 ;
        RECT 139.775 107.495 141.125 107.725 ;
        RECT 133.815 106.815 141.125 107.495 ;
        RECT 141.635 106.815 143.005 107.625 ;
        RECT 73.695 106.605 73.865 106.815 ;
        RECT 75.530 106.605 75.700 106.795 ;
        RECT 75.995 106.605 76.165 106.795 ;
        RECT 77.375 106.625 77.545 106.815 ;
        RECT 81.240 106.625 81.410 106.815 ;
        RECT 81.515 106.605 81.685 106.795 ;
        RECT 82.435 106.625 82.605 106.815 ;
        RECT 87.030 106.655 87.150 106.765 ;
        RECT 87.495 106.605 87.665 106.795 ;
        RECT 90.250 106.655 90.370 106.765 ;
        RECT 93.015 106.625 93.185 106.815 ;
        RECT 93.475 106.625 93.645 106.815 ;
        RECT 95.305 106.605 95.475 106.795 ;
        RECT 97.155 106.625 97.325 106.815 ;
        RECT 98.535 106.605 98.705 106.795 ;
        RECT 100.370 106.625 100.540 106.815 ;
        RECT 100.840 106.625 101.010 106.815 ;
        RECT 103.135 106.625 103.305 106.815 ;
        RECT 105.455 106.795 105.605 106.815 ;
        RECT 104.055 106.605 104.225 106.795 ;
        RECT 104.525 106.660 104.685 106.770 ;
        RECT 105.435 106.625 105.605 106.795 ;
        RECT 105.890 106.655 106.010 106.765 ;
        RECT 106.360 106.605 106.530 106.795 ;
        RECT 108.200 106.625 108.370 106.815 ;
        RECT 110.495 106.625 110.665 106.815 ;
        RECT 111.875 106.625 112.045 106.795 ;
        RECT 111.875 106.605 112.040 106.625 ;
        RECT 112.335 106.605 112.505 106.795 ;
        RECT 113.715 106.625 113.885 106.795 ;
        RECT 114.175 106.625 114.345 106.815 ;
        RECT 115.555 106.625 115.725 106.815 ;
        RECT 113.720 106.605 113.885 106.625 ;
        RECT 116.020 106.605 116.190 106.795 ;
        RECT 119.705 106.650 119.865 106.760 ;
        RECT 121.075 106.605 121.245 106.795 ;
        RECT 122.915 106.625 123.085 106.815 ;
        RECT 126.135 106.605 126.305 106.795 ;
        RECT 131.190 106.605 131.360 106.815 ;
        RECT 131.655 106.605 131.825 106.815 ;
        RECT 133.955 106.625 134.125 106.815 ;
        RECT 139.025 106.650 139.185 106.760 ;
        RECT 139.935 106.605 140.105 106.795 ;
        RECT 141.310 106.655 141.430 106.765 ;
        RECT 142.695 106.605 142.865 106.815 ;
        RECT 51.935 105.895 55.605 106.575 ;
        RECT 55.760 105.925 57.595 106.605 ;
        RECT 51.935 105.695 52.885 105.895 ;
        RECT 56.665 105.695 57.595 105.925 ;
        RECT 57.915 105.795 63.425 106.605 ;
        RECT 63.895 105.695 65.725 106.605 ;
        RECT 65.835 105.695 68.945 106.605 ;
        RECT 68.965 105.735 69.395 106.520 ;
        RECT 69.415 105.695 70.765 106.605 ;
        RECT 72.165 106.575 74.005 106.605 ;
        RECT 70.840 105.925 74.005 106.575 ;
        RECT 70.840 105.895 73.520 105.925 ;
        RECT 72.165 105.695 73.520 105.895 ;
        RECT 74.015 105.695 75.845 106.605 ;
        RECT 75.855 105.795 81.365 106.605 ;
        RECT 81.375 105.795 86.885 106.605 ;
        RECT 87.355 105.925 94.665 106.605 ;
        RECT 90.870 105.705 91.780 105.925 ;
        RECT 93.315 105.695 94.665 105.925 ;
        RECT 94.725 105.735 95.155 106.520 ;
        RECT 95.175 105.695 98.385 106.605 ;
        RECT 98.395 105.795 103.905 106.605 ;
        RECT 103.915 105.795 105.745 106.605 ;
        RECT 106.215 105.695 109.690 106.605 ;
        RECT 110.205 105.925 112.040 106.605 ;
        RECT 110.205 105.695 111.135 105.925 ;
        RECT 112.195 105.795 113.565 106.605 ;
        RECT 113.720 105.925 115.555 106.605 ;
        RECT 114.625 105.695 115.555 105.925 ;
        RECT 115.875 105.695 119.350 106.605 ;
        RECT 120.485 105.735 120.915 106.520 ;
        RECT 120.935 105.925 125.750 106.605 ;
        RECT 125.995 105.795 127.825 106.605 ;
        RECT 128.030 105.695 131.505 106.605 ;
        RECT 131.515 105.925 138.825 106.605 ;
        RECT 139.795 105.925 141.625 106.605 ;
        RECT 135.030 105.705 135.940 105.925 ;
        RECT 137.475 105.695 138.825 105.925 ;
        RECT 140.280 105.695 141.625 105.925 ;
        RECT 141.635 105.795 143.005 106.605 ;
      LAYER nwell ;
        RECT 17.240 102.575 143.200 105.405 ;
      LAYER pwell ;
        RECT 17.435 101.375 18.805 102.185 ;
        RECT 18.815 101.375 21.565 102.185 ;
        RECT 25.090 102.055 26.000 102.275 ;
        RECT 27.535 102.055 28.885 102.285 ;
        RECT 21.575 101.375 28.885 102.055 ;
        RECT 28.935 101.375 30.305 102.185 ;
        RECT 30.325 101.460 30.755 102.245 ;
        RECT 32.850 102.055 33.985 102.285 ;
        RECT 30.775 101.375 33.985 102.055 ;
        RECT 33.995 101.375 39.505 102.185 ;
        RECT 39.515 101.375 45.025 102.185 ;
        RECT 45.035 101.375 46.865 102.185 ;
        RECT 48.755 102.055 50.105 102.285 ;
        RECT 51.640 102.055 52.550 102.275 ;
        RECT 46.875 101.375 48.705 102.055 ;
        RECT 48.755 101.375 56.065 102.055 ;
        RECT 56.085 101.460 56.515 102.245 ;
        RECT 59.190 102.055 60.110 102.285 ;
        RECT 56.645 101.375 60.110 102.055 ;
        RECT 60.225 101.375 61.575 102.285 ;
        RECT 61.595 101.375 65.265 102.185 ;
        RECT 65.275 101.375 67.105 102.285 ;
        RECT 70.630 102.055 71.540 102.275 ;
        RECT 73.075 102.055 74.425 102.285 ;
        RECT 67.115 101.375 74.425 102.055 ;
        RECT 74.475 101.375 79.985 102.185 ;
        RECT 79.995 101.375 81.825 102.185 ;
        RECT 81.845 101.460 82.275 102.245 ;
        RECT 83.345 102.055 84.275 102.285 ;
        RECT 82.440 101.375 84.275 102.055 ;
        RECT 84.595 101.375 86.425 102.185 ;
        RECT 86.435 101.375 89.645 102.285 ;
        RECT 95.945 102.055 96.875 102.285 ;
        RECT 90.810 101.375 95.625 102.055 ;
        RECT 95.945 101.375 97.780 102.055 ;
        RECT 97.935 101.375 101.605 102.185 ;
        RECT 101.925 102.055 102.855 102.285 ;
        RECT 101.925 101.375 103.760 102.055 ;
        RECT 104.110 101.375 107.585 102.285 ;
        RECT 107.605 101.460 108.035 102.245 ;
        RECT 111.570 102.055 112.480 102.275 ;
        RECT 114.015 102.055 115.365 102.285 ;
        RECT 108.055 101.375 115.365 102.055 ;
        RECT 115.610 101.375 119.085 102.285 ;
        RECT 123.915 102.195 124.865 102.285 ;
        RECT 119.095 101.375 122.765 102.185 ;
        RECT 122.935 101.375 124.865 102.195 ;
        RECT 125.385 102.055 126.315 102.285 ;
        RECT 125.385 101.375 127.220 102.055 ;
        RECT 127.375 101.375 129.205 102.185 ;
        RECT 129.525 102.055 130.455 102.285 ;
        RECT 129.525 101.375 131.360 102.055 ;
        RECT 131.515 101.375 133.345 102.185 ;
        RECT 133.365 101.460 133.795 102.245 ;
        RECT 133.815 101.375 137.025 102.285 ;
        RECT 138.440 102.055 139.785 102.285 ;
        RECT 140.280 102.055 141.625 102.285 ;
        RECT 137.955 101.375 139.785 102.055 ;
        RECT 139.795 101.375 141.625 102.055 ;
        RECT 141.635 101.375 143.005 102.185 ;
        RECT 17.575 101.165 17.745 101.375 ;
        RECT 18.955 101.165 19.125 101.375 ;
        RECT 21.715 101.355 21.885 101.375 ;
        RECT 21.715 101.185 21.890 101.355 ;
        RECT 21.720 101.165 21.890 101.185 ;
        RECT 25.395 101.165 25.565 101.355 ;
        RECT 25.860 101.165 26.030 101.355 ;
        RECT 29.075 101.185 29.245 101.375 ;
        RECT 30.915 101.185 31.085 101.375 ;
        RECT 31.375 101.165 31.545 101.355 ;
        RECT 31.835 101.165 32.005 101.355 ;
        RECT 34.135 101.185 34.305 101.375 ;
        RECT 37.350 101.215 37.470 101.325 ;
        RECT 37.815 101.165 37.985 101.355 ;
        RECT 39.655 101.185 39.825 101.375 ;
        RECT 40.115 101.165 40.285 101.355 ;
        RECT 42.870 101.215 42.990 101.325 ;
        RECT 44.720 101.165 44.890 101.355 ;
        RECT 45.175 101.165 45.345 101.375 ;
        RECT 47.015 101.185 47.185 101.375 ;
        RECT 47.930 101.215 48.050 101.325 ;
        RECT 48.395 101.185 48.565 101.355 ;
        RECT 50.695 101.185 50.865 101.355 ;
        RECT 48.415 101.165 48.565 101.185 ;
        RECT 50.845 101.165 50.865 101.185 ;
        RECT 53.455 101.165 53.625 101.355 ;
        RECT 55.755 101.185 55.925 101.375 ;
        RECT 56.675 101.185 56.845 101.375 ;
        RECT 57.135 101.185 57.305 101.355 ;
        RECT 60.355 101.185 60.525 101.375 ;
        RECT 57.140 101.165 57.305 101.185 ;
        RECT 61.275 101.165 61.445 101.355 ;
        RECT 61.735 101.165 61.905 101.375 ;
        RECT 65.420 101.165 65.590 101.375 ;
        RECT 67.255 101.185 67.425 101.375 ;
        RECT 69.555 101.165 69.725 101.355 ;
        RECT 74.155 101.165 74.325 101.355 ;
        RECT 74.615 101.165 74.785 101.375 ;
        RECT 78.295 101.165 78.465 101.355 ;
        RECT 80.135 101.185 80.305 101.375 ;
        RECT 82.440 101.355 82.605 101.375 ;
        RECT 82.435 101.185 82.605 101.355 ;
        RECT 84.735 101.185 84.905 101.375 ;
        RECT 85.655 101.165 85.825 101.355 ;
        RECT 86.565 101.185 86.735 101.375 ;
        RECT 89.330 101.215 89.450 101.325 ;
        RECT 89.800 101.165 89.970 101.355 ;
        RECT 93.475 101.165 93.645 101.355 ;
        RECT 95.315 101.185 95.485 101.375 ;
        RECT 97.615 101.355 97.780 101.375 ;
        RECT 97.615 101.185 97.785 101.355 ;
        RECT 98.075 101.165 98.245 101.375 ;
        RECT 103.595 101.355 103.760 101.375 ;
        RECT 107.270 101.355 107.440 101.375 ;
        RECT 98.535 101.165 98.705 101.355 ;
        RECT 103.595 101.185 103.765 101.355 ;
        RECT 104.055 101.165 104.225 101.355 ;
        RECT 106.810 101.215 106.930 101.325 ;
        RECT 107.270 101.185 107.445 101.355 ;
        RECT 108.195 101.185 108.365 101.375 ;
        RECT 107.275 101.165 107.445 101.185 ;
        RECT 114.635 101.165 114.805 101.355 ;
        RECT 117.390 101.215 117.510 101.325 ;
        RECT 117.855 101.185 118.025 101.355 ;
        RECT 118.770 101.185 118.940 101.375 ;
        RECT 119.235 101.185 119.405 101.375 ;
        RECT 122.935 101.355 123.085 101.375 ;
        RECT 120.150 101.215 120.270 101.325 ;
        RECT 117.875 101.165 118.025 101.185 ;
        RECT 121.075 101.165 121.245 101.355 ;
        RECT 122.915 101.185 123.085 101.355 ;
        RECT 127.055 101.355 127.220 101.375 ;
        RECT 127.055 101.185 127.225 101.355 ;
        RECT 127.515 101.185 127.685 101.375 ;
        RECT 131.195 101.355 131.360 101.375 ;
        RECT 129.810 101.165 129.980 101.355 ;
        RECT 130.275 101.165 130.445 101.355 ;
        RECT 131.195 101.185 131.365 101.355 ;
        RECT 131.655 101.185 131.825 101.375 ;
        RECT 136.715 101.185 136.885 101.375 ;
        RECT 137.185 101.220 137.345 101.330 ;
        RECT 138.095 101.185 138.265 101.375 ;
        RECT 139.935 101.185 140.105 101.375 ;
        RECT 140.395 101.165 140.565 101.355 ;
        RECT 140.865 101.210 141.025 101.320 ;
        RECT 142.695 101.165 142.865 101.375 ;
        RECT 17.435 100.355 18.805 101.165 ;
        RECT 18.815 100.355 21.565 101.165 ;
        RECT 21.575 100.255 23.405 101.165 ;
        RECT 23.415 100.485 25.705 101.165 ;
        RECT 23.415 100.255 24.335 100.485 ;
        RECT 25.715 100.255 28.635 101.165 ;
        RECT 28.945 100.255 31.675 101.165 ;
        RECT 31.695 100.355 37.205 101.165 ;
        RECT 37.675 100.485 39.965 101.165 ;
        RECT 39.045 100.255 39.965 100.485 ;
        RECT 39.985 100.255 42.715 101.165 ;
        RECT 43.205 100.295 43.635 101.080 ;
        RECT 43.655 100.255 45.005 101.165 ;
        RECT 45.035 100.355 47.785 101.165 ;
        RECT 48.415 100.345 50.345 101.165 ;
        RECT 50.845 100.485 53.295 101.165 ;
        RECT 53.425 100.485 56.890 101.165 ;
        RECT 57.140 100.485 58.975 101.165 ;
        RECT 49.395 100.255 50.345 100.345 ;
        RECT 51.335 100.255 53.295 100.485 ;
        RECT 55.970 100.255 56.890 100.485 ;
        RECT 58.045 100.255 58.975 100.485 ;
        RECT 59.295 100.485 61.585 101.165 ;
        RECT 59.295 100.255 60.215 100.485 ;
        RECT 61.595 100.355 65.265 101.165 ;
        RECT 65.275 100.255 68.945 101.165 ;
        RECT 68.965 100.295 69.395 101.080 ;
        RECT 69.415 100.355 70.785 101.165 ;
        RECT 70.890 100.485 74.355 101.165 ;
        RECT 70.890 100.255 71.810 100.485 ;
        RECT 74.475 100.355 78.145 101.165 ;
        RECT 78.155 100.485 85.465 101.165 ;
        RECT 81.670 100.265 82.580 100.485 ;
        RECT 84.115 100.255 85.465 100.485 ;
        RECT 85.515 100.355 89.185 101.165 ;
        RECT 89.655 100.255 93.130 101.165 ;
        RECT 93.335 100.355 94.705 101.165 ;
        RECT 94.725 100.295 95.155 101.080 ;
        RECT 95.175 100.255 98.385 101.165 ;
        RECT 98.395 100.355 103.905 101.165 ;
        RECT 103.915 100.355 106.665 101.165 ;
        RECT 107.135 100.485 114.445 101.165 ;
        RECT 110.650 100.265 111.560 100.485 ;
        RECT 113.095 100.255 114.445 100.485 ;
        RECT 114.495 100.355 117.245 101.165 ;
        RECT 117.875 100.345 119.805 101.165 ;
        RECT 118.855 100.255 119.805 100.345 ;
        RECT 120.485 100.295 120.915 101.080 ;
        RECT 120.935 100.355 126.445 101.165 ;
        RECT 126.650 100.255 130.125 101.165 ;
        RECT 130.135 100.485 137.445 101.165 ;
        RECT 133.650 100.265 134.560 100.485 ;
        RECT 136.095 100.255 137.445 100.485 ;
        RECT 137.495 100.255 140.705 101.165 ;
        RECT 141.635 100.355 143.005 101.165 ;
      LAYER nwell ;
        RECT 17.240 97.135 143.200 99.965 ;
      LAYER pwell ;
        RECT 17.435 95.935 18.805 96.745 ;
        RECT 18.815 95.935 24.325 96.745 ;
        RECT 24.335 95.935 26.165 96.745 ;
        RECT 27.225 96.615 28.155 96.845 ;
        RECT 26.320 95.935 28.155 96.615 ;
        RECT 28.475 95.935 30.305 96.745 ;
        RECT 30.325 96.020 30.755 96.805 ;
        RECT 30.775 95.935 34.445 96.745 ;
        RECT 34.455 95.935 35.825 96.745 ;
        RECT 36.145 96.615 37.075 96.845 ;
        RECT 41.650 96.615 42.560 96.835 ;
        RECT 44.095 96.615 45.445 96.845 ;
        RECT 36.145 95.935 37.980 96.615 ;
        RECT 38.135 95.935 45.445 96.615 ;
        RECT 45.535 96.615 46.885 96.845 ;
        RECT 48.420 96.615 49.330 96.835 ;
        RECT 52.855 96.645 53.785 96.845 ;
        RECT 55.115 96.645 56.065 96.845 ;
        RECT 45.535 95.935 52.845 96.615 ;
        RECT 52.855 96.165 56.065 96.645 ;
        RECT 53.000 95.965 56.065 96.165 ;
        RECT 56.085 96.020 56.515 96.805 ;
        RECT 56.575 96.615 57.925 96.845 ;
        RECT 59.460 96.615 60.370 96.835 ;
        RECT 67.870 96.615 68.780 96.835 ;
        RECT 70.315 96.615 71.665 96.845 ;
        RECT 17.575 95.725 17.745 95.935 ;
        RECT 18.955 95.725 19.125 95.935 ;
        RECT 21.710 95.725 21.880 95.915 ;
        RECT 24.475 95.745 24.645 95.935 ;
        RECT 26.320 95.915 26.485 95.935 ;
        RECT 25.395 95.725 25.565 95.915 ;
        RECT 26.315 95.745 26.485 95.915 ;
        RECT 28.615 95.745 28.785 95.935 ;
        RECT 30.915 95.745 31.085 95.935 ;
        RECT 32.755 95.725 32.925 95.915 ;
        RECT 34.595 95.745 34.765 95.935 ;
        RECT 37.815 95.915 37.980 95.935 ;
        RECT 35.055 95.725 35.225 95.915 ;
        RECT 35.515 95.725 35.685 95.915 ;
        RECT 37.815 95.745 37.985 95.915 ;
        RECT 38.275 95.745 38.445 95.935 ;
        RECT 39.190 95.775 39.310 95.885 ;
        RECT 17.435 94.915 18.805 95.725 ;
        RECT 18.815 94.915 21.565 95.725 ;
        RECT 21.595 94.815 22.945 95.725 ;
        RECT 22.955 95.045 25.705 95.725 ;
        RECT 25.755 95.045 33.065 95.725 ;
        RECT 33.075 95.045 35.365 95.725 ;
        RECT 22.955 94.815 23.885 95.045 ;
        RECT 25.755 94.815 27.105 95.045 ;
        RECT 28.640 94.825 29.550 95.045 ;
        RECT 33.075 94.815 33.995 95.045 ;
        RECT 35.375 94.915 39.045 95.725 ;
        RECT 39.515 95.695 40.450 95.725 ;
        RECT 42.410 95.695 42.580 95.915 ;
        RECT 42.870 95.775 42.990 95.885 ;
        RECT 43.795 95.725 43.965 95.915 ;
        RECT 46.095 95.725 46.265 95.915 ;
        RECT 48.850 95.775 48.970 95.885 ;
        RECT 49.315 95.745 49.485 95.915 ;
        RECT 52.535 95.745 52.705 95.935 ;
        RECT 53.000 95.745 53.170 95.965 ;
        RECT 55.130 95.935 56.065 95.965 ;
        RECT 56.575 95.935 63.885 96.615 ;
        RECT 64.355 95.935 71.665 96.615 ;
        RECT 71.715 95.935 77.225 96.745 ;
        RECT 77.235 95.935 79.065 96.745 ;
        RECT 79.845 96.615 80.775 96.845 ;
        RECT 79.845 95.935 81.680 96.615 ;
        RECT 81.845 96.020 82.275 96.805 ;
        RECT 82.295 95.935 85.770 96.845 ;
        RECT 86.435 95.935 89.645 96.845 ;
        RECT 93.170 96.615 94.080 96.835 ;
        RECT 95.615 96.615 96.965 96.845 ;
        RECT 89.655 95.935 96.965 96.615 ;
        RECT 97.325 96.615 98.255 96.845 ;
        RECT 97.325 95.935 99.160 96.615 ;
        RECT 99.775 95.935 101.965 96.845 ;
        RECT 102.275 96.755 103.225 96.845 ;
        RECT 102.275 95.935 104.205 96.755 ;
        RECT 104.375 95.935 107.125 96.745 ;
        RECT 107.605 96.020 108.035 96.805 ;
        RECT 108.055 95.935 111.725 96.745 ;
        RECT 111.735 95.935 113.105 96.745 ;
        RECT 113.115 95.935 115.305 96.845 ;
        RECT 118.930 96.615 119.840 96.835 ;
        RECT 121.375 96.615 122.725 96.845 ;
        RECT 115.415 95.935 122.725 96.615 ;
        RECT 122.775 95.935 128.285 96.745 ;
        RECT 129.065 96.615 129.995 96.845 ;
        RECT 131.365 96.615 132.295 96.845 ;
        RECT 129.065 95.935 130.900 96.615 ;
        RECT 131.365 95.935 133.200 96.615 ;
        RECT 133.365 96.020 133.795 96.805 ;
        RECT 133.815 95.935 137.025 96.845 ;
        RECT 138.085 96.615 139.015 96.845 ;
        RECT 140.280 96.615 141.625 96.845 ;
        RECT 137.180 95.935 139.015 96.615 ;
        RECT 139.795 95.935 141.625 96.615 ;
        RECT 141.635 95.935 143.005 96.745 ;
        RECT 49.320 95.725 49.485 95.745 ;
        RECT 58.515 95.725 58.685 95.915 ;
        RECT 58.975 95.725 59.145 95.915 ;
        RECT 63.575 95.745 63.745 95.935 ;
        RECT 64.030 95.775 64.150 95.885 ;
        RECT 64.495 95.725 64.665 95.935 ;
        RECT 68.185 95.770 68.345 95.880 ;
        RECT 69.555 95.725 69.725 95.915 ;
        RECT 71.855 95.745 72.025 95.935 ;
        RECT 75.075 95.725 75.245 95.915 ;
        RECT 77.375 95.745 77.545 95.935 ;
        RECT 81.515 95.915 81.680 95.935 ;
        RECT 77.830 95.775 77.950 95.885 ;
        RECT 78.300 95.725 78.470 95.915 ;
        RECT 79.210 95.775 79.330 95.885 ;
        RECT 81.515 95.745 81.685 95.915 ;
        RECT 82.440 95.745 82.610 95.935 ;
        RECT 83.815 95.745 83.985 95.915 ;
        RECT 83.815 95.725 83.980 95.745 ;
        RECT 84.275 95.725 84.445 95.915 ;
        RECT 86.110 95.775 86.230 95.885 ;
        RECT 86.565 95.745 86.735 95.935 ;
        RECT 87.025 95.725 87.195 95.915 ;
        RECT 89.795 95.745 89.965 95.935 ;
        RECT 98.995 95.915 99.160 95.935 ;
        RECT 90.250 95.775 90.370 95.885 ;
        RECT 90.720 95.725 90.890 95.915 ;
        RECT 94.390 95.775 94.510 95.885 ;
        RECT 95.315 95.725 95.485 95.915 ;
        RECT 98.995 95.745 99.165 95.915 ;
        RECT 99.450 95.775 99.570 95.885 ;
        RECT 99.920 95.745 100.090 95.935 ;
        RECT 104.055 95.915 104.205 95.935 ;
        RECT 100.835 95.725 101.005 95.915 ;
        RECT 102.675 95.725 102.845 95.915 ;
        RECT 104.055 95.745 104.225 95.915 ;
        RECT 104.515 95.745 104.685 95.935 ;
        RECT 107.270 95.775 107.390 95.885 ;
        RECT 108.195 95.745 108.365 95.935 ;
        RECT 110.035 95.725 110.205 95.915 ;
        RECT 111.875 95.745 112.045 95.935 ;
        RECT 113.260 95.745 113.430 95.935 ;
        RECT 114.635 95.725 114.805 95.915 ;
        RECT 115.095 95.725 115.265 95.915 ;
        RECT 115.555 95.745 115.725 95.935 ;
        RECT 116.940 95.725 117.110 95.915 ;
        RECT 121.075 95.725 121.245 95.915 ;
        RECT 122.915 95.745 123.085 95.935 ;
        RECT 130.735 95.915 130.900 95.935 ;
        RECT 133.035 95.915 133.200 95.935 ;
        RECT 128.430 95.775 128.550 95.885 ;
        RECT 130.735 95.745 130.905 95.915 ;
        RECT 132.110 95.725 132.280 95.915 ;
        RECT 132.575 95.725 132.745 95.915 ;
        RECT 133.035 95.745 133.205 95.915 ;
        RECT 136.715 95.745 136.885 95.935 ;
        RECT 137.180 95.915 137.345 95.935 ;
        RECT 137.175 95.745 137.345 95.915 ;
        RECT 139.470 95.775 139.590 95.885 ;
        RECT 139.935 95.725 140.105 95.935 ;
        RECT 142.695 95.725 142.865 95.935 ;
        RECT 39.515 95.495 42.580 95.695 ;
        RECT 39.515 95.015 42.725 95.495 ;
        RECT 39.515 94.815 40.465 95.015 ;
        RECT 41.795 94.815 42.725 95.015 ;
        RECT 43.205 94.855 43.635 95.640 ;
        RECT 43.655 95.045 45.945 95.725 ;
        RECT 45.025 94.815 45.945 95.045 ;
        RECT 45.955 94.915 48.705 95.725 ;
        RECT 49.320 95.045 51.155 95.725 ;
        RECT 50.225 94.815 51.155 95.045 ;
        RECT 51.515 95.045 58.825 95.725 ;
        RECT 51.515 94.815 52.865 95.045 ;
        RECT 54.400 94.825 55.310 95.045 ;
        RECT 58.835 94.915 64.345 95.725 ;
        RECT 64.355 94.915 68.025 95.725 ;
        RECT 68.965 94.855 69.395 95.640 ;
        RECT 69.415 94.915 74.925 95.725 ;
        RECT 74.935 94.915 77.685 95.725 ;
        RECT 78.155 94.815 81.630 95.725 ;
        RECT 82.145 95.045 83.980 95.725 ;
        RECT 82.145 94.815 83.075 95.045 ;
        RECT 84.135 94.915 86.885 95.725 ;
        RECT 86.895 94.815 90.105 95.725 ;
        RECT 90.575 94.815 94.050 95.725 ;
        RECT 94.725 94.855 95.155 95.640 ;
        RECT 95.175 94.915 100.685 95.725 ;
        RECT 100.695 94.915 102.525 95.725 ;
        RECT 102.535 95.045 109.845 95.725 ;
        RECT 106.050 94.825 106.960 95.045 ;
        RECT 108.495 94.815 109.845 95.045 ;
        RECT 109.895 94.915 111.725 95.725 ;
        RECT 111.735 94.815 114.945 95.725 ;
        RECT 114.955 94.915 116.785 95.725 ;
        RECT 116.795 94.815 120.270 95.725 ;
        RECT 120.485 94.855 120.915 95.640 ;
        RECT 120.935 95.045 128.245 95.725 ;
        RECT 124.450 94.825 125.360 95.045 ;
        RECT 126.895 94.815 128.245 95.045 ;
        RECT 128.950 94.815 132.425 95.725 ;
        RECT 132.435 95.045 139.745 95.725 ;
        RECT 139.795 95.045 141.625 95.725 ;
        RECT 135.950 94.825 136.860 95.045 ;
        RECT 138.395 94.815 139.745 95.045 ;
        RECT 140.280 94.815 141.625 95.045 ;
        RECT 141.635 94.915 143.005 95.725 ;
      LAYER nwell ;
        RECT 17.240 91.695 143.200 94.525 ;
      LAYER pwell ;
        RECT 17.435 90.495 18.805 91.305 ;
        RECT 18.815 90.495 22.485 91.305 ;
        RECT 26.010 91.175 26.920 91.395 ;
        RECT 28.455 91.175 29.805 91.405 ;
        RECT 22.495 90.495 29.805 91.175 ;
        RECT 30.325 90.580 30.755 91.365 ;
        RECT 30.775 90.495 36.285 91.305 ;
        RECT 36.295 90.495 41.805 91.305 ;
        RECT 41.815 90.495 47.325 91.305 ;
        RECT 47.335 90.495 52.845 91.305 ;
        RECT 52.855 90.495 54.205 91.405 ;
        RECT 54.235 90.495 56.065 91.305 ;
        RECT 56.085 90.580 56.515 91.365 ;
        RECT 56.535 90.495 62.045 91.305 ;
        RECT 62.055 90.495 67.565 91.305 ;
        RECT 67.575 90.495 73.085 91.305 ;
        RECT 73.095 90.495 74.465 91.305 ;
        RECT 77.990 91.175 78.900 91.395 ;
        RECT 80.435 91.175 81.785 91.405 ;
        RECT 74.475 90.495 81.785 91.175 ;
        RECT 81.845 90.580 82.275 91.365 ;
        RECT 82.295 90.495 85.770 91.405 ;
        RECT 86.920 91.175 88.265 91.405 ;
        RECT 86.435 90.495 88.265 91.175 ;
        RECT 88.275 90.495 91.025 91.305 ;
        RECT 91.035 90.495 94.245 91.405 ;
        RECT 94.255 90.495 99.765 91.305 ;
        RECT 99.775 90.495 101.605 91.305 ;
        RECT 102.075 90.495 105.550 91.405 ;
        RECT 105.755 91.175 107.100 91.405 ;
        RECT 105.755 90.495 107.585 91.175 ;
        RECT 107.605 90.580 108.035 91.365 ;
        RECT 108.365 91.175 109.295 91.405 ;
        RECT 108.365 90.495 110.200 91.175 ;
        RECT 110.355 90.495 115.865 91.305 ;
        RECT 115.875 90.495 117.705 91.305 ;
        RECT 119.225 91.175 120.155 91.405 ;
        RECT 120.960 91.175 122.305 91.405 ;
        RECT 118.320 90.495 120.155 91.175 ;
        RECT 120.475 90.495 122.305 91.175 ;
        RECT 122.315 90.495 127.825 91.305 ;
        RECT 127.835 90.495 129.665 91.305 ;
        RECT 129.870 90.495 133.345 91.405 ;
        RECT 133.365 90.580 133.795 91.365 ;
        RECT 137.330 91.175 138.240 91.395 ;
        RECT 139.775 91.175 141.125 91.405 ;
        RECT 133.815 90.495 141.125 91.175 ;
        RECT 141.635 90.495 143.005 91.305 ;
        RECT 17.575 90.285 17.745 90.495 ;
        RECT 18.955 90.285 19.125 90.495 ;
        RECT 22.635 90.305 22.805 90.495 ;
        RECT 24.475 90.285 24.645 90.475 ;
        RECT 29.995 90.445 30.165 90.475 ;
        RECT 29.990 90.335 30.165 90.445 ;
        RECT 29.995 90.285 30.165 90.335 ;
        RECT 30.915 90.305 31.085 90.495 ;
        RECT 35.515 90.285 35.685 90.475 ;
        RECT 36.435 90.305 36.605 90.495 ;
        RECT 41.035 90.285 41.205 90.475 ;
        RECT 41.955 90.305 42.125 90.495 ;
        RECT 42.870 90.335 42.990 90.445 ;
        RECT 43.795 90.285 43.965 90.475 ;
        RECT 47.475 90.305 47.645 90.495 ;
        RECT 49.315 90.285 49.485 90.475 ;
        RECT 53.920 90.305 54.090 90.495 ;
        RECT 54.375 90.305 54.545 90.495 ;
        RECT 54.835 90.285 55.005 90.475 ;
        RECT 56.675 90.305 56.845 90.495 ;
        RECT 60.355 90.285 60.525 90.475 ;
        RECT 62.195 90.305 62.365 90.495 ;
        RECT 65.875 90.285 66.045 90.475 ;
        RECT 67.715 90.305 67.885 90.495 ;
        RECT 68.630 90.335 68.750 90.445 ;
        RECT 69.555 90.285 69.725 90.475 ;
        RECT 73.235 90.305 73.405 90.495 ;
        RECT 74.615 90.305 74.785 90.495 ;
        RECT 82.440 90.475 82.610 90.495 ;
        RECT 75.075 90.285 75.245 90.475 ;
        RECT 82.435 90.305 82.610 90.475 ;
        RECT 82.435 90.285 82.605 90.305 ;
        RECT 83.820 90.285 83.990 90.475 ;
        RECT 86.110 90.335 86.230 90.445 ;
        RECT 86.575 90.305 86.745 90.495 ;
        RECT 87.500 90.285 87.670 90.475 ;
        RECT 88.415 90.305 88.585 90.495 ;
        RECT 93.935 90.285 94.105 90.495 ;
        RECT 94.395 90.445 94.565 90.495 ;
        RECT 94.390 90.335 94.565 90.445 ;
        RECT 94.395 90.305 94.565 90.335 ;
        RECT 95.315 90.305 95.485 90.475 ;
        RECT 99.915 90.305 100.085 90.495 ;
        RECT 95.320 90.285 95.485 90.305 ;
        RECT 100.830 90.285 101.000 90.475 ;
        RECT 101.295 90.285 101.465 90.475 ;
        RECT 101.750 90.335 101.870 90.445 ;
        RECT 102.220 90.305 102.390 90.495 ;
        RECT 102.675 90.285 102.845 90.475 ;
        RECT 107.275 90.305 107.445 90.495 ;
        RECT 110.035 90.475 110.200 90.495 ;
        RECT 110.035 90.305 110.210 90.475 ;
        RECT 110.495 90.305 110.665 90.495 ;
        RECT 110.040 90.285 110.210 90.305 ;
        RECT 113.715 90.285 113.885 90.475 ;
        RECT 116.015 90.305 116.185 90.495 ;
        RECT 118.320 90.475 118.485 90.495 ;
        RECT 116.935 90.285 117.105 90.475 ;
        RECT 117.850 90.335 117.970 90.445 ;
        RECT 118.315 90.305 118.485 90.475 ;
        RECT 120.615 90.305 120.785 90.495 ;
        RECT 122.455 90.305 122.625 90.495 ;
        RECT 118.320 90.285 118.485 90.305 ;
        RECT 124.290 90.285 124.460 90.475 ;
        RECT 124.750 90.335 124.870 90.445 ;
        RECT 125.220 90.285 125.390 90.475 ;
        RECT 127.975 90.305 128.145 90.495 ;
        RECT 128.890 90.335 129.010 90.445 ;
        RECT 133.030 90.305 133.200 90.495 ;
        RECT 133.955 90.305 134.125 90.495 ;
        RECT 136.255 90.285 136.425 90.475 ;
        RECT 136.715 90.285 136.885 90.475 ;
        RECT 138.095 90.285 138.265 90.475 ;
        RECT 139.935 90.285 140.105 90.475 ;
        RECT 141.310 90.335 141.430 90.445 ;
        RECT 142.695 90.285 142.865 90.495 ;
        RECT 17.435 89.475 18.805 90.285 ;
        RECT 18.815 89.475 24.325 90.285 ;
        RECT 24.335 89.475 29.845 90.285 ;
        RECT 29.855 89.475 35.365 90.285 ;
        RECT 35.375 89.475 40.885 90.285 ;
        RECT 40.895 89.475 42.725 90.285 ;
        RECT 43.205 89.415 43.635 90.200 ;
        RECT 43.655 89.475 49.165 90.285 ;
        RECT 49.175 89.475 54.685 90.285 ;
        RECT 54.695 89.475 60.205 90.285 ;
        RECT 60.215 89.475 65.725 90.285 ;
        RECT 65.735 89.475 68.485 90.285 ;
        RECT 68.965 89.415 69.395 90.200 ;
        RECT 69.415 89.475 74.925 90.285 ;
        RECT 74.935 89.605 82.245 90.285 ;
        RECT 78.450 89.385 79.360 89.605 ;
        RECT 80.895 89.375 82.245 89.605 ;
        RECT 82.295 89.475 83.665 90.285 ;
        RECT 83.675 89.375 87.150 90.285 ;
        RECT 87.355 89.375 90.830 90.285 ;
        RECT 91.035 89.375 94.245 90.285 ;
        RECT 94.725 89.415 95.155 90.200 ;
        RECT 95.320 89.605 97.155 90.285 ;
        RECT 96.225 89.375 97.155 89.605 ;
        RECT 97.670 89.375 101.145 90.285 ;
        RECT 101.155 89.475 102.525 90.285 ;
        RECT 102.535 89.605 109.845 90.285 ;
        RECT 106.050 89.385 106.960 89.605 ;
        RECT 108.495 89.375 109.845 89.605 ;
        RECT 109.895 89.375 113.370 90.285 ;
        RECT 113.575 89.375 116.785 90.285 ;
        RECT 116.795 89.475 118.165 90.285 ;
        RECT 118.320 89.605 120.155 90.285 ;
        RECT 119.225 89.375 120.155 89.605 ;
        RECT 120.485 89.415 120.915 90.200 ;
        RECT 121.130 89.375 124.605 90.285 ;
        RECT 125.075 89.375 128.550 90.285 ;
        RECT 129.255 89.605 136.565 90.285 ;
        RECT 129.255 89.375 130.605 89.605 ;
        RECT 132.140 89.385 133.050 89.605 ;
        RECT 136.575 89.475 137.945 90.285 ;
        RECT 137.955 89.605 139.785 90.285 ;
        RECT 139.795 89.605 141.625 90.285 ;
        RECT 138.440 89.375 139.785 89.605 ;
        RECT 140.280 89.375 141.625 89.605 ;
        RECT 141.635 89.475 143.005 90.285 ;
      LAYER nwell ;
        RECT 17.240 86.255 143.200 89.085 ;
      LAYER pwell ;
        RECT 17.435 85.055 18.805 85.865 ;
        RECT 18.815 85.055 24.325 85.865 ;
        RECT 24.335 85.055 29.845 85.865 ;
        RECT 30.325 85.140 30.755 85.925 ;
        RECT 30.775 85.055 36.285 85.865 ;
        RECT 36.295 85.055 41.805 85.865 ;
        RECT 41.815 85.055 47.325 85.865 ;
        RECT 47.335 85.055 52.845 85.865 ;
        RECT 52.855 85.055 55.605 85.865 ;
        RECT 56.085 85.140 56.515 85.925 ;
        RECT 56.535 85.055 62.045 85.865 ;
        RECT 62.055 85.055 67.565 85.865 ;
        RECT 67.575 85.055 73.085 85.865 ;
        RECT 73.095 85.055 78.605 85.865 ;
        RECT 78.615 85.055 81.365 85.865 ;
        RECT 81.845 85.140 82.275 85.925 ;
        RECT 85.810 85.735 86.720 85.955 ;
        RECT 88.255 85.735 89.605 85.965 ;
        RECT 82.295 85.055 89.605 85.735 ;
        RECT 89.655 85.055 91.025 85.865 ;
        RECT 94.550 85.735 95.460 85.955 ;
        RECT 96.995 85.735 98.345 85.965 ;
        RECT 101.910 85.735 102.820 85.955 ;
        RECT 104.355 85.735 105.705 85.965 ;
        RECT 91.035 85.055 98.345 85.735 ;
        RECT 98.395 85.055 105.705 85.735 ;
        RECT 105.755 85.055 107.585 85.735 ;
        RECT 107.605 85.140 108.035 85.925 ;
        RECT 108.055 85.055 111.530 85.965 ;
        RECT 111.735 85.055 114.945 85.965 ;
        RECT 115.455 85.735 116.805 85.965 ;
        RECT 118.340 85.735 119.250 85.955 ;
        RECT 126.290 85.735 127.200 85.955 ;
        RECT 128.735 85.735 130.085 85.965 ;
        RECT 115.455 85.055 122.765 85.735 ;
        RECT 122.775 85.055 130.085 85.735 ;
        RECT 130.445 85.735 131.375 85.965 ;
        RECT 130.445 85.055 132.280 85.735 ;
        RECT 133.365 85.140 133.795 85.925 ;
        RECT 134.010 85.055 137.485 85.965 ;
        RECT 137.495 85.055 139.325 85.865 ;
        RECT 140.280 85.735 141.625 85.965 ;
        RECT 139.795 85.055 141.625 85.735 ;
        RECT 141.635 85.055 143.005 85.865 ;
        RECT 17.575 84.845 17.745 85.055 ;
        RECT 18.955 84.845 19.125 85.055 ;
        RECT 24.475 84.845 24.645 85.055 ;
        RECT 29.995 85.005 30.165 85.035 ;
        RECT 29.990 84.895 30.165 85.005 ;
        RECT 29.995 84.845 30.165 84.895 ;
        RECT 30.915 84.865 31.085 85.055 ;
        RECT 35.515 84.845 35.685 85.035 ;
        RECT 36.435 84.865 36.605 85.055 ;
        RECT 41.035 84.845 41.205 85.035 ;
        RECT 41.955 84.865 42.125 85.055 ;
        RECT 42.870 84.895 42.990 85.005 ;
        RECT 43.795 84.845 43.965 85.035 ;
        RECT 47.475 84.865 47.645 85.055 ;
        RECT 49.315 84.845 49.485 85.035 ;
        RECT 52.995 84.865 53.165 85.055 ;
        RECT 54.835 84.845 55.005 85.035 ;
        RECT 55.750 84.895 55.870 85.005 ;
        RECT 56.675 84.865 56.845 85.055 ;
        RECT 60.355 84.845 60.525 85.035 ;
        RECT 62.195 84.865 62.365 85.055 ;
        RECT 65.875 84.845 66.045 85.035 ;
        RECT 67.715 84.865 67.885 85.055 ;
        RECT 68.630 84.895 68.750 85.005 ;
        RECT 69.555 84.845 69.725 85.035 ;
        RECT 73.235 84.865 73.405 85.055 ;
        RECT 75.075 84.845 75.245 85.035 ;
        RECT 78.755 84.865 78.925 85.055 ;
        RECT 80.595 84.845 80.765 85.035 ;
        RECT 81.510 84.895 81.630 85.005 ;
        RECT 82.435 84.865 82.605 85.055 ;
        RECT 89.795 84.865 89.965 85.055 ;
        RECT 91.175 84.865 91.345 85.055 ;
        RECT 92.095 84.865 92.265 85.035 ;
        RECT 89.795 84.845 89.960 84.865 ;
        RECT 92.095 84.845 92.260 84.865 ;
        RECT 92.555 84.845 92.725 85.035 ;
        RECT 94.390 84.895 94.510 85.005 ;
        RECT 95.320 84.845 95.490 85.035 ;
        RECT 98.535 84.865 98.705 85.055 ;
        RECT 98.990 84.895 99.110 85.005 ;
        RECT 101.295 84.865 101.465 85.035 ;
        RECT 105.895 84.865 106.065 85.055 ;
        RECT 108.200 84.865 108.370 85.055 ;
        RECT 101.295 84.845 101.460 84.865 ;
        RECT 108.655 84.845 108.825 85.035 ;
        RECT 109.115 84.865 109.285 85.035 ;
        RECT 109.120 84.845 109.285 84.865 ;
        RECT 111.415 84.845 111.585 85.035 ;
        RECT 111.875 84.865 112.045 85.055 ;
        RECT 115.090 84.895 115.210 85.005 ;
        RECT 116.015 84.845 116.185 85.035 ;
        RECT 116.475 84.845 116.645 85.035 ;
        RECT 119.705 84.890 119.865 85.000 ;
        RECT 121.080 84.845 121.250 85.035 ;
        RECT 122.455 84.865 122.625 85.055 ;
        RECT 122.915 84.865 123.085 85.055 ;
        RECT 132.115 85.035 132.280 85.055 ;
        RECT 124.750 84.895 124.870 85.005 ;
        RECT 125.215 84.845 125.385 85.035 ;
        RECT 132.115 84.865 132.285 85.035 ;
        RECT 132.575 84.865 132.745 85.035 ;
        RECT 132.580 84.845 132.745 84.865 ;
        RECT 134.875 84.845 135.045 85.035 ;
        RECT 137.170 84.865 137.340 85.055 ;
        RECT 137.635 84.865 137.805 85.055 ;
        RECT 138.555 84.845 138.725 85.035 ;
        RECT 139.470 84.895 139.590 85.005 ;
        RECT 139.935 84.845 140.105 85.055 ;
        RECT 142.695 84.845 142.865 85.055 ;
        RECT 17.435 84.035 18.805 84.845 ;
        RECT 18.815 84.035 24.325 84.845 ;
        RECT 24.335 84.035 29.845 84.845 ;
        RECT 29.855 84.035 35.365 84.845 ;
        RECT 35.375 84.035 40.885 84.845 ;
        RECT 40.895 84.035 42.725 84.845 ;
        RECT 43.205 83.975 43.635 84.760 ;
        RECT 43.655 84.035 49.165 84.845 ;
        RECT 49.175 84.035 54.685 84.845 ;
        RECT 54.695 84.035 60.205 84.845 ;
        RECT 60.215 84.035 65.725 84.845 ;
        RECT 65.735 84.035 68.485 84.845 ;
        RECT 68.965 83.975 69.395 84.760 ;
        RECT 69.415 84.035 74.925 84.845 ;
        RECT 74.935 84.035 80.445 84.845 ;
        RECT 80.455 84.165 87.765 84.845 ;
        RECT 83.970 83.945 84.880 84.165 ;
        RECT 86.415 83.935 87.765 84.165 ;
        RECT 88.125 84.165 89.960 84.845 ;
        RECT 90.425 84.165 92.260 84.845 ;
        RECT 88.125 83.935 89.055 84.165 ;
        RECT 90.425 83.935 91.355 84.165 ;
        RECT 92.415 84.035 94.245 84.845 ;
        RECT 94.725 83.975 95.155 84.760 ;
        RECT 95.175 83.935 98.650 84.845 ;
        RECT 99.625 84.165 101.460 84.845 ;
        RECT 101.655 84.165 108.965 84.845 ;
        RECT 109.120 84.165 110.955 84.845 ;
        RECT 99.625 83.935 100.555 84.165 ;
        RECT 101.655 83.935 103.005 84.165 ;
        RECT 104.540 83.945 105.450 84.165 ;
        RECT 110.025 83.935 110.955 84.165 ;
        RECT 111.275 84.035 113.105 84.845 ;
        RECT 113.115 83.935 116.325 84.845 ;
        RECT 116.335 83.935 119.545 84.845 ;
        RECT 120.485 83.975 120.915 84.760 ;
        RECT 120.935 83.935 124.410 84.845 ;
        RECT 125.075 84.165 132.385 84.845 ;
        RECT 132.580 84.165 134.415 84.845 ;
        RECT 128.590 83.945 129.500 84.165 ;
        RECT 131.035 83.935 132.385 84.165 ;
        RECT 133.485 83.935 134.415 84.165 ;
        RECT 134.735 84.035 138.405 84.845 ;
        RECT 138.415 84.035 139.785 84.845 ;
        RECT 139.795 84.165 141.625 84.845 ;
        RECT 140.280 83.935 141.625 84.165 ;
        RECT 141.635 84.035 143.005 84.845 ;
      LAYER nwell ;
        RECT 17.240 80.815 143.200 83.645 ;
      LAYER pwell ;
        RECT 17.435 79.615 18.805 80.425 ;
        RECT 18.815 79.615 24.325 80.425 ;
        RECT 24.335 79.615 29.845 80.425 ;
        RECT 30.325 79.700 30.755 80.485 ;
        RECT 30.775 79.615 36.285 80.425 ;
        RECT 36.295 79.615 41.805 80.425 ;
        RECT 41.815 79.615 43.185 80.425 ;
        RECT 43.205 79.700 43.635 80.485 ;
        RECT 43.655 79.615 49.165 80.425 ;
        RECT 49.175 79.615 54.685 80.425 ;
        RECT 54.695 79.615 56.065 80.425 ;
        RECT 56.085 79.700 56.515 80.485 ;
        RECT 56.535 79.615 62.045 80.425 ;
        RECT 62.055 79.615 63.885 80.425 ;
        RECT 64.380 80.295 65.725 80.525 ;
        RECT 63.895 79.615 65.725 80.295 ;
        RECT 65.735 79.615 68.485 80.425 ;
        RECT 68.965 79.700 69.395 80.485 ;
        RECT 70.335 80.295 71.680 80.525 ;
        RECT 70.335 79.615 72.165 80.295 ;
        RECT 72.175 79.615 73.545 80.425 ;
        RECT 74.215 80.295 78.145 80.525 ;
        RECT 73.730 79.615 78.145 80.295 ;
        RECT 78.155 80.295 79.500 80.525 ;
        RECT 79.995 80.295 81.340 80.525 ;
        RECT 78.155 79.615 79.985 80.295 ;
        RECT 79.995 79.615 81.825 80.295 ;
        RECT 81.845 79.700 82.275 80.485 ;
        RECT 83.215 80.295 84.560 80.525 ;
        RECT 83.215 79.615 85.045 80.295 ;
        RECT 85.055 79.615 86.425 80.425 ;
        RECT 86.435 80.295 87.780 80.525 ;
        RECT 86.435 79.615 88.265 80.295 ;
        RECT 88.275 79.615 89.645 80.425 ;
        RECT 89.655 80.295 91.000 80.525 ;
        RECT 89.655 79.615 91.485 80.295 ;
        RECT 91.495 79.615 92.865 80.425 ;
        RECT 92.875 80.295 94.220 80.525 ;
        RECT 92.875 79.615 94.705 80.295 ;
        RECT 94.725 79.700 95.155 80.485 ;
        RECT 96.095 80.295 97.440 80.525 ;
        RECT 96.095 79.615 97.925 80.295 ;
        RECT 97.935 79.615 99.305 80.425 ;
        RECT 99.315 80.295 100.660 80.525 ;
        RECT 102.075 80.295 103.420 80.525 ;
        RECT 104.965 80.295 105.895 80.525 ;
        RECT 99.315 79.615 101.145 80.295 ;
        RECT 102.075 79.615 103.905 80.295 ;
        RECT 104.060 79.615 105.895 80.295 ;
        RECT 106.215 79.615 107.585 80.425 ;
        RECT 107.605 79.700 108.035 80.485 ;
        RECT 108.055 80.295 109.400 80.525 ;
        RECT 109.895 80.295 111.240 80.525 ;
        RECT 112.195 80.295 113.540 80.525 ;
        RECT 108.055 79.615 109.885 80.295 ;
        RECT 109.895 79.615 111.725 80.295 ;
        RECT 112.195 79.615 114.025 80.295 ;
        RECT 114.035 79.615 115.405 80.425 ;
        RECT 115.900 80.295 117.245 80.525 ;
        RECT 118.765 80.295 119.695 80.525 ;
        RECT 115.415 79.615 117.245 80.295 ;
        RECT 117.860 79.615 119.695 80.295 ;
        RECT 120.485 79.700 120.915 80.485 ;
        RECT 121.420 80.295 122.765 80.525 ;
        RECT 123.260 80.295 124.605 80.525 ;
        RECT 120.935 79.615 122.765 80.295 ;
        RECT 122.775 79.615 124.605 80.295 ;
        RECT 125.075 80.295 126.420 80.525 ;
        RECT 125.075 79.615 126.905 80.295 ;
        RECT 126.915 79.615 128.285 80.425 ;
        RECT 128.780 80.295 130.125 80.525 ;
        RECT 128.295 79.615 130.125 80.295 ;
        RECT 130.135 79.615 131.505 80.425 ;
        RECT 132.000 80.295 133.345 80.525 ;
        RECT 131.515 79.615 133.345 80.295 ;
        RECT 133.365 79.700 133.795 80.485 ;
        RECT 134.735 80.295 136.080 80.525 ;
        RECT 134.735 79.615 136.565 80.295 ;
        RECT 136.575 79.615 140.245 80.425 ;
        RECT 140.255 79.615 141.625 80.425 ;
        RECT 141.635 79.615 143.005 80.425 ;
        RECT 17.575 79.425 17.745 79.615 ;
        RECT 18.955 79.425 19.125 79.615 ;
        RECT 24.475 79.425 24.645 79.615 ;
        RECT 29.990 79.455 30.110 79.565 ;
        RECT 30.915 79.425 31.085 79.615 ;
        RECT 36.435 79.425 36.605 79.615 ;
        RECT 41.955 79.425 42.125 79.615 ;
        RECT 43.795 79.425 43.965 79.615 ;
        RECT 49.315 79.425 49.485 79.615 ;
        RECT 54.835 79.425 55.005 79.615 ;
        RECT 56.675 79.425 56.845 79.615 ;
        RECT 62.195 79.425 62.365 79.615 ;
        RECT 64.035 79.425 64.205 79.615 ;
        RECT 65.875 79.425 66.045 79.615 ;
        RECT 68.630 79.455 68.750 79.565 ;
        RECT 69.565 79.460 69.725 79.570 ;
        RECT 71.855 79.425 72.025 79.615 ;
        RECT 72.315 79.425 72.485 79.615 ;
        RECT 73.730 79.595 73.840 79.615 ;
        RECT 73.670 79.425 73.840 79.595 ;
        RECT 79.675 79.425 79.845 79.615 ;
        RECT 81.515 79.425 81.685 79.615 ;
        RECT 82.445 79.460 82.605 79.570 ;
        RECT 84.735 79.425 84.905 79.615 ;
        RECT 85.195 79.425 85.365 79.615 ;
        RECT 87.955 79.425 88.125 79.615 ;
        RECT 88.415 79.425 88.585 79.615 ;
        RECT 91.175 79.425 91.345 79.615 ;
        RECT 91.635 79.425 91.805 79.615 ;
        RECT 94.395 79.425 94.565 79.615 ;
        RECT 95.325 79.460 95.485 79.570 ;
        RECT 97.615 79.425 97.785 79.615 ;
        RECT 98.075 79.425 98.245 79.615 ;
        RECT 100.835 79.425 101.005 79.615 ;
        RECT 101.305 79.460 101.465 79.570 ;
        RECT 103.595 79.425 103.765 79.615 ;
        RECT 104.060 79.595 104.225 79.615 ;
        RECT 104.055 79.425 104.225 79.595 ;
        RECT 106.355 79.425 106.525 79.615 ;
        RECT 109.575 79.425 109.745 79.615 ;
        RECT 111.415 79.425 111.585 79.615 ;
        RECT 111.870 79.455 111.990 79.565 ;
        RECT 113.715 79.425 113.885 79.615 ;
        RECT 114.175 79.425 114.345 79.615 ;
        RECT 115.555 79.425 115.725 79.615 ;
        RECT 117.860 79.595 118.025 79.615 ;
        RECT 117.390 79.455 117.510 79.565 ;
        RECT 117.855 79.425 118.025 79.595 ;
        RECT 120.150 79.455 120.270 79.565 ;
        RECT 121.075 79.425 121.245 79.615 ;
        RECT 122.915 79.425 123.085 79.615 ;
        RECT 124.750 79.455 124.870 79.565 ;
        RECT 126.595 79.425 126.765 79.615 ;
        RECT 127.055 79.425 127.225 79.615 ;
        RECT 128.435 79.425 128.605 79.615 ;
        RECT 130.275 79.425 130.445 79.615 ;
        RECT 131.655 79.425 131.825 79.615 ;
        RECT 133.965 79.460 134.125 79.570 ;
        RECT 136.255 79.425 136.425 79.615 ;
        RECT 136.715 79.425 136.885 79.615 ;
        RECT 140.395 79.425 140.565 79.615 ;
        RECT 142.695 79.425 142.865 79.615 ;
      LAYER nwell ;
        RECT 12.560 47.315 48.820 48.920 ;
      LAYER pwell ;
        RECT 12.755 46.115 14.125 46.925 ;
        RECT 14.135 46.115 19.645 46.925 ;
        RECT 21.060 46.795 22.405 47.025 ;
        RECT 20.575 46.115 22.405 46.795 ;
        RECT 22.545 46.115 25.545 47.025 ;
        RECT 25.645 46.200 26.075 46.985 ;
        RECT 29.670 46.795 30.590 47.025 ;
        RECT 27.125 46.115 30.590 46.795 ;
        RECT 31.615 46.795 32.960 47.025 ;
        RECT 36.110 46.795 37.030 47.025 ;
        RECT 31.615 46.115 33.445 46.795 ;
        RECT 33.565 46.115 37.030 46.795 ;
        RECT 37.135 46.115 38.505 46.895 ;
        RECT 38.525 46.200 38.955 46.985 ;
        RECT 39.895 46.795 41.240 47.025 ;
        RECT 39.895 46.115 41.725 46.795 ;
        RECT 41.735 46.115 43.105 46.925 ;
        RECT 43.115 46.115 44.485 46.895 ;
        RECT 44.495 46.115 45.865 46.895 ;
        RECT 45.875 46.115 47.245 46.895 ;
        RECT 47.255 46.115 48.625 46.925 ;
        RECT 12.895 45.905 13.065 46.115 ;
        RECT 14.275 45.905 14.445 46.115 ;
        RECT 17.950 45.955 18.070 46.065 ;
        RECT 19.805 45.960 19.965 46.070 ;
        RECT 20.715 45.925 20.885 46.115 ;
        RECT 25.315 45.905 25.485 46.115 ;
        RECT 25.775 45.905 25.945 46.095 ;
        RECT 26.245 45.960 26.405 46.070 ;
        RECT 27.155 45.925 27.325 46.115 ;
        RECT 30.845 45.960 31.005 46.070 ;
        RECT 33.135 45.925 33.305 46.115 ;
        RECT 33.595 45.925 33.765 46.115 ;
        RECT 37.285 46.095 37.455 46.115 ;
        RECT 34.975 45.925 35.145 46.095 ;
        RECT 34.975 45.905 35.140 45.925 ;
        RECT 35.435 45.905 35.605 46.095 ;
        RECT 37.275 45.925 37.455 46.095 ;
        RECT 37.275 45.905 37.445 45.925 ;
        RECT 39.115 45.905 39.285 46.095 ;
        RECT 41.415 45.925 41.585 46.115 ;
        RECT 41.875 45.925 42.045 46.115 ;
        RECT 42.335 45.905 42.505 46.095 ;
        RECT 44.175 45.925 44.345 46.115 ;
        RECT 45.555 45.925 45.725 46.115 ;
        RECT 46.925 45.905 47.095 46.115 ;
        RECT 48.315 45.905 48.485 46.115 ;
        RECT 12.755 45.095 14.125 45.905 ;
        RECT 14.135 45.095 17.805 45.905 ;
        RECT 18.315 45.225 25.625 45.905 ;
        RECT 25.635 45.225 32.945 45.905 ;
        RECT 18.315 44.995 19.665 45.225 ;
        RECT 21.200 45.005 22.110 45.225 ;
        RECT 29.150 45.005 30.060 45.225 ;
        RECT 31.595 44.995 32.945 45.225 ;
        RECT 33.305 45.225 35.140 45.905 ;
        RECT 35.295 45.225 37.125 45.905 ;
        RECT 33.305 44.995 34.235 45.225 ;
        RECT 35.780 44.995 37.125 45.225 ;
        RECT 37.145 44.995 38.495 45.905 ;
        RECT 38.525 45.035 38.955 45.820 ;
        RECT 39.055 44.995 42.055 45.905 ;
        RECT 42.305 45.225 45.770 45.905 ;
        RECT 44.850 44.995 45.770 45.225 ;
        RECT 45.875 45.125 47.245 45.905 ;
        RECT 47.255 45.095 48.625 45.905 ;
      LAYER nwell ;
        RECT 12.560 41.875 48.820 44.705 ;
      LAYER pwell ;
        RECT 12.755 40.675 14.125 41.485 ;
        RECT 17.650 41.355 18.560 41.575 ;
        RECT 20.095 41.355 21.445 41.585 ;
        RECT 14.135 40.675 21.445 41.355 ;
        RECT 21.590 41.355 22.510 41.585 ;
        RECT 21.590 40.675 25.055 41.355 ;
        RECT 25.645 40.760 26.075 41.545 ;
        RECT 26.095 41.355 27.025 41.585 ;
        RECT 31.745 41.355 32.675 41.585 ;
        RECT 26.095 40.675 29.995 41.355 ;
        RECT 30.840 40.675 32.675 41.355 ;
        RECT 33.005 40.675 34.355 41.585 ;
        RECT 37.890 41.355 38.800 41.575 ;
        RECT 40.335 41.355 41.685 41.585 ;
        RECT 43.245 41.355 44.175 41.585 ;
        RECT 34.375 40.675 41.685 41.355 ;
        RECT 42.340 40.675 44.175 41.355 ;
        RECT 44.495 40.675 45.865 41.455 ;
        RECT 45.875 40.675 47.245 41.455 ;
        RECT 47.255 40.675 48.625 41.485 ;
        RECT 12.895 40.465 13.065 40.675 ;
        RECT 14.275 40.485 14.445 40.675 ;
        RECT 15.655 40.465 15.825 40.655 ;
        RECT 16.390 40.465 16.560 40.655 ;
        RECT 20.255 40.465 20.425 40.655 ;
        RECT 24.855 40.485 25.025 40.675 ;
        RECT 25.310 40.515 25.430 40.625 ;
        RECT 26.510 40.485 26.680 40.675 ;
        RECT 30.840 40.655 31.005 40.675 ;
        RECT 30.375 40.625 30.545 40.655 ;
        RECT 30.370 40.515 30.545 40.625 ;
        RECT 30.375 40.465 30.545 40.515 ;
        RECT 30.835 40.485 31.005 40.655 ;
        RECT 34.055 40.465 34.225 40.675 ;
        RECT 34.515 40.465 34.685 40.675 ;
        RECT 42.340 40.655 42.505 40.675 ;
        RECT 12.755 39.655 14.125 40.465 ;
        RECT 14.135 39.785 15.965 40.465 ;
        RECT 15.975 39.785 19.875 40.465 ;
        RECT 14.135 39.555 15.480 39.785 ;
        RECT 15.975 39.555 16.905 39.785 ;
        RECT 20.115 39.655 21.485 40.465 ;
        RECT 21.580 39.785 30.685 40.465 ;
        RECT 30.790 39.785 34.255 40.465 ;
        RECT 30.790 39.555 31.710 39.785 ;
        RECT 34.375 39.655 35.745 40.465 ;
        RECT 35.900 40.435 36.070 40.655 ;
        RECT 39.115 40.465 39.285 40.655 ;
        RECT 41.870 40.515 41.990 40.625 ;
        RECT 42.335 40.485 42.505 40.655 ;
        RECT 42.795 40.465 42.965 40.655 ;
        RECT 44.635 40.485 44.805 40.675 ;
        RECT 46.485 40.510 46.645 40.620 ;
        RECT 46.925 40.485 47.095 40.675 ;
        RECT 48.315 40.465 48.485 40.675 ;
        RECT 37.560 40.435 38.505 40.465 ;
        RECT 35.755 39.755 38.505 40.435 ;
        RECT 37.560 39.555 38.505 39.755 ;
        RECT 38.525 39.595 38.955 40.380 ;
        RECT 39.055 39.555 42.505 40.465 ;
        RECT 42.735 39.555 46.185 40.465 ;
        RECT 47.255 39.655 48.625 40.465 ;
      LAYER nwell ;
        RECT 12.560 36.435 48.820 39.265 ;
      LAYER pwell ;
        RECT 12.755 35.235 14.125 36.045 ;
        RECT 14.135 35.915 15.065 36.145 ;
        RECT 21.790 35.915 22.700 36.135 ;
        RECT 24.235 35.915 25.585 36.145 ;
        RECT 14.135 35.235 18.035 35.915 ;
        RECT 18.275 35.235 25.585 35.915 ;
        RECT 25.645 35.320 26.075 36.105 ;
        RECT 29.610 35.915 30.520 36.135 ;
        RECT 32.055 35.915 33.405 36.145 ;
        RECT 26.095 35.235 33.405 35.915 ;
        RECT 33.915 35.915 35.280 36.145 ;
        RECT 33.915 35.235 37.125 35.915 ;
        RECT 38.135 35.235 41.135 36.145 ;
        RECT 41.275 35.235 42.625 36.145 ;
        RECT 43.195 35.235 46.645 36.145 ;
        RECT 47.255 35.235 48.625 36.045 ;
        RECT 12.895 35.025 13.065 35.235 ;
        RECT 14.550 35.045 14.720 35.235 ;
        RECT 18.415 35.045 18.585 35.235 ;
        RECT 21.175 35.025 21.345 35.215 ;
        RECT 21.635 35.025 21.805 35.215 ;
        RECT 24.390 35.075 24.510 35.185 ;
        RECT 24.855 35.025 25.025 35.215 ;
        RECT 26.235 35.045 26.405 35.235 ;
        RECT 33.590 35.075 33.710 35.185 ;
        RECT 36.810 35.045 36.980 35.235 ;
        RECT 37.275 35.025 37.445 35.215 ;
        RECT 37.745 35.070 37.905 35.180 ;
        RECT 38.195 35.045 38.365 35.235 ;
        RECT 41.420 35.215 41.590 35.235 ;
        RECT 12.755 34.215 14.125 35.025 ;
        RECT 14.175 34.345 21.485 35.025 ;
        RECT 14.175 34.115 15.525 34.345 ;
        RECT 17.060 34.125 17.970 34.345 ;
        RECT 21.495 34.215 24.245 35.025 ;
        RECT 24.715 34.345 33.820 35.025 ;
        RECT 34.010 34.345 37.475 35.025 ;
        RECT 39.110 34.995 39.280 35.215 ;
        RECT 41.415 35.045 41.590 35.215 ;
        RECT 42.790 35.075 42.910 35.185 ;
        RECT 43.255 35.045 43.425 35.235 ;
        RECT 44.170 35.075 44.290 35.185 ;
        RECT 41.415 35.025 41.585 35.045 ;
        RECT 45.550 35.025 45.720 35.215 ;
        RECT 46.935 35.185 47.105 35.215 ;
        RECT 46.930 35.075 47.105 35.185 ;
        RECT 46.935 35.025 47.105 35.075 ;
        RECT 48.315 35.025 48.485 35.235 ;
        RECT 40.310 34.995 41.265 35.025 ;
        RECT 34.010 34.115 34.930 34.345 ;
        RECT 38.525 34.155 38.955 34.940 ;
        RECT 38.985 34.315 41.265 34.995 ;
        RECT 40.310 34.115 41.265 34.315 ;
        RECT 41.275 34.215 44.025 35.025 ;
        RECT 44.515 34.115 45.865 35.025 ;
        RECT 45.875 34.245 47.245 35.025 ;
        RECT 47.255 34.215 48.625 35.025 ;
      LAYER nwell ;
        RECT 12.560 30.995 48.820 33.825 ;
      LAYER pwell ;
        RECT 12.755 29.795 14.125 30.605 ;
        RECT 14.135 29.795 15.505 30.605 ;
        RECT 18.170 30.475 19.090 30.705 ;
        RECT 15.625 29.795 19.090 30.475 ;
        RECT 19.290 30.475 20.210 30.705 ;
        RECT 19.290 29.795 22.755 30.475 ;
        RECT 22.875 29.795 25.625 30.605 ;
        RECT 25.645 29.880 26.075 30.665 ;
        RECT 26.115 29.795 27.465 30.705 ;
        RECT 27.545 29.795 31.605 30.705 ;
        RECT 31.710 30.475 32.630 30.705 ;
        RECT 31.710 29.795 35.175 30.475 ;
        RECT 35.295 29.795 36.665 30.605 ;
        RECT 36.675 30.505 37.625 30.705 ;
        RECT 36.675 29.825 40.345 30.505 ;
        RECT 36.675 29.795 37.625 29.825 ;
        RECT 12.895 29.585 13.065 29.795 ;
        RECT 14.275 29.605 14.445 29.795 ;
        RECT 15.655 29.585 15.825 29.795 ;
        RECT 16.110 29.635 16.230 29.745 ;
        RECT 16.850 29.585 17.020 29.775 ;
        RECT 20.715 29.585 20.885 29.775 ;
        RECT 22.555 29.605 22.725 29.795 ;
        RECT 23.015 29.605 23.185 29.795 ;
        RECT 27.150 29.605 27.320 29.795 ;
        RECT 28.350 29.585 28.520 29.775 ;
        RECT 31.295 29.605 31.465 29.795 ;
        RECT 34.975 29.605 35.145 29.795 ;
        RECT 35.435 29.585 35.605 29.795 ;
        RECT 35.895 29.585 36.065 29.775 ;
        RECT 40.030 29.605 40.200 29.825 ;
        RECT 40.355 29.795 41.705 30.705 ;
        RECT 41.735 29.795 43.105 30.575 ;
        RECT 43.255 29.795 46.705 30.705 ;
        RECT 47.255 29.795 48.625 30.605 ;
        RECT 40.500 29.605 40.670 29.795 ;
        RECT 41.885 29.775 42.055 29.795 ;
        RECT 41.870 29.605 42.055 29.775 ;
        RECT 42.345 29.630 42.505 29.740 ;
        RECT 41.870 29.585 42.040 29.605 ;
        RECT 46.475 29.585 46.645 29.795 ;
        RECT 46.930 29.635 47.050 29.745 ;
        RECT 48.315 29.585 48.485 29.795 ;
        RECT 12.755 28.775 14.125 29.585 ;
        RECT 14.135 28.905 15.965 29.585 ;
        RECT 16.435 28.905 20.335 29.585 ;
        RECT 20.575 28.905 27.885 29.585 ;
        RECT 14.135 28.675 15.480 28.905 ;
        RECT 16.435 28.675 17.365 28.905 ;
        RECT 24.090 28.685 25.000 28.905 ;
        RECT 26.535 28.675 27.885 28.905 ;
        RECT 27.935 28.905 31.835 29.585 ;
        RECT 32.170 28.905 35.635 29.585 ;
        RECT 27.935 28.675 28.865 28.905 ;
        RECT 32.170 28.675 33.090 28.905 ;
        RECT 35.755 28.775 38.505 29.585 ;
        RECT 38.525 28.715 38.955 29.500 ;
        RECT 39.265 28.675 42.185 29.585 ;
        RECT 43.255 28.675 46.705 29.585 ;
        RECT 47.255 28.775 48.625 29.585 ;
      LAYER nwell ;
        RECT 12.560 25.555 48.820 28.385 ;
      LAYER pwell ;
        RECT 12.755 24.355 14.125 25.165 ;
        RECT 17.650 25.035 18.560 25.255 ;
        RECT 20.095 25.035 21.445 25.265 ;
        RECT 14.135 24.355 21.445 25.035 ;
        RECT 21.495 24.355 25.165 25.165 ;
        RECT 25.645 24.440 26.075 25.225 ;
        RECT 29.610 25.035 30.520 25.255 ;
        RECT 32.055 25.035 33.405 25.265 ;
        RECT 35.300 25.035 36.665 25.265 ;
        RECT 26.095 24.355 33.405 25.035 ;
        RECT 33.455 24.355 36.665 25.035 ;
        RECT 36.675 24.355 39.425 25.165 ;
        RECT 42.550 25.035 43.470 25.265 ;
        RECT 40.005 24.355 43.470 25.035 ;
        RECT 43.655 24.355 46.655 25.265 ;
        RECT 47.255 24.355 48.625 25.165 ;
        RECT 12.895 24.145 13.065 24.355 ;
        RECT 14.275 24.165 14.445 24.355 ;
        RECT 15.655 24.145 15.825 24.335 ;
        RECT 16.125 24.190 16.285 24.300 ;
        RECT 17.035 24.145 17.205 24.335 ;
        RECT 20.725 24.190 20.885 24.300 ;
        RECT 21.635 24.145 21.805 24.355 ;
        RECT 25.310 24.195 25.430 24.305 ;
        RECT 26.235 24.165 26.405 24.355 ;
        RECT 28.720 24.145 28.890 24.335 ;
        RECT 29.455 24.145 29.625 24.335 ;
        RECT 31.295 24.145 31.465 24.335 ;
        RECT 33.600 24.165 33.770 24.355 ;
        RECT 36.815 24.165 36.985 24.355 ;
        RECT 39.390 24.145 39.560 24.335 ;
        RECT 39.570 24.195 39.690 24.305 ;
        RECT 40.035 24.165 40.205 24.355 ;
        RECT 43.255 24.145 43.425 24.335 ;
        RECT 43.715 24.165 43.885 24.355 ;
        RECT 12.755 23.335 14.125 24.145 ;
        RECT 14.135 23.465 15.965 24.145 ;
        RECT 17.005 23.465 20.470 24.145 ;
        RECT 21.605 23.465 25.070 24.145 ;
        RECT 25.405 23.465 29.305 24.145 ;
        RECT 14.135 23.235 15.480 23.465 ;
        RECT 19.550 23.235 20.470 23.465 ;
        RECT 24.150 23.235 25.070 23.465 ;
        RECT 28.375 23.235 29.305 23.465 ;
        RECT 29.315 23.335 31.145 24.145 ;
        RECT 31.155 23.465 38.465 24.145 ;
        RECT 34.670 23.245 35.580 23.465 ;
        RECT 37.115 23.235 38.465 23.465 ;
        RECT 38.525 23.275 38.955 24.060 ;
        RECT 38.975 23.465 42.875 24.145 ;
        RECT 38.975 23.235 39.905 23.465 ;
        RECT 43.115 23.365 44.485 24.145 ;
        RECT 44.495 24.115 45.440 24.145 ;
        RECT 46.930 24.115 47.100 24.335 ;
        RECT 48.315 24.145 48.485 24.355 ;
        RECT 44.495 23.435 47.245 24.115 ;
        RECT 44.495 23.235 45.440 23.435 ;
        RECT 47.255 23.335 48.625 24.145 ;
      LAYER nwell ;
        RECT 12.560 20.115 48.820 22.945 ;
      LAYER pwell ;
        RECT 12.755 18.915 14.125 19.725 ;
        RECT 14.175 19.595 15.525 19.825 ;
        RECT 17.060 19.595 17.970 19.815 ;
        RECT 14.175 18.915 21.485 19.595 ;
        RECT 21.495 18.915 25.165 19.725 ;
        RECT 25.645 19.000 26.075 19.785 ;
        RECT 26.095 18.915 35.200 19.595 ;
        RECT 35.295 18.915 36.665 19.725 ;
        RECT 36.675 18.915 38.045 19.695 ;
        RECT 38.055 18.915 39.425 19.695 ;
        RECT 39.435 18.915 40.805 19.695 ;
        RECT 40.815 18.915 42.185 19.695 ;
        RECT 42.215 18.915 43.565 19.825 ;
        RECT 43.655 18.915 47.105 19.825 ;
        RECT 47.255 18.915 48.625 19.725 ;
        RECT 12.895 18.705 13.065 18.915 ;
        RECT 15.655 18.705 15.825 18.895 ;
        RECT 16.125 18.750 16.285 18.860 ;
        RECT 17.310 18.705 17.480 18.895 ;
        RECT 21.175 18.705 21.345 18.915 ;
        RECT 21.635 18.725 21.805 18.915 ;
        RECT 24.855 18.705 25.025 18.895 ;
        RECT 25.310 18.755 25.430 18.865 ;
        RECT 26.235 18.725 26.405 18.915 ;
        RECT 33.135 18.705 33.305 18.895 ;
        RECT 33.870 18.705 34.040 18.895 ;
        RECT 35.435 18.725 35.605 18.915 ;
        RECT 36.815 18.725 36.985 18.915 ;
        RECT 37.745 18.750 37.905 18.860 ;
        RECT 38.195 18.725 38.365 18.915 ;
        RECT 39.575 18.725 39.745 18.915 ;
        RECT 40.955 18.725 41.125 18.915 ;
        RECT 42.335 18.705 42.505 18.895 ;
        RECT 42.805 18.750 42.965 18.860 ;
        RECT 43.250 18.725 43.420 18.915 ;
        RECT 43.715 18.725 43.885 18.915 ;
        RECT 46.015 18.705 46.185 18.895 ;
        RECT 46.485 18.750 46.645 18.860 ;
        RECT 48.315 18.705 48.485 18.915 ;
        RECT 12.755 17.895 14.125 18.705 ;
        RECT 14.135 18.025 15.965 18.705 ;
        RECT 16.895 18.025 20.795 18.705 ;
        RECT 14.135 17.795 15.480 18.025 ;
        RECT 16.895 17.795 17.825 18.025 ;
        RECT 21.035 17.895 24.705 18.705 ;
        RECT 24.715 17.895 26.085 18.705 ;
        RECT 26.135 18.025 33.445 18.705 ;
        RECT 33.455 18.025 37.355 18.705 ;
        RECT 26.135 17.795 27.485 18.025 ;
        RECT 29.020 17.805 29.930 18.025 ;
        RECT 33.455 17.795 34.385 18.025 ;
        RECT 38.525 17.835 38.955 18.620 ;
        RECT 39.070 18.025 42.535 18.705 ;
        RECT 39.070 17.795 39.990 18.025 ;
        RECT 43.575 17.795 46.325 18.705 ;
        RECT 47.255 17.895 48.625 18.705 ;
      LAYER nwell ;
        RECT 12.560 14.675 48.820 17.505 ;
      LAYER pwell ;
        RECT 12.755 13.475 14.125 14.285 ;
        RECT 14.135 13.475 19.645 14.285 ;
        RECT 19.655 13.475 23.325 14.285 ;
        RECT 24.280 14.155 25.625 14.385 ;
        RECT 23.795 13.475 25.625 14.155 ;
        RECT 25.645 13.560 26.075 14.345 ;
        RECT 26.555 14.155 27.900 14.385 ;
        RECT 31.910 14.155 32.820 14.375 ;
        RECT 34.355 14.155 35.705 14.385 ;
        RECT 26.555 13.475 28.385 14.155 ;
        RECT 28.395 13.475 35.705 14.155 ;
        RECT 35.755 14.155 37.100 14.385 ;
        RECT 35.755 13.475 37.585 14.155 ;
        RECT 38.525 13.560 38.955 14.345 ;
        RECT 40.380 14.155 41.725 14.385 ;
        RECT 39.895 13.475 41.725 14.155 ;
        RECT 41.735 13.475 43.105 14.255 ;
        RECT 45.855 14.155 46.785 14.385 ;
        RECT 44.035 13.475 46.785 14.155 ;
        RECT 47.255 13.475 48.625 14.285 ;
        RECT 12.895 13.285 13.065 13.475 ;
        RECT 14.275 13.285 14.445 13.475 ;
        RECT 19.795 13.285 19.965 13.475 ;
        RECT 23.470 13.315 23.590 13.425 ;
        RECT 23.935 13.285 24.105 13.475 ;
        RECT 26.230 13.315 26.350 13.425 ;
        RECT 28.075 13.285 28.245 13.475 ;
        RECT 28.535 13.285 28.705 13.475 ;
        RECT 37.275 13.285 37.445 13.475 ;
        RECT 37.745 13.320 37.905 13.430 ;
        RECT 39.125 13.320 39.285 13.430 ;
        RECT 40.035 13.285 40.205 13.475 ;
        RECT 42.785 13.285 42.955 13.475 ;
        RECT 43.265 13.320 43.425 13.430 ;
        RECT 44.175 13.285 44.345 13.475 ;
        RECT 46.930 13.315 47.050 13.425 ;
        RECT 48.315 13.285 48.485 13.475 ;
      LAYER li1 ;
        RECT 17.430 204.545 143.010 204.715 ;
        RECT 17.515 203.795 18.725 204.545 ;
        RECT 18.895 204.000 24.240 204.545 ;
        RECT 24.415 204.000 29.760 204.545 ;
        RECT 17.515 203.255 18.035 203.795 ;
        RECT 18.205 203.085 18.725 203.625 ;
        RECT 20.480 203.170 20.820 204.000 ;
        RECT 17.515 201.995 18.725 203.085 ;
        RECT 22.300 202.430 22.650 203.680 ;
        RECT 26.000 203.170 26.340 204.000 ;
        RECT 30.395 203.820 30.685 204.545 ;
        RECT 30.855 204.000 36.200 204.545 ;
        RECT 36.375 204.000 41.720 204.545 ;
        RECT 27.820 202.430 28.170 203.680 ;
        RECT 32.440 203.170 32.780 204.000 ;
        RECT 18.895 201.995 24.240 202.430 ;
        RECT 24.415 201.995 29.760 202.430 ;
        RECT 30.395 201.995 30.685 203.160 ;
        RECT 34.260 202.430 34.610 203.680 ;
        RECT 37.960 203.170 38.300 204.000 ;
        RECT 41.895 203.795 43.105 204.545 ;
        RECT 43.275 203.820 43.565 204.545 ;
        RECT 43.735 204.000 49.080 204.545 ;
        RECT 49.255 204.000 54.600 204.545 ;
        RECT 39.780 202.430 40.130 203.680 ;
        RECT 41.895 203.255 42.415 203.795 ;
        RECT 42.585 203.085 43.105 203.625 ;
        RECT 45.320 203.170 45.660 204.000 ;
        RECT 30.855 201.995 36.200 202.430 ;
        RECT 36.375 201.995 41.720 202.430 ;
        RECT 41.895 201.995 43.105 203.085 ;
        RECT 43.275 201.995 43.565 203.160 ;
        RECT 47.140 202.430 47.490 203.680 ;
        RECT 50.840 203.170 51.180 204.000 ;
        RECT 54.775 203.795 55.985 204.545 ;
        RECT 56.155 203.820 56.445 204.545 ;
        RECT 56.615 204.000 61.960 204.545 ;
        RECT 62.135 204.000 67.480 204.545 ;
        RECT 52.660 202.430 53.010 203.680 ;
        RECT 54.775 203.255 55.295 203.795 ;
        RECT 55.465 203.085 55.985 203.625 ;
        RECT 58.200 203.170 58.540 204.000 ;
        RECT 43.735 201.995 49.080 202.430 ;
        RECT 49.255 201.995 54.600 202.430 ;
        RECT 54.775 201.995 55.985 203.085 ;
        RECT 56.155 201.995 56.445 203.160 ;
        RECT 60.020 202.430 60.370 203.680 ;
        RECT 63.720 203.170 64.060 204.000 ;
        RECT 67.655 203.795 68.865 204.545 ;
        RECT 69.035 203.820 69.325 204.545 ;
        RECT 69.495 204.000 74.840 204.545 ;
        RECT 65.540 202.430 65.890 203.680 ;
        RECT 67.655 203.255 68.175 203.795 ;
        RECT 68.345 203.085 68.865 203.625 ;
        RECT 71.080 203.170 71.420 204.000 ;
        RECT 75.015 203.775 76.685 204.545 ;
        RECT 56.615 201.995 61.960 202.430 ;
        RECT 62.135 201.995 67.480 202.430 ;
        RECT 67.655 201.995 68.865 203.085 ;
        RECT 69.035 201.995 69.325 203.160 ;
        RECT 72.900 202.430 73.250 203.680 ;
        RECT 75.015 203.255 75.765 203.775 ;
        RECT 76.860 203.705 77.120 204.545 ;
        RECT 77.295 203.800 77.550 204.375 ;
        RECT 77.720 204.165 78.050 204.545 ;
        RECT 78.265 203.995 78.435 204.375 ;
        RECT 77.720 203.825 78.435 203.995 ;
        RECT 75.935 203.085 76.685 203.605 ;
        RECT 69.495 201.995 74.840 202.430 ;
        RECT 75.015 201.995 76.685 203.085 ;
        RECT 76.860 201.995 77.120 203.145 ;
        RECT 77.295 203.070 77.465 203.800 ;
        RECT 77.720 203.635 77.890 203.825 ;
        RECT 78.695 203.775 81.285 204.545 ;
        RECT 81.915 203.820 82.205 204.545 ;
        RECT 82.375 204.000 87.720 204.545 ;
        RECT 87.895 204.000 93.240 204.545 ;
        RECT 77.635 203.305 77.890 203.635 ;
        RECT 77.720 203.095 77.890 203.305 ;
        RECT 78.170 203.275 78.525 203.645 ;
        RECT 78.695 203.255 79.905 203.775 ;
        RECT 77.295 202.165 77.550 203.070 ;
        RECT 77.720 202.925 78.435 203.095 ;
        RECT 80.075 203.085 81.285 203.605 ;
        RECT 83.960 203.170 84.300 204.000 ;
        RECT 77.720 201.995 78.050 202.755 ;
        RECT 78.265 202.165 78.435 202.925 ;
        RECT 78.695 201.995 81.285 203.085 ;
        RECT 81.915 201.995 82.205 203.160 ;
        RECT 85.780 202.430 86.130 203.680 ;
        RECT 89.480 203.170 89.820 204.000 ;
        RECT 93.415 203.795 94.625 204.545 ;
        RECT 94.795 203.820 95.085 204.545 ;
        RECT 95.255 204.000 100.600 204.545 ;
        RECT 100.775 204.000 106.120 204.545 ;
        RECT 91.300 202.430 91.650 203.680 ;
        RECT 93.415 203.255 93.935 203.795 ;
        RECT 94.105 203.085 94.625 203.625 ;
        RECT 96.840 203.170 97.180 204.000 ;
        RECT 82.375 201.995 87.720 202.430 ;
        RECT 87.895 201.995 93.240 202.430 ;
        RECT 93.415 201.995 94.625 203.085 ;
        RECT 94.795 201.995 95.085 203.160 ;
        RECT 98.660 202.430 99.010 203.680 ;
        RECT 102.360 203.170 102.700 204.000 ;
        RECT 106.295 203.795 107.505 204.545 ;
        RECT 107.675 203.820 107.965 204.545 ;
        RECT 108.135 204.000 113.480 204.545 ;
        RECT 113.655 204.000 119.000 204.545 ;
        RECT 104.180 202.430 104.530 203.680 ;
        RECT 106.295 203.255 106.815 203.795 ;
        RECT 106.985 203.085 107.505 203.625 ;
        RECT 109.720 203.170 110.060 204.000 ;
        RECT 95.255 201.995 100.600 202.430 ;
        RECT 100.775 201.995 106.120 202.430 ;
        RECT 106.295 201.995 107.505 203.085 ;
        RECT 107.675 201.995 107.965 203.160 ;
        RECT 111.540 202.430 111.890 203.680 ;
        RECT 115.240 203.170 115.580 204.000 ;
        RECT 119.175 203.795 120.385 204.545 ;
        RECT 120.555 203.820 120.845 204.545 ;
        RECT 121.015 204.000 126.360 204.545 ;
        RECT 126.535 204.000 131.880 204.545 ;
        RECT 117.060 202.430 117.410 203.680 ;
        RECT 119.175 203.255 119.695 203.795 ;
        RECT 119.865 203.085 120.385 203.625 ;
        RECT 122.600 203.170 122.940 204.000 ;
        RECT 108.135 201.995 113.480 202.430 ;
        RECT 113.655 201.995 119.000 202.430 ;
        RECT 119.175 201.995 120.385 203.085 ;
        RECT 120.555 201.995 120.845 203.160 ;
        RECT 124.420 202.430 124.770 203.680 ;
        RECT 128.120 203.170 128.460 204.000 ;
        RECT 132.055 203.795 133.265 204.545 ;
        RECT 133.435 203.820 133.725 204.545 ;
        RECT 133.895 204.000 139.240 204.545 ;
        RECT 129.940 202.430 130.290 203.680 ;
        RECT 132.055 203.255 132.575 203.795 ;
        RECT 132.745 203.085 133.265 203.625 ;
        RECT 135.480 203.170 135.820 204.000 ;
        RECT 139.415 203.775 141.085 204.545 ;
        RECT 141.715 203.795 142.925 204.545 ;
        RECT 121.015 201.995 126.360 202.430 ;
        RECT 126.535 201.995 131.880 202.430 ;
        RECT 132.055 201.995 133.265 203.085 ;
        RECT 133.435 201.995 133.725 203.160 ;
        RECT 137.300 202.430 137.650 203.680 ;
        RECT 139.415 203.255 140.165 203.775 ;
        RECT 140.335 203.085 141.085 203.605 ;
        RECT 133.895 201.995 139.240 202.430 ;
        RECT 139.415 201.995 141.085 203.085 ;
        RECT 141.715 203.085 142.235 203.625 ;
        RECT 142.405 203.255 142.925 203.795 ;
        RECT 141.715 201.995 142.925 203.085 ;
        RECT 17.430 201.825 143.010 201.995 ;
        RECT 17.515 200.735 18.725 201.825 ;
        RECT 18.895 201.390 24.240 201.825 ;
        RECT 24.415 201.390 29.760 201.825 ;
        RECT 17.515 200.025 18.035 200.565 ;
        RECT 18.205 200.195 18.725 200.735 ;
        RECT 17.515 199.275 18.725 200.025 ;
        RECT 20.480 199.820 20.820 200.650 ;
        RECT 22.300 200.140 22.650 201.390 ;
        RECT 26.000 199.820 26.340 200.650 ;
        RECT 27.820 200.140 28.170 201.390 ;
        RECT 30.395 200.660 30.685 201.825 ;
        RECT 30.855 201.390 36.200 201.825 ;
        RECT 36.375 201.390 41.720 201.825 ;
        RECT 41.895 201.390 47.240 201.825 ;
        RECT 47.415 201.390 52.760 201.825 ;
        RECT 18.895 199.275 24.240 199.820 ;
        RECT 24.415 199.275 29.760 199.820 ;
        RECT 30.395 199.275 30.685 200.000 ;
        RECT 32.440 199.820 32.780 200.650 ;
        RECT 34.260 200.140 34.610 201.390 ;
        RECT 37.960 199.820 38.300 200.650 ;
        RECT 39.780 200.140 40.130 201.390 ;
        RECT 43.480 199.820 43.820 200.650 ;
        RECT 45.300 200.140 45.650 201.390 ;
        RECT 49.000 199.820 49.340 200.650 ;
        RECT 50.820 200.140 51.170 201.390 ;
        RECT 52.935 200.735 55.525 201.825 ;
        RECT 52.935 200.045 54.145 200.565 ;
        RECT 54.315 200.215 55.525 200.735 ;
        RECT 56.155 200.660 56.445 201.825 ;
        RECT 56.615 201.390 61.960 201.825 ;
        RECT 62.135 201.390 67.480 201.825 ;
        RECT 67.655 201.390 73.000 201.825 ;
        RECT 73.175 201.390 78.520 201.825 ;
        RECT 30.855 199.275 36.200 199.820 ;
        RECT 36.375 199.275 41.720 199.820 ;
        RECT 41.895 199.275 47.240 199.820 ;
        RECT 47.415 199.275 52.760 199.820 ;
        RECT 52.935 199.275 55.525 200.045 ;
        RECT 56.155 199.275 56.445 200.000 ;
        RECT 58.200 199.820 58.540 200.650 ;
        RECT 60.020 200.140 60.370 201.390 ;
        RECT 63.720 199.820 64.060 200.650 ;
        RECT 65.540 200.140 65.890 201.390 ;
        RECT 69.240 199.820 69.580 200.650 ;
        RECT 71.060 200.140 71.410 201.390 ;
        RECT 74.760 199.820 75.100 200.650 ;
        RECT 76.580 200.140 76.930 201.390 ;
        RECT 78.695 200.735 81.285 201.825 ;
        RECT 78.695 200.045 79.905 200.565 ;
        RECT 80.075 200.215 81.285 200.735 ;
        RECT 81.915 200.660 82.205 201.825 ;
        RECT 82.375 201.390 87.720 201.825 ;
        RECT 87.895 201.390 93.240 201.825 ;
        RECT 93.415 201.390 98.760 201.825 ;
        RECT 98.935 201.390 104.280 201.825 ;
        RECT 56.615 199.275 61.960 199.820 ;
        RECT 62.135 199.275 67.480 199.820 ;
        RECT 67.655 199.275 73.000 199.820 ;
        RECT 73.175 199.275 78.520 199.820 ;
        RECT 78.695 199.275 81.285 200.045 ;
        RECT 81.915 199.275 82.205 200.000 ;
        RECT 83.960 199.820 84.300 200.650 ;
        RECT 85.780 200.140 86.130 201.390 ;
        RECT 89.480 199.820 89.820 200.650 ;
        RECT 91.300 200.140 91.650 201.390 ;
        RECT 95.000 199.820 95.340 200.650 ;
        RECT 96.820 200.140 97.170 201.390 ;
        RECT 100.520 199.820 100.860 200.650 ;
        RECT 102.340 200.140 102.690 201.390 ;
        RECT 104.455 200.735 107.045 201.825 ;
        RECT 104.455 200.045 105.665 200.565 ;
        RECT 105.835 200.215 107.045 200.735 ;
        RECT 107.675 200.660 107.965 201.825 ;
        RECT 108.135 201.390 113.480 201.825 ;
        RECT 113.655 201.390 119.000 201.825 ;
        RECT 119.175 201.390 124.520 201.825 ;
        RECT 124.695 201.390 130.040 201.825 ;
        RECT 82.375 199.275 87.720 199.820 ;
        RECT 87.895 199.275 93.240 199.820 ;
        RECT 93.415 199.275 98.760 199.820 ;
        RECT 98.935 199.275 104.280 199.820 ;
        RECT 104.455 199.275 107.045 200.045 ;
        RECT 107.675 199.275 107.965 200.000 ;
        RECT 109.720 199.820 110.060 200.650 ;
        RECT 111.540 200.140 111.890 201.390 ;
        RECT 115.240 199.820 115.580 200.650 ;
        RECT 117.060 200.140 117.410 201.390 ;
        RECT 120.760 199.820 121.100 200.650 ;
        RECT 122.580 200.140 122.930 201.390 ;
        RECT 126.280 199.820 126.620 200.650 ;
        RECT 128.100 200.140 128.450 201.390 ;
        RECT 130.215 200.735 132.805 201.825 ;
        RECT 130.215 200.045 131.425 200.565 ;
        RECT 131.595 200.215 132.805 200.735 ;
        RECT 133.435 200.660 133.725 201.825 ;
        RECT 133.895 201.390 139.240 201.825 ;
        RECT 108.135 199.275 113.480 199.820 ;
        RECT 113.655 199.275 119.000 199.820 ;
        RECT 119.175 199.275 124.520 199.820 ;
        RECT 124.695 199.275 130.040 199.820 ;
        RECT 130.215 199.275 132.805 200.045 ;
        RECT 133.435 199.275 133.725 200.000 ;
        RECT 135.480 199.820 135.820 200.650 ;
        RECT 137.300 200.140 137.650 201.390 ;
        RECT 139.415 200.735 141.085 201.825 ;
        RECT 139.415 200.045 140.165 200.565 ;
        RECT 140.335 200.215 141.085 200.735 ;
        RECT 141.715 200.735 142.925 201.825 ;
        RECT 141.715 200.195 142.235 200.735 ;
        RECT 133.895 199.275 139.240 199.820 ;
        RECT 139.415 199.275 141.085 200.045 ;
        RECT 142.405 200.025 142.925 200.565 ;
        RECT 141.715 199.275 142.925 200.025 ;
        RECT 17.430 199.105 143.010 199.275 ;
        RECT 17.515 198.355 18.725 199.105 ;
        RECT 18.895 198.560 24.240 199.105 ;
        RECT 24.415 198.560 29.760 199.105 ;
        RECT 29.935 198.560 35.280 199.105 ;
        RECT 35.455 198.560 40.800 199.105 ;
        RECT 17.515 197.815 18.035 198.355 ;
        RECT 18.205 197.645 18.725 198.185 ;
        RECT 20.480 197.730 20.820 198.560 ;
        RECT 17.515 196.555 18.725 197.645 ;
        RECT 22.300 196.990 22.650 198.240 ;
        RECT 26.000 197.730 26.340 198.560 ;
        RECT 27.820 196.990 28.170 198.240 ;
        RECT 31.520 197.730 31.860 198.560 ;
        RECT 33.340 196.990 33.690 198.240 ;
        RECT 37.040 197.730 37.380 198.560 ;
        RECT 40.975 198.335 42.645 199.105 ;
        RECT 43.275 198.380 43.565 199.105 ;
        RECT 43.735 198.560 49.080 199.105 ;
        RECT 49.255 198.560 54.600 199.105 ;
        RECT 54.775 198.560 60.120 199.105 ;
        RECT 60.295 198.560 65.640 199.105 ;
        RECT 38.860 196.990 39.210 198.240 ;
        RECT 40.975 197.815 41.725 198.335 ;
        RECT 41.895 197.645 42.645 198.165 ;
        RECT 45.320 197.730 45.660 198.560 ;
        RECT 18.895 196.555 24.240 196.990 ;
        RECT 24.415 196.555 29.760 196.990 ;
        RECT 29.935 196.555 35.280 196.990 ;
        RECT 35.455 196.555 40.800 196.990 ;
        RECT 40.975 196.555 42.645 197.645 ;
        RECT 43.275 196.555 43.565 197.720 ;
        RECT 47.140 196.990 47.490 198.240 ;
        RECT 50.840 197.730 51.180 198.560 ;
        RECT 52.660 196.990 53.010 198.240 ;
        RECT 56.360 197.730 56.700 198.560 ;
        RECT 58.180 196.990 58.530 198.240 ;
        RECT 61.880 197.730 62.220 198.560 ;
        RECT 65.815 198.335 68.405 199.105 ;
        RECT 69.035 198.380 69.325 199.105 ;
        RECT 69.495 198.560 74.840 199.105 ;
        RECT 75.015 198.560 80.360 199.105 ;
        RECT 80.535 198.560 85.880 199.105 ;
        RECT 86.055 198.560 91.400 199.105 ;
        RECT 63.700 196.990 64.050 198.240 ;
        RECT 65.815 197.815 67.025 198.335 ;
        RECT 67.195 197.645 68.405 198.165 ;
        RECT 71.080 197.730 71.420 198.560 ;
        RECT 43.735 196.555 49.080 196.990 ;
        RECT 49.255 196.555 54.600 196.990 ;
        RECT 54.775 196.555 60.120 196.990 ;
        RECT 60.295 196.555 65.640 196.990 ;
        RECT 65.815 196.555 68.405 197.645 ;
        RECT 69.035 196.555 69.325 197.720 ;
        RECT 72.900 196.990 73.250 198.240 ;
        RECT 76.600 197.730 76.940 198.560 ;
        RECT 78.420 196.990 78.770 198.240 ;
        RECT 82.120 197.730 82.460 198.560 ;
        RECT 83.940 196.990 84.290 198.240 ;
        RECT 87.640 197.730 87.980 198.560 ;
        RECT 91.575 198.335 94.165 199.105 ;
        RECT 94.795 198.380 95.085 199.105 ;
        RECT 95.255 198.560 100.600 199.105 ;
        RECT 100.775 198.560 106.120 199.105 ;
        RECT 106.295 198.560 111.640 199.105 ;
        RECT 111.815 198.560 117.160 199.105 ;
        RECT 89.460 196.990 89.810 198.240 ;
        RECT 91.575 197.815 92.785 198.335 ;
        RECT 92.955 197.645 94.165 198.165 ;
        RECT 96.840 197.730 97.180 198.560 ;
        RECT 69.495 196.555 74.840 196.990 ;
        RECT 75.015 196.555 80.360 196.990 ;
        RECT 80.535 196.555 85.880 196.990 ;
        RECT 86.055 196.555 91.400 196.990 ;
        RECT 91.575 196.555 94.165 197.645 ;
        RECT 94.795 196.555 95.085 197.720 ;
        RECT 98.660 196.990 99.010 198.240 ;
        RECT 102.360 197.730 102.700 198.560 ;
        RECT 104.180 196.990 104.530 198.240 ;
        RECT 107.880 197.730 108.220 198.560 ;
        RECT 109.700 196.990 110.050 198.240 ;
        RECT 113.400 197.730 113.740 198.560 ;
        RECT 117.335 198.335 119.925 199.105 ;
        RECT 120.555 198.380 120.845 199.105 ;
        RECT 121.015 198.560 126.360 199.105 ;
        RECT 126.535 198.560 131.880 199.105 ;
        RECT 132.055 198.560 137.400 199.105 ;
        RECT 115.220 196.990 115.570 198.240 ;
        RECT 117.335 197.815 118.545 198.335 ;
        RECT 118.715 197.645 119.925 198.165 ;
        RECT 122.600 197.730 122.940 198.560 ;
        RECT 95.255 196.555 100.600 196.990 ;
        RECT 100.775 196.555 106.120 196.990 ;
        RECT 106.295 196.555 111.640 196.990 ;
        RECT 111.815 196.555 117.160 196.990 ;
        RECT 117.335 196.555 119.925 197.645 ;
        RECT 120.555 196.555 120.845 197.720 ;
        RECT 124.420 196.990 124.770 198.240 ;
        RECT 128.120 197.730 128.460 198.560 ;
        RECT 129.940 196.990 130.290 198.240 ;
        RECT 133.640 197.730 133.980 198.560 ;
        RECT 137.575 198.335 141.085 199.105 ;
        RECT 141.715 198.355 142.925 199.105 ;
        RECT 135.460 196.990 135.810 198.240 ;
        RECT 137.575 197.815 139.225 198.335 ;
        RECT 139.395 197.645 141.085 198.165 ;
        RECT 121.015 196.555 126.360 196.990 ;
        RECT 126.535 196.555 131.880 196.990 ;
        RECT 132.055 196.555 137.400 196.990 ;
        RECT 137.575 196.555 141.085 197.645 ;
        RECT 141.715 197.645 142.235 198.185 ;
        RECT 142.405 197.815 142.925 198.355 ;
        RECT 141.715 196.555 142.925 197.645 ;
        RECT 17.430 196.385 143.010 196.555 ;
        RECT 17.515 195.295 18.725 196.385 ;
        RECT 18.895 195.950 24.240 196.385 ;
        RECT 24.415 195.950 29.760 196.385 ;
        RECT 17.515 194.585 18.035 195.125 ;
        RECT 18.205 194.755 18.725 195.295 ;
        RECT 17.515 193.835 18.725 194.585 ;
        RECT 20.480 194.380 20.820 195.210 ;
        RECT 22.300 194.700 22.650 195.950 ;
        RECT 26.000 194.380 26.340 195.210 ;
        RECT 27.820 194.700 28.170 195.950 ;
        RECT 30.395 195.220 30.685 196.385 ;
        RECT 30.855 195.950 36.200 196.385 ;
        RECT 36.375 195.950 41.720 196.385 ;
        RECT 41.895 195.950 47.240 196.385 ;
        RECT 47.415 195.950 52.760 196.385 ;
        RECT 18.895 193.835 24.240 194.380 ;
        RECT 24.415 193.835 29.760 194.380 ;
        RECT 30.395 193.835 30.685 194.560 ;
        RECT 32.440 194.380 32.780 195.210 ;
        RECT 34.260 194.700 34.610 195.950 ;
        RECT 37.960 194.380 38.300 195.210 ;
        RECT 39.780 194.700 40.130 195.950 ;
        RECT 43.480 194.380 43.820 195.210 ;
        RECT 45.300 194.700 45.650 195.950 ;
        RECT 49.000 194.380 49.340 195.210 ;
        RECT 50.820 194.700 51.170 195.950 ;
        RECT 52.935 195.295 55.525 196.385 ;
        RECT 52.935 194.605 54.145 195.125 ;
        RECT 54.315 194.775 55.525 195.295 ;
        RECT 56.155 195.220 56.445 196.385 ;
        RECT 56.615 195.950 61.960 196.385 ;
        RECT 62.135 195.950 67.480 196.385 ;
        RECT 67.655 195.950 73.000 196.385 ;
        RECT 73.175 195.950 78.520 196.385 ;
        RECT 30.855 193.835 36.200 194.380 ;
        RECT 36.375 193.835 41.720 194.380 ;
        RECT 41.895 193.835 47.240 194.380 ;
        RECT 47.415 193.835 52.760 194.380 ;
        RECT 52.935 193.835 55.525 194.605 ;
        RECT 56.155 193.835 56.445 194.560 ;
        RECT 58.200 194.380 58.540 195.210 ;
        RECT 60.020 194.700 60.370 195.950 ;
        RECT 63.720 194.380 64.060 195.210 ;
        RECT 65.540 194.700 65.890 195.950 ;
        RECT 69.240 194.380 69.580 195.210 ;
        RECT 71.060 194.700 71.410 195.950 ;
        RECT 74.760 194.380 75.100 195.210 ;
        RECT 76.580 194.700 76.930 195.950 ;
        RECT 78.695 195.295 81.285 196.385 ;
        RECT 78.695 194.605 79.905 195.125 ;
        RECT 80.075 194.775 81.285 195.295 ;
        RECT 81.915 195.220 82.205 196.385 ;
        RECT 82.375 195.950 87.720 196.385 ;
        RECT 87.895 195.950 93.240 196.385 ;
        RECT 93.415 195.950 98.760 196.385 ;
        RECT 98.935 195.950 104.280 196.385 ;
        RECT 56.615 193.835 61.960 194.380 ;
        RECT 62.135 193.835 67.480 194.380 ;
        RECT 67.655 193.835 73.000 194.380 ;
        RECT 73.175 193.835 78.520 194.380 ;
        RECT 78.695 193.835 81.285 194.605 ;
        RECT 81.915 193.835 82.205 194.560 ;
        RECT 83.960 194.380 84.300 195.210 ;
        RECT 85.780 194.700 86.130 195.950 ;
        RECT 89.480 194.380 89.820 195.210 ;
        RECT 91.300 194.700 91.650 195.950 ;
        RECT 95.000 194.380 95.340 195.210 ;
        RECT 96.820 194.700 97.170 195.950 ;
        RECT 100.520 194.380 100.860 195.210 ;
        RECT 102.340 194.700 102.690 195.950 ;
        RECT 104.455 195.295 107.045 196.385 ;
        RECT 104.455 194.605 105.665 195.125 ;
        RECT 105.835 194.775 107.045 195.295 ;
        RECT 107.675 195.220 107.965 196.385 ;
        RECT 108.135 195.950 113.480 196.385 ;
        RECT 113.655 195.950 119.000 196.385 ;
        RECT 119.175 195.950 124.520 196.385 ;
        RECT 124.695 195.950 130.040 196.385 ;
        RECT 82.375 193.835 87.720 194.380 ;
        RECT 87.895 193.835 93.240 194.380 ;
        RECT 93.415 193.835 98.760 194.380 ;
        RECT 98.935 193.835 104.280 194.380 ;
        RECT 104.455 193.835 107.045 194.605 ;
        RECT 107.675 193.835 107.965 194.560 ;
        RECT 109.720 194.380 110.060 195.210 ;
        RECT 111.540 194.700 111.890 195.950 ;
        RECT 115.240 194.380 115.580 195.210 ;
        RECT 117.060 194.700 117.410 195.950 ;
        RECT 120.760 194.380 121.100 195.210 ;
        RECT 122.580 194.700 122.930 195.950 ;
        RECT 126.280 194.380 126.620 195.210 ;
        RECT 128.100 194.700 128.450 195.950 ;
        RECT 130.215 195.295 132.805 196.385 ;
        RECT 130.215 194.605 131.425 195.125 ;
        RECT 131.595 194.775 132.805 195.295 ;
        RECT 133.435 195.220 133.725 196.385 ;
        RECT 133.895 195.950 139.240 196.385 ;
        RECT 108.135 193.835 113.480 194.380 ;
        RECT 113.655 193.835 119.000 194.380 ;
        RECT 119.175 193.835 124.520 194.380 ;
        RECT 124.695 193.835 130.040 194.380 ;
        RECT 130.215 193.835 132.805 194.605 ;
        RECT 133.435 193.835 133.725 194.560 ;
        RECT 135.480 194.380 135.820 195.210 ;
        RECT 137.300 194.700 137.650 195.950 ;
        RECT 139.415 195.295 141.085 196.385 ;
        RECT 139.415 194.605 140.165 195.125 ;
        RECT 140.335 194.775 141.085 195.295 ;
        RECT 141.715 195.295 142.925 196.385 ;
        RECT 141.715 194.755 142.235 195.295 ;
        RECT 133.895 193.835 139.240 194.380 ;
        RECT 139.415 193.835 141.085 194.605 ;
        RECT 142.405 194.585 142.925 195.125 ;
        RECT 141.715 193.835 142.925 194.585 ;
        RECT 17.430 193.665 143.010 193.835 ;
        RECT 17.515 192.915 18.725 193.665 ;
        RECT 18.895 193.120 24.240 193.665 ;
        RECT 24.415 193.120 29.760 193.665 ;
        RECT 29.935 193.120 35.280 193.665 ;
        RECT 35.455 193.120 40.800 193.665 ;
        RECT 17.515 192.375 18.035 192.915 ;
        RECT 18.205 192.205 18.725 192.745 ;
        RECT 20.480 192.290 20.820 193.120 ;
        RECT 17.515 191.115 18.725 192.205 ;
        RECT 22.300 191.550 22.650 192.800 ;
        RECT 26.000 192.290 26.340 193.120 ;
        RECT 27.820 191.550 28.170 192.800 ;
        RECT 31.520 192.290 31.860 193.120 ;
        RECT 33.340 191.550 33.690 192.800 ;
        RECT 37.040 192.290 37.380 193.120 ;
        RECT 40.975 192.895 42.645 193.665 ;
        RECT 43.275 192.940 43.565 193.665 ;
        RECT 43.735 193.120 49.080 193.665 ;
        RECT 49.255 193.120 54.600 193.665 ;
        RECT 54.775 193.120 60.120 193.665 ;
        RECT 60.295 193.120 65.640 193.665 ;
        RECT 38.860 191.550 39.210 192.800 ;
        RECT 40.975 192.375 41.725 192.895 ;
        RECT 41.895 192.205 42.645 192.725 ;
        RECT 45.320 192.290 45.660 193.120 ;
        RECT 18.895 191.115 24.240 191.550 ;
        RECT 24.415 191.115 29.760 191.550 ;
        RECT 29.935 191.115 35.280 191.550 ;
        RECT 35.455 191.115 40.800 191.550 ;
        RECT 40.975 191.115 42.645 192.205 ;
        RECT 43.275 191.115 43.565 192.280 ;
        RECT 47.140 191.550 47.490 192.800 ;
        RECT 50.840 192.290 51.180 193.120 ;
        RECT 52.660 191.550 53.010 192.800 ;
        RECT 56.360 192.290 56.700 193.120 ;
        RECT 58.180 191.550 58.530 192.800 ;
        RECT 61.880 192.290 62.220 193.120 ;
        RECT 65.815 192.915 67.025 193.665 ;
        RECT 67.195 192.990 67.455 193.495 ;
        RECT 67.635 193.285 67.965 193.665 ;
        RECT 68.145 193.115 68.315 193.495 ;
        RECT 63.700 191.550 64.050 192.800 ;
        RECT 65.815 192.375 66.335 192.915 ;
        RECT 66.505 192.205 67.025 192.745 ;
        RECT 43.735 191.115 49.080 191.550 ;
        RECT 49.255 191.115 54.600 191.550 ;
        RECT 54.775 191.115 60.120 191.550 ;
        RECT 60.295 191.115 65.640 191.550 ;
        RECT 65.815 191.115 67.025 192.205 ;
        RECT 67.195 192.190 67.365 192.990 ;
        RECT 67.650 192.945 68.315 193.115 ;
        RECT 67.650 192.690 67.820 192.945 ;
        RECT 69.035 192.940 69.325 193.665 ;
        RECT 69.555 192.845 69.765 193.665 ;
        RECT 69.935 192.865 70.265 193.495 ;
        RECT 67.535 192.360 67.820 192.690 ;
        RECT 68.055 192.395 68.385 192.765 ;
        RECT 67.650 192.215 67.820 192.360 ;
        RECT 67.195 191.285 67.465 192.190 ;
        RECT 67.650 192.045 68.315 192.215 ;
        RECT 67.635 191.115 67.965 191.875 ;
        RECT 68.145 191.285 68.315 192.045 ;
        RECT 69.035 191.115 69.325 192.280 ;
        RECT 69.935 192.265 70.185 192.865 ;
        RECT 70.435 192.845 70.665 193.665 ;
        RECT 70.965 193.115 71.135 193.405 ;
        RECT 71.305 193.285 71.635 193.665 ;
        RECT 70.965 192.945 71.630 193.115 ;
        RECT 70.355 192.425 70.685 192.675 ;
        RECT 69.555 191.115 69.765 192.255 ;
        RECT 69.935 191.285 70.265 192.265 ;
        RECT 70.435 191.115 70.665 192.255 ;
        RECT 70.880 192.125 71.230 192.775 ;
        RECT 71.400 191.955 71.630 192.945 ;
        RECT 70.965 191.785 71.630 191.955 ;
        RECT 70.965 191.285 71.135 191.785 ;
        RECT 71.305 191.115 71.635 191.615 ;
        RECT 71.805 191.285 71.990 193.405 ;
        RECT 72.245 193.205 72.495 193.665 ;
        RECT 72.665 193.215 73.000 193.385 ;
        RECT 73.195 193.215 73.870 193.385 ;
        RECT 72.665 193.075 72.835 193.215 ;
        RECT 72.160 192.085 72.440 193.035 ;
        RECT 72.610 192.945 72.835 193.075 ;
        RECT 72.610 191.840 72.780 192.945 ;
        RECT 73.005 192.795 73.530 193.015 ;
        RECT 72.950 192.030 73.190 192.625 ;
        RECT 73.360 192.095 73.530 192.795 ;
        RECT 73.700 192.435 73.870 193.215 ;
        RECT 74.190 193.165 74.560 193.665 ;
        RECT 74.740 193.215 75.145 193.385 ;
        RECT 75.315 193.215 76.100 193.385 ;
        RECT 74.740 192.985 74.910 193.215 ;
        RECT 74.080 192.685 74.910 192.985 ;
        RECT 75.295 192.715 75.760 193.045 ;
        RECT 74.080 192.655 74.280 192.685 ;
        RECT 74.400 192.435 74.570 192.505 ;
        RECT 73.700 192.265 74.570 192.435 ;
        RECT 74.060 192.175 74.570 192.265 ;
        RECT 72.610 191.710 72.915 191.840 ;
        RECT 73.360 191.730 73.890 192.095 ;
        RECT 72.230 191.115 72.495 191.575 ;
        RECT 72.665 191.285 72.915 191.710 ;
        RECT 74.060 191.560 74.230 192.175 ;
        RECT 73.125 191.390 74.230 191.560 ;
        RECT 74.400 191.115 74.570 191.915 ;
        RECT 74.740 191.615 74.910 192.685 ;
        RECT 75.080 191.785 75.270 192.505 ;
        RECT 75.440 191.755 75.760 192.715 ;
        RECT 75.930 192.755 76.100 193.215 ;
        RECT 76.375 193.135 76.585 193.665 ;
        RECT 76.845 192.925 77.175 193.450 ;
        RECT 77.345 193.055 77.515 193.665 ;
        RECT 77.685 193.010 78.015 193.445 ;
        RECT 77.685 192.925 78.065 193.010 ;
        RECT 76.975 192.755 77.175 192.925 ;
        RECT 77.840 192.885 78.065 192.925 ;
        RECT 75.930 192.425 76.805 192.755 ;
        RECT 76.975 192.425 77.725 192.755 ;
        RECT 74.740 191.285 74.990 191.615 ;
        RECT 75.930 191.585 76.100 192.425 ;
        RECT 76.975 192.220 77.165 192.425 ;
        RECT 77.895 192.305 78.065 192.885 ;
        RECT 77.850 192.255 78.065 192.305 ;
        RECT 76.270 191.845 77.165 192.220 ;
        RECT 77.675 192.175 78.065 192.255 ;
        RECT 78.235 192.925 78.620 193.495 ;
        RECT 78.790 193.205 79.115 193.665 ;
        RECT 79.635 193.035 79.915 193.495 ;
        RECT 78.235 192.255 78.515 192.925 ;
        RECT 78.790 192.865 79.915 193.035 ;
        RECT 78.790 192.755 79.240 192.865 ;
        RECT 78.685 192.425 79.240 192.755 ;
        RECT 80.105 192.695 80.505 193.495 ;
        RECT 80.905 193.205 81.175 193.665 ;
        RECT 81.345 193.035 81.630 193.495 ;
        RECT 81.975 193.185 82.255 193.665 ;
        RECT 75.215 191.415 76.100 191.585 ;
        RECT 76.280 191.115 76.595 191.615 ;
        RECT 76.825 191.285 77.165 191.845 ;
        RECT 77.335 191.115 77.505 192.125 ;
        RECT 77.675 191.330 78.005 192.175 ;
        RECT 78.235 191.285 78.620 192.255 ;
        RECT 78.790 191.965 79.240 192.425 ;
        RECT 79.410 192.135 80.505 192.695 ;
        RECT 78.790 191.745 79.915 191.965 ;
        RECT 78.790 191.115 79.115 191.575 ;
        RECT 79.635 191.285 79.915 191.745 ;
        RECT 80.105 191.285 80.505 192.135 ;
        RECT 80.675 192.865 81.630 193.035 ;
        RECT 82.425 193.015 82.685 193.405 ;
        RECT 82.860 193.185 83.115 193.665 ;
        RECT 83.285 193.015 83.580 193.405 ;
        RECT 83.760 193.185 84.035 193.665 ;
        RECT 84.205 193.165 84.505 193.495 ;
        RECT 80.675 191.965 80.885 192.865 ;
        RECT 81.930 192.845 83.580 193.015 ;
        RECT 81.055 192.135 81.745 192.695 ;
        RECT 81.930 192.335 82.335 192.845 ;
        RECT 82.505 192.505 83.645 192.675 ;
        RECT 81.930 192.165 82.685 192.335 ;
        RECT 80.675 191.745 81.630 191.965 ;
        RECT 80.905 191.115 81.175 191.575 ;
        RECT 81.345 191.285 81.630 191.745 ;
        RECT 81.970 191.115 82.255 191.985 ;
        RECT 82.425 191.915 82.685 192.165 ;
        RECT 83.475 192.255 83.645 192.505 ;
        RECT 83.815 192.425 84.165 192.995 ;
        RECT 84.335 192.255 84.505 193.165 ;
        RECT 84.675 193.120 90.020 193.665 ;
        RECT 86.260 192.290 86.600 193.120 ;
        RECT 90.195 192.895 93.705 193.665 ;
        RECT 94.795 192.940 95.085 193.665 ;
        RECT 95.255 193.120 100.600 193.665 ;
        RECT 100.775 193.120 106.120 193.665 ;
        RECT 106.295 193.120 111.640 193.665 ;
        RECT 111.815 193.120 117.160 193.665 ;
        RECT 83.475 192.085 84.505 192.255 ;
        RECT 82.425 191.745 83.545 191.915 ;
        RECT 82.425 191.285 82.685 191.745 ;
        RECT 82.860 191.115 83.115 191.575 ;
        RECT 83.285 191.285 83.545 191.745 ;
        RECT 83.715 191.115 84.025 191.915 ;
        RECT 84.195 191.285 84.505 192.085 ;
        RECT 88.080 191.550 88.430 192.800 ;
        RECT 90.195 192.375 91.845 192.895 ;
        RECT 92.015 192.205 93.705 192.725 ;
        RECT 96.840 192.290 97.180 193.120 ;
        RECT 84.675 191.115 90.020 191.550 ;
        RECT 90.195 191.115 93.705 192.205 ;
        RECT 94.795 191.115 95.085 192.280 ;
        RECT 98.660 191.550 99.010 192.800 ;
        RECT 102.360 192.290 102.700 193.120 ;
        RECT 104.180 191.550 104.530 192.800 ;
        RECT 107.880 192.290 108.220 193.120 ;
        RECT 109.700 191.550 110.050 192.800 ;
        RECT 113.400 192.290 113.740 193.120 ;
        RECT 117.340 192.825 117.600 193.665 ;
        RECT 117.775 192.920 118.030 193.495 ;
        RECT 118.200 193.285 118.530 193.665 ;
        RECT 118.745 193.115 118.915 193.495 ;
        RECT 118.200 192.945 118.915 193.115 ;
        RECT 115.220 191.550 115.570 192.800 ;
        RECT 95.255 191.115 100.600 191.550 ;
        RECT 100.775 191.115 106.120 191.550 ;
        RECT 106.295 191.115 111.640 191.550 ;
        RECT 111.815 191.115 117.160 191.550 ;
        RECT 117.340 191.115 117.600 192.265 ;
        RECT 117.775 192.190 117.945 192.920 ;
        RECT 118.200 192.755 118.370 192.945 ;
        RECT 119.175 192.915 120.385 193.665 ;
        RECT 120.555 192.940 120.845 193.665 ;
        RECT 121.015 193.120 126.360 193.665 ;
        RECT 126.535 193.120 131.880 193.665 ;
        RECT 132.055 193.120 137.400 193.665 ;
        RECT 118.115 192.425 118.370 192.755 ;
        RECT 118.200 192.215 118.370 192.425 ;
        RECT 118.650 192.395 119.005 192.765 ;
        RECT 119.175 192.375 119.695 192.915 ;
        RECT 117.775 191.285 118.030 192.190 ;
        RECT 118.200 192.045 118.915 192.215 ;
        RECT 119.865 192.205 120.385 192.745 ;
        RECT 122.600 192.290 122.940 193.120 ;
        RECT 118.200 191.115 118.530 191.875 ;
        RECT 118.745 191.285 118.915 192.045 ;
        RECT 119.175 191.115 120.385 192.205 ;
        RECT 120.555 191.115 120.845 192.280 ;
        RECT 124.420 191.550 124.770 192.800 ;
        RECT 128.120 192.290 128.460 193.120 ;
        RECT 129.940 191.550 130.290 192.800 ;
        RECT 133.640 192.290 133.980 193.120 ;
        RECT 137.575 192.895 141.085 193.665 ;
        RECT 141.715 192.915 142.925 193.665 ;
        RECT 135.460 191.550 135.810 192.800 ;
        RECT 137.575 192.375 139.225 192.895 ;
        RECT 139.395 192.205 141.085 192.725 ;
        RECT 121.015 191.115 126.360 191.550 ;
        RECT 126.535 191.115 131.880 191.550 ;
        RECT 132.055 191.115 137.400 191.550 ;
        RECT 137.575 191.115 141.085 192.205 ;
        RECT 141.715 192.205 142.235 192.745 ;
        RECT 142.405 192.375 142.925 192.915 ;
        RECT 141.715 191.115 142.925 192.205 ;
        RECT 17.430 190.945 143.010 191.115 ;
        RECT 17.515 189.855 18.725 190.945 ;
        RECT 18.895 190.510 24.240 190.945 ;
        RECT 24.415 190.510 29.760 190.945 ;
        RECT 17.515 189.145 18.035 189.685 ;
        RECT 18.205 189.315 18.725 189.855 ;
        RECT 17.515 188.395 18.725 189.145 ;
        RECT 20.480 188.940 20.820 189.770 ;
        RECT 22.300 189.260 22.650 190.510 ;
        RECT 26.000 188.940 26.340 189.770 ;
        RECT 27.820 189.260 28.170 190.510 ;
        RECT 30.395 189.780 30.685 190.945 ;
        RECT 30.855 190.510 36.200 190.945 ;
        RECT 36.375 190.510 41.720 190.945 ;
        RECT 41.895 190.510 47.240 190.945 ;
        RECT 47.415 190.510 52.760 190.945 ;
        RECT 18.895 188.395 24.240 188.940 ;
        RECT 24.415 188.395 29.760 188.940 ;
        RECT 30.395 188.395 30.685 189.120 ;
        RECT 32.440 188.940 32.780 189.770 ;
        RECT 34.260 189.260 34.610 190.510 ;
        RECT 37.960 188.940 38.300 189.770 ;
        RECT 39.780 189.260 40.130 190.510 ;
        RECT 43.480 188.940 43.820 189.770 ;
        RECT 45.300 189.260 45.650 190.510 ;
        RECT 49.000 188.940 49.340 189.770 ;
        RECT 50.820 189.260 51.170 190.510 ;
        RECT 52.935 189.855 55.525 190.945 ;
        RECT 52.935 189.165 54.145 189.685 ;
        RECT 54.315 189.335 55.525 189.855 ;
        RECT 56.155 189.780 56.445 190.945 ;
        RECT 56.615 190.510 61.960 190.945 ;
        RECT 30.855 188.395 36.200 188.940 ;
        RECT 36.375 188.395 41.720 188.940 ;
        RECT 41.895 188.395 47.240 188.940 ;
        RECT 47.415 188.395 52.760 188.940 ;
        RECT 52.935 188.395 55.525 189.165 ;
        RECT 56.155 188.395 56.445 189.120 ;
        RECT 58.200 188.940 58.540 189.770 ;
        RECT 60.020 189.260 60.370 190.510 ;
        RECT 62.135 189.855 64.725 190.945 ;
        RECT 62.135 189.165 63.345 189.685 ;
        RECT 63.515 189.335 64.725 189.855 ;
        RECT 65.355 189.805 65.740 190.775 ;
        RECT 65.910 190.485 66.235 190.945 ;
        RECT 66.755 190.315 67.035 190.775 ;
        RECT 65.910 190.095 67.035 190.315 ;
        RECT 56.615 188.395 61.960 188.940 ;
        RECT 62.135 188.395 64.725 189.165 ;
        RECT 65.355 189.135 65.635 189.805 ;
        RECT 65.910 189.635 66.360 190.095 ;
        RECT 67.225 189.925 67.625 190.775 ;
        RECT 68.025 190.485 68.295 190.945 ;
        RECT 68.465 190.315 68.750 190.775 ;
        RECT 65.805 189.305 66.360 189.635 ;
        RECT 66.530 189.365 67.625 189.925 ;
        RECT 65.910 189.195 66.360 189.305 ;
        RECT 65.355 188.565 65.740 189.135 ;
        RECT 65.910 189.025 67.035 189.195 ;
        RECT 65.910 188.395 66.235 188.855 ;
        RECT 66.755 188.565 67.035 189.025 ;
        RECT 67.225 188.565 67.625 189.365 ;
        RECT 67.795 190.095 68.750 190.315 ;
        RECT 67.795 189.195 68.005 190.095 ;
        RECT 68.175 189.365 68.865 189.925 ;
        RECT 69.965 189.805 70.295 190.945 ;
        RECT 70.825 189.975 71.155 190.760 ;
        RECT 71.335 190.435 71.635 190.945 ;
        RECT 71.805 190.265 72.135 190.775 ;
        RECT 72.305 190.435 72.935 190.945 ;
        RECT 73.515 190.435 73.895 190.605 ;
        RECT 74.065 190.435 74.365 190.945 ;
        RECT 73.725 190.265 73.895 190.435 ;
        RECT 74.645 190.275 74.815 190.775 ;
        RECT 74.985 190.445 75.315 190.945 ;
        RECT 70.475 189.805 71.155 189.975 ;
        RECT 71.335 190.095 73.555 190.265 ;
        RECT 69.955 189.385 70.305 189.635 ;
        RECT 70.475 189.205 70.645 189.805 ;
        RECT 70.815 189.385 71.165 189.635 ;
        RECT 67.795 189.025 68.750 189.195 ;
        RECT 68.025 188.395 68.295 188.855 ;
        RECT 68.465 188.565 68.750 189.025 ;
        RECT 69.965 188.395 70.235 189.205 ;
        RECT 70.405 188.565 70.735 189.205 ;
        RECT 70.905 188.395 71.145 189.205 ;
        RECT 71.335 189.135 71.505 190.095 ;
        RECT 71.675 189.755 73.215 189.925 ;
        RECT 71.675 189.305 71.920 189.755 ;
        RECT 72.180 189.385 72.875 189.585 ;
        RECT 73.045 189.555 73.215 189.755 ;
        RECT 73.385 189.895 73.555 190.095 ;
        RECT 73.725 190.065 74.385 190.265 ;
        RECT 74.645 190.105 75.310 190.275 ;
        RECT 73.385 189.725 74.045 189.895 ;
        RECT 73.045 189.385 73.645 189.555 ;
        RECT 73.875 189.305 74.045 189.725 ;
        RECT 71.335 188.590 71.800 189.135 ;
        RECT 72.305 188.395 72.475 189.215 ;
        RECT 72.645 189.135 73.555 189.215 ;
        RECT 74.215 189.135 74.385 190.065 ;
        RECT 74.560 189.285 74.910 189.935 ;
        RECT 72.645 189.045 73.895 189.135 ;
        RECT 72.645 188.565 72.975 189.045 ;
        RECT 73.385 188.965 73.895 189.045 ;
        RECT 73.145 188.395 73.495 188.785 ;
        RECT 73.665 188.565 73.895 188.965 ;
        RECT 74.065 188.655 74.385 189.135 ;
        RECT 75.080 189.115 75.310 190.105 ;
        RECT 74.645 188.945 75.310 189.115 ;
        RECT 74.645 188.655 74.815 188.945 ;
        RECT 74.985 188.395 75.315 188.775 ;
        RECT 75.485 188.655 75.670 190.775 ;
        RECT 75.910 190.485 76.175 190.945 ;
        RECT 76.345 190.350 76.595 190.775 ;
        RECT 76.805 190.500 77.910 190.670 ;
        RECT 76.290 190.220 76.595 190.350 ;
        RECT 75.840 189.025 76.120 189.975 ;
        RECT 76.290 189.115 76.460 190.220 ;
        RECT 76.630 189.435 76.870 190.030 ;
        RECT 77.040 189.965 77.570 190.330 ;
        RECT 77.040 189.265 77.210 189.965 ;
        RECT 77.740 189.885 77.910 190.500 ;
        RECT 78.080 190.145 78.250 190.945 ;
        RECT 78.420 190.445 78.670 190.775 ;
        RECT 78.895 190.475 79.780 190.645 ;
        RECT 77.740 189.795 78.250 189.885 ;
        RECT 76.290 188.985 76.515 189.115 ;
        RECT 76.685 189.045 77.210 189.265 ;
        RECT 77.380 189.625 78.250 189.795 ;
        RECT 75.925 188.395 76.175 188.855 ;
        RECT 76.345 188.845 76.515 188.985 ;
        RECT 77.380 188.845 77.550 189.625 ;
        RECT 78.080 189.555 78.250 189.625 ;
        RECT 77.760 189.375 77.960 189.405 ;
        RECT 78.420 189.375 78.590 190.445 ;
        RECT 78.760 189.555 78.950 190.275 ;
        RECT 77.760 189.075 78.590 189.375 ;
        RECT 79.120 189.345 79.440 190.305 ;
        RECT 76.345 188.675 76.680 188.845 ;
        RECT 76.875 188.675 77.550 188.845 ;
        RECT 77.870 188.395 78.240 188.895 ;
        RECT 78.420 188.845 78.590 189.075 ;
        RECT 78.975 189.015 79.440 189.345 ;
        RECT 79.610 189.635 79.780 190.475 ;
        RECT 79.960 190.445 80.275 190.945 ;
        RECT 80.505 190.215 80.845 190.775 ;
        RECT 79.950 189.840 80.845 190.215 ;
        RECT 81.015 189.935 81.185 190.945 ;
        RECT 80.655 189.635 80.845 189.840 ;
        RECT 81.355 189.885 81.685 190.730 ;
        RECT 81.355 189.805 81.745 189.885 ;
        RECT 81.530 189.755 81.745 189.805 ;
        RECT 81.915 189.780 82.205 190.945 ;
        RECT 82.560 189.975 82.950 190.150 ;
        RECT 83.435 190.145 83.765 190.945 ;
        RECT 83.935 190.155 84.470 190.775 ;
        RECT 84.675 190.510 90.020 190.945 ;
        RECT 82.560 189.805 83.985 189.975 ;
        RECT 79.610 189.305 80.485 189.635 ;
        RECT 80.655 189.305 81.405 189.635 ;
        RECT 79.610 188.845 79.780 189.305 ;
        RECT 80.655 189.135 80.855 189.305 ;
        RECT 81.575 189.175 81.745 189.755 ;
        RECT 81.520 189.135 81.745 189.175 ;
        RECT 78.420 188.675 78.825 188.845 ;
        RECT 78.995 188.675 79.780 188.845 ;
        RECT 80.055 188.395 80.265 188.925 ;
        RECT 80.525 188.610 80.855 189.135 ;
        RECT 81.365 189.050 81.745 189.135 ;
        RECT 81.025 188.395 81.195 189.005 ;
        RECT 81.365 188.615 81.695 189.050 ;
        RECT 81.915 188.395 82.205 189.120 ;
        RECT 82.435 189.075 82.790 189.635 ;
        RECT 82.960 188.905 83.130 189.805 ;
        RECT 83.300 189.075 83.565 189.635 ;
        RECT 83.815 189.305 83.985 189.805 ;
        RECT 84.155 189.135 84.470 190.155 ;
        RECT 82.540 188.395 82.780 188.905 ;
        RECT 82.960 188.575 83.240 188.905 ;
        RECT 83.470 188.395 83.685 188.905 ;
        RECT 83.855 188.565 84.470 189.135 ;
        RECT 86.260 188.940 86.600 189.770 ;
        RECT 88.080 189.260 88.430 190.510 ;
        RECT 90.195 189.855 92.785 190.945 ;
        RECT 90.195 189.165 91.405 189.685 ;
        RECT 91.575 189.335 92.785 189.855 ;
        RECT 93.425 189.805 93.755 190.945 ;
        RECT 94.285 189.975 94.615 190.760 ;
        RECT 93.935 189.805 94.615 189.975 ;
        RECT 95.775 189.885 96.105 190.730 ;
        RECT 96.275 189.935 96.445 190.945 ;
        RECT 96.615 190.215 96.955 190.775 ;
        RECT 97.185 190.445 97.500 190.945 ;
        RECT 97.680 190.475 98.565 190.645 ;
        RECT 95.715 189.805 96.105 189.885 ;
        RECT 96.615 189.840 97.510 190.215 ;
        RECT 93.415 189.385 93.765 189.635 ;
        RECT 93.935 189.205 94.105 189.805 ;
        RECT 95.715 189.755 95.930 189.805 ;
        RECT 94.275 189.385 94.625 189.635 ;
        RECT 84.675 188.395 90.020 188.940 ;
        RECT 90.195 188.395 92.785 189.165 ;
        RECT 93.425 188.395 93.695 189.205 ;
        RECT 93.865 188.565 94.195 189.205 ;
        RECT 94.365 188.395 94.605 189.205 ;
        RECT 95.715 189.175 95.885 189.755 ;
        RECT 96.615 189.635 96.805 189.840 ;
        RECT 97.680 189.635 97.850 190.475 ;
        RECT 98.790 190.445 99.040 190.775 ;
        RECT 96.055 189.305 96.805 189.635 ;
        RECT 96.975 189.305 97.850 189.635 ;
        RECT 95.715 189.135 95.940 189.175 ;
        RECT 96.605 189.135 96.805 189.305 ;
        RECT 95.715 189.050 96.095 189.135 ;
        RECT 95.765 188.615 96.095 189.050 ;
        RECT 96.265 188.395 96.435 189.005 ;
        RECT 96.605 188.610 96.935 189.135 ;
        RECT 97.195 188.395 97.405 188.925 ;
        RECT 97.680 188.845 97.850 189.305 ;
        RECT 98.020 189.345 98.340 190.305 ;
        RECT 98.510 189.555 98.700 190.275 ;
        RECT 98.870 189.375 99.040 190.445 ;
        RECT 99.210 190.145 99.380 190.945 ;
        RECT 99.550 190.500 100.655 190.670 ;
        RECT 99.550 189.885 99.720 190.500 ;
        RECT 100.865 190.350 101.115 190.775 ;
        RECT 101.285 190.485 101.550 190.945 ;
        RECT 99.890 189.965 100.420 190.330 ;
        RECT 100.865 190.220 101.170 190.350 ;
        RECT 99.210 189.795 99.720 189.885 ;
        RECT 99.210 189.625 100.080 189.795 ;
        RECT 99.210 189.555 99.380 189.625 ;
        RECT 99.500 189.375 99.700 189.405 ;
        RECT 98.020 189.015 98.485 189.345 ;
        RECT 98.870 189.075 99.700 189.375 ;
        RECT 98.870 188.845 99.040 189.075 ;
        RECT 97.680 188.675 98.465 188.845 ;
        RECT 98.635 188.675 99.040 188.845 ;
        RECT 99.220 188.395 99.590 188.895 ;
        RECT 99.910 188.845 100.080 189.625 ;
        RECT 100.250 189.265 100.420 189.965 ;
        RECT 100.590 189.435 100.830 190.030 ;
        RECT 100.250 189.045 100.775 189.265 ;
        RECT 101.000 189.115 101.170 190.220 ;
        RECT 100.945 188.985 101.170 189.115 ;
        RECT 101.340 189.025 101.620 189.975 ;
        RECT 100.945 188.845 101.115 188.985 ;
        RECT 99.910 188.675 100.585 188.845 ;
        RECT 100.780 188.675 101.115 188.845 ;
        RECT 101.285 188.395 101.535 188.855 ;
        RECT 101.790 188.655 101.975 190.775 ;
        RECT 102.145 190.445 102.475 190.945 ;
        RECT 102.645 190.275 102.815 190.775 ;
        RECT 103.125 190.485 103.335 190.945 ;
        RECT 103.825 190.355 104.325 190.775 ;
        RECT 102.150 190.105 102.815 190.275 ;
        RECT 102.150 189.115 102.380 190.105 ;
        RECT 102.550 189.285 102.900 189.935 ;
        RECT 102.150 188.945 102.815 189.115 ;
        RECT 103.075 188.975 103.315 190.300 ;
        RECT 103.485 190.145 104.325 190.355 ;
        RECT 103.485 189.135 103.655 190.145 ;
        RECT 103.825 189.725 104.225 189.975 ;
        RECT 104.515 189.925 104.715 190.715 ;
        RECT 104.395 189.755 104.715 189.925 ;
        RECT 104.885 189.765 105.205 190.945 ;
        RECT 105.380 189.805 105.700 190.945 ;
        RECT 103.825 189.305 103.995 189.725 ;
        RECT 104.395 189.555 104.575 189.755 ;
        RECT 105.880 189.635 106.075 190.685 ;
        RECT 106.255 190.095 106.585 190.775 ;
        RECT 106.785 190.145 107.040 190.945 ;
        RECT 106.255 189.815 106.605 190.095 ;
        RECT 105.440 189.585 105.700 189.635 ;
        RECT 104.210 189.385 104.575 189.555 ;
        RECT 104.745 189.385 105.205 189.585 ;
        RECT 105.435 189.415 105.700 189.585 ;
        RECT 105.440 189.305 105.700 189.415 ;
        RECT 105.880 189.305 106.265 189.635 ;
        RECT 106.435 189.435 106.605 189.815 ;
        RECT 106.795 189.605 107.040 189.965 ;
        RECT 107.675 189.780 107.965 190.945 ;
        RECT 108.135 189.855 111.645 190.945 ;
        RECT 112.795 189.885 113.125 190.730 ;
        RECT 113.295 189.935 113.465 190.945 ;
        RECT 113.635 190.215 113.975 190.775 ;
        RECT 114.205 190.445 114.520 190.945 ;
        RECT 114.700 190.475 115.585 190.645 ;
        RECT 106.435 189.265 106.955 189.435 ;
        RECT 104.175 189.135 105.205 189.175 ;
        RECT 103.485 188.955 103.835 189.135 ;
        RECT 104.005 189.005 105.205 189.135 ;
        RECT 102.145 188.395 102.475 188.775 ;
        RECT 102.645 188.655 102.815 188.945 ;
        RECT 104.005 188.785 104.335 189.005 ;
        RECT 103.075 188.605 104.335 188.785 ;
        RECT 104.525 188.395 104.695 188.835 ;
        RECT 104.865 188.590 105.205 189.005 ;
        RECT 105.380 188.925 106.595 189.095 ;
        RECT 105.380 188.575 105.670 188.925 ;
        RECT 105.865 188.395 106.195 188.755 ;
        RECT 106.365 188.620 106.595 188.925 ;
        RECT 106.785 188.905 106.955 189.265 ;
        RECT 108.135 189.165 109.785 189.685 ;
        RECT 109.955 189.335 111.645 189.855 ;
        RECT 112.735 189.805 113.125 189.885 ;
        RECT 113.635 189.840 114.530 190.215 ;
        RECT 112.735 189.755 112.950 189.805 ;
        RECT 112.735 189.175 112.905 189.755 ;
        RECT 113.635 189.635 113.825 189.840 ;
        RECT 114.700 189.635 114.870 190.475 ;
        RECT 115.810 190.445 116.060 190.775 ;
        RECT 113.075 189.305 113.825 189.635 ;
        RECT 113.995 189.305 114.870 189.635 ;
        RECT 106.785 188.735 106.985 188.905 ;
        RECT 106.785 188.700 106.955 188.735 ;
        RECT 107.675 188.395 107.965 189.120 ;
        RECT 108.135 188.395 111.645 189.165 ;
        RECT 112.735 189.135 112.960 189.175 ;
        RECT 113.625 189.135 113.825 189.305 ;
        RECT 112.735 189.050 113.115 189.135 ;
        RECT 112.785 188.615 113.115 189.050 ;
        RECT 113.285 188.395 113.455 189.005 ;
        RECT 113.625 188.610 113.955 189.135 ;
        RECT 114.215 188.395 114.425 188.925 ;
        RECT 114.700 188.845 114.870 189.305 ;
        RECT 115.040 189.345 115.360 190.305 ;
        RECT 115.530 189.555 115.720 190.275 ;
        RECT 115.890 189.375 116.060 190.445 ;
        RECT 116.230 190.145 116.400 190.945 ;
        RECT 116.570 190.500 117.675 190.670 ;
        RECT 116.570 189.885 116.740 190.500 ;
        RECT 117.885 190.350 118.135 190.775 ;
        RECT 118.305 190.485 118.570 190.945 ;
        RECT 116.910 189.965 117.440 190.330 ;
        RECT 117.885 190.220 118.190 190.350 ;
        RECT 116.230 189.795 116.740 189.885 ;
        RECT 116.230 189.625 117.100 189.795 ;
        RECT 116.230 189.555 116.400 189.625 ;
        RECT 116.520 189.375 116.720 189.405 ;
        RECT 115.040 189.015 115.505 189.345 ;
        RECT 115.890 189.075 116.720 189.375 ;
        RECT 115.890 188.845 116.060 189.075 ;
        RECT 114.700 188.675 115.485 188.845 ;
        RECT 115.655 188.675 116.060 188.845 ;
        RECT 116.240 188.395 116.610 188.895 ;
        RECT 116.930 188.845 117.100 189.625 ;
        RECT 117.270 189.265 117.440 189.965 ;
        RECT 117.610 189.435 117.850 190.030 ;
        RECT 117.270 189.045 117.795 189.265 ;
        RECT 118.020 189.115 118.190 190.220 ;
        RECT 117.965 188.985 118.190 189.115 ;
        RECT 118.360 189.025 118.640 189.975 ;
        RECT 117.965 188.845 118.135 188.985 ;
        RECT 116.930 188.675 117.605 188.845 ;
        RECT 117.800 188.675 118.135 188.845 ;
        RECT 118.305 188.395 118.555 188.855 ;
        RECT 118.810 188.655 118.995 190.775 ;
        RECT 119.165 190.445 119.495 190.945 ;
        RECT 119.665 190.275 119.835 190.775 ;
        RECT 119.170 190.105 119.835 190.275 ;
        RECT 119.170 189.115 119.400 190.105 ;
        RECT 119.570 189.285 119.920 189.935 ;
        RECT 120.155 189.885 120.485 190.730 ;
        RECT 120.655 189.935 120.825 190.945 ;
        RECT 120.995 190.215 121.335 190.775 ;
        RECT 121.565 190.445 121.880 190.945 ;
        RECT 122.060 190.475 122.945 190.645 ;
        RECT 120.095 189.805 120.485 189.885 ;
        RECT 120.995 189.840 121.890 190.215 ;
        RECT 120.095 189.755 120.310 189.805 ;
        RECT 120.095 189.175 120.265 189.755 ;
        RECT 120.995 189.635 121.185 189.840 ;
        RECT 122.060 189.635 122.230 190.475 ;
        RECT 123.170 190.445 123.420 190.775 ;
        RECT 120.435 189.305 121.185 189.635 ;
        RECT 121.355 189.305 122.230 189.635 ;
        RECT 120.095 189.135 120.320 189.175 ;
        RECT 120.985 189.135 121.185 189.305 ;
        RECT 119.170 188.945 119.835 189.115 ;
        RECT 120.095 189.050 120.475 189.135 ;
        RECT 119.165 188.395 119.495 188.775 ;
        RECT 119.665 188.655 119.835 188.945 ;
        RECT 120.145 188.615 120.475 189.050 ;
        RECT 120.645 188.395 120.815 189.005 ;
        RECT 120.985 188.610 121.315 189.135 ;
        RECT 121.575 188.395 121.785 188.925 ;
        RECT 122.060 188.845 122.230 189.305 ;
        RECT 122.400 189.345 122.720 190.305 ;
        RECT 122.890 189.555 123.080 190.275 ;
        RECT 123.250 189.375 123.420 190.445 ;
        RECT 123.590 190.145 123.760 190.945 ;
        RECT 123.930 190.500 125.035 190.670 ;
        RECT 123.930 189.885 124.100 190.500 ;
        RECT 125.245 190.350 125.495 190.775 ;
        RECT 125.665 190.485 125.930 190.945 ;
        RECT 124.270 189.965 124.800 190.330 ;
        RECT 125.245 190.220 125.550 190.350 ;
        RECT 123.590 189.795 124.100 189.885 ;
        RECT 123.590 189.625 124.460 189.795 ;
        RECT 123.590 189.555 123.760 189.625 ;
        RECT 123.880 189.375 124.080 189.405 ;
        RECT 122.400 189.015 122.865 189.345 ;
        RECT 123.250 189.075 124.080 189.375 ;
        RECT 123.250 188.845 123.420 189.075 ;
        RECT 122.060 188.675 122.845 188.845 ;
        RECT 123.015 188.675 123.420 188.845 ;
        RECT 123.600 188.395 123.970 188.895 ;
        RECT 124.290 188.845 124.460 189.625 ;
        RECT 124.630 189.265 124.800 189.965 ;
        RECT 124.970 189.435 125.210 190.030 ;
        RECT 124.630 189.045 125.155 189.265 ;
        RECT 125.380 189.115 125.550 190.220 ;
        RECT 125.325 188.985 125.550 189.115 ;
        RECT 125.720 189.025 126.000 189.975 ;
        RECT 125.325 188.845 125.495 188.985 ;
        RECT 124.290 188.675 124.965 188.845 ;
        RECT 125.160 188.675 125.495 188.845 ;
        RECT 125.665 188.395 125.915 188.855 ;
        RECT 126.170 188.655 126.355 190.775 ;
        RECT 126.525 190.445 126.855 190.945 ;
        RECT 127.025 190.275 127.195 190.775 ;
        RECT 127.455 190.510 132.800 190.945 ;
        RECT 126.530 190.105 127.195 190.275 ;
        RECT 126.530 189.115 126.760 190.105 ;
        RECT 126.930 189.285 127.280 189.935 ;
        RECT 126.530 188.945 127.195 189.115 ;
        RECT 126.525 188.395 126.855 188.775 ;
        RECT 127.025 188.655 127.195 188.945 ;
        RECT 129.040 188.940 129.380 189.770 ;
        RECT 130.860 189.260 131.210 190.510 ;
        RECT 133.435 189.780 133.725 190.945 ;
        RECT 133.895 190.510 139.240 190.945 ;
        RECT 127.455 188.395 132.800 188.940 ;
        RECT 133.435 188.395 133.725 189.120 ;
        RECT 135.480 188.940 135.820 189.770 ;
        RECT 137.300 189.260 137.650 190.510 ;
        RECT 139.415 189.855 141.085 190.945 ;
        RECT 139.415 189.165 140.165 189.685 ;
        RECT 140.335 189.335 141.085 189.855 ;
        RECT 141.715 189.855 142.925 190.945 ;
        RECT 141.715 189.315 142.235 189.855 ;
        RECT 133.895 188.395 139.240 188.940 ;
        RECT 139.415 188.395 141.085 189.165 ;
        RECT 142.405 189.145 142.925 189.685 ;
        RECT 141.715 188.395 142.925 189.145 ;
        RECT 17.430 188.225 143.010 188.395 ;
        RECT 17.515 187.475 18.725 188.225 ;
        RECT 18.895 187.680 24.240 188.225 ;
        RECT 24.415 187.680 29.760 188.225 ;
        RECT 29.935 187.680 35.280 188.225 ;
        RECT 17.515 186.935 18.035 187.475 ;
        RECT 18.205 186.765 18.725 187.305 ;
        RECT 20.480 186.850 20.820 187.680 ;
        RECT 17.515 185.675 18.725 186.765 ;
        RECT 22.300 186.110 22.650 187.360 ;
        RECT 26.000 186.850 26.340 187.680 ;
        RECT 27.820 186.110 28.170 187.360 ;
        RECT 31.520 186.850 31.860 187.680 ;
        RECT 36.460 187.655 36.635 188.055 ;
        RECT 36.805 187.845 37.135 188.225 ;
        RECT 37.380 187.725 37.610 188.055 ;
        RECT 36.460 187.485 37.090 187.655 ;
        RECT 33.340 186.110 33.690 187.360 ;
        RECT 36.920 187.315 37.090 187.485 ;
        RECT 36.375 186.635 36.740 187.315 ;
        RECT 36.920 186.985 37.270 187.315 ;
        RECT 36.920 186.465 37.090 186.985 ;
        RECT 36.460 186.295 37.090 186.465 ;
        RECT 37.440 186.435 37.610 187.725 ;
        RECT 37.810 186.615 38.090 187.890 ;
        RECT 38.315 186.865 38.585 187.890 ;
        RECT 39.045 187.845 39.375 188.225 ;
        RECT 39.545 187.970 39.880 188.015 ;
        RECT 38.275 186.695 38.585 186.865 ;
        RECT 38.315 186.615 38.585 186.695 ;
        RECT 38.775 186.615 39.115 187.645 ;
        RECT 39.545 187.505 39.885 187.970 ;
        RECT 39.285 186.985 39.545 187.315 ;
        RECT 39.285 186.435 39.455 186.985 ;
        RECT 39.715 186.815 39.885 187.505 ;
        RECT 40.055 187.455 42.645 188.225 ;
        RECT 43.275 187.500 43.565 188.225 ;
        RECT 43.735 187.680 49.080 188.225 ;
        RECT 49.255 187.680 54.600 188.225 ;
        RECT 54.780 187.825 55.115 188.225 ;
        RECT 40.055 186.935 41.265 187.455 ;
        RECT 18.895 185.675 24.240 186.110 ;
        RECT 24.415 185.675 29.760 186.110 ;
        RECT 29.935 185.675 35.280 186.110 ;
        RECT 36.460 185.845 36.635 186.295 ;
        RECT 37.440 186.265 39.455 186.435 ;
        RECT 36.805 185.675 37.135 186.115 ;
        RECT 37.440 185.845 37.610 186.265 ;
        RECT 37.845 185.675 38.515 186.085 ;
        RECT 38.730 185.845 38.900 186.265 ;
        RECT 39.100 185.675 39.430 186.085 ;
        RECT 39.625 185.845 39.885 186.815 ;
        RECT 41.435 186.765 42.645 187.285 ;
        RECT 45.320 186.850 45.660 187.680 ;
        RECT 40.055 185.675 42.645 186.765 ;
        RECT 43.275 185.675 43.565 186.840 ;
        RECT 47.140 186.110 47.490 187.360 ;
        RECT 50.840 186.850 51.180 187.680 ;
        RECT 55.285 187.655 55.490 188.055 ;
        RECT 55.700 187.745 55.975 188.225 ;
        RECT 56.185 187.725 56.445 188.055 ;
        RECT 54.805 187.485 55.490 187.655 ;
        RECT 52.660 186.110 53.010 187.360 ;
        RECT 54.805 186.455 55.145 187.485 ;
        RECT 55.315 186.815 55.565 187.315 ;
        RECT 55.745 186.985 56.105 187.565 ;
        RECT 56.275 186.815 56.445 187.725 ;
        RECT 56.615 187.455 58.285 188.225 ;
        RECT 58.965 187.570 59.295 188.005 ;
        RECT 59.465 187.615 59.635 188.225 ;
        RECT 58.915 187.485 59.295 187.570 ;
        RECT 59.805 187.485 60.135 188.010 ;
        RECT 60.395 187.695 60.605 188.225 ;
        RECT 60.880 187.775 61.665 187.945 ;
        RECT 61.835 187.775 62.240 187.945 ;
        RECT 56.615 186.935 57.365 187.455 ;
        RECT 58.915 187.445 59.140 187.485 ;
        RECT 55.315 186.645 56.445 186.815 ;
        RECT 57.535 186.765 58.285 187.285 ;
        RECT 54.805 186.280 55.470 186.455 ;
        RECT 43.735 185.675 49.080 186.110 ;
        RECT 49.255 185.675 54.600 186.110 ;
        RECT 54.780 185.675 55.115 186.100 ;
        RECT 55.285 185.875 55.470 186.280 ;
        RECT 55.675 185.675 56.005 186.455 ;
        RECT 56.175 185.875 56.445 186.645 ;
        RECT 56.615 185.675 58.285 186.765 ;
        RECT 58.915 186.865 59.085 187.445 ;
        RECT 59.805 187.315 60.005 187.485 ;
        RECT 60.880 187.315 61.050 187.775 ;
        RECT 59.255 186.985 60.005 187.315 ;
        RECT 60.175 186.985 61.050 187.315 ;
        RECT 58.915 186.815 59.130 186.865 ;
        RECT 58.915 186.735 59.305 186.815 ;
        RECT 58.975 185.890 59.305 186.735 ;
        RECT 59.815 186.780 60.005 186.985 ;
        RECT 59.475 185.675 59.645 186.685 ;
        RECT 59.815 186.405 60.710 186.780 ;
        RECT 59.815 185.845 60.155 186.405 ;
        RECT 60.385 185.675 60.700 186.175 ;
        RECT 60.880 186.145 61.050 186.985 ;
        RECT 61.220 187.275 61.685 187.605 ;
        RECT 62.070 187.545 62.240 187.775 ;
        RECT 62.420 187.725 62.790 188.225 ;
        RECT 63.110 187.775 63.785 187.945 ;
        RECT 63.980 187.775 64.315 187.945 ;
        RECT 61.220 186.315 61.540 187.275 ;
        RECT 62.070 187.245 62.900 187.545 ;
        RECT 61.710 186.345 61.900 187.065 ;
        RECT 62.070 186.175 62.240 187.245 ;
        RECT 62.700 187.215 62.900 187.245 ;
        RECT 62.410 186.995 62.580 187.065 ;
        RECT 63.110 186.995 63.280 187.775 ;
        RECT 64.145 187.635 64.315 187.775 ;
        RECT 64.485 187.765 64.735 188.225 ;
        RECT 62.410 186.825 63.280 186.995 ;
        RECT 63.450 187.355 63.975 187.575 ;
        RECT 64.145 187.505 64.370 187.635 ;
        RECT 62.410 186.735 62.920 186.825 ;
        RECT 60.880 185.975 61.765 186.145 ;
        RECT 61.990 185.845 62.240 186.175 ;
        RECT 62.410 185.675 62.580 186.475 ;
        RECT 62.750 186.120 62.920 186.735 ;
        RECT 63.450 186.655 63.620 187.355 ;
        RECT 63.090 186.290 63.620 186.655 ;
        RECT 63.790 186.590 64.030 187.185 ;
        RECT 64.200 186.400 64.370 187.505 ;
        RECT 64.540 186.645 64.820 187.595 ;
        RECT 64.065 186.270 64.370 186.400 ;
        RECT 62.750 185.950 63.855 186.120 ;
        RECT 64.065 185.845 64.315 186.270 ;
        RECT 64.485 185.675 64.750 186.135 ;
        RECT 64.990 185.845 65.175 187.965 ;
        RECT 65.345 187.845 65.675 188.225 ;
        RECT 65.845 187.675 66.015 187.965 ;
        RECT 65.350 187.505 66.015 187.675 ;
        RECT 66.285 187.695 66.615 188.055 ;
        RECT 66.785 187.865 67.115 188.225 ;
        RECT 67.315 187.695 67.645 188.055 ;
        RECT 65.350 186.515 65.580 187.505 ;
        RECT 66.285 187.485 67.645 187.695 ;
        RECT 68.155 187.465 68.865 188.055 ;
        RECT 69.035 187.500 69.325 188.225 ;
        RECT 69.585 187.675 69.755 187.965 ;
        RECT 69.925 187.845 70.255 188.225 ;
        RECT 69.585 187.505 70.250 187.675 ;
        RECT 65.750 186.685 66.100 187.335 ;
        RECT 66.275 186.985 66.585 187.315 ;
        RECT 66.795 186.985 67.170 187.315 ;
        RECT 67.490 186.985 67.985 187.315 ;
        RECT 65.350 186.345 66.015 186.515 ;
        RECT 65.345 185.675 65.675 186.175 ;
        RECT 65.845 185.845 66.015 186.345 ;
        RECT 66.285 185.675 66.615 186.735 ;
        RECT 66.795 186.060 66.965 186.985 ;
        RECT 67.135 186.495 67.465 186.715 ;
        RECT 67.660 186.695 67.985 186.985 ;
        RECT 68.160 186.695 68.490 187.235 ;
        RECT 68.660 186.495 68.865 187.465 ;
        RECT 67.135 186.265 68.865 186.495 ;
        RECT 67.135 185.865 67.465 186.265 ;
        RECT 67.635 185.675 67.965 186.035 ;
        RECT 68.165 185.845 68.865 186.265 ;
        RECT 69.035 185.675 69.325 186.840 ;
        RECT 69.500 186.685 69.850 187.335 ;
        RECT 70.020 186.515 70.250 187.505 ;
        RECT 69.585 186.345 70.250 186.515 ;
        RECT 69.585 185.845 69.755 186.345 ;
        RECT 69.925 185.675 70.255 186.175 ;
        RECT 70.425 185.845 70.610 187.965 ;
        RECT 70.865 187.765 71.115 188.225 ;
        RECT 71.285 187.775 71.620 187.945 ;
        RECT 71.815 187.775 72.490 187.945 ;
        RECT 71.285 187.635 71.455 187.775 ;
        RECT 70.780 186.645 71.060 187.595 ;
        RECT 71.230 187.505 71.455 187.635 ;
        RECT 71.230 186.400 71.400 187.505 ;
        RECT 71.625 187.355 72.150 187.575 ;
        RECT 71.570 186.590 71.810 187.185 ;
        RECT 71.980 186.655 72.150 187.355 ;
        RECT 72.320 186.995 72.490 187.775 ;
        RECT 72.810 187.725 73.180 188.225 ;
        RECT 73.360 187.775 73.765 187.945 ;
        RECT 73.935 187.775 74.720 187.945 ;
        RECT 73.360 187.545 73.530 187.775 ;
        RECT 72.700 187.245 73.530 187.545 ;
        RECT 73.915 187.275 74.380 187.605 ;
        RECT 72.700 187.215 72.900 187.245 ;
        RECT 73.020 186.995 73.190 187.065 ;
        RECT 72.320 186.825 73.190 186.995 ;
        RECT 72.680 186.735 73.190 186.825 ;
        RECT 71.230 186.270 71.535 186.400 ;
        RECT 71.980 186.290 72.510 186.655 ;
        RECT 70.850 185.675 71.115 186.135 ;
        RECT 71.285 185.845 71.535 186.270 ;
        RECT 72.680 186.120 72.850 186.735 ;
        RECT 71.745 185.950 72.850 186.120 ;
        RECT 73.020 185.675 73.190 186.475 ;
        RECT 73.360 186.175 73.530 187.245 ;
        RECT 73.700 186.345 73.890 187.065 ;
        RECT 74.060 186.315 74.380 187.275 ;
        RECT 74.550 187.315 74.720 187.775 ;
        RECT 74.995 187.695 75.205 188.225 ;
        RECT 75.465 187.485 75.795 188.010 ;
        RECT 75.965 187.615 76.135 188.225 ;
        RECT 76.305 187.570 76.635 188.005 ;
        RECT 76.305 187.485 76.685 187.570 ;
        RECT 75.595 187.315 75.795 187.485 ;
        RECT 76.460 187.445 76.685 187.485 ;
        RECT 74.550 186.985 75.425 187.315 ;
        RECT 75.595 186.985 76.345 187.315 ;
        RECT 73.360 185.845 73.610 186.175 ;
        RECT 74.550 186.145 74.720 186.985 ;
        RECT 75.595 186.780 75.785 186.985 ;
        RECT 76.515 186.865 76.685 187.445 ;
        RECT 76.470 186.815 76.685 186.865 ;
        RECT 74.890 186.405 75.785 186.780 ;
        RECT 76.295 186.735 76.685 186.815 ;
        RECT 76.855 187.500 77.115 188.055 ;
        RECT 77.285 187.780 77.715 188.225 ;
        RECT 77.950 187.655 78.120 188.055 ;
        RECT 78.290 187.825 79.010 188.225 ;
        RECT 76.855 186.785 77.030 187.500 ;
        RECT 77.950 187.485 78.830 187.655 ;
        RECT 79.180 187.610 79.350 188.055 ;
        RECT 79.925 187.715 80.325 188.225 ;
        RECT 77.200 186.985 77.455 187.315 ;
        RECT 73.835 185.975 74.720 186.145 ;
        RECT 74.900 185.675 75.215 186.175 ;
        RECT 75.445 185.845 75.785 186.405 ;
        RECT 75.955 185.675 76.125 186.685 ;
        RECT 76.295 185.890 76.625 186.735 ;
        RECT 76.855 185.845 77.115 186.785 ;
        RECT 77.285 186.505 77.455 186.985 ;
        RECT 77.680 186.695 78.010 187.315 ;
        RECT 78.180 186.935 78.470 187.315 ;
        RECT 78.660 186.765 78.830 187.485 ;
        RECT 78.310 186.595 78.830 186.765 ;
        RECT 79.000 187.440 79.350 187.610 ;
        RECT 77.285 186.335 78.045 186.505 ;
        RECT 78.310 186.405 78.480 186.595 ;
        RECT 79.000 186.415 79.170 187.440 ;
        RECT 79.590 186.955 79.850 187.545 ;
        RECT 79.370 186.655 79.850 186.955 ;
        RECT 80.050 186.655 80.310 187.545 ;
        RECT 80.535 187.485 80.920 188.055 ;
        RECT 81.090 187.765 81.415 188.225 ;
        RECT 81.935 187.595 82.215 188.055 ;
        RECT 80.535 186.815 80.815 187.485 ;
        RECT 81.090 187.425 82.215 187.595 ;
        RECT 81.090 187.315 81.540 187.425 ;
        RECT 80.985 186.985 81.540 187.315 ;
        RECT 82.405 187.255 82.805 188.055 ;
        RECT 83.205 187.765 83.475 188.225 ;
        RECT 83.645 187.595 83.930 188.055 ;
        RECT 77.875 186.110 78.045 186.335 ;
        RECT 78.760 186.245 79.170 186.415 ;
        RECT 79.345 186.305 80.285 186.475 ;
        RECT 78.760 186.110 79.015 186.245 ;
        RECT 77.285 185.675 77.615 186.075 ;
        RECT 77.875 185.940 79.015 186.110 ;
        RECT 79.345 186.055 79.515 186.305 ;
        RECT 78.760 185.845 79.015 185.940 ;
        RECT 79.185 185.885 79.515 186.055 ;
        RECT 79.685 185.675 79.935 186.135 ;
        RECT 80.105 185.845 80.285 186.305 ;
        RECT 80.535 185.845 80.920 186.815 ;
        RECT 81.090 186.525 81.540 186.985 ;
        RECT 81.710 186.695 82.805 187.255 ;
        RECT 81.090 186.305 82.215 186.525 ;
        RECT 81.090 185.675 81.415 186.135 ;
        RECT 81.935 185.845 82.215 186.305 ;
        RECT 82.405 185.845 82.805 186.695 ;
        RECT 82.975 187.425 83.930 187.595 ;
        RECT 82.975 186.525 83.185 187.425 ;
        RECT 84.685 187.415 84.955 188.225 ;
        RECT 85.125 187.415 85.455 188.055 ;
        RECT 85.625 187.415 85.865 188.225 ;
        RECT 86.055 187.455 89.565 188.225 ;
        RECT 90.195 187.485 90.580 188.055 ;
        RECT 90.750 187.765 91.075 188.225 ;
        RECT 91.595 187.595 91.875 188.055 ;
        RECT 83.355 186.695 84.045 187.255 ;
        RECT 84.675 186.985 85.025 187.235 ;
        RECT 85.195 186.815 85.365 187.415 ;
        RECT 85.535 186.985 85.885 187.235 ;
        RECT 86.055 186.935 87.705 187.455 ;
        RECT 82.975 186.305 83.930 186.525 ;
        RECT 83.205 185.675 83.475 186.135 ;
        RECT 83.645 185.845 83.930 186.305 ;
        RECT 84.685 185.675 85.015 186.815 ;
        RECT 85.195 186.645 85.875 186.815 ;
        RECT 87.875 186.765 89.565 187.285 ;
        RECT 85.545 185.860 85.875 186.645 ;
        RECT 86.055 185.675 89.565 186.765 ;
        RECT 90.195 186.815 90.475 187.485 ;
        RECT 90.750 187.425 91.875 187.595 ;
        RECT 90.750 187.315 91.200 187.425 ;
        RECT 90.645 186.985 91.200 187.315 ;
        RECT 92.065 187.255 92.465 188.055 ;
        RECT 92.865 187.765 93.135 188.225 ;
        RECT 93.305 187.595 93.590 188.055 ;
        RECT 90.195 185.845 90.580 186.815 ;
        RECT 90.750 186.525 91.200 186.985 ;
        RECT 91.370 186.695 92.465 187.255 ;
        RECT 90.750 186.305 91.875 186.525 ;
        RECT 90.750 185.675 91.075 186.135 ;
        RECT 91.595 185.845 91.875 186.305 ;
        RECT 92.065 185.845 92.465 186.695 ;
        RECT 92.635 187.425 93.590 187.595 ;
        RECT 94.795 187.500 95.085 188.225 ;
        RECT 95.305 187.570 95.635 188.005 ;
        RECT 95.805 187.615 95.975 188.225 ;
        RECT 95.255 187.485 95.635 187.570 ;
        RECT 96.145 187.485 96.475 188.010 ;
        RECT 96.735 187.695 96.945 188.225 ;
        RECT 97.220 187.775 98.005 187.945 ;
        RECT 98.175 187.775 98.580 187.945 ;
        RECT 95.255 187.445 95.480 187.485 ;
        RECT 92.635 186.525 92.845 187.425 ;
        RECT 93.015 186.695 93.705 187.255 ;
        RECT 95.255 186.865 95.425 187.445 ;
        RECT 96.145 187.315 96.345 187.485 ;
        RECT 97.220 187.315 97.390 187.775 ;
        RECT 95.595 186.985 96.345 187.315 ;
        RECT 96.515 186.985 97.390 187.315 ;
        RECT 92.635 186.305 93.590 186.525 ;
        RECT 92.865 185.675 93.135 186.135 ;
        RECT 93.305 185.845 93.590 186.305 ;
        RECT 94.795 185.675 95.085 186.840 ;
        RECT 95.255 186.815 95.470 186.865 ;
        RECT 95.255 186.735 95.645 186.815 ;
        RECT 95.315 185.890 95.645 186.735 ;
        RECT 96.155 186.780 96.345 186.985 ;
        RECT 95.815 185.675 95.985 186.685 ;
        RECT 96.155 186.405 97.050 186.780 ;
        RECT 96.155 185.845 96.495 186.405 ;
        RECT 96.725 185.675 97.040 186.175 ;
        RECT 97.220 186.145 97.390 186.985 ;
        RECT 97.560 187.275 98.025 187.605 ;
        RECT 98.410 187.545 98.580 187.775 ;
        RECT 98.760 187.725 99.130 188.225 ;
        RECT 99.450 187.775 100.125 187.945 ;
        RECT 100.320 187.775 100.655 187.945 ;
        RECT 97.560 186.315 97.880 187.275 ;
        RECT 98.410 187.245 99.240 187.545 ;
        RECT 98.050 186.345 98.240 187.065 ;
        RECT 98.410 186.175 98.580 187.245 ;
        RECT 99.040 187.215 99.240 187.245 ;
        RECT 98.750 186.995 98.920 187.065 ;
        RECT 99.450 186.995 99.620 187.775 ;
        RECT 100.485 187.635 100.655 187.775 ;
        RECT 100.825 187.765 101.075 188.225 ;
        RECT 98.750 186.825 99.620 186.995 ;
        RECT 99.790 187.355 100.315 187.575 ;
        RECT 100.485 187.505 100.710 187.635 ;
        RECT 98.750 186.735 99.260 186.825 ;
        RECT 97.220 185.975 98.105 186.145 ;
        RECT 98.330 185.845 98.580 186.175 ;
        RECT 98.750 185.675 98.920 186.475 ;
        RECT 99.090 186.120 99.260 186.735 ;
        RECT 99.790 186.655 99.960 187.355 ;
        RECT 99.430 186.290 99.960 186.655 ;
        RECT 100.130 186.590 100.370 187.185 ;
        RECT 100.540 186.400 100.710 187.505 ;
        RECT 100.880 186.645 101.160 187.595 ;
        RECT 100.405 186.270 100.710 186.400 ;
        RECT 99.090 185.950 100.195 186.120 ;
        RECT 100.405 185.845 100.655 186.270 ;
        RECT 100.825 185.675 101.090 186.135 ;
        RECT 101.330 185.845 101.515 187.965 ;
        RECT 101.685 187.845 102.015 188.225 ;
        RECT 102.185 187.675 102.355 187.965 ;
        RECT 101.690 187.505 102.355 187.675 ;
        RECT 102.730 187.595 103.015 188.055 ;
        RECT 103.185 187.765 103.455 188.225 ;
        RECT 101.690 186.515 101.920 187.505 ;
        RECT 102.730 187.425 103.685 187.595 ;
        RECT 102.090 186.685 102.440 187.335 ;
        RECT 102.615 186.695 103.305 187.255 ;
        RECT 103.475 186.525 103.685 187.425 ;
        RECT 101.690 186.345 102.355 186.515 ;
        RECT 101.685 185.675 102.015 186.175 ;
        RECT 102.185 185.845 102.355 186.345 ;
        RECT 102.730 186.305 103.685 186.525 ;
        RECT 103.855 187.255 104.255 188.055 ;
        RECT 104.445 187.595 104.725 188.055 ;
        RECT 105.245 187.765 105.570 188.225 ;
        RECT 104.445 187.425 105.570 187.595 ;
        RECT 105.740 187.485 106.125 188.055 ;
        RECT 107.305 187.675 107.475 187.965 ;
        RECT 107.645 187.845 107.975 188.225 ;
        RECT 107.305 187.505 107.970 187.675 ;
        RECT 105.120 187.315 105.570 187.425 ;
        RECT 103.855 186.695 104.950 187.255 ;
        RECT 105.120 186.985 105.675 187.315 ;
        RECT 102.730 185.845 103.015 186.305 ;
        RECT 103.185 185.675 103.455 186.135 ;
        RECT 103.855 185.845 104.255 186.695 ;
        RECT 105.120 186.525 105.570 186.985 ;
        RECT 105.845 186.815 106.125 187.485 ;
        RECT 104.445 186.305 105.570 186.525 ;
        RECT 104.445 185.845 104.725 186.305 ;
        RECT 105.245 185.675 105.570 186.135 ;
        RECT 105.740 185.845 106.125 186.815 ;
        RECT 107.220 186.685 107.570 187.335 ;
        RECT 107.740 186.515 107.970 187.505 ;
        RECT 107.305 186.345 107.970 186.515 ;
        RECT 107.305 185.845 107.475 186.345 ;
        RECT 107.645 185.675 107.975 186.175 ;
        RECT 108.145 185.845 108.330 187.965 ;
        RECT 108.585 187.765 108.835 188.225 ;
        RECT 109.005 187.775 109.340 187.945 ;
        RECT 109.535 187.775 110.210 187.945 ;
        RECT 109.005 187.635 109.175 187.775 ;
        RECT 108.500 186.645 108.780 187.595 ;
        RECT 108.950 187.505 109.175 187.635 ;
        RECT 108.950 186.400 109.120 187.505 ;
        RECT 109.345 187.355 109.870 187.575 ;
        RECT 109.290 186.590 109.530 187.185 ;
        RECT 109.700 186.655 109.870 187.355 ;
        RECT 110.040 186.995 110.210 187.775 ;
        RECT 110.530 187.725 110.900 188.225 ;
        RECT 111.080 187.775 111.485 187.945 ;
        RECT 111.655 187.775 112.440 187.945 ;
        RECT 111.080 187.545 111.250 187.775 ;
        RECT 110.420 187.245 111.250 187.545 ;
        RECT 111.635 187.275 112.100 187.605 ;
        RECT 110.420 187.215 110.620 187.245 ;
        RECT 110.740 186.995 110.910 187.065 ;
        RECT 110.040 186.825 110.910 186.995 ;
        RECT 110.400 186.735 110.910 186.825 ;
        RECT 108.950 186.270 109.255 186.400 ;
        RECT 109.700 186.290 110.230 186.655 ;
        RECT 108.570 185.675 108.835 186.135 ;
        RECT 109.005 185.845 109.255 186.270 ;
        RECT 110.400 186.120 110.570 186.735 ;
        RECT 109.465 185.950 110.570 186.120 ;
        RECT 110.740 185.675 110.910 186.475 ;
        RECT 111.080 186.175 111.250 187.245 ;
        RECT 111.420 186.345 111.610 187.065 ;
        RECT 111.780 186.315 112.100 187.275 ;
        RECT 112.270 187.315 112.440 187.775 ;
        RECT 112.715 187.695 112.925 188.225 ;
        RECT 113.185 187.485 113.515 188.010 ;
        RECT 113.685 187.615 113.855 188.225 ;
        RECT 114.025 187.570 114.355 188.005 ;
        RECT 114.025 187.485 114.405 187.570 ;
        RECT 113.315 187.315 113.515 187.485 ;
        RECT 114.180 187.445 114.405 187.485 ;
        RECT 112.270 186.985 113.145 187.315 ;
        RECT 113.315 186.985 114.065 187.315 ;
        RECT 111.080 185.845 111.330 186.175 ;
        RECT 112.270 186.145 112.440 186.985 ;
        RECT 113.315 186.780 113.505 186.985 ;
        RECT 114.235 186.865 114.405 187.445 ;
        RECT 115.310 187.415 115.555 188.020 ;
        RECT 115.775 187.690 116.285 188.225 ;
        RECT 114.190 186.815 114.405 186.865 ;
        RECT 112.610 186.405 113.505 186.780 ;
        RECT 114.015 186.735 114.405 186.815 ;
        RECT 115.035 187.245 116.265 187.415 ;
        RECT 111.555 185.975 112.440 186.145 ;
        RECT 112.620 185.675 112.935 186.175 ;
        RECT 113.165 185.845 113.505 186.405 ;
        RECT 113.675 185.675 113.845 186.685 ;
        RECT 114.015 185.890 114.345 186.735 ;
        RECT 115.035 186.435 115.375 187.245 ;
        RECT 115.545 186.680 116.295 186.870 ;
        RECT 115.035 186.025 115.550 186.435 ;
        RECT 115.785 185.675 115.955 186.435 ;
        RECT 116.125 186.015 116.295 186.680 ;
        RECT 116.465 186.695 116.655 188.055 ;
        RECT 116.825 187.205 117.100 188.055 ;
        RECT 117.290 187.690 117.820 188.055 ;
        RECT 118.245 187.825 118.575 188.225 ;
        RECT 117.645 187.655 117.820 187.690 ;
        RECT 116.825 187.035 117.105 187.205 ;
        RECT 116.825 186.895 117.100 187.035 ;
        RECT 117.305 186.695 117.475 187.495 ;
        RECT 116.465 186.525 117.475 186.695 ;
        RECT 117.645 187.485 118.575 187.655 ;
        RECT 118.745 187.485 119.000 188.055 ;
        RECT 117.645 186.355 117.815 187.485 ;
        RECT 118.405 187.315 118.575 187.485 ;
        RECT 116.690 186.185 117.815 186.355 ;
        RECT 117.985 186.985 118.180 187.315 ;
        RECT 118.405 186.985 118.660 187.315 ;
        RECT 117.985 186.015 118.155 186.985 ;
        RECT 118.830 186.815 119.000 187.485 ;
        RECT 119.175 187.475 120.385 188.225 ;
        RECT 120.555 187.500 120.845 188.225 ;
        RECT 121.015 187.680 126.360 188.225 ;
        RECT 126.535 187.680 131.880 188.225 ;
        RECT 132.055 187.680 137.400 188.225 ;
        RECT 119.175 186.935 119.695 187.475 ;
        RECT 116.125 185.845 118.155 186.015 ;
        RECT 118.325 185.675 118.495 186.815 ;
        RECT 118.665 185.845 119.000 186.815 ;
        RECT 119.865 186.765 120.385 187.305 ;
        RECT 122.600 186.850 122.940 187.680 ;
        RECT 119.175 185.675 120.385 186.765 ;
        RECT 120.555 185.675 120.845 186.840 ;
        RECT 124.420 186.110 124.770 187.360 ;
        RECT 128.120 186.850 128.460 187.680 ;
        RECT 129.940 186.110 130.290 187.360 ;
        RECT 133.640 186.850 133.980 187.680 ;
        RECT 137.575 187.455 141.085 188.225 ;
        RECT 141.715 187.475 142.925 188.225 ;
        RECT 135.460 186.110 135.810 187.360 ;
        RECT 137.575 186.935 139.225 187.455 ;
        RECT 139.395 186.765 141.085 187.285 ;
        RECT 121.015 185.675 126.360 186.110 ;
        RECT 126.535 185.675 131.880 186.110 ;
        RECT 132.055 185.675 137.400 186.110 ;
        RECT 137.575 185.675 141.085 186.765 ;
        RECT 141.715 186.765 142.235 187.305 ;
        RECT 142.405 186.935 142.925 187.475 ;
        RECT 141.715 185.675 142.925 186.765 ;
        RECT 17.430 185.505 143.010 185.675 ;
        RECT 17.515 184.415 18.725 185.505 ;
        RECT 18.895 184.415 22.405 185.505 ;
        RECT 23.125 184.835 23.295 185.335 ;
        RECT 23.465 185.005 23.795 185.505 ;
        RECT 23.125 184.665 23.790 184.835 ;
        RECT 17.515 183.705 18.035 184.245 ;
        RECT 18.205 183.875 18.725 184.415 ;
        RECT 18.895 183.725 20.545 184.245 ;
        RECT 20.715 183.895 22.405 184.415 ;
        RECT 23.040 183.845 23.390 184.495 ;
        RECT 17.515 182.955 18.725 183.705 ;
        RECT 18.895 182.955 22.405 183.725 ;
        RECT 23.560 183.675 23.790 184.665 ;
        RECT 23.125 183.505 23.790 183.675 ;
        RECT 23.125 183.215 23.295 183.505 ;
        RECT 23.465 182.955 23.795 183.335 ;
        RECT 23.965 183.215 24.150 185.335 ;
        RECT 24.390 185.045 24.655 185.505 ;
        RECT 24.825 184.910 25.075 185.335 ;
        RECT 25.285 185.060 26.390 185.230 ;
        RECT 24.770 184.780 25.075 184.910 ;
        RECT 24.320 183.585 24.600 184.535 ;
        RECT 24.770 183.675 24.940 184.780 ;
        RECT 25.110 183.995 25.350 184.590 ;
        RECT 25.520 184.525 26.050 184.890 ;
        RECT 25.520 183.825 25.690 184.525 ;
        RECT 26.220 184.445 26.390 185.060 ;
        RECT 26.560 184.705 26.730 185.505 ;
        RECT 26.900 185.005 27.150 185.335 ;
        RECT 27.375 185.035 28.260 185.205 ;
        RECT 26.220 184.355 26.730 184.445 ;
        RECT 24.770 183.545 24.995 183.675 ;
        RECT 25.165 183.605 25.690 183.825 ;
        RECT 25.860 184.185 26.730 184.355 ;
        RECT 24.405 182.955 24.655 183.415 ;
        RECT 24.825 183.405 24.995 183.545 ;
        RECT 25.860 183.405 26.030 184.185 ;
        RECT 26.560 184.115 26.730 184.185 ;
        RECT 26.240 183.935 26.440 183.965 ;
        RECT 26.900 183.935 27.070 185.005 ;
        RECT 27.240 184.115 27.430 184.835 ;
        RECT 26.240 183.635 27.070 183.935 ;
        RECT 27.600 183.905 27.920 184.865 ;
        RECT 24.825 183.235 25.160 183.405 ;
        RECT 25.355 183.235 26.030 183.405 ;
        RECT 26.350 182.955 26.720 183.455 ;
        RECT 26.900 183.405 27.070 183.635 ;
        RECT 27.455 183.575 27.920 183.905 ;
        RECT 28.090 184.195 28.260 185.035 ;
        RECT 28.440 185.005 28.755 185.505 ;
        RECT 28.985 184.775 29.325 185.335 ;
        RECT 28.430 184.400 29.325 184.775 ;
        RECT 29.495 184.495 29.665 185.505 ;
        RECT 29.135 184.195 29.325 184.400 ;
        RECT 29.835 184.445 30.165 185.290 ;
        RECT 29.835 184.365 30.225 184.445 ;
        RECT 30.010 184.315 30.225 184.365 ;
        RECT 30.395 184.340 30.685 185.505 ;
        RECT 30.855 184.415 32.525 185.505 ;
        RECT 33.240 184.885 33.415 185.335 ;
        RECT 33.585 185.065 33.915 185.505 ;
        RECT 34.220 184.915 34.390 185.335 ;
        RECT 34.625 185.095 35.295 185.505 ;
        RECT 35.510 184.915 35.680 185.335 ;
        RECT 35.880 185.095 36.210 185.505 ;
        RECT 33.240 184.715 33.870 184.885 ;
        RECT 28.090 183.865 28.965 184.195 ;
        RECT 29.135 183.865 29.885 184.195 ;
        RECT 28.090 183.405 28.260 183.865 ;
        RECT 29.135 183.695 29.335 183.865 ;
        RECT 30.055 183.735 30.225 184.315 ;
        RECT 30.000 183.695 30.225 183.735 ;
        RECT 26.900 183.235 27.305 183.405 ;
        RECT 27.475 183.235 28.260 183.405 ;
        RECT 28.535 182.955 28.745 183.485 ;
        RECT 29.005 183.170 29.335 183.695 ;
        RECT 29.845 183.610 30.225 183.695 ;
        RECT 30.855 183.725 31.605 184.245 ;
        RECT 31.775 183.895 32.525 184.415 ;
        RECT 33.155 183.865 33.520 184.545 ;
        RECT 33.700 184.195 33.870 184.715 ;
        RECT 34.220 184.745 36.235 184.915 ;
        RECT 33.700 183.865 34.050 184.195 ;
        RECT 29.505 182.955 29.675 183.565 ;
        RECT 29.845 183.175 30.175 183.610 ;
        RECT 30.395 182.955 30.685 183.680 ;
        RECT 30.855 182.955 32.525 183.725 ;
        RECT 33.700 183.695 33.870 183.865 ;
        RECT 33.240 183.525 33.870 183.695 ;
        RECT 33.240 183.125 33.415 183.525 ;
        RECT 34.220 183.455 34.390 184.745 ;
        RECT 33.585 182.955 33.915 183.335 ;
        RECT 34.160 183.125 34.390 183.455 ;
        RECT 34.590 183.290 34.870 184.565 ;
        RECT 35.095 184.485 35.365 184.565 ;
        RECT 35.055 184.315 35.365 184.485 ;
        RECT 35.095 183.290 35.365 184.315 ;
        RECT 35.555 183.535 35.895 184.565 ;
        RECT 36.065 184.195 36.235 184.745 ;
        RECT 36.405 184.365 36.665 185.335 ;
        RECT 36.925 184.835 37.095 185.335 ;
        RECT 37.265 185.005 37.595 185.505 ;
        RECT 36.925 184.665 37.590 184.835 ;
        RECT 36.065 183.865 36.325 184.195 ;
        RECT 36.495 183.675 36.665 184.365 ;
        RECT 36.840 183.845 37.190 184.495 ;
        RECT 37.360 183.675 37.590 184.665 ;
        RECT 35.825 182.955 36.155 183.335 ;
        RECT 36.325 183.210 36.665 183.675 ;
        RECT 36.925 183.505 37.590 183.675 ;
        RECT 36.925 183.215 37.095 183.505 ;
        RECT 36.325 183.165 36.660 183.210 ;
        RECT 37.265 182.955 37.595 183.335 ;
        RECT 37.765 183.215 37.950 185.335 ;
        RECT 38.190 185.045 38.455 185.505 ;
        RECT 38.625 184.910 38.875 185.335 ;
        RECT 39.085 185.060 40.190 185.230 ;
        RECT 38.570 184.780 38.875 184.910 ;
        RECT 38.120 183.585 38.400 184.535 ;
        RECT 38.570 183.675 38.740 184.780 ;
        RECT 38.910 183.995 39.150 184.590 ;
        RECT 39.320 184.525 39.850 184.890 ;
        RECT 39.320 183.825 39.490 184.525 ;
        RECT 40.020 184.445 40.190 185.060 ;
        RECT 40.360 184.705 40.530 185.505 ;
        RECT 40.700 185.005 40.950 185.335 ;
        RECT 41.175 185.035 42.060 185.205 ;
        RECT 40.020 184.355 40.530 184.445 ;
        RECT 38.570 183.545 38.795 183.675 ;
        RECT 38.965 183.605 39.490 183.825 ;
        RECT 39.660 184.185 40.530 184.355 ;
        RECT 38.205 182.955 38.455 183.415 ;
        RECT 38.625 183.405 38.795 183.545 ;
        RECT 39.660 183.405 39.830 184.185 ;
        RECT 40.360 184.115 40.530 184.185 ;
        RECT 40.040 183.935 40.240 183.965 ;
        RECT 40.700 183.935 40.870 185.005 ;
        RECT 41.040 184.115 41.230 184.835 ;
        RECT 40.040 183.635 40.870 183.935 ;
        RECT 41.400 183.905 41.720 184.865 ;
        RECT 38.625 183.235 38.960 183.405 ;
        RECT 39.155 183.235 39.830 183.405 ;
        RECT 40.150 182.955 40.520 183.455 ;
        RECT 40.700 183.405 40.870 183.635 ;
        RECT 41.255 183.575 41.720 183.905 ;
        RECT 41.890 184.195 42.060 185.035 ;
        RECT 42.240 185.005 42.555 185.505 ;
        RECT 42.785 184.775 43.125 185.335 ;
        RECT 42.230 184.400 43.125 184.775 ;
        RECT 43.295 184.495 43.465 185.505 ;
        RECT 42.935 184.195 43.125 184.400 ;
        RECT 43.635 184.445 43.965 185.290 ;
        RECT 43.635 184.365 44.025 184.445 ;
        RECT 44.195 184.415 47.705 185.505 ;
        RECT 47.965 184.835 48.135 185.335 ;
        RECT 48.305 185.005 48.635 185.505 ;
        RECT 47.965 184.665 48.630 184.835 ;
        RECT 43.810 184.315 44.025 184.365 ;
        RECT 41.890 183.865 42.765 184.195 ;
        RECT 42.935 183.865 43.685 184.195 ;
        RECT 41.890 183.405 42.060 183.865 ;
        RECT 42.935 183.695 43.135 183.865 ;
        RECT 43.855 183.735 44.025 184.315 ;
        RECT 43.800 183.695 44.025 183.735 ;
        RECT 40.700 183.235 41.105 183.405 ;
        RECT 41.275 183.235 42.060 183.405 ;
        RECT 42.335 182.955 42.545 183.485 ;
        RECT 42.805 183.170 43.135 183.695 ;
        RECT 43.645 183.610 44.025 183.695 ;
        RECT 44.195 183.725 45.845 184.245 ;
        RECT 46.015 183.895 47.705 184.415 ;
        RECT 47.880 183.845 48.230 184.495 ;
        RECT 43.305 182.955 43.475 183.565 ;
        RECT 43.645 183.175 43.975 183.610 ;
        RECT 44.195 182.955 47.705 183.725 ;
        RECT 48.400 183.675 48.630 184.665 ;
        RECT 47.965 183.505 48.630 183.675 ;
        RECT 47.965 183.215 48.135 183.505 ;
        RECT 48.305 182.955 48.635 183.335 ;
        RECT 48.805 183.215 48.990 185.335 ;
        RECT 49.230 185.045 49.495 185.505 ;
        RECT 49.665 184.910 49.915 185.335 ;
        RECT 50.125 185.060 51.230 185.230 ;
        RECT 49.610 184.780 49.915 184.910 ;
        RECT 49.160 183.585 49.440 184.535 ;
        RECT 49.610 183.675 49.780 184.780 ;
        RECT 49.950 183.995 50.190 184.590 ;
        RECT 50.360 184.525 50.890 184.890 ;
        RECT 50.360 183.825 50.530 184.525 ;
        RECT 51.060 184.445 51.230 185.060 ;
        RECT 51.400 184.705 51.570 185.505 ;
        RECT 51.740 185.005 51.990 185.335 ;
        RECT 52.215 185.035 53.100 185.205 ;
        RECT 51.060 184.355 51.570 184.445 ;
        RECT 49.610 183.545 49.835 183.675 ;
        RECT 50.005 183.605 50.530 183.825 ;
        RECT 50.700 184.185 51.570 184.355 ;
        RECT 49.245 182.955 49.495 183.415 ;
        RECT 49.665 183.405 49.835 183.545 ;
        RECT 50.700 183.405 50.870 184.185 ;
        RECT 51.400 184.115 51.570 184.185 ;
        RECT 51.080 183.935 51.280 183.965 ;
        RECT 51.740 183.935 51.910 185.005 ;
        RECT 52.080 184.115 52.270 184.835 ;
        RECT 51.080 183.635 51.910 183.935 ;
        RECT 52.440 183.905 52.760 184.865 ;
        RECT 49.665 183.235 50.000 183.405 ;
        RECT 50.195 183.235 50.870 183.405 ;
        RECT 51.190 182.955 51.560 183.455 ;
        RECT 51.740 183.405 51.910 183.635 ;
        RECT 52.295 183.575 52.760 183.905 ;
        RECT 52.930 184.195 53.100 185.035 ;
        RECT 53.280 185.005 53.595 185.505 ;
        RECT 53.825 184.775 54.165 185.335 ;
        RECT 53.270 184.400 54.165 184.775 ;
        RECT 54.335 184.495 54.505 185.505 ;
        RECT 53.975 184.195 54.165 184.400 ;
        RECT 54.675 184.445 55.005 185.290 ;
        RECT 54.675 184.365 55.065 184.445 ;
        RECT 54.850 184.315 55.065 184.365 ;
        RECT 56.155 184.340 56.445 185.505 ;
        RECT 56.705 184.835 56.875 185.335 ;
        RECT 57.045 185.005 57.375 185.505 ;
        RECT 56.705 184.665 57.370 184.835 ;
        RECT 52.930 183.865 53.805 184.195 ;
        RECT 53.975 183.865 54.725 184.195 ;
        RECT 52.930 183.405 53.100 183.865 ;
        RECT 53.975 183.695 54.175 183.865 ;
        RECT 54.895 183.735 55.065 184.315 ;
        RECT 56.620 183.845 56.970 184.495 ;
        RECT 54.840 183.695 55.065 183.735 ;
        RECT 51.740 183.235 52.145 183.405 ;
        RECT 52.315 183.235 53.100 183.405 ;
        RECT 53.375 182.955 53.585 183.485 ;
        RECT 53.845 183.170 54.175 183.695 ;
        RECT 54.685 183.610 55.065 183.695 ;
        RECT 54.345 182.955 54.515 183.565 ;
        RECT 54.685 183.175 55.015 183.610 ;
        RECT 56.155 182.955 56.445 183.680 ;
        RECT 57.140 183.675 57.370 184.665 ;
        RECT 56.705 183.505 57.370 183.675 ;
        RECT 56.705 183.215 56.875 183.505 ;
        RECT 57.045 182.955 57.375 183.335 ;
        RECT 57.545 183.215 57.730 185.335 ;
        RECT 57.970 185.045 58.235 185.505 ;
        RECT 58.405 184.910 58.655 185.335 ;
        RECT 58.865 185.060 59.970 185.230 ;
        RECT 58.350 184.780 58.655 184.910 ;
        RECT 57.900 183.585 58.180 184.535 ;
        RECT 58.350 183.675 58.520 184.780 ;
        RECT 58.690 183.995 58.930 184.590 ;
        RECT 59.100 184.525 59.630 184.890 ;
        RECT 59.100 183.825 59.270 184.525 ;
        RECT 59.800 184.445 59.970 185.060 ;
        RECT 60.140 184.705 60.310 185.505 ;
        RECT 60.480 185.005 60.730 185.335 ;
        RECT 60.955 185.035 61.840 185.205 ;
        RECT 59.800 184.355 60.310 184.445 ;
        RECT 58.350 183.545 58.575 183.675 ;
        RECT 58.745 183.605 59.270 183.825 ;
        RECT 59.440 184.185 60.310 184.355 ;
        RECT 57.985 182.955 58.235 183.415 ;
        RECT 58.405 183.405 58.575 183.545 ;
        RECT 59.440 183.405 59.610 184.185 ;
        RECT 60.140 184.115 60.310 184.185 ;
        RECT 59.820 183.935 60.020 183.965 ;
        RECT 60.480 183.935 60.650 185.005 ;
        RECT 60.820 184.115 61.010 184.835 ;
        RECT 59.820 183.635 60.650 183.935 ;
        RECT 61.180 183.905 61.500 184.865 ;
        RECT 58.405 183.235 58.740 183.405 ;
        RECT 58.935 183.235 59.610 183.405 ;
        RECT 59.930 182.955 60.300 183.455 ;
        RECT 60.480 183.405 60.650 183.635 ;
        RECT 61.035 183.575 61.500 183.905 ;
        RECT 61.670 184.195 61.840 185.035 ;
        RECT 62.020 185.005 62.335 185.505 ;
        RECT 62.565 184.775 62.905 185.335 ;
        RECT 62.010 184.400 62.905 184.775 ;
        RECT 63.075 184.495 63.245 185.505 ;
        RECT 62.715 184.195 62.905 184.400 ;
        RECT 63.415 184.445 63.745 185.290 ;
        RECT 63.415 184.365 63.805 184.445 ;
        RECT 63.590 184.315 63.805 184.365 ;
        RECT 61.670 183.865 62.545 184.195 ;
        RECT 62.715 183.865 63.465 184.195 ;
        RECT 61.670 183.405 61.840 183.865 ;
        RECT 62.715 183.695 62.915 183.865 ;
        RECT 63.635 183.735 63.805 184.315 ;
        RECT 63.580 183.695 63.805 183.735 ;
        RECT 60.480 183.235 60.885 183.405 ;
        RECT 61.055 183.235 61.840 183.405 ;
        RECT 62.115 182.955 62.325 183.485 ;
        RECT 62.585 183.170 62.915 183.695 ;
        RECT 63.425 183.610 63.805 183.695 ;
        RECT 64.435 184.395 64.695 185.335 ;
        RECT 64.865 185.105 65.195 185.505 ;
        RECT 66.340 185.240 66.595 185.335 ;
        RECT 65.455 185.070 66.595 185.240 ;
        RECT 66.765 185.125 67.095 185.295 ;
        RECT 65.455 184.845 65.625 185.070 ;
        RECT 64.865 184.675 65.625 184.845 ;
        RECT 66.340 184.935 66.595 185.070 ;
        RECT 64.435 183.680 64.610 184.395 ;
        RECT 64.865 184.195 65.035 184.675 ;
        RECT 65.890 184.585 66.060 184.775 ;
        RECT 66.340 184.765 66.750 184.935 ;
        RECT 64.780 183.865 65.035 184.195 ;
        RECT 65.260 183.865 65.590 184.485 ;
        RECT 65.890 184.415 66.410 184.585 ;
        RECT 65.760 183.865 66.050 184.245 ;
        RECT 66.240 183.695 66.410 184.415 ;
        RECT 63.085 182.955 63.255 183.565 ;
        RECT 63.425 183.175 63.755 183.610 ;
        RECT 64.435 183.125 64.695 183.680 ;
        RECT 65.530 183.525 66.410 183.695 ;
        RECT 66.580 183.740 66.750 184.765 ;
        RECT 66.925 184.875 67.095 185.125 ;
        RECT 67.265 185.045 67.515 185.505 ;
        RECT 67.685 184.875 67.865 185.335 ;
        RECT 66.925 184.705 67.865 184.875 ;
        RECT 66.950 184.225 67.430 184.525 ;
        RECT 66.580 183.570 66.930 183.740 ;
        RECT 67.170 183.635 67.430 184.225 ;
        RECT 67.630 183.635 67.890 184.525 ;
        RECT 68.115 184.365 68.395 185.505 ;
        RECT 68.565 184.355 68.895 185.335 ;
        RECT 69.065 184.365 69.325 185.505 ;
        RECT 69.610 184.875 69.895 185.335 ;
        RECT 70.065 185.045 70.335 185.505 ;
        RECT 69.610 184.655 70.565 184.875 ;
        RECT 68.125 183.925 68.460 184.195 ;
        RECT 68.630 183.755 68.800 184.355 ;
        RECT 68.970 183.945 69.305 184.195 ;
        RECT 69.495 183.925 70.185 184.485 ;
        RECT 70.355 183.755 70.565 184.655 ;
        RECT 64.865 182.955 65.295 183.400 ;
        RECT 65.530 183.125 65.700 183.525 ;
        RECT 65.870 182.955 66.590 183.355 ;
        RECT 66.760 183.125 66.930 183.570 ;
        RECT 67.505 182.955 67.905 183.465 ;
        RECT 68.115 182.955 68.425 183.755 ;
        RECT 68.630 183.125 69.325 183.755 ;
        RECT 69.610 183.585 70.565 183.755 ;
        RECT 70.735 184.485 71.135 185.335 ;
        RECT 71.325 184.875 71.605 185.335 ;
        RECT 72.125 185.045 72.450 185.505 ;
        RECT 71.325 184.655 72.450 184.875 ;
        RECT 70.735 183.925 71.830 184.485 ;
        RECT 72.000 184.195 72.450 184.655 ;
        RECT 72.620 184.365 73.005 185.335 ;
        RECT 69.610 183.125 69.895 183.585 ;
        RECT 70.065 182.955 70.335 183.415 ;
        RECT 70.735 183.125 71.135 183.925 ;
        RECT 72.000 183.865 72.555 184.195 ;
        RECT 72.000 183.755 72.450 183.865 ;
        RECT 71.325 183.585 72.450 183.755 ;
        RECT 72.725 183.695 73.005 184.365 ;
        RECT 71.325 183.125 71.605 183.585 ;
        RECT 72.125 182.955 72.450 183.415 ;
        RECT 72.620 183.125 73.005 183.695 ;
        RECT 73.175 183.940 73.525 185.335 ;
        RECT 73.695 184.705 74.100 185.505 ;
        RECT 74.270 185.165 75.805 185.335 ;
        RECT 74.270 184.535 74.440 185.165 ;
        RECT 73.695 184.365 74.440 184.535 ;
        RECT 73.175 183.125 73.445 183.940 ;
        RECT 73.695 183.865 73.865 184.365 ;
        RECT 74.610 184.195 74.880 184.940 ;
        RECT 74.035 183.865 74.370 184.195 ;
        RECT 74.540 183.865 74.880 184.195 ;
        RECT 75.070 184.195 75.305 184.940 ;
        RECT 75.475 184.535 75.805 185.165 ;
        RECT 75.990 184.705 76.225 185.505 ;
        RECT 76.395 184.535 76.685 185.335 ;
        RECT 75.475 184.365 76.685 184.535 ;
        RECT 76.855 184.415 78.065 185.505 ;
        RECT 78.235 184.995 79.425 185.285 ;
        RECT 75.070 183.865 75.360 184.195 ;
        RECT 75.530 183.865 75.930 184.195 ;
        RECT 76.100 183.695 76.270 184.365 ;
        RECT 76.440 183.865 76.685 184.195 ;
        RECT 76.855 183.705 77.375 184.245 ;
        RECT 77.545 183.875 78.065 184.415 ;
        RECT 78.255 184.655 79.425 184.825 ;
        RECT 79.595 184.705 79.875 185.505 ;
        RECT 78.255 184.365 78.580 184.655 ;
        RECT 79.255 184.535 79.425 184.655 ;
        RECT 78.750 184.195 78.945 184.485 ;
        RECT 79.255 184.365 79.915 184.535 ;
        RECT 80.085 184.365 80.360 185.335 ;
        RECT 80.535 184.365 80.795 185.505 ;
        RECT 79.745 184.195 79.915 184.365 ;
        RECT 78.235 183.865 78.580 184.195 ;
        RECT 78.750 183.865 79.575 184.195 ;
        RECT 79.745 183.865 80.020 184.195 ;
        RECT 73.615 182.955 74.285 183.695 ;
        RECT 74.455 183.525 75.850 183.695 ;
        RECT 74.455 183.180 74.750 183.525 ;
        RECT 74.930 182.955 75.305 183.355 ;
        RECT 75.520 183.180 75.850 183.525 ;
        RECT 76.100 183.125 76.685 183.695 ;
        RECT 76.855 182.955 78.065 183.705 ;
        RECT 79.745 183.695 79.915 183.865 ;
        RECT 78.250 183.525 79.915 183.695 ;
        RECT 80.190 183.630 80.360 184.365 ;
        RECT 80.965 184.355 81.295 185.335 ;
        RECT 81.465 184.365 81.745 185.505 ;
        RECT 80.555 183.945 80.890 184.195 ;
        RECT 81.060 183.755 81.230 184.355 ;
        RECT 81.915 184.340 82.205 185.505 ;
        RECT 83.355 184.445 83.685 185.290 ;
        RECT 83.855 184.495 84.025 185.505 ;
        RECT 84.195 184.775 84.535 185.335 ;
        RECT 84.765 185.005 85.080 185.505 ;
        RECT 85.260 185.035 86.145 185.205 ;
        RECT 83.295 184.365 83.685 184.445 ;
        RECT 84.195 184.400 85.090 184.775 ;
        RECT 83.295 184.315 83.510 184.365 ;
        RECT 81.400 183.925 81.735 184.195 ;
        RECT 78.250 183.175 78.505 183.525 ;
        RECT 78.675 182.955 79.005 183.355 ;
        RECT 79.175 183.175 79.345 183.525 ;
        RECT 79.515 182.955 79.895 183.355 ;
        RECT 80.085 183.285 80.360 183.630 ;
        RECT 80.535 183.125 81.230 183.755 ;
        RECT 81.435 182.955 81.745 183.755 ;
        RECT 83.295 183.735 83.465 184.315 ;
        RECT 84.195 184.195 84.385 184.400 ;
        RECT 85.260 184.195 85.430 185.035 ;
        RECT 86.370 185.005 86.620 185.335 ;
        RECT 83.635 183.865 84.385 184.195 ;
        RECT 84.555 183.865 85.430 184.195 ;
        RECT 83.295 183.695 83.520 183.735 ;
        RECT 84.185 183.695 84.385 183.865 ;
        RECT 81.915 182.955 82.205 183.680 ;
        RECT 83.295 183.610 83.675 183.695 ;
        RECT 83.345 183.175 83.675 183.610 ;
        RECT 83.845 182.955 84.015 183.565 ;
        RECT 84.185 183.170 84.515 183.695 ;
        RECT 84.775 182.955 84.985 183.485 ;
        RECT 85.260 183.405 85.430 183.865 ;
        RECT 85.600 183.905 85.920 184.865 ;
        RECT 86.090 184.115 86.280 184.835 ;
        RECT 86.450 183.935 86.620 185.005 ;
        RECT 86.790 184.705 86.960 185.505 ;
        RECT 87.130 185.060 88.235 185.230 ;
        RECT 87.130 184.445 87.300 185.060 ;
        RECT 88.445 184.910 88.695 185.335 ;
        RECT 88.865 185.045 89.130 185.505 ;
        RECT 87.470 184.525 88.000 184.890 ;
        RECT 88.445 184.780 88.750 184.910 ;
        RECT 86.790 184.355 87.300 184.445 ;
        RECT 86.790 184.185 87.660 184.355 ;
        RECT 86.790 184.115 86.960 184.185 ;
        RECT 87.080 183.935 87.280 183.965 ;
        RECT 85.600 183.575 86.065 183.905 ;
        RECT 86.450 183.635 87.280 183.935 ;
        RECT 86.450 183.405 86.620 183.635 ;
        RECT 85.260 183.235 86.045 183.405 ;
        RECT 86.215 183.235 86.620 183.405 ;
        RECT 86.800 182.955 87.170 183.455 ;
        RECT 87.490 183.405 87.660 184.185 ;
        RECT 87.830 183.825 88.000 184.525 ;
        RECT 88.170 183.995 88.410 184.590 ;
        RECT 87.830 183.605 88.355 183.825 ;
        RECT 88.580 183.675 88.750 184.780 ;
        RECT 88.525 183.545 88.750 183.675 ;
        RECT 88.920 183.585 89.200 184.535 ;
        RECT 88.525 183.405 88.695 183.545 ;
        RECT 87.490 183.235 88.165 183.405 ;
        RECT 88.360 183.235 88.695 183.405 ;
        RECT 88.865 182.955 89.115 183.415 ;
        RECT 89.370 183.215 89.555 185.335 ;
        RECT 89.725 185.005 90.055 185.505 ;
        RECT 90.225 184.835 90.395 185.335 ;
        RECT 89.730 184.665 90.395 184.835 ;
        RECT 90.770 184.875 91.055 185.335 ;
        RECT 91.225 185.045 91.495 185.505 ;
        RECT 89.730 183.675 89.960 184.665 ;
        RECT 90.770 184.655 91.725 184.875 ;
        RECT 90.130 183.845 90.480 184.495 ;
        RECT 90.655 183.925 91.345 184.485 ;
        RECT 91.515 183.755 91.725 184.655 ;
        RECT 89.730 183.505 90.395 183.675 ;
        RECT 89.725 182.955 90.055 183.335 ;
        RECT 90.225 183.215 90.395 183.505 ;
        RECT 90.770 183.585 91.725 183.755 ;
        RECT 91.895 184.485 92.295 185.335 ;
        RECT 92.485 184.875 92.765 185.335 ;
        RECT 93.285 185.045 93.610 185.505 ;
        RECT 92.485 184.655 93.610 184.875 ;
        RECT 91.895 183.925 92.990 184.485 ;
        RECT 93.160 184.195 93.610 184.655 ;
        RECT 93.780 184.365 94.165 185.335 ;
        RECT 94.425 184.835 94.595 185.335 ;
        RECT 94.765 185.005 95.095 185.505 ;
        RECT 94.425 184.665 95.090 184.835 ;
        RECT 90.770 183.125 91.055 183.585 ;
        RECT 91.225 182.955 91.495 183.415 ;
        RECT 91.895 183.125 92.295 183.925 ;
        RECT 93.160 183.865 93.715 184.195 ;
        RECT 93.160 183.755 93.610 183.865 ;
        RECT 92.485 183.585 93.610 183.755 ;
        RECT 93.885 183.695 94.165 184.365 ;
        RECT 94.340 183.845 94.690 184.495 ;
        RECT 92.485 183.125 92.765 183.585 ;
        RECT 93.285 182.955 93.610 183.415 ;
        RECT 93.780 183.125 94.165 183.695 ;
        RECT 94.860 183.675 95.090 184.665 ;
        RECT 94.425 183.505 95.090 183.675 ;
        RECT 94.425 183.215 94.595 183.505 ;
        RECT 94.765 182.955 95.095 183.335 ;
        RECT 95.265 183.215 95.450 185.335 ;
        RECT 95.690 185.045 95.955 185.505 ;
        RECT 96.125 184.910 96.375 185.335 ;
        RECT 96.585 185.060 97.690 185.230 ;
        RECT 96.070 184.780 96.375 184.910 ;
        RECT 95.620 183.585 95.900 184.535 ;
        RECT 96.070 183.675 96.240 184.780 ;
        RECT 96.410 183.995 96.650 184.590 ;
        RECT 96.820 184.525 97.350 184.890 ;
        RECT 96.820 183.825 96.990 184.525 ;
        RECT 97.520 184.445 97.690 185.060 ;
        RECT 97.860 184.705 98.030 185.505 ;
        RECT 98.200 185.005 98.450 185.335 ;
        RECT 98.675 185.035 99.560 185.205 ;
        RECT 97.520 184.355 98.030 184.445 ;
        RECT 96.070 183.545 96.295 183.675 ;
        RECT 96.465 183.605 96.990 183.825 ;
        RECT 97.160 184.185 98.030 184.355 ;
        RECT 95.705 182.955 95.955 183.415 ;
        RECT 96.125 183.405 96.295 183.545 ;
        RECT 97.160 183.405 97.330 184.185 ;
        RECT 97.860 184.115 98.030 184.185 ;
        RECT 97.540 183.935 97.740 183.965 ;
        RECT 98.200 183.935 98.370 185.005 ;
        RECT 98.540 184.115 98.730 184.835 ;
        RECT 97.540 183.635 98.370 183.935 ;
        RECT 98.900 183.905 99.220 184.865 ;
        RECT 96.125 183.235 96.460 183.405 ;
        RECT 96.655 183.235 97.330 183.405 ;
        RECT 97.650 182.955 98.020 183.455 ;
        RECT 98.200 183.405 98.370 183.635 ;
        RECT 98.755 183.575 99.220 183.905 ;
        RECT 99.390 184.195 99.560 185.035 ;
        RECT 99.740 185.005 100.055 185.505 ;
        RECT 100.285 184.775 100.625 185.335 ;
        RECT 99.730 184.400 100.625 184.775 ;
        RECT 100.795 184.495 100.965 185.505 ;
        RECT 100.435 184.195 100.625 184.400 ;
        RECT 101.135 184.445 101.465 185.290 ;
        RECT 101.135 184.365 101.525 184.445 ;
        RECT 101.310 184.315 101.525 184.365 ;
        RECT 99.390 183.865 100.265 184.195 ;
        RECT 100.435 183.865 101.185 184.195 ;
        RECT 99.390 183.405 99.560 183.865 ;
        RECT 100.435 183.695 100.635 183.865 ;
        RECT 101.355 183.735 101.525 184.315 ;
        RECT 101.300 183.695 101.525 183.735 ;
        RECT 98.200 183.235 98.605 183.405 ;
        RECT 98.775 183.235 99.560 183.405 ;
        RECT 99.835 182.955 100.045 183.485 ;
        RECT 100.305 183.170 100.635 183.695 ;
        RECT 101.145 183.610 101.525 183.695 ;
        RECT 101.695 184.365 102.080 185.335 ;
        RECT 102.250 185.045 102.575 185.505 ;
        RECT 103.095 184.875 103.375 185.335 ;
        RECT 102.250 184.655 103.375 184.875 ;
        RECT 101.695 183.695 101.975 184.365 ;
        RECT 102.250 184.195 102.700 184.655 ;
        RECT 103.565 184.485 103.965 185.335 ;
        RECT 104.365 185.045 104.635 185.505 ;
        RECT 104.805 184.875 105.090 185.335 ;
        RECT 105.375 184.995 106.565 185.285 ;
        RECT 102.145 183.865 102.700 184.195 ;
        RECT 102.870 183.925 103.965 184.485 ;
        RECT 102.250 183.755 102.700 183.865 ;
        RECT 100.805 182.955 100.975 183.565 ;
        RECT 101.145 183.175 101.475 183.610 ;
        RECT 101.695 183.125 102.080 183.695 ;
        RECT 102.250 183.585 103.375 183.755 ;
        RECT 102.250 182.955 102.575 183.415 ;
        RECT 103.095 183.125 103.375 183.585 ;
        RECT 103.565 183.125 103.965 183.925 ;
        RECT 104.135 184.655 105.090 184.875 ;
        RECT 105.395 184.655 106.565 184.825 ;
        RECT 106.735 184.705 107.015 185.505 ;
        RECT 104.135 183.755 104.345 184.655 ;
        RECT 104.515 183.925 105.205 184.485 ;
        RECT 105.395 184.365 105.720 184.655 ;
        RECT 106.395 184.535 106.565 184.655 ;
        RECT 105.890 184.195 106.085 184.485 ;
        RECT 106.395 184.365 107.055 184.535 ;
        RECT 107.225 184.365 107.500 185.335 ;
        RECT 106.885 184.195 107.055 184.365 ;
        RECT 105.375 183.865 105.720 184.195 ;
        RECT 105.890 183.865 106.715 184.195 ;
        RECT 106.885 183.865 107.160 184.195 ;
        RECT 104.135 183.585 105.090 183.755 ;
        RECT 106.885 183.695 107.055 183.865 ;
        RECT 104.365 182.955 104.635 183.415 ;
        RECT 104.805 183.125 105.090 183.585 ;
        RECT 105.390 183.525 107.055 183.695 ;
        RECT 107.330 183.630 107.500 184.365 ;
        RECT 107.675 184.340 107.965 185.505 ;
        RECT 108.140 184.555 108.405 185.325 ;
        RECT 108.575 184.785 108.905 185.505 ;
        RECT 109.095 184.965 109.355 185.325 ;
        RECT 109.525 185.135 109.855 185.505 ;
        RECT 110.025 184.965 110.285 185.325 ;
        RECT 109.095 184.735 110.285 184.965 ;
        RECT 110.855 184.555 111.145 185.325 ;
        RECT 105.390 183.175 105.645 183.525 ;
        RECT 105.815 182.955 106.145 183.355 ;
        RECT 106.315 183.175 106.485 183.525 ;
        RECT 106.655 182.955 107.035 183.355 ;
        RECT 107.225 183.285 107.500 183.630 ;
        RECT 107.675 182.955 107.965 183.680 ;
        RECT 108.140 183.135 108.475 184.555 ;
        RECT 108.650 184.375 111.145 184.555 ;
        RECT 108.650 183.685 108.875 184.375 ;
        RECT 111.355 184.365 111.615 185.505 ;
        RECT 111.785 184.535 112.115 185.335 ;
        RECT 112.285 184.705 112.455 185.505 ;
        RECT 112.625 184.535 112.955 185.335 ;
        RECT 113.125 184.705 113.380 185.505 ;
        RECT 114.205 185.165 115.365 185.335 ;
        RECT 114.205 184.665 114.375 185.165 ;
        RECT 114.635 184.535 114.805 184.995 ;
        RECT 115.035 184.915 115.365 185.165 ;
        RECT 115.590 185.085 115.920 185.505 ;
        RECT 116.175 184.915 116.460 185.335 ;
        RECT 115.035 184.745 116.460 184.915 ;
        RECT 116.705 184.705 117.035 185.505 ;
        RECT 117.285 184.785 117.620 185.295 ;
        RECT 111.785 184.365 113.485 184.535 ;
        RECT 109.075 183.865 109.355 184.195 ;
        RECT 109.535 183.865 110.110 184.195 ;
        RECT 110.290 183.865 110.725 184.195 ;
        RECT 110.905 183.865 111.175 184.195 ;
        RECT 111.355 183.945 112.115 184.195 ;
        RECT 112.285 183.945 113.035 184.195 ;
        RECT 113.205 183.775 113.485 184.365 ;
        RECT 114.180 184.195 114.385 184.485 ;
        RECT 114.635 184.365 117.005 184.535 ;
        RECT 116.835 184.195 117.005 184.365 ;
        RECT 114.180 184.145 114.530 184.195 ;
        RECT 114.175 183.975 114.530 184.145 ;
        RECT 114.180 183.865 114.530 183.975 ;
        RECT 108.650 183.495 111.135 183.685 ;
        RECT 108.655 182.955 109.400 183.325 ;
        RECT 109.965 183.135 110.220 183.495 ;
        RECT 110.400 182.955 110.730 183.325 ;
        RECT 110.910 183.135 111.135 183.495 ;
        RECT 111.355 183.585 112.455 183.755 ;
        RECT 111.355 183.125 111.695 183.585 ;
        RECT 111.865 182.955 112.035 183.415 ;
        RECT 112.205 183.335 112.455 183.585 ;
        RECT 112.625 183.525 113.485 183.775 ;
        RECT 113.045 183.335 113.375 183.355 ;
        RECT 112.205 183.125 113.375 183.335 ;
        RECT 114.125 182.955 114.455 183.675 ;
        RECT 114.840 183.530 115.260 184.195 ;
        RECT 115.430 183.805 115.720 184.195 ;
        RECT 115.910 183.805 116.180 184.195 ;
        RECT 116.390 184.145 116.640 184.195 ;
        RECT 116.390 183.975 116.645 184.145 ;
        RECT 116.390 183.865 116.640 183.975 ;
        RECT 116.835 183.865 117.140 184.195 ;
        RECT 115.430 183.635 115.725 183.805 ;
        RECT 115.910 183.635 116.185 183.805 ;
        RECT 116.835 183.695 117.005 183.865 ;
        RECT 115.430 183.535 115.720 183.635 ;
        RECT 115.910 183.535 116.180 183.635 ;
        RECT 116.445 183.525 117.005 183.695 ;
        RECT 116.445 183.355 116.615 183.525 ;
        RECT 117.365 183.430 117.620 184.785 ;
        RECT 115.000 183.185 116.615 183.355 ;
        RECT 116.785 182.955 117.115 183.355 ;
        RECT 117.285 183.170 117.620 183.430 ;
        RECT 117.830 184.715 118.365 185.335 ;
        RECT 117.830 183.695 118.145 184.715 ;
        RECT 118.535 184.705 118.865 185.505 ;
        RECT 119.350 184.535 119.740 184.710 ;
        RECT 118.315 184.365 119.740 184.535 ;
        RECT 120.105 184.535 120.435 185.320 ;
        RECT 120.105 184.365 120.785 184.535 ;
        RECT 120.965 184.365 121.295 185.505 ;
        RECT 121.475 184.365 121.735 185.505 ;
        RECT 118.315 183.865 118.485 184.365 ;
        RECT 117.830 183.125 118.445 183.695 ;
        RECT 118.735 183.635 119.000 184.195 ;
        RECT 119.170 183.465 119.340 184.365 ;
        RECT 119.510 183.635 119.865 184.195 ;
        RECT 120.095 183.945 120.445 184.195 ;
        RECT 120.615 183.765 120.785 184.365 ;
        RECT 121.905 184.355 122.235 185.335 ;
        RECT 122.405 184.365 122.685 185.505 ;
        RECT 122.855 185.070 128.200 185.505 ;
        RECT 120.955 183.945 121.305 184.195 ;
        RECT 121.495 183.945 121.830 184.195 ;
        RECT 118.615 182.955 118.830 183.465 ;
        RECT 119.060 183.135 119.340 183.465 ;
        RECT 119.520 182.955 119.760 183.465 ;
        RECT 120.115 182.955 120.355 183.765 ;
        RECT 120.525 183.125 120.855 183.765 ;
        RECT 121.025 182.955 121.295 183.765 ;
        RECT 122.000 183.755 122.170 184.355 ;
        RECT 122.340 183.925 122.675 184.195 ;
        RECT 121.475 183.125 122.170 183.755 ;
        RECT 122.375 182.955 122.685 183.755 ;
        RECT 124.440 183.500 124.780 184.330 ;
        RECT 126.260 183.820 126.610 185.070 ;
        RECT 128.375 184.415 131.885 185.505 ;
        RECT 132.055 184.415 133.265 185.505 ;
        RECT 128.375 183.725 130.025 184.245 ;
        RECT 130.195 183.895 131.885 184.415 ;
        RECT 122.855 182.955 128.200 183.500 ;
        RECT 128.375 182.955 131.885 183.725 ;
        RECT 132.055 183.705 132.575 184.245 ;
        RECT 132.745 183.875 133.265 184.415 ;
        RECT 133.435 184.340 133.725 185.505 ;
        RECT 133.895 184.415 137.405 185.505 ;
        RECT 133.895 183.725 135.545 184.245 ;
        RECT 135.715 183.895 137.405 184.415 ;
        RECT 138.125 184.575 138.295 185.335 ;
        RECT 138.475 184.745 138.805 185.505 ;
        RECT 138.125 184.405 138.790 184.575 ;
        RECT 138.975 184.430 139.245 185.335 ;
        RECT 138.620 184.260 138.790 184.405 ;
        RECT 138.055 183.855 138.385 184.225 ;
        RECT 138.620 183.930 138.905 184.260 ;
        RECT 132.055 182.955 133.265 183.705 ;
        RECT 133.435 182.955 133.725 183.680 ;
        RECT 133.895 182.955 137.405 183.725 ;
        RECT 138.620 183.675 138.790 183.930 ;
        RECT 138.125 183.505 138.790 183.675 ;
        RECT 139.075 183.630 139.245 184.430 ;
        RECT 138.125 183.125 138.295 183.505 ;
        RECT 138.475 182.955 138.805 183.335 ;
        RECT 138.985 183.125 139.245 183.630 ;
        RECT 140.335 184.430 140.605 185.335 ;
        RECT 140.775 184.745 141.105 185.505 ;
        RECT 141.285 184.575 141.465 185.335 ;
        RECT 140.335 183.630 140.515 184.430 ;
        RECT 140.790 184.405 141.465 184.575 ;
        RECT 141.715 184.415 142.925 185.505 ;
        RECT 140.790 184.260 140.960 184.405 ;
        RECT 140.685 183.930 140.960 184.260 ;
        RECT 140.790 183.675 140.960 183.930 ;
        RECT 141.185 183.855 141.525 184.225 ;
        RECT 141.715 183.875 142.235 184.415 ;
        RECT 142.405 183.705 142.925 184.245 ;
        RECT 140.335 183.125 140.595 183.630 ;
        RECT 140.790 183.505 141.455 183.675 ;
        RECT 140.775 182.955 141.105 183.335 ;
        RECT 141.285 183.125 141.455 183.505 ;
        RECT 141.715 182.955 142.925 183.705 ;
        RECT 17.430 182.785 143.010 182.955 ;
        RECT 17.515 182.035 18.725 182.785 ;
        RECT 18.895 182.240 24.240 182.785 ;
        RECT 24.420 182.530 24.755 182.575 ;
        RECT 17.515 181.495 18.035 182.035 ;
        RECT 18.205 181.325 18.725 181.865 ;
        RECT 20.480 181.410 20.820 182.240 ;
        RECT 24.415 182.065 24.755 182.530 ;
        RECT 24.925 182.405 25.255 182.785 ;
        RECT 17.515 180.235 18.725 181.325 ;
        RECT 22.300 180.670 22.650 181.920 ;
        RECT 24.415 181.375 24.585 182.065 ;
        RECT 24.755 181.545 25.015 181.875 ;
        RECT 18.895 180.235 24.240 180.670 ;
        RECT 24.415 180.405 24.675 181.375 ;
        RECT 24.845 180.995 25.015 181.545 ;
        RECT 25.185 181.175 25.525 182.205 ;
        RECT 25.715 181.425 25.985 182.450 ;
        RECT 25.715 181.255 26.025 181.425 ;
        RECT 25.715 181.175 25.985 181.255 ;
        RECT 26.210 181.175 26.490 182.450 ;
        RECT 26.690 182.285 26.920 182.615 ;
        RECT 27.165 182.405 27.495 182.785 ;
        RECT 26.690 180.995 26.860 182.285 ;
        RECT 27.665 182.215 27.840 182.615 ;
        RECT 27.210 182.045 27.840 182.215 ;
        RECT 27.210 181.875 27.380 182.045 ;
        RECT 28.095 181.950 28.385 182.785 ;
        RECT 28.555 182.385 29.510 182.555 ;
        RECT 29.925 182.395 30.255 182.785 ;
        RECT 27.030 181.545 27.380 181.875 ;
        RECT 24.845 180.825 26.860 180.995 ;
        RECT 27.210 181.025 27.380 181.545 ;
        RECT 27.560 181.195 27.925 181.875 ;
        RECT 28.555 181.505 28.725 182.385 ;
        RECT 30.425 182.215 30.595 182.535 ;
        RECT 30.765 182.395 31.095 182.785 ;
        RECT 28.895 182.045 31.145 182.215 ;
        RECT 28.895 181.545 29.125 182.045 ;
        RECT 29.295 181.625 29.670 181.795 ;
        RECT 28.095 181.335 28.725 181.505 ;
        RECT 29.500 181.425 29.670 181.625 ;
        RECT 29.840 181.595 30.390 181.795 ;
        RECT 30.560 181.425 30.805 181.875 ;
        RECT 27.210 180.855 27.840 181.025 ;
        RECT 24.870 180.235 25.200 180.645 ;
        RECT 25.400 180.405 25.570 180.825 ;
        RECT 25.785 180.235 26.455 180.645 ;
        RECT 26.690 180.405 26.860 180.825 ;
        RECT 27.165 180.235 27.495 180.675 ;
        RECT 27.665 180.405 27.840 180.855 ;
        RECT 28.095 180.405 28.415 181.335 ;
        RECT 29.500 181.255 30.805 181.425 ;
        RECT 30.975 181.085 31.145 182.045 ;
        RECT 31.315 182.035 32.525 182.785 ;
        RECT 32.695 182.405 33.585 182.575 ;
        RECT 31.315 181.495 31.835 182.035 ;
        RECT 32.005 181.325 32.525 181.865 ;
        RECT 32.695 181.850 33.245 182.235 ;
        RECT 33.415 181.680 33.585 182.405 ;
        RECT 28.595 180.915 29.835 181.085 ;
        RECT 28.595 180.405 28.995 180.915 ;
        RECT 29.165 180.235 29.335 180.745 ;
        RECT 29.505 180.405 29.835 180.915 ;
        RECT 30.005 180.235 30.175 181.085 ;
        RECT 30.765 180.405 31.145 181.085 ;
        RECT 31.315 180.235 32.525 181.325 ;
        RECT 32.695 181.610 33.585 181.680 ;
        RECT 33.755 182.080 33.975 182.565 ;
        RECT 34.145 182.245 34.395 182.785 ;
        RECT 34.565 182.135 34.825 182.615 ;
        RECT 33.755 181.655 34.085 182.080 ;
        RECT 32.695 181.585 33.590 181.610 ;
        RECT 32.695 181.570 33.600 181.585 ;
        RECT 32.695 181.555 33.605 181.570 ;
        RECT 32.695 181.550 33.615 181.555 ;
        RECT 32.695 181.540 33.620 181.550 ;
        RECT 32.695 181.530 33.625 181.540 ;
        RECT 32.695 181.525 33.635 181.530 ;
        RECT 32.695 181.515 33.645 181.525 ;
        RECT 32.695 181.510 33.655 181.515 ;
        RECT 32.695 181.060 32.955 181.510 ;
        RECT 33.320 181.505 33.655 181.510 ;
        RECT 33.320 181.500 33.670 181.505 ;
        RECT 33.320 181.490 33.685 181.500 ;
        RECT 33.320 181.485 33.710 181.490 ;
        RECT 34.255 181.485 34.485 181.880 ;
        RECT 33.320 181.480 34.485 181.485 ;
        RECT 33.350 181.445 34.485 181.480 ;
        RECT 33.385 181.420 34.485 181.445 ;
        RECT 33.415 181.390 34.485 181.420 ;
        RECT 33.435 181.360 34.485 181.390 ;
        RECT 33.455 181.330 34.485 181.360 ;
        RECT 33.525 181.320 34.485 181.330 ;
        RECT 33.550 181.310 34.485 181.320 ;
        RECT 33.570 181.295 34.485 181.310 ;
        RECT 33.590 181.280 34.485 181.295 ;
        RECT 33.595 181.270 34.380 181.280 ;
        RECT 33.610 181.235 34.380 181.270 ;
        RECT 33.125 180.915 33.455 181.160 ;
        RECT 33.625 180.985 34.380 181.235 ;
        RECT 34.655 181.105 34.825 182.135 ;
        RECT 35.085 182.235 35.255 182.525 ;
        RECT 35.425 182.405 35.755 182.785 ;
        RECT 35.085 182.065 35.750 182.235 ;
        RECT 35.000 181.245 35.350 181.895 ;
        RECT 33.125 180.890 33.310 180.915 ;
        RECT 32.695 180.790 33.310 180.890 ;
        RECT 32.695 180.235 33.300 180.790 ;
        RECT 33.475 180.405 33.955 180.745 ;
        RECT 34.125 180.235 34.380 180.780 ;
        RECT 34.550 180.405 34.825 181.105 ;
        RECT 35.520 181.075 35.750 182.065 ;
        RECT 35.085 180.905 35.750 181.075 ;
        RECT 35.085 180.405 35.255 180.905 ;
        RECT 35.425 180.235 35.755 180.735 ;
        RECT 35.925 180.405 36.110 182.525 ;
        RECT 36.365 182.325 36.615 182.785 ;
        RECT 36.785 182.335 37.120 182.505 ;
        RECT 37.315 182.335 37.990 182.505 ;
        RECT 36.785 182.195 36.955 182.335 ;
        RECT 36.280 181.205 36.560 182.155 ;
        RECT 36.730 182.065 36.955 182.195 ;
        RECT 36.730 180.960 36.900 182.065 ;
        RECT 37.125 181.915 37.650 182.135 ;
        RECT 37.070 181.150 37.310 181.745 ;
        RECT 37.480 181.215 37.650 181.915 ;
        RECT 37.820 181.555 37.990 182.335 ;
        RECT 38.310 182.285 38.680 182.785 ;
        RECT 38.860 182.335 39.265 182.505 ;
        RECT 39.435 182.335 40.220 182.505 ;
        RECT 38.860 182.105 39.030 182.335 ;
        RECT 38.200 181.805 39.030 182.105 ;
        RECT 39.415 181.835 39.880 182.165 ;
        RECT 38.200 181.775 38.400 181.805 ;
        RECT 38.520 181.555 38.690 181.625 ;
        RECT 37.820 181.385 38.690 181.555 ;
        RECT 38.180 181.295 38.690 181.385 ;
        RECT 36.730 180.830 37.035 180.960 ;
        RECT 37.480 180.850 38.010 181.215 ;
        RECT 36.350 180.235 36.615 180.695 ;
        RECT 36.785 180.405 37.035 180.830 ;
        RECT 38.180 180.680 38.350 181.295 ;
        RECT 37.245 180.510 38.350 180.680 ;
        RECT 38.520 180.235 38.690 181.035 ;
        RECT 38.860 180.735 39.030 181.805 ;
        RECT 39.200 180.905 39.390 181.625 ;
        RECT 39.560 180.875 39.880 181.835 ;
        RECT 40.050 181.875 40.220 182.335 ;
        RECT 40.495 182.255 40.705 182.785 ;
        RECT 40.965 182.045 41.295 182.570 ;
        RECT 41.465 182.175 41.635 182.785 ;
        RECT 41.805 182.130 42.135 182.565 ;
        RECT 41.805 182.045 42.185 182.130 ;
        RECT 43.275 182.060 43.565 182.785 ;
        RECT 43.785 182.395 44.115 182.785 ;
        RECT 44.285 182.215 44.455 182.535 ;
        RECT 44.625 182.395 44.955 182.785 ;
        RECT 45.370 182.385 46.325 182.555 ;
        RECT 41.095 181.875 41.295 182.045 ;
        RECT 41.960 182.005 42.185 182.045 ;
        RECT 40.050 181.545 40.925 181.875 ;
        RECT 41.095 181.545 41.845 181.875 ;
        RECT 38.860 180.405 39.110 180.735 ;
        RECT 40.050 180.705 40.220 181.545 ;
        RECT 41.095 181.340 41.285 181.545 ;
        RECT 42.015 181.425 42.185 182.005 ;
        RECT 41.970 181.375 42.185 181.425 ;
        RECT 43.735 182.045 45.985 182.215 ;
        RECT 40.390 180.965 41.285 181.340 ;
        RECT 41.795 181.295 42.185 181.375 ;
        RECT 39.335 180.535 40.220 180.705 ;
        RECT 40.400 180.235 40.715 180.735 ;
        RECT 40.945 180.405 41.285 180.965 ;
        RECT 41.455 180.235 41.625 181.245 ;
        RECT 41.795 180.450 42.125 181.295 ;
        RECT 43.275 180.235 43.565 181.400 ;
        RECT 43.735 181.085 43.905 182.045 ;
        RECT 44.075 181.425 44.320 181.875 ;
        RECT 44.490 181.595 45.040 181.795 ;
        RECT 45.210 181.625 45.585 181.795 ;
        RECT 45.210 181.425 45.380 181.625 ;
        RECT 45.755 181.545 45.985 182.045 ;
        RECT 44.075 181.255 45.380 181.425 ;
        RECT 46.155 181.505 46.325 182.385 ;
        RECT 46.495 181.950 46.785 182.785 ;
        RECT 46.960 182.530 47.295 182.575 ;
        RECT 46.955 182.065 47.295 182.530 ;
        RECT 47.465 182.405 47.795 182.785 ;
        RECT 46.155 181.335 46.785 181.505 ;
        RECT 43.735 180.405 44.115 181.085 ;
        RECT 44.705 180.235 44.875 181.085 ;
        RECT 45.045 180.915 46.285 181.085 ;
        RECT 45.045 180.405 45.375 180.915 ;
        RECT 45.545 180.235 45.715 180.745 ;
        RECT 45.885 180.405 46.285 180.915 ;
        RECT 46.465 180.405 46.785 181.335 ;
        RECT 46.955 181.375 47.125 182.065 ;
        RECT 47.295 181.545 47.555 181.875 ;
        RECT 46.955 180.405 47.215 181.375 ;
        RECT 47.385 180.995 47.555 181.545 ;
        RECT 47.725 181.175 48.065 182.205 ;
        RECT 48.255 182.105 48.525 182.450 ;
        RECT 48.255 181.935 48.565 182.105 ;
        RECT 48.255 181.175 48.525 181.935 ;
        RECT 48.750 181.175 49.030 182.450 ;
        RECT 49.230 182.285 49.460 182.615 ;
        RECT 49.705 182.405 50.035 182.785 ;
        RECT 49.230 180.995 49.400 182.285 ;
        RECT 50.205 182.215 50.380 182.615 ;
        RECT 49.750 182.045 50.380 182.215 ;
        RECT 49.750 181.875 49.920 182.045 ;
        RECT 50.635 182.015 54.145 182.785 ;
        RECT 54.325 182.055 54.625 182.785 ;
        RECT 49.570 181.545 49.920 181.875 ;
        RECT 47.385 180.825 49.400 180.995 ;
        RECT 49.750 181.025 49.920 181.545 ;
        RECT 50.100 181.195 50.465 181.875 ;
        RECT 50.635 181.495 52.285 182.015 ;
        RECT 54.805 181.875 55.035 182.495 ;
        RECT 55.235 182.225 55.460 182.605 ;
        RECT 55.630 182.395 55.960 182.785 ;
        RECT 56.155 182.240 61.500 182.785 ;
        RECT 61.675 182.240 67.020 182.785 ;
        RECT 55.235 182.045 55.565 182.225 ;
        RECT 52.455 181.325 54.145 181.845 ;
        RECT 54.330 181.545 54.625 181.875 ;
        RECT 54.805 181.545 55.220 181.875 ;
        RECT 55.390 181.375 55.565 182.045 ;
        RECT 55.735 181.545 55.975 182.195 ;
        RECT 57.740 181.410 58.080 182.240 ;
        RECT 49.750 180.855 50.380 181.025 ;
        RECT 47.410 180.235 47.740 180.645 ;
        RECT 47.940 180.405 48.110 180.825 ;
        RECT 48.325 180.235 48.995 180.645 ;
        RECT 49.230 180.405 49.400 180.825 ;
        RECT 49.705 180.235 50.035 180.675 ;
        RECT 50.205 180.405 50.380 180.855 ;
        RECT 50.635 180.235 54.145 181.325 ;
        RECT 54.325 181.015 55.220 181.345 ;
        RECT 55.390 181.185 55.975 181.375 ;
        RECT 54.325 180.845 55.530 181.015 ;
        RECT 54.325 180.415 54.655 180.845 ;
        RECT 54.835 180.235 55.030 180.675 ;
        RECT 55.200 180.415 55.530 180.845 ;
        RECT 55.700 180.415 55.975 181.185 ;
        RECT 59.560 180.670 59.910 181.920 ;
        RECT 63.260 181.410 63.600 182.240 ;
        RECT 67.715 181.965 67.925 182.785 ;
        RECT 68.095 181.985 68.425 182.615 ;
        RECT 65.080 180.670 65.430 181.920 ;
        RECT 68.095 181.385 68.345 181.985 ;
        RECT 68.595 181.965 68.825 182.785 ;
        RECT 69.035 182.060 69.325 182.785 ;
        RECT 69.500 182.110 69.775 182.455 ;
        RECT 69.965 182.385 70.345 182.785 ;
        RECT 70.515 182.215 70.685 182.565 ;
        RECT 70.855 182.385 71.185 182.785 ;
        RECT 71.355 182.215 71.610 182.565 ;
        RECT 71.960 182.275 72.200 182.785 ;
        RECT 72.380 182.275 72.660 182.605 ;
        RECT 72.890 182.275 73.105 182.785 ;
        RECT 68.515 181.545 68.845 181.795 ;
        RECT 56.155 180.235 61.500 180.670 ;
        RECT 61.675 180.235 67.020 180.670 ;
        RECT 67.715 180.235 67.925 181.375 ;
        RECT 68.095 180.405 68.425 181.385 ;
        RECT 68.595 180.235 68.825 181.375 ;
        RECT 69.035 180.235 69.325 181.400 ;
        RECT 69.500 181.375 69.670 182.110 ;
        RECT 69.945 182.045 71.610 182.215 ;
        RECT 69.945 181.875 70.115 182.045 ;
        RECT 69.840 181.545 70.115 181.875 ;
        RECT 70.285 181.545 71.110 181.875 ;
        RECT 71.280 181.545 71.625 181.875 ;
        RECT 71.855 181.545 72.210 182.105 ;
        RECT 69.945 181.375 70.115 181.545 ;
        RECT 69.500 180.405 69.775 181.375 ;
        RECT 69.945 181.205 70.605 181.375 ;
        RECT 70.915 181.255 71.110 181.545 ;
        RECT 72.380 181.375 72.550 182.275 ;
        RECT 72.720 181.545 72.985 182.105 ;
        RECT 73.275 182.045 73.890 182.615 ;
        RECT 74.095 182.240 79.440 182.785 ;
        RECT 73.235 181.375 73.405 181.875 ;
        RECT 70.435 181.085 70.605 181.205 ;
        RECT 71.280 181.085 71.605 181.375 ;
        RECT 69.985 180.235 70.265 181.035 ;
        RECT 70.435 180.915 71.605 181.085 ;
        RECT 71.980 181.205 73.405 181.375 ;
        RECT 71.980 181.030 72.370 181.205 ;
        RECT 70.435 180.455 71.625 180.745 ;
        RECT 72.855 180.235 73.185 181.035 ;
        RECT 73.575 181.025 73.890 182.045 ;
        RECT 75.680 181.410 76.020 182.240 ;
        RECT 79.705 182.235 79.875 182.525 ;
        RECT 80.045 182.405 80.375 182.785 ;
        RECT 79.705 182.065 80.370 182.235 ;
        RECT 73.355 180.405 73.890 181.025 ;
        RECT 77.500 180.670 77.850 181.920 ;
        RECT 79.620 181.245 79.970 181.895 ;
        RECT 80.140 181.075 80.370 182.065 ;
        RECT 79.705 180.905 80.370 181.075 ;
        RECT 74.095 180.235 79.440 180.670 ;
        RECT 79.705 180.405 79.875 180.905 ;
        RECT 80.045 180.235 80.375 180.735 ;
        RECT 80.545 180.405 80.730 182.525 ;
        RECT 80.985 182.325 81.235 182.785 ;
        RECT 81.405 182.335 81.740 182.505 ;
        RECT 81.935 182.335 82.610 182.505 ;
        RECT 81.405 182.195 81.575 182.335 ;
        RECT 80.900 181.205 81.180 182.155 ;
        RECT 81.350 182.065 81.575 182.195 ;
        RECT 81.350 180.960 81.520 182.065 ;
        RECT 81.745 181.915 82.270 182.135 ;
        RECT 81.690 181.150 81.930 181.745 ;
        RECT 82.100 181.215 82.270 181.915 ;
        RECT 82.440 181.555 82.610 182.335 ;
        RECT 82.930 182.285 83.300 182.785 ;
        RECT 83.480 182.335 83.885 182.505 ;
        RECT 84.055 182.335 84.840 182.505 ;
        RECT 83.480 182.105 83.650 182.335 ;
        RECT 82.820 181.805 83.650 182.105 ;
        RECT 84.035 181.835 84.500 182.165 ;
        RECT 82.820 181.775 83.020 181.805 ;
        RECT 83.140 181.555 83.310 181.625 ;
        RECT 82.440 181.385 83.310 181.555 ;
        RECT 82.800 181.295 83.310 181.385 ;
        RECT 81.350 180.830 81.655 180.960 ;
        RECT 82.100 180.850 82.630 181.215 ;
        RECT 80.970 180.235 81.235 180.695 ;
        RECT 81.405 180.405 81.655 180.830 ;
        RECT 82.800 180.680 82.970 181.295 ;
        RECT 81.865 180.510 82.970 180.680 ;
        RECT 83.140 180.235 83.310 181.035 ;
        RECT 83.480 180.735 83.650 181.805 ;
        RECT 83.820 180.905 84.010 181.625 ;
        RECT 84.180 180.875 84.500 181.835 ;
        RECT 84.670 181.875 84.840 182.335 ;
        RECT 85.115 182.255 85.325 182.785 ;
        RECT 85.585 182.045 85.915 182.570 ;
        RECT 86.085 182.175 86.255 182.785 ;
        RECT 86.425 182.130 86.755 182.565 ;
        RECT 86.425 182.045 86.805 182.130 ;
        RECT 85.715 181.875 85.915 182.045 ;
        RECT 86.580 182.005 86.805 182.045 ;
        RECT 84.670 181.545 85.545 181.875 ;
        RECT 85.715 181.545 86.465 181.875 ;
        RECT 83.480 180.405 83.730 180.735 ;
        RECT 84.670 180.705 84.840 181.545 ;
        RECT 85.715 181.340 85.905 181.545 ;
        RECT 86.635 181.425 86.805 182.005 ;
        RECT 86.975 182.015 90.485 182.785 ;
        RECT 86.975 181.495 88.625 182.015 ;
        RECT 90.655 181.985 90.995 182.615 ;
        RECT 91.165 181.985 91.415 182.785 ;
        RECT 91.605 182.135 91.935 182.615 ;
        RECT 92.105 182.325 92.330 182.785 ;
        RECT 92.500 182.135 92.830 182.615 ;
        RECT 86.590 181.375 86.805 181.425 ;
        RECT 85.010 180.965 85.905 181.340 ;
        RECT 86.415 181.295 86.805 181.375 ;
        RECT 88.795 181.325 90.485 181.845 ;
        RECT 83.955 180.535 84.840 180.705 ;
        RECT 85.020 180.235 85.335 180.735 ;
        RECT 85.565 180.405 85.905 180.965 ;
        RECT 86.075 180.235 86.245 181.245 ;
        RECT 86.415 180.450 86.745 181.295 ;
        RECT 86.975 180.235 90.485 181.325 ;
        RECT 90.655 181.375 90.830 181.985 ;
        RECT 91.605 181.965 92.830 182.135 ;
        RECT 93.460 182.005 93.960 182.615 ;
        RECT 94.795 182.060 95.085 182.785 ;
        RECT 95.800 182.215 95.975 182.615 ;
        RECT 96.145 182.405 96.475 182.785 ;
        RECT 96.720 182.285 96.950 182.615 ;
        RECT 95.800 182.045 96.430 182.215 ;
        RECT 91.000 181.625 91.695 181.795 ;
        RECT 91.525 181.375 91.695 181.625 ;
        RECT 91.870 181.595 92.290 181.795 ;
        RECT 92.460 181.595 92.790 181.795 ;
        RECT 92.960 181.595 93.290 181.795 ;
        RECT 93.460 181.375 93.630 182.005 ;
        RECT 96.260 181.875 96.430 182.045 ;
        RECT 93.815 181.545 94.165 181.795 ;
        RECT 90.655 180.405 90.995 181.375 ;
        RECT 91.165 180.235 91.335 181.375 ;
        RECT 91.525 181.205 93.960 181.375 ;
        RECT 91.605 180.235 91.855 181.035 ;
        RECT 92.500 180.405 92.830 181.205 ;
        RECT 93.130 180.235 93.460 181.035 ;
        RECT 93.630 180.405 93.960 181.205 ;
        RECT 94.795 180.235 95.085 181.400 ;
        RECT 95.715 181.195 96.080 181.875 ;
        RECT 96.260 181.545 96.610 181.875 ;
        RECT 96.260 181.025 96.430 181.545 ;
        RECT 95.800 180.855 96.430 181.025 ;
        RECT 96.780 180.995 96.950 182.285 ;
        RECT 97.150 181.175 97.430 182.450 ;
        RECT 97.655 182.105 97.925 182.450 ;
        RECT 98.385 182.405 98.715 182.785 ;
        RECT 98.885 182.530 99.220 182.575 ;
        RECT 97.615 181.935 97.925 182.105 ;
        RECT 97.655 181.175 97.925 181.935 ;
        RECT 98.115 181.175 98.455 182.205 ;
        RECT 98.885 182.065 99.225 182.530 ;
        RECT 98.625 181.545 98.885 181.875 ;
        RECT 98.625 180.995 98.795 181.545 ;
        RECT 99.055 181.375 99.225 182.065 ;
        RECT 99.395 181.965 99.655 182.785 ;
        RECT 99.825 181.965 100.155 182.385 ;
        RECT 100.335 182.300 101.125 182.565 ;
        RECT 99.905 181.875 100.155 181.965 ;
        RECT 95.800 180.405 95.975 180.855 ;
        RECT 96.780 180.825 98.795 180.995 ;
        RECT 96.145 180.235 96.475 180.675 ;
        RECT 96.780 180.405 96.950 180.825 ;
        RECT 97.185 180.235 97.855 180.645 ;
        RECT 98.070 180.405 98.240 180.825 ;
        RECT 98.440 180.235 98.770 180.645 ;
        RECT 98.965 180.405 99.225 181.375 ;
        RECT 99.395 180.915 99.735 181.795 ;
        RECT 99.905 181.625 100.700 181.875 ;
        RECT 99.395 180.235 99.655 180.745 ;
        RECT 99.905 180.405 100.075 181.625 ;
        RECT 100.870 181.445 101.125 182.300 ;
        RECT 101.295 182.145 101.495 182.565 ;
        RECT 101.685 182.325 102.015 182.785 ;
        RECT 101.295 181.625 101.705 182.145 ;
        RECT 102.185 182.135 102.445 182.615 ;
        RECT 101.875 181.445 102.105 181.875 ;
        RECT 100.315 181.275 102.105 181.445 ;
        RECT 100.315 180.910 100.565 181.275 ;
        RECT 100.735 180.915 101.065 181.105 ;
        RECT 101.285 180.980 102.000 181.275 ;
        RECT 102.275 181.105 102.445 182.135 ;
        RECT 100.735 180.740 100.930 180.915 ;
        RECT 100.315 180.235 100.930 180.740 ;
        RECT 101.100 180.405 101.575 180.745 ;
        RECT 101.745 180.235 101.960 180.780 ;
        RECT 102.170 180.405 102.445 181.105 ;
        RECT 102.615 182.285 102.875 182.615 ;
        RECT 103.045 182.425 103.375 182.785 ;
        RECT 103.630 182.405 104.930 182.615 ;
        RECT 102.615 182.275 102.845 182.285 ;
        RECT 102.615 181.085 102.785 182.275 ;
        RECT 103.630 182.255 103.800 182.405 ;
        RECT 103.045 182.130 103.800 182.255 ;
        RECT 102.955 182.085 103.800 182.130 ;
        RECT 102.955 181.965 103.225 182.085 ;
        RECT 102.955 181.390 103.125 181.965 ;
        RECT 103.355 181.525 103.765 181.830 ;
        RECT 104.055 181.795 104.265 182.195 ;
        RECT 103.935 181.585 104.265 181.795 ;
        RECT 104.510 181.795 104.730 182.195 ;
        RECT 105.205 182.020 105.660 182.785 ;
        RECT 105.835 181.840 106.175 182.615 ;
        RECT 106.345 182.325 106.515 182.785 ;
        RECT 106.755 182.350 107.115 182.615 ;
        RECT 106.755 182.345 107.110 182.350 ;
        RECT 106.755 182.335 107.105 182.345 ;
        RECT 106.755 182.330 107.100 182.335 ;
        RECT 106.755 182.320 107.095 182.330 ;
        RECT 107.745 182.325 107.915 182.785 ;
        RECT 106.755 182.315 107.090 182.320 ;
        RECT 106.755 182.305 107.080 182.315 ;
        RECT 106.755 182.295 107.070 182.305 ;
        RECT 106.755 182.155 107.055 182.295 ;
        RECT 106.345 181.965 107.055 182.155 ;
        RECT 107.245 182.155 107.575 182.235 ;
        RECT 108.085 182.155 108.425 182.615 ;
        RECT 107.245 181.965 108.425 182.155 ;
        RECT 108.595 182.155 108.935 182.615 ;
        RECT 109.105 182.325 109.275 182.785 ;
        RECT 109.445 182.405 110.615 182.615 ;
        RECT 109.445 182.155 109.695 182.405 ;
        RECT 110.285 182.385 110.615 182.405 ;
        RECT 108.595 181.985 109.695 182.155 ;
        RECT 109.865 181.965 110.725 182.215 ;
        RECT 104.510 181.585 104.985 181.795 ;
        RECT 105.175 181.595 105.665 181.795 ;
        RECT 102.955 181.355 103.155 181.390 ;
        RECT 104.485 181.355 105.660 181.415 ;
        RECT 102.955 181.245 105.660 181.355 ;
        RECT 103.015 181.185 104.815 181.245 ;
        RECT 104.485 181.155 104.815 181.185 ;
        RECT 102.615 180.405 102.875 181.085 ;
        RECT 103.045 180.235 103.295 181.015 ;
        RECT 103.545 180.985 104.380 180.995 ;
        RECT 104.970 180.985 105.155 181.075 ;
        RECT 103.545 180.785 105.155 180.985 ;
        RECT 103.545 180.405 103.795 180.785 ;
        RECT 104.925 180.745 105.155 180.785 ;
        RECT 105.405 180.625 105.660 181.245 ;
        RECT 103.965 180.235 104.320 180.615 ;
        RECT 105.325 180.405 105.660 180.625 ;
        RECT 105.835 180.405 106.115 181.840 ;
        RECT 106.345 181.395 106.630 181.965 ;
        RECT 106.815 181.565 107.285 181.795 ;
        RECT 107.455 181.775 107.785 181.795 ;
        RECT 107.455 181.595 107.905 181.775 ;
        RECT 108.095 181.595 108.425 181.795 ;
        RECT 106.345 181.180 107.495 181.395 ;
        RECT 106.285 180.235 106.995 181.010 ;
        RECT 107.165 180.405 107.495 181.180 ;
        RECT 107.690 180.480 107.905 181.595 ;
        RECT 108.195 181.255 108.425 181.595 ;
        RECT 108.595 181.545 109.355 181.795 ;
        RECT 109.525 181.545 110.275 181.795 ;
        RECT 110.445 181.375 110.725 181.965 ;
        RECT 108.085 180.235 108.415 180.955 ;
        RECT 108.595 180.235 108.855 181.375 ;
        RECT 109.025 181.205 110.725 181.375 ;
        RECT 110.895 182.135 111.155 182.615 ;
        RECT 111.325 182.245 111.575 182.785 ;
        RECT 109.025 180.405 109.355 181.205 ;
        RECT 109.525 180.235 109.695 181.035 ;
        RECT 109.865 180.405 110.195 181.205 ;
        RECT 110.895 181.105 111.065 182.135 ;
        RECT 111.745 182.080 111.965 182.565 ;
        RECT 111.235 181.485 111.465 181.880 ;
        RECT 111.635 181.655 111.965 182.080 ;
        RECT 112.135 182.405 113.025 182.575 ;
        RECT 114.115 182.405 115.005 182.575 ;
        RECT 112.135 181.680 112.305 182.405 ;
        RECT 112.475 181.850 113.025 182.235 ;
        RECT 114.115 181.850 114.665 182.235 ;
        RECT 114.835 181.680 115.005 182.405 ;
        RECT 112.135 181.610 113.025 181.680 ;
        RECT 112.130 181.585 113.025 181.610 ;
        RECT 112.120 181.570 113.025 181.585 ;
        RECT 112.115 181.555 113.025 181.570 ;
        RECT 112.105 181.550 113.025 181.555 ;
        RECT 112.100 181.540 113.025 181.550 ;
        RECT 112.095 181.530 113.025 181.540 ;
        RECT 112.085 181.525 113.025 181.530 ;
        RECT 112.075 181.515 113.025 181.525 ;
        RECT 112.065 181.510 113.025 181.515 ;
        RECT 112.065 181.505 112.400 181.510 ;
        RECT 112.050 181.500 112.400 181.505 ;
        RECT 112.035 181.490 112.400 181.500 ;
        RECT 112.010 181.485 112.400 181.490 ;
        RECT 111.235 181.480 112.400 181.485 ;
        RECT 111.235 181.445 112.370 181.480 ;
        RECT 111.235 181.420 112.335 181.445 ;
        RECT 111.235 181.390 112.305 181.420 ;
        RECT 111.235 181.360 112.285 181.390 ;
        RECT 111.235 181.330 112.265 181.360 ;
        RECT 111.235 181.320 112.195 181.330 ;
        RECT 111.235 181.310 112.170 181.320 ;
        RECT 111.235 181.295 112.150 181.310 ;
        RECT 111.235 181.280 112.130 181.295 ;
        RECT 111.340 181.270 112.125 181.280 ;
        RECT 111.340 181.235 112.110 181.270 ;
        RECT 110.365 180.235 110.620 181.035 ;
        RECT 110.895 180.405 111.170 181.105 ;
        RECT 111.340 180.985 112.095 181.235 ;
        RECT 112.265 180.915 112.595 181.160 ;
        RECT 112.765 181.060 113.025 181.510 ;
        RECT 114.115 181.610 115.005 181.680 ;
        RECT 115.175 182.080 115.395 182.565 ;
        RECT 115.565 182.245 115.815 182.785 ;
        RECT 115.985 182.135 116.245 182.615 ;
        RECT 115.175 181.655 115.505 182.080 ;
        RECT 114.115 181.585 115.010 181.610 ;
        RECT 114.115 181.570 115.020 181.585 ;
        RECT 114.115 181.555 115.025 181.570 ;
        RECT 114.115 181.550 115.035 181.555 ;
        RECT 114.115 181.540 115.040 181.550 ;
        RECT 114.115 181.530 115.045 181.540 ;
        RECT 114.115 181.525 115.055 181.530 ;
        RECT 114.115 181.515 115.065 181.525 ;
        RECT 114.115 181.510 115.075 181.515 ;
        RECT 114.115 181.060 114.375 181.510 ;
        RECT 114.740 181.505 115.075 181.510 ;
        RECT 114.740 181.500 115.090 181.505 ;
        RECT 114.740 181.490 115.105 181.500 ;
        RECT 114.740 181.485 115.130 181.490 ;
        RECT 115.675 181.485 115.905 181.880 ;
        RECT 114.740 181.480 115.905 181.485 ;
        RECT 114.770 181.445 115.905 181.480 ;
        RECT 114.805 181.420 115.905 181.445 ;
        RECT 114.835 181.390 115.905 181.420 ;
        RECT 114.855 181.360 115.905 181.390 ;
        RECT 114.875 181.330 115.905 181.360 ;
        RECT 114.945 181.320 115.905 181.330 ;
        RECT 114.970 181.310 115.905 181.320 ;
        RECT 114.990 181.295 115.905 181.310 ;
        RECT 115.010 181.280 115.905 181.295 ;
        RECT 115.015 181.270 115.800 181.280 ;
        RECT 115.030 181.235 115.800 181.270 ;
        RECT 112.410 180.890 112.595 180.915 ;
        RECT 114.545 180.915 114.875 181.160 ;
        RECT 115.045 180.985 115.800 181.235 ;
        RECT 116.075 181.105 116.245 182.135 ;
        RECT 116.415 181.965 116.675 182.785 ;
        RECT 116.845 181.965 117.175 182.385 ;
        RECT 117.355 182.300 118.145 182.565 ;
        RECT 116.925 181.875 117.175 181.965 ;
        RECT 114.545 180.890 114.730 180.915 ;
        RECT 112.410 180.790 113.025 180.890 ;
        RECT 111.340 180.235 111.595 180.780 ;
        RECT 111.765 180.405 112.245 180.745 ;
        RECT 112.420 180.235 113.025 180.790 ;
        RECT 114.115 180.790 114.730 180.890 ;
        RECT 114.115 180.235 114.720 180.790 ;
        RECT 114.895 180.405 115.375 180.745 ;
        RECT 115.545 180.235 115.800 180.780 ;
        RECT 115.970 180.405 116.245 181.105 ;
        RECT 116.415 180.915 116.755 181.795 ;
        RECT 116.925 181.625 117.720 181.875 ;
        RECT 116.415 180.235 116.675 180.745 ;
        RECT 116.925 180.405 117.095 181.625 ;
        RECT 117.890 181.445 118.145 182.300 ;
        RECT 118.315 182.145 118.515 182.565 ;
        RECT 118.705 182.325 119.035 182.785 ;
        RECT 118.315 181.625 118.725 182.145 ;
        RECT 119.205 182.135 119.465 182.615 ;
        RECT 118.895 181.445 119.125 181.875 ;
        RECT 117.335 181.275 119.125 181.445 ;
        RECT 117.335 180.910 117.585 181.275 ;
        RECT 117.755 180.915 118.085 181.105 ;
        RECT 118.305 180.980 119.020 181.275 ;
        RECT 119.295 181.105 119.465 182.135 ;
        RECT 120.555 182.060 120.845 182.785 ;
        RECT 121.015 182.240 126.360 182.785 ;
        RECT 122.600 181.410 122.940 182.240 ;
        RECT 126.535 182.015 128.205 182.785 ;
        RECT 128.925 182.235 129.095 182.525 ;
        RECT 129.265 182.405 129.595 182.785 ;
        RECT 128.925 182.065 129.590 182.235 ;
        RECT 117.755 180.740 117.950 180.915 ;
        RECT 117.335 180.235 117.950 180.740 ;
        RECT 118.120 180.405 118.595 180.745 ;
        RECT 118.765 180.235 118.980 180.780 ;
        RECT 119.190 180.405 119.465 181.105 ;
        RECT 120.555 180.235 120.845 181.400 ;
        RECT 124.420 180.670 124.770 181.920 ;
        RECT 126.535 181.495 127.285 182.015 ;
        RECT 127.455 181.325 128.205 181.845 ;
        RECT 121.015 180.235 126.360 180.670 ;
        RECT 126.535 180.235 128.205 181.325 ;
        RECT 128.840 181.245 129.190 181.895 ;
        RECT 129.360 181.075 129.590 182.065 ;
        RECT 128.925 180.905 129.590 181.075 ;
        RECT 128.925 180.405 129.095 180.905 ;
        RECT 129.265 180.235 129.595 180.735 ;
        RECT 129.765 180.405 129.950 182.525 ;
        RECT 130.205 182.325 130.455 182.785 ;
        RECT 130.625 182.335 130.960 182.505 ;
        RECT 131.155 182.335 131.830 182.505 ;
        RECT 130.625 182.195 130.795 182.335 ;
        RECT 130.120 181.205 130.400 182.155 ;
        RECT 130.570 182.065 130.795 182.195 ;
        RECT 130.570 180.960 130.740 182.065 ;
        RECT 130.965 181.915 131.490 182.135 ;
        RECT 130.910 181.150 131.150 181.745 ;
        RECT 131.320 181.215 131.490 181.915 ;
        RECT 131.660 181.555 131.830 182.335 ;
        RECT 132.150 182.285 132.520 182.785 ;
        RECT 132.700 182.335 133.105 182.505 ;
        RECT 133.275 182.335 134.060 182.505 ;
        RECT 132.700 182.105 132.870 182.335 ;
        RECT 132.040 181.805 132.870 182.105 ;
        RECT 133.255 181.835 133.720 182.165 ;
        RECT 132.040 181.775 132.240 181.805 ;
        RECT 132.360 181.555 132.530 181.625 ;
        RECT 131.660 181.385 132.530 181.555 ;
        RECT 132.020 181.295 132.530 181.385 ;
        RECT 130.570 180.830 130.875 180.960 ;
        RECT 131.320 180.850 131.850 181.215 ;
        RECT 130.190 180.235 130.455 180.695 ;
        RECT 130.625 180.405 130.875 180.830 ;
        RECT 132.020 180.680 132.190 181.295 ;
        RECT 131.085 180.510 132.190 180.680 ;
        RECT 132.360 180.235 132.530 181.035 ;
        RECT 132.700 180.735 132.870 181.805 ;
        RECT 133.040 180.905 133.230 181.625 ;
        RECT 133.400 180.875 133.720 181.835 ;
        RECT 133.890 181.875 134.060 182.335 ;
        RECT 134.335 182.255 134.545 182.785 ;
        RECT 134.805 182.045 135.135 182.570 ;
        RECT 135.305 182.175 135.475 182.785 ;
        RECT 135.645 182.130 135.975 182.565 ;
        RECT 135.645 182.045 136.025 182.130 ;
        RECT 134.935 181.875 135.135 182.045 ;
        RECT 135.800 182.005 136.025 182.045 ;
        RECT 133.890 181.545 134.765 181.875 ;
        RECT 134.935 181.545 135.685 181.875 ;
        RECT 132.700 180.405 132.950 180.735 ;
        RECT 133.890 180.705 134.060 181.545 ;
        RECT 134.935 181.340 135.125 181.545 ;
        RECT 135.855 181.425 136.025 182.005 ;
        RECT 135.810 181.375 136.025 181.425 ;
        RECT 134.230 180.965 135.125 181.340 ;
        RECT 135.635 181.295 136.025 181.375 ;
        RECT 136.195 182.045 136.580 182.615 ;
        RECT 136.750 182.325 137.075 182.785 ;
        RECT 137.595 182.155 137.875 182.615 ;
        RECT 136.195 181.375 136.475 182.045 ;
        RECT 136.750 181.985 137.875 182.155 ;
        RECT 136.750 181.875 137.200 181.985 ;
        RECT 136.645 181.545 137.200 181.875 ;
        RECT 138.065 181.815 138.465 182.615 ;
        RECT 138.865 182.325 139.135 182.785 ;
        RECT 139.305 182.155 139.590 182.615 ;
        RECT 133.175 180.535 134.060 180.705 ;
        RECT 134.240 180.235 134.555 180.735 ;
        RECT 134.785 180.405 135.125 180.965 ;
        RECT 135.295 180.235 135.465 181.245 ;
        RECT 135.635 180.450 135.965 181.295 ;
        RECT 136.195 180.405 136.580 181.375 ;
        RECT 136.750 181.085 137.200 181.545 ;
        RECT 137.370 181.255 138.465 181.815 ;
        RECT 136.750 180.865 137.875 181.085 ;
        RECT 136.750 180.235 137.075 180.695 ;
        RECT 137.595 180.405 137.875 180.865 ;
        RECT 138.065 180.405 138.465 181.255 ;
        RECT 138.635 181.985 139.590 182.155 ;
        RECT 139.965 182.235 140.135 182.615 ;
        RECT 140.350 182.405 140.680 182.785 ;
        RECT 139.965 182.065 140.680 182.235 ;
        RECT 138.635 181.085 138.845 181.985 ;
        RECT 139.015 181.255 139.705 181.815 ;
        RECT 139.875 181.515 140.230 181.885 ;
        RECT 140.510 181.875 140.680 182.065 ;
        RECT 140.850 182.040 141.105 182.615 ;
        RECT 140.510 181.545 140.765 181.875 ;
        RECT 140.510 181.335 140.680 181.545 ;
        RECT 139.965 181.165 140.680 181.335 ;
        RECT 140.935 181.310 141.105 182.040 ;
        RECT 141.280 181.945 141.540 182.785 ;
        RECT 141.715 182.035 142.925 182.785 ;
        RECT 138.635 180.865 139.590 181.085 ;
        RECT 138.865 180.235 139.135 180.695 ;
        RECT 139.305 180.405 139.590 180.865 ;
        RECT 139.965 180.405 140.135 181.165 ;
        RECT 140.350 180.235 140.680 180.995 ;
        RECT 140.850 180.405 141.105 181.310 ;
        RECT 141.280 180.235 141.540 181.385 ;
        RECT 141.715 181.325 142.235 181.865 ;
        RECT 142.405 181.495 142.925 182.035 ;
        RECT 141.715 180.235 142.925 181.325 ;
        RECT 17.430 180.065 143.010 180.235 ;
        RECT 17.515 178.975 18.725 180.065 ;
        RECT 18.895 178.975 22.405 180.065 ;
        RECT 17.515 178.265 18.035 178.805 ;
        RECT 18.205 178.435 18.725 178.975 ;
        RECT 18.895 178.285 20.545 178.805 ;
        RECT 20.715 178.455 22.405 178.975 ;
        RECT 22.575 178.925 22.835 179.895 ;
        RECT 23.030 179.655 23.360 180.065 ;
        RECT 23.560 179.475 23.730 179.895 ;
        RECT 23.945 179.655 24.615 180.065 ;
        RECT 24.850 179.475 25.020 179.895 ;
        RECT 25.325 179.625 25.655 180.065 ;
        RECT 23.005 179.305 25.020 179.475 ;
        RECT 25.825 179.445 26.000 179.895 ;
        RECT 17.515 177.515 18.725 178.265 ;
        RECT 18.895 177.515 22.405 178.285 ;
        RECT 22.575 178.235 22.745 178.925 ;
        RECT 23.005 178.755 23.175 179.305 ;
        RECT 22.915 178.425 23.175 178.755 ;
        RECT 22.575 177.770 22.915 178.235 ;
        RECT 23.345 178.095 23.685 179.125 ;
        RECT 23.875 178.705 24.145 179.125 ;
        RECT 23.875 178.535 24.185 178.705 ;
        RECT 22.580 177.725 22.915 177.770 ;
        RECT 23.085 177.515 23.415 177.895 ;
        RECT 23.875 177.850 24.145 178.535 ;
        RECT 24.370 177.850 24.650 179.125 ;
        RECT 24.850 178.015 25.020 179.305 ;
        RECT 25.370 179.275 26.000 179.445 ;
        RECT 25.370 178.755 25.540 179.275 ;
        RECT 25.190 178.425 25.540 178.755 ;
        RECT 25.720 178.425 26.085 179.105 ;
        RECT 26.255 178.975 29.765 180.065 ;
        RECT 25.370 178.255 25.540 178.425 ;
        RECT 26.255 178.285 27.905 178.805 ;
        RECT 28.075 178.455 29.765 178.975 ;
        RECT 30.395 178.900 30.685 180.065 ;
        RECT 30.855 178.975 34.365 180.065 ;
        RECT 30.855 178.285 32.505 178.805 ;
        RECT 32.675 178.455 34.365 178.975 ;
        RECT 35.005 178.925 35.335 180.065 ;
        RECT 35.865 179.095 36.195 179.880 ;
        RECT 35.515 178.925 36.195 179.095 ;
        RECT 36.385 179.115 36.660 179.885 ;
        RECT 36.830 179.455 37.160 179.885 ;
        RECT 37.330 179.625 37.525 180.065 ;
        RECT 37.705 179.455 38.035 179.885 ;
        RECT 38.220 179.685 38.555 180.065 ;
        RECT 36.830 179.285 38.035 179.455 ;
        RECT 36.385 178.925 36.970 179.115 ;
        RECT 37.140 178.955 38.035 179.285 ;
        RECT 34.995 178.505 35.345 178.755 ;
        RECT 35.515 178.325 35.685 178.925 ;
        RECT 35.855 178.505 36.205 178.755 ;
        RECT 25.370 178.085 26.000 178.255 ;
        RECT 24.850 177.685 25.080 178.015 ;
        RECT 25.325 177.515 25.655 177.895 ;
        RECT 25.825 177.685 26.000 178.085 ;
        RECT 26.255 177.515 29.765 178.285 ;
        RECT 30.395 177.515 30.685 178.240 ;
        RECT 30.855 177.515 34.365 178.285 ;
        RECT 35.005 177.515 35.275 178.325 ;
        RECT 35.445 177.685 35.775 178.325 ;
        RECT 35.945 177.515 36.185 178.325 ;
        RECT 36.385 178.105 36.625 178.755 ;
        RECT 36.795 178.255 36.970 178.925 ;
        RECT 37.140 178.425 37.555 178.755 ;
        RECT 37.735 178.425 38.030 178.755 ;
        RECT 36.795 178.075 37.125 178.255 ;
        RECT 36.400 177.515 36.730 177.905 ;
        RECT 36.900 177.695 37.125 178.075 ;
        RECT 37.325 177.805 37.555 178.425 ;
        RECT 37.735 177.515 38.035 178.245 ;
        RECT 38.215 178.195 38.455 179.505 ;
        RECT 38.725 179.095 38.975 179.895 ;
        RECT 39.195 179.345 39.525 180.065 ;
        RECT 39.710 179.095 39.960 179.895 ;
        RECT 40.425 179.265 40.755 180.065 ;
        RECT 40.925 179.635 41.265 179.895 ;
        RECT 38.625 178.925 40.815 179.095 ;
        RECT 38.625 178.015 38.795 178.925 ;
        RECT 40.500 178.755 40.815 178.925 ;
        RECT 38.300 177.685 38.795 178.015 ;
        RECT 39.015 177.790 39.365 178.755 ;
        RECT 39.545 177.785 39.845 178.755 ;
        RECT 40.025 177.785 40.305 178.755 ;
        RECT 40.500 178.505 40.830 178.755 ;
        RECT 40.485 177.515 40.755 178.315 ;
        RECT 41.005 178.235 41.265 179.635 ;
        RECT 41.445 178.925 41.775 180.065 ;
        RECT 42.305 179.095 42.635 179.880 ;
        RECT 41.955 178.925 42.635 179.095 ;
        RECT 42.825 179.095 43.155 179.880 ;
        RECT 42.825 178.925 43.505 179.095 ;
        RECT 43.685 178.925 44.015 180.065 ;
        RECT 44.195 179.630 49.540 180.065 ;
        RECT 41.435 178.505 41.785 178.755 ;
        RECT 41.955 178.325 42.125 178.925 ;
        RECT 42.295 178.505 42.645 178.755 ;
        RECT 42.815 178.505 43.165 178.755 ;
        RECT 43.335 178.325 43.505 178.925 ;
        RECT 43.675 178.505 44.025 178.755 ;
        RECT 40.925 177.725 41.265 178.235 ;
        RECT 41.445 177.515 41.715 178.325 ;
        RECT 41.885 177.685 42.215 178.325 ;
        RECT 42.385 177.515 42.625 178.325 ;
        RECT 42.835 177.515 43.075 178.325 ;
        RECT 43.245 177.685 43.575 178.325 ;
        RECT 43.745 177.515 44.015 178.325 ;
        RECT 45.780 178.060 46.120 178.890 ;
        RECT 47.600 178.380 47.950 179.630 ;
        RECT 49.800 179.445 49.975 179.895 ;
        RECT 50.145 179.625 50.475 180.065 ;
        RECT 50.780 179.475 50.950 179.895 ;
        RECT 51.185 179.655 51.855 180.065 ;
        RECT 52.070 179.475 52.240 179.895 ;
        RECT 52.440 179.655 52.770 180.065 ;
        RECT 49.800 179.275 50.430 179.445 ;
        RECT 49.715 178.425 50.080 179.105 ;
        RECT 50.260 178.755 50.430 179.275 ;
        RECT 50.780 179.305 52.795 179.475 ;
        RECT 50.260 178.425 50.610 178.755 ;
        RECT 50.260 178.255 50.430 178.425 ;
        RECT 49.800 178.085 50.430 178.255 ;
        RECT 44.195 177.515 49.540 178.060 ;
        RECT 49.800 177.685 49.975 178.085 ;
        RECT 50.780 178.015 50.950 179.305 ;
        RECT 50.145 177.515 50.475 177.895 ;
        RECT 50.720 177.685 50.950 178.015 ;
        RECT 51.150 177.850 51.430 179.125 ;
        RECT 51.655 178.025 51.925 179.125 ;
        RECT 52.115 178.095 52.455 179.125 ;
        RECT 52.625 178.755 52.795 179.305 ;
        RECT 52.965 178.925 53.225 179.895 ;
        RECT 53.405 179.095 53.735 179.880 ;
        RECT 53.405 178.925 54.085 179.095 ;
        RECT 54.265 178.925 54.595 180.065 ;
        RECT 54.775 178.975 55.985 180.065 ;
        RECT 52.625 178.425 52.885 178.755 ;
        RECT 53.055 178.235 53.225 178.925 ;
        RECT 53.395 178.505 53.745 178.755 ;
        RECT 53.915 178.325 54.085 178.925 ;
        RECT 54.255 178.505 54.605 178.755 ;
        RECT 51.615 177.855 51.925 178.025 ;
        RECT 51.655 177.850 51.925 177.855 ;
        RECT 52.385 177.515 52.715 177.895 ;
        RECT 52.885 177.770 53.225 178.235 ;
        RECT 52.885 177.725 53.220 177.770 ;
        RECT 53.415 177.515 53.655 178.325 ;
        RECT 53.825 177.685 54.155 178.325 ;
        RECT 54.325 177.515 54.595 178.325 ;
        RECT 54.775 178.265 55.295 178.805 ;
        RECT 55.465 178.435 55.985 178.975 ;
        RECT 56.155 178.900 56.445 180.065 ;
        RECT 56.615 179.630 61.960 180.065 ;
        RECT 54.775 177.515 55.985 178.265 ;
        RECT 56.155 177.515 56.445 178.240 ;
        RECT 58.200 178.060 58.540 178.890 ;
        RECT 60.020 178.380 60.370 179.630 ;
        RECT 63.065 179.005 63.395 179.855 ;
        RECT 63.065 178.240 63.255 179.005 ;
        RECT 63.565 178.925 63.815 180.065 ;
        RECT 64.005 179.425 64.255 179.845 ;
        RECT 64.485 179.595 64.815 180.065 ;
        RECT 65.045 179.425 65.295 179.845 ;
        RECT 64.005 179.255 65.295 179.425 ;
        RECT 65.475 179.425 65.805 179.855 ;
        RECT 65.475 179.255 65.930 179.425 ;
        RECT 63.995 178.755 64.210 179.085 ;
        RECT 63.425 178.425 63.735 178.755 ;
        RECT 63.905 178.425 64.210 178.755 ;
        RECT 64.385 178.425 64.670 179.085 ;
        RECT 64.865 178.425 65.130 179.085 ;
        RECT 65.345 178.425 65.590 179.085 ;
        RECT 63.565 178.255 63.735 178.425 ;
        RECT 65.760 178.255 65.930 179.255 ;
        RECT 56.615 177.515 61.960 178.060 ;
        RECT 63.065 177.730 63.395 178.240 ;
        RECT 63.565 178.085 65.930 178.255 ;
        RECT 66.275 178.925 66.660 179.895 ;
        RECT 66.830 179.605 67.155 180.065 ;
        RECT 67.675 179.435 67.955 179.895 ;
        RECT 66.830 179.215 67.955 179.435 ;
        RECT 66.275 178.255 66.555 178.925 ;
        RECT 66.830 178.755 67.280 179.215 ;
        RECT 68.145 179.045 68.545 179.895 ;
        RECT 68.945 179.605 69.215 180.065 ;
        RECT 69.385 179.435 69.670 179.895 ;
        RECT 66.725 178.425 67.280 178.755 ;
        RECT 67.450 178.485 68.545 179.045 ;
        RECT 66.830 178.315 67.280 178.425 ;
        RECT 63.565 177.515 63.895 177.915 ;
        RECT 64.945 177.745 65.275 178.085 ;
        RECT 65.445 177.515 65.775 177.915 ;
        RECT 66.275 177.685 66.660 178.255 ;
        RECT 66.830 178.145 67.955 178.315 ;
        RECT 66.830 177.515 67.155 177.975 ;
        RECT 67.675 177.685 67.955 178.145 ;
        RECT 68.145 177.685 68.545 178.485 ;
        RECT 68.715 179.215 69.670 179.435 ;
        RECT 68.715 178.315 68.925 179.215 ;
        RECT 69.095 178.485 69.785 179.045 ;
        RECT 69.955 178.925 70.340 179.895 ;
        RECT 70.510 179.605 70.835 180.065 ;
        RECT 71.355 179.435 71.635 179.895 ;
        RECT 70.510 179.215 71.635 179.435 ;
        RECT 68.715 178.145 69.670 178.315 ;
        RECT 68.945 177.515 69.215 177.975 ;
        RECT 69.385 177.685 69.670 178.145 ;
        RECT 69.955 178.255 70.235 178.925 ;
        RECT 70.510 178.755 70.960 179.215 ;
        RECT 71.825 179.045 72.225 179.895 ;
        RECT 72.625 179.605 72.895 180.065 ;
        RECT 73.065 179.435 73.350 179.895 ;
        RECT 70.405 178.425 70.960 178.755 ;
        RECT 71.130 178.485 72.225 179.045 ;
        RECT 70.510 178.315 70.960 178.425 ;
        RECT 69.955 177.685 70.340 178.255 ;
        RECT 70.510 178.145 71.635 178.315 ;
        RECT 70.510 177.515 70.835 177.975 ;
        RECT 71.355 177.685 71.635 178.145 ;
        RECT 71.825 177.685 72.225 178.485 ;
        RECT 72.395 179.215 73.350 179.435 ;
        RECT 72.395 178.315 72.605 179.215 ;
        RECT 72.775 178.485 73.465 179.045 ;
        RECT 73.635 178.925 73.915 180.065 ;
        RECT 74.085 178.915 74.415 179.895 ;
        RECT 74.585 178.925 74.845 180.065 ;
        RECT 75.015 178.925 75.275 180.065 ;
        RECT 75.445 178.915 75.775 179.895 ;
        RECT 75.945 178.925 76.225 180.065 ;
        RECT 76.395 179.630 81.740 180.065 ;
        RECT 73.645 178.485 73.980 178.755 ;
        RECT 74.150 178.365 74.320 178.915 ;
        RECT 74.490 178.505 74.825 178.755 ;
        RECT 75.035 178.505 75.370 178.755 ;
        RECT 74.150 178.315 74.325 178.365 ;
        RECT 75.540 178.315 75.710 178.915 ;
        RECT 75.880 178.485 76.215 178.755 ;
        RECT 72.395 178.145 73.350 178.315 ;
        RECT 72.625 177.515 72.895 177.975 ;
        RECT 73.065 177.685 73.350 178.145 ;
        RECT 73.635 177.515 73.945 178.315 ;
        RECT 74.150 177.685 74.845 178.315 ;
        RECT 75.015 177.685 75.710 178.315 ;
        RECT 75.915 177.515 76.225 178.315 ;
        RECT 77.980 178.060 78.320 178.890 ;
        RECT 79.800 178.380 80.150 179.630 ;
        RECT 81.915 178.900 82.205 180.065 ;
        RECT 82.490 179.435 82.775 179.895 ;
        RECT 82.945 179.605 83.215 180.065 ;
        RECT 82.490 179.215 83.445 179.435 ;
        RECT 82.375 178.485 83.065 179.045 ;
        RECT 83.235 178.315 83.445 179.215 ;
        RECT 76.395 177.515 81.740 178.060 ;
        RECT 81.915 177.515 82.205 178.240 ;
        RECT 82.490 178.145 83.445 178.315 ;
        RECT 83.615 179.045 84.015 179.895 ;
        RECT 84.205 179.435 84.485 179.895 ;
        RECT 85.005 179.605 85.330 180.065 ;
        RECT 84.205 179.215 85.330 179.435 ;
        RECT 83.615 178.485 84.710 179.045 ;
        RECT 84.880 178.755 85.330 179.215 ;
        RECT 85.500 178.925 85.885 179.895 ;
        RECT 86.055 179.630 91.400 180.065 ;
        RECT 82.490 177.685 82.775 178.145 ;
        RECT 82.945 177.515 83.215 177.975 ;
        RECT 83.615 177.685 84.015 178.485 ;
        RECT 84.880 178.425 85.435 178.755 ;
        RECT 84.880 178.315 85.330 178.425 ;
        RECT 84.205 178.145 85.330 178.315 ;
        RECT 85.605 178.255 85.885 178.925 ;
        RECT 84.205 177.685 84.485 178.145 ;
        RECT 85.005 177.515 85.330 177.975 ;
        RECT 85.500 177.685 85.885 178.255 ;
        RECT 87.640 178.060 87.980 178.890 ;
        RECT 89.460 178.380 89.810 179.630 ;
        RECT 92.035 178.925 92.295 180.065 ;
        RECT 92.465 178.915 92.795 179.895 ;
        RECT 92.965 178.925 93.245 180.065 ;
        RECT 93.425 178.925 93.755 180.065 ;
        RECT 94.285 179.095 94.615 179.880 ;
        RECT 93.935 178.925 94.615 179.095 ;
        RECT 94.795 178.975 96.465 180.065 ;
        RECT 96.725 179.445 96.895 179.875 ;
        RECT 97.065 179.615 97.395 180.065 ;
        RECT 96.725 179.215 97.400 179.445 ;
        RECT 92.055 178.505 92.390 178.755 ;
        RECT 92.560 178.315 92.730 178.915 ;
        RECT 92.900 178.485 93.235 178.755 ;
        RECT 93.415 178.505 93.765 178.755 ;
        RECT 93.935 178.325 94.105 178.925 ;
        RECT 94.275 178.505 94.625 178.755 ;
        RECT 86.055 177.515 91.400 178.060 ;
        RECT 92.035 177.685 92.730 178.315 ;
        RECT 92.935 177.515 93.245 178.315 ;
        RECT 93.425 177.515 93.695 178.325 ;
        RECT 93.865 177.685 94.195 178.325 ;
        RECT 94.365 177.515 94.605 178.325 ;
        RECT 94.795 178.285 95.545 178.805 ;
        RECT 95.715 178.455 96.465 178.975 ;
        RECT 94.795 177.515 96.465 178.285 ;
        RECT 96.695 178.195 96.995 179.045 ;
        RECT 97.165 178.565 97.400 179.215 ;
        RECT 97.570 178.905 97.855 179.850 ;
        RECT 98.035 179.595 98.720 180.065 ;
        RECT 98.030 179.075 98.725 179.385 ;
        RECT 98.900 179.010 99.205 179.795 ;
        RECT 97.570 178.755 98.430 178.905 ;
        RECT 97.570 178.735 98.855 178.755 ;
        RECT 97.165 178.235 97.700 178.565 ;
        RECT 97.870 178.375 98.855 178.735 ;
        RECT 97.165 178.085 97.385 178.235 ;
        RECT 96.640 177.515 96.975 178.020 ;
        RECT 97.145 177.710 97.385 178.085 ;
        RECT 97.870 178.040 98.040 178.375 ;
        RECT 99.030 178.205 99.205 179.010 ;
        RECT 99.455 178.925 99.665 180.065 ;
        RECT 99.835 178.915 100.165 179.895 ;
        RECT 100.335 178.925 100.565 180.065 ;
        RECT 101.275 178.925 101.505 180.065 ;
        RECT 101.675 178.915 102.005 179.895 ;
        RECT 102.175 178.925 102.385 180.065 ;
        RECT 102.615 178.975 103.825 180.065 ;
        RECT 104.495 179.605 104.710 180.065 ;
        RECT 104.880 179.435 105.210 179.895 ;
        RECT 97.665 177.845 98.040 178.040 ;
        RECT 97.665 177.700 97.835 177.845 ;
        RECT 98.400 177.515 98.795 178.010 ;
        RECT 98.965 177.685 99.205 178.205 ;
        RECT 99.455 177.515 99.665 178.335 ;
        RECT 99.835 178.315 100.085 178.915 ;
        RECT 100.255 178.505 100.585 178.755 ;
        RECT 101.255 178.505 101.585 178.755 ;
        RECT 99.835 177.685 100.165 178.315 ;
        RECT 100.335 177.515 100.565 178.335 ;
        RECT 101.275 177.515 101.505 178.335 ;
        RECT 101.755 178.315 102.005 178.915 ;
        RECT 101.675 177.685 102.005 178.315 ;
        RECT 102.175 177.515 102.385 178.335 ;
        RECT 102.615 178.265 103.135 178.805 ;
        RECT 103.305 178.435 103.825 178.975 ;
        RECT 104.040 179.265 105.210 179.435 ;
        RECT 105.380 179.265 105.630 180.065 ;
        RECT 102.615 177.515 103.825 178.265 ;
        RECT 104.040 177.975 104.410 179.265 ;
        RECT 105.840 179.095 106.120 179.255 ;
        RECT 104.785 178.925 106.120 179.095 ;
        RECT 106.295 178.975 107.505 180.065 ;
        RECT 104.785 178.755 104.955 178.925 ;
        RECT 104.580 178.505 104.955 178.755 ;
        RECT 105.125 178.505 105.600 178.745 ;
        RECT 105.770 178.505 106.120 178.745 ;
        RECT 104.785 178.335 104.955 178.505 ;
        RECT 104.785 178.165 106.120 178.335 ;
        RECT 104.040 177.685 104.790 177.975 ;
        RECT 105.300 177.515 105.630 177.975 ;
        RECT 105.850 177.955 106.120 178.165 ;
        RECT 106.295 178.265 106.815 178.805 ;
        RECT 106.985 178.435 107.505 178.975 ;
        RECT 107.675 178.900 107.965 180.065 ;
        RECT 108.135 178.975 110.725 180.065 ;
        RECT 108.135 178.285 109.345 178.805 ;
        RECT 109.515 178.455 110.725 178.975 ;
        RECT 111.355 179.195 111.630 179.895 ;
        RECT 111.800 179.520 112.055 180.065 ;
        RECT 112.225 179.555 112.705 179.895 ;
        RECT 112.880 179.510 113.485 180.065 ;
        RECT 112.870 179.410 113.485 179.510 ;
        RECT 113.745 179.445 113.915 179.875 ;
        RECT 114.085 179.615 114.415 180.065 ;
        RECT 112.870 179.385 113.055 179.410 ;
        RECT 106.295 177.515 107.505 178.265 ;
        RECT 107.675 177.515 107.965 178.240 ;
        RECT 108.135 177.515 110.725 178.285 ;
        RECT 111.355 178.165 111.525 179.195 ;
        RECT 111.800 179.065 112.555 179.315 ;
        RECT 112.725 179.140 113.055 179.385 ;
        RECT 111.800 179.030 112.570 179.065 ;
        RECT 111.800 179.020 112.585 179.030 ;
        RECT 111.695 179.005 112.590 179.020 ;
        RECT 111.695 178.990 112.610 179.005 ;
        RECT 111.695 178.980 112.630 178.990 ;
        RECT 111.695 178.970 112.655 178.980 ;
        RECT 111.695 178.940 112.725 178.970 ;
        RECT 111.695 178.910 112.745 178.940 ;
        RECT 111.695 178.880 112.765 178.910 ;
        RECT 111.695 178.855 112.795 178.880 ;
        RECT 111.695 178.820 112.830 178.855 ;
        RECT 111.695 178.815 112.860 178.820 ;
        RECT 111.695 178.420 111.925 178.815 ;
        RECT 112.470 178.810 112.860 178.815 ;
        RECT 112.495 178.800 112.860 178.810 ;
        RECT 112.510 178.795 112.860 178.800 ;
        RECT 112.525 178.790 112.860 178.795 ;
        RECT 113.225 178.790 113.485 179.240 ;
        RECT 113.745 179.215 114.420 179.445 ;
        RECT 112.525 178.785 113.485 178.790 ;
        RECT 112.535 178.775 113.485 178.785 ;
        RECT 112.545 178.770 113.485 178.775 ;
        RECT 112.555 178.760 113.485 178.770 ;
        RECT 112.560 178.750 113.485 178.760 ;
        RECT 112.565 178.745 113.485 178.750 ;
        RECT 112.575 178.730 113.485 178.745 ;
        RECT 112.580 178.715 113.485 178.730 ;
        RECT 112.590 178.690 113.485 178.715 ;
        RECT 112.095 178.220 112.425 178.645 ;
        RECT 111.355 177.685 111.615 178.165 ;
        RECT 111.785 177.515 112.035 178.055 ;
        RECT 112.205 177.735 112.425 178.220 ;
        RECT 112.595 178.620 113.485 178.690 ;
        RECT 112.595 177.895 112.765 178.620 ;
        RECT 112.935 178.065 113.485 178.450 ;
        RECT 113.715 178.195 114.015 179.045 ;
        RECT 114.185 178.565 114.420 179.215 ;
        RECT 114.590 178.905 114.875 179.850 ;
        RECT 115.055 179.595 115.740 180.065 ;
        RECT 115.050 179.075 115.745 179.385 ;
        RECT 115.920 179.010 116.225 179.795 ;
        RECT 114.590 178.755 115.450 178.905 ;
        RECT 114.590 178.735 115.875 178.755 ;
        RECT 114.185 178.235 114.720 178.565 ;
        RECT 114.890 178.375 115.875 178.735 ;
        RECT 114.185 178.085 114.405 178.235 ;
        RECT 112.595 177.725 113.485 177.895 ;
        RECT 113.660 177.515 113.995 178.020 ;
        RECT 114.165 177.710 114.405 178.085 ;
        RECT 114.890 178.040 115.060 178.375 ;
        RECT 116.050 178.205 116.225 179.010 ;
        RECT 114.685 177.845 115.060 178.040 ;
        RECT 114.685 177.700 114.855 177.845 ;
        RECT 115.420 177.515 115.815 178.010 ;
        RECT 115.985 177.685 116.225 178.205 ;
        RECT 116.435 179.010 116.740 179.795 ;
        RECT 116.920 179.595 117.605 180.065 ;
        RECT 116.915 179.075 117.610 179.385 ;
        RECT 116.435 178.205 116.610 179.010 ;
        RECT 117.785 178.905 118.070 179.850 ;
        RECT 118.245 179.615 118.575 180.065 ;
        RECT 118.745 179.445 118.915 179.875 ;
        RECT 119.175 179.555 120.365 179.845 ;
        RECT 117.210 178.755 118.070 178.905 ;
        RECT 116.785 178.735 118.070 178.755 ;
        RECT 118.240 179.215 118.915 179.445 ;
        RECT 119.195 179.215 120.365 179.385 ;
        RECT 120.535 179.265 120.815 180.065 ;
        RECT 116.785 178.375 117.770 178.735 ;
        RECT 118.240 178.565 118.475 179.215 ;
        RECT 116.435 177.685 116.675 178.205 ;
        RECT 117.600 178.040 117.770 178.375 ;
        RECT 117.940 178.235 118.475 178.565 ;
        RECT 118.255 178.085 118.475 178.235 ;
        RECT 118.645 178.195 118.945 179.045 ;
        RECT 119.195 178.925 119.520 179.215 ;
        RECT 120.195 179.095 120.365 179.215 ;
        RECT 119.690 178.755 119.885 179.045 ;
        RECT 120.195 178.925 120.855 179.095 ;
        RECT 121.025 178.925 121.300 179.895 ;
        RECT 121.480 178.925 121.800 180.065 ;
        RECT 120.685 178.755 120.855 178.925 ;
        RECT 119.175 178.425 119.520 178.755 ;
        RECT 119.690 178.425 120.515 178.755 ;
        RECT 120.685 178.425 120.960 178.755 ;
        RECT 120.685 178.255 120.855 178.425 ;
        RECT 119.190 178.085 120.855 178.255 ;
        RECT 121.130 178.190 121.300 178.925 ;
        RECT 121.980 178.755 122.175 179.805 ;
        RECT 122.355 179.215 122.685 179.895 ;
        RECT 122.885 179.265 123.140 180.065 ;
        RECT 122.355 178.935 122.705 179.215 ;
        RECT 123.405 179.135 123.575 179.895 ;
        RECT 123.790 179.305 124.120 180.065 ;
        RECT 121.540 178.705 121.800 178.755 ;
        RECT 121.535 178.535 121.800 178.705 ;
        RECT 121.540 178.425 121.800 178.535 ;
        RECT 121.980 178.425 122.365 178.755 ;
        RECT 122.535 178.555 122.705 178.935 ;
        RECT 122.895 178.725 123.140 179.085 ;
        RECT 123.405 178.965 124.120 179.135 ;
        RECT 124.290 178.990 124.545 179.895 ;
        RECT 122.535 178.385 123.055 178.555 ;
        RECT 123.315 178.415 123.670 178.785 ;
        RECT 123.950 178.755 124.120 178.965 ;
        RECT 123.950 178.425 124.205 178.755 ;
        RECT 116.845 177.515 117.240 178.010 ;
        RECT 117.600 177.845 117.975 178.040 ;
        RECT 117.805 177.700 117.975 177.845 ;
        RECT 118.255 177.710 118.495 178.085 ;
        RECT 118.665 177.515 119.000 178.020 ;
        RECT 119.190 177.735 119.445 178.085 ;
        RECT 119.615 177.515 119.945 177.915 ;
        RECT 120.115 177.735 120.285 178.085 ;
        RECT 120.455 177.515 120.835 177.915 ;
        RECT 121.025 177.845 121.300 178.190 ;
        RECT 121.480 178.045 122.695 178.215 ;
        RECT 121.480 177.695 121.770 178.045 ;
        RECT 121.965 177.515 122.295 177.875 ;
        RECT 122.465 177.740 122.695 178.045 ;
        RECT 122.885 178.025 123.055 178.385 ;
        RECT 123.950 178.235 124.120 178.425 ;
        RECT 124.375 178.260 124.545 178.990 ;
        RECT 124.720 178.915 124.980 180.065 ;
        RECT 125.155 179.630 130.500 180.065 ;
        RECT 123.405 178.065 124.120 178.235 ;
        RECT 122.885 177.855 123.085 178.025 ;
        RECT 122.885 177.820 123.055 177.855 ;
        RECT 123.405 177.685 123.575 178.065 ;
        RECT 123.790 177.515 124.120 177.895 ;
        RECT 124.290 177.685 124.545 178.260 ;
        RECT 124.720 177.515 124.980 178.355 ;
        RECT 126.740 178.060 127.080 178.890 ;
        RECT 128.560 178.380 128.910 179.630 ;
        RECT 130.675 178.975 133.265 180.065 ;
        RECT 130.675 178.285 131.885 178.805 ;
        RECT 132.055 178.455 133.265 178.975 ;
        RECT 133.435 178.900 133.725 180.065 ;
        RECT 133.900 178.925 134.235 179.895 ;
        RECT 134.405 178.925 134.575 180.065 ;
        RECT 134.745 179.725 136.775 179.895 ;
        RECT 125.155 177.515 130.500 178.060 ;
        RECT 130.675 177.515 133.265 178.285 ;
        RECT 133.900 178.255 134.070 178.925 ;
        RECT 134.745 178.755 134.915 179.725 ;
        RECT 134.240 178.425 134.495 178.755 ;
        RECT 134.720 178.425 134.915 178.755 ;
        RECT 135.085 179.385 136.210 179.555 ;
        RECT 134.325 178.255 134.495 178.425 ;
        RECT 135.085 178.255 135.255 179.385 ;
        RECT 133.435 177.515 133.725 178.240 ;
        RECT 133.900 177.685 134.155 178.255 ;
        RECT 134.325 178.085 135.255 178.255 ;
        RECT 135.425 179.045 136.435 179.215 ;
        RECT 135.425 178.245 135.595 179.045 ;
        RECT 135.800 178.705 136.075 178.845 ;
        RECT 135.795 178.535 136.075 178.705 ;
        RECT 135.080 178.050 135.255 178.085 ;
        RECT 134.325 177.515 134.655 177.915 ;
        RECT 135.080 177.685 135.610 178.050 ;
        RECT 135.800 177.685 136.075 178.535 ;
        RECT 136.245 177.685 136.435 179.045 ;
        RECT 136.605 179.060 136.775 179.725 ;
        RECT 136.945 179.305 137.115 180.065 ;
        RECT 137.350 179.305 137.865 179.715 ;
        RECT 136.605 178.870 137.355 179.060 ;
        RECT 137.525 178.495 137.865 179.305 ;
        RECT 138.125 179.135 138.295 179.895 ;
        RECT 138.510 179.305 138.840 180.065 ;
        RECT 138.125 178.965 138.840 179.135 ;
        RECT 139.010 178.990 139.265 179.895 ;
        RECT 136.635 178.325 137.865 178.495 ;
        RECT 138.035 178.415 138.390 178.785 ;
        RECT 138.670 178.755 138.840 178.965 ;
        RECT 138.670 178.425 138.925 178.755 ;
        RECT 136.615 177.515 137.125 178.050 ;
        RECT 137.345 177.720 137.590 178.325 ;
        RECT 138.670 178.235 138.840 178.425 ;
        RECT 139.095 178.260 139.265 178.990 ;
        RECT 139.440 178.915 139.700 180.065 ;
        RECT 139.965 179.135 140.135 179.895 ;
        RECT 140.350 179.305 140.680 180.065 ;
        RECT 139.965 178.965 140.680 179.135 ;
        RECT 140.850 178.990 141.105 179.895 ;
        RECT 139.875 178.415 140.230 178.785 ;
        RECT 140.510 178.755 140.680 178.965 ;
        RECT 140.510 178.425 140.765 178.755 ;
        RECT 138.125 178.065 138.840 178.235 ;
        RECT 138.125 177.685 138.295 178.065 ;
        RECT 138.510 177.515 138.840 177.895 ;
        RECT 139.010 177.685 139.265 178.260 ;
        RECT 139.440 177.515 139.700 178.355 ;
        RECT 140.510 178.235 140.680 178.425 ;
        RECT 140.935 178.260 141.105 178.990 ;
        RECT 141.280 178.915 141.540 180.065 ;
        RECT 141.715 178.975 142.925 180.065 ;
        RECT 141.715 178.435 142.235 178.975 ;
        RECT 139.965 178.065 140.680 178.235 ;
        RECT 139.965 177.685 140.135 178.065 ;
        RECT 140.350 177.515 140.680 177.895 ;
        RECT 140.850 177.685 141.105 178.260 ;
        RECT 141.280 177.515 141.540 178.355 ;
        RECT 142.405 178.265 142.925 178.805 ;
        RECT 141.715 177.515 142.925 178.265 ;
        RECT 17.430 177.345 143.010 177.515 ;
        RECT 17.515 176.595 18.725 177.345 ;
        RECT 18.985 176.795 19.155 177.175 ;
        RECT 19.335 176.965 19.665 177.345 ;
        RECT 18.985 176.625 19.650 176.795 ;
        RECT 19.845 176.670 20.105 177.175 ;
        RECT 17.515 176.055 18.035 176.595 ;
        RECT 18.205 175.885 18.725 176.425 ;
        RECT 18.915 176.075 19.245 176.445 ;
        RECT 19.480 176.370 19.650 176.625 ;
        RECT 19.480 176.040 19.765 176.370 ;
        RECT 19.480 175.895 19.650 176.040 ;
        RECT 17.515 174.795 18.725 175.885 ;
        RECT 18.985 175.725 19.650 175.895 ;
        RECT 19.935 175.870 20.105 176.670 ;
        RECT 20.275 176.575 21.945 177.345 ;
        RECT 22.205 176.795 22.375 177.085 ;
        RECT 22.545 176.965 22.875 177.345 ;
        RECT 22.205 176.625 22.870 176.795 ;
        RECT 20.275 176.055 21.025 176.575 ;
        RECT 21.195 175.885 21.945 176.405 ;
        RECT 18.985 174.965 19.155 175.725 ;
        RECT 19.335 174.795 19.665 175.555 ;
        RECT 19.835 174.965 20.105 175.870 ;
        RECT 20.275 174.795 21.945 175.885 ;
        RECT 22.120 175.805 22.470 176.455 ;
        RECT 22.640 175.635 22.870 176.625 ;
        RECT 22.205 175.465 22.870 175.635 ;
        RECT 22.205 174.965 22.375 175.465 ;
        RECT 22.545 174.795 22.875 175.295 ;
        RECT 23.045 174.965 23.230 177.085 ;
        RECT 23.485 176.885 23.735 177.345 ;
        RECT 23.905 176.895 24.240 177.065 ;
        RECT 24.435 176.895 25.110 177.065 ;
        RECT 23.905 176.755 24.075 176.895 ;
        RECT 23.400 175.765 23.680 176.715 ;
        RECT 23.850 176.625 24.075 176.755 ;
        RECT 23.850 175.520 24.020 176.625 ;
        RECT 24.245 176.475 24.770 176.695 ;
        RECT 24.190 175.710 24.430 176.305 ;
        RECT 24.600 175.775 24.770 176.475 ;
        RECT 24.940 176.115 25.110 176.895 ;
        RECT 25.430 176.845 25.800 177.345 ;
        RECT 25.980 176.895 26.385 177.065 ;
        RECT 26.555 176.895 27.340 177.065 ;
        RECT 25.980 176.665 26.150 176.895 ;
        RECT 25.320 176.365 26.150 176.665 ;
        RECT 26.535 176.395 27.000 176.725 ;
        RECT 25.320 176.335 25.520 176.365 ;
        RECT 25.640 176.115 25.810 176.185 ;
        RECT 24.940 175.945 25.810 176.115 ;
        RECT 25.300 175.855 25.810 175.945 ;
        RECT 23.850 175.390 24.155 175.520 ;
        RECT 24.600 175.410 25.130 175.775 ;
        RECT 23.470 174.795 23.735 175.255 ;
        RECT 23.905 174.965 24.155 175.390 ;
        RECT 25.300 175.240 25.470 175.855 ;
        RECT 24.365 175.070 25.470 175.240 ;
        RECT 25.640 174.795 25.810 175.595 ;
        RECT 25.980 175.295 26.150 176.365 ;
        RECT 26.320 175.465 26.510 176.185 ;
        RECT 26.680 175.435 27.000 176.395 ;
        RECT 27.170 176.435 27.340 176.895 ;
        RECT 27.615 176.815 27.825 177.345 ;
        RECT 28.085 176.605 28.415 177.130 ;
        RECT 28.585 176.735 28.755 177.345 ;
        RECT 28.925 176.690 29.255 177.125 ;
        RECT 28.925 176.605 29.305 176.690 ;
        RECT 28.215 176.435 28.415 176.605 ;
        RECT 29.080 176.565 29.305 176.605 ;
        RECT 27.170 176.105 28.045 176.435 ;
        RECT 28.215 176.105 28.965 176.435 ;
        RECT 25.980 174.965 26.230 175.295 ;
        RECT 27.170 175.265 27.340 176.105 ;
        RECT 28.215 175.900 28.405 176.105 ;
        RECT 29.135 175.985 29.305 176.565 ;
        RECT 29.495 176.535 29.735 177.345 ;
        RECT 29.905 176.535 30.235 177.175 ;
        RECT 30.405 176.535 30.675 177.345 ;
        RECT 30.855 176.800 36.200 177.345 ;
        RECT 36.375 176.800 41.720 177.345 ;
        RECT 29.475 176.105 29.825 176.355 ;
        RECT 29.090 175.935 29.305 175.985 ;
        RECT 29.995 175.935 30.165 176.535 ;
        RECT 30.335 176.105 30.685 176.355 ;
        RECT 32.440 175.970 32.780 176.800 ;
        RECT 27.510 175.525 28.405 175.900 ;
        RECT 28.915 175.855 29.305 175.935 ;
        RECT 26.455 175.095 27.340 175.265 ;
        RECT 27.520 174.795 27.835 175.295 ;
        RECT 28.065 174.965 28.405 175.525 ;
        RECT 28.575 174.795 28.745 175.805 ;
        RECT 28.915 175.010 29.245 175.855 ;
        RECT 29.485 175.765 30.165 175.935 ;
        RECT 29.485 174.980 29.815 175.765 ;
        RECT 30.345 174.795 30.675 175.935 ;
        RECT 34.260 175.230 34.610 176.480 ;
        RECT 37.960 175.970 38.300 176.800 ;
        RECT 41.895 176.595 43.105 177.345 ;
        RECT 43.275 176.620 43.565 177.345 ;
        RECT 39.780 175.230 40.130 176.480 ;
        RECT 41.895 176.055 42.415 176.595 ;
        RECT 43.735 176.575 45.405 177.345 ;
        RECT 46.045 176.615 46.345 177.345 ;
        RECT 42.585 175.885 43.105 176.425 ;
        RECT 43.735 176.055 44.485 176.575 ;
        RECT 46.525 176.435 46.755 177.055 ;
        RECT 46.955 176.785 47.180 177.165 ;
        RECT 47.350 176.955 47.680 177.345 ;
        RECT 47.875 176.965 48.765 177.135 ;
        RECT 46.955 176.605 47.285 176.785 ;
        RECT 30.855 174.795 36.200 175.230 ;
        RECT 36.375 174.795 41.720 175.230 ;
        RECT 41.895 174.795 43.105 175.885 ;
        RECT 43.275 174.795 43.565 175.960 ;
        RECT 44.655 175.885 45.405 176.405 ;
        RECT 46.050 176.105 46.345 176.435 ;
        RECT 46.525 176.105 46.940 176.435 ;
        RECT 47.110 175.935 47.285 176.605 ;
        RECT 47.455 176.105 47.695 176.755 ;
        RECT 47.875 176.410 48.425 176.795 ;
        RECT 48.595 176.240 48.765 176.965 ;
        RECT 47.875 176.170 48.765 176.240 ;
        RECT 48.935 176.640 49.155 177.125 ;
        RECT 49.325 176.805 49.575 177.345 ;
        RECT 49.745 176.695 50.005 177.175 ;
        RECT 48.935 176.215 49.265 176.640 ;
        RECT 47.875 176.145 48.770 176.170 ;
        RECT 47.875 176.130 48.780 176.145 ;
        RECT 47.875 176.115 48.785 176.130 ;
        RECT 47.875 176.110 48.795 176.115 ;
        RECT 47.875 176.100 48.800 176.110 ;
        RECT 47.875 176.090 48.805 176.100 ;
        RECT 47.875 176.085 48.815 176.090 ;
        RECT 47.875 176.075 48.825 176.085 ;
        RECT 47.875 176.070 48.835 176.075 ;
        RECT 43.735 174.795 45.405 175.885 ;
        RECT 46.045 175.575 46.940 175.905 ;
        RECT 47.110 175.745 47.695 175.935 ;
        RECT 46.045 175.405 47.250 175.575 ;
        RECT 46.045 174.975 46.375 175.405 ;
        RECT 46.555 174.795 46.750 175.235 ;
        RECT 46.920 174.975 47.250 175.405 ;
        RECT 47.420 174.975 47.695 175.745 ;
        RECT 47.875 175.620 48.135 176.070 ;
        RECT 48.500 176.065 48.835 176.070 ;
        RECT 48.500 176.060 48.850 176.065 ;
        RECT 48.500 176.050 48.865 176.060 ;
        RECT 48.500 176.045 48.890 176.050 ;
        RECT 49.435 176.045 49.665 176.440 ;
        RECT 48.500 176.040 49.665 176.045 ;
        RECT 48.530 176.005 49.665 176.040 ;
        RECT 48.565 175.980 49.665 176.005 ;
        RECT 48.595 175.950 49.665 175.980 ;
        RECT 48.615 175.920 49.665 175.950 ;
        RECT 48.635 175.890 49.665 175.920 ;
        RECT 48.705 175.880 49.665 175.890 ;
        RECT 48.730 175.870 49.665 175.880 ;
        RECT 48.750 175.855 49.665 175.870 ;
        RECT 48.770 175.840 49.665 175.855 ;
        RECT 48.775 175.830 49.560 175.840 ;
        RECT 48.790 175.795 49.560 175.830 ;
        RECT 48.305 175.475 48.635 175.720 ;
        RECT 48.805 175.545 49.560 175.795 ;
        RECT 49.835 175.665 50.005 176.695 ;
        RECT 50.265 176.795 50.435 177.085 ;
        RECT 50.605 176.965 50.935 177.345 ;
        RECT 50.265 176.625 50.930 176.795 ;
        RECT 50.180 175.805 50.530 176.455 ;
        RECT 48.305 175.450 48.490 175.475 ;
        RECT 47.875 175.350 48.490 175.450 ;
        RECT 47.875 174.795 48.480 175.350 ;
        RECT 48.655 174.965 49.135 175.305 ;
        RECT 49.305 174.795 49.560 175.340 ;
        RECT 49.730 174.965 50.005 175.665 ;
        RECT 50.700 175.635 50.930 176.625 ;
        RECT 50.265 175.465 50.930 175.635 ;
        RECT 50.265 174.965 50.435 175.465 ;
        RECT 50.605 174.795 50.935 175.295 ;
        RECT 51.105 174.965 51.290 177.085 ;
        RECT 51.545 176.885 51.795 177.345 ;
        RECT 51.965 176.895 52.300 177.065 ;
        RECT 52.495 176.895 53.170 177.065 ;
        RECT 51.965 176.755 52.135 176.895 ;
        RECT 51.460 175.765 51.740 176.715 ;
        RECT 51.910 176.625 52.135 176.755 ;
        RECT 51.910 175.520 52.080 176.625 ;
        RECT 52.305 176.475 52.830 176.695 ;
        RECT 52.250 175.710 52.490 176.305 ;
        RECT 52.660 175.775 52.830 176.475 ;
        RECT 53.000 176.115 53.170 176.895 ;
        RECT 53.490 176.845 53.860 177.345 ;
        RECT 54.040 176.895 54.445 177.065 ;
        RECT 54.615 176.895 55.400 177.065 ;
        RECT 54.040 176.665 54.210 176.895 ;
        RECT 53.380 176.365 54.210 176.665 ;
        RECT 54.595 176.395 55.060 176.725 ;
        RECT 53.380 176.335 53.580 176.365 ;
        RECT 53.700 176.115 53.870 176.185 ;
        RECT 53.000 175.945 53.870 176.115 ;
        RECT 53.360 175.855 53.870 175.945 ;
        RECT 51.910 175.390 52.215 175.520 ;
        RECT 52.660 175.410 53.190 175.775 ;
        RECT 51.530 174.795 51.795 175.255 ;
        RECT 51.965 174.965 52.215 175.390 ;
        RECT 53.360 175.240 53.530 175.855 ;
        RECT 52.425 175.070 53.530 175.240 ;
        RECT 53.700 174.795 53.870 175.595 ;
        RECT 54.040 175.295 54.210 176.365 ;
        RECT 54.380 175.465 54.570 176.185 ;
        RECT 54.740 175.435 55.060 176.395 ;
        RECT 55.230 176.435 55.400 176.895 ;
        RECT 55.675 176.815 55.885 177.345 ;
        RECT 56.145 176.605 56.475 177.130 ;
        RECT 56.645 176.735 56.815 177.345 ;
        RECT 56.985 176.690 57.315 177.125 ;
        RECT 56.985 176.605 57.365 176.690 ;
        RECT 56.275 176.435 56.475 176.605 ;
        RECT 57.140 176.565 57.365 176.605 ;
        RECT 55.230 176.105 56.105 176.435 ;
        RECT 56.275 176.105 57.025 176.435 ;
        RECT 54.040 174.965 54.290 175.295 ;
        RECT 55.230 175.265 55.400 176.105 ;
        RECT 56.275 175.900 56.465 176.105 ;
        RECT 57.195 175.985 57.365 176.565 ;
        RECT 57.535 176.575 61.045 177.345 ;
        RECT 61.765 176.795 61.935 177.085 ;
        RECT 62.105 176.965 62.435 177.345 ;
        RECT 61.765 176.625 62.430 176.795 ;
        RECT 57.535 176.055 59.185 176.575 ;
        RECT 57.150 175.935 57.365 175.985 ;
        RECT 55.570 175.525 56.465 175.900 ;
        RECT 56.975 175.855 57.365 175.935 ;
        RECT 59.355 175.885 61.045 176.405 ;
        RECT 54.515 175.095 55.400 175.265 ;
        RECT 55.580 174.795 55.895 175.295 ;
        RECT 56.125 174.965 56.465 175.525 ;
        RECT 56.635 174.795 56.805 175.805 ;
        RECT 56.975 175.010 57.305 175.855 ;
        RECT 57.535 174.795 61.045 175.885 ;
        RECT 61.680 175.805 62.030 176.455 ;
        RECT 62.200 175.635 62.430 176.625 ;
        RECT 61.765 175.465 62.430 175.635 ;
        RECT 61.765 174.965 61.935 175.465 ;
        RECT 62.105 174.795 62.435 175.295 ;
        RECT 62.605 174.965 62.790 177.085 ;
        RECT 63.045 176.885 63.295 177.345 ;
        RECT 63.465 176.895 63.800 177.065 ;
        RECT 63.995 176.895 64.670 177.065 ;
        RECT 63.465 176.755 63.635 176.895 ;
        RECT 62.960 175.765 63.240 176.715 ;
        RECT 63.410 176.625 63.635 176.755 ;
        RECT 63.410 175.520 63.580 176.625 ;
        RECT 63.805 176.475 64.330 176.695 ;
        RECT 63.750 175.710 63.990 176.305 ;
        RECT 64.160 175.775 64.330 176.475 ;
        RECT 64.500 176.115 64.670 176.895 ;
        RECT 64.990 176.845 65.360 177.345 ;
        RECT 65.540 176.895 65.945 177.065 ;
        RECT 66.115 176.895 66.900 177.065 ;
        RECT 65.540 176.665 65.710 176.895 ;
        RECT 64.880 176.365 65.710 176.665 ;
        RECT 66.095 176.395 66.560 176.725 ;
        RECT 64.880 176.335 65.080 176.365 ;
        RECT 65.200 176.115 65.370 176.185 ;
        RECT 64.500 175.945 65.370 176.115 ;
        RECT 64.860 175.855 65.370 175.945 ;
        RECT 63.410 175.390 63.715 175.520 ;
        RECT 64.160 175.410 64.690 175.775 ;
        RECT 63.030 174.795 63.295 175.255 ;
        RECT 63.465 174.965 63.715 175.390 ;
        RECT 64.860 175.240 65.030 175.855 ;
        RECT 63.925 175.070 65.030 175.240 ;
        RECT 65.200 174.795 65.370 175.595 ;
        RECT 65.540 175.295 65.710 176.365 ;
        RECT 65.880 175.465 66.070 176.185 ;
        RECT 66.240 175.435 66.560 176.395 ;
        RECT 66.730 176.435 66.900 176.895 ;
        RECT 67.175 176.815 67.385 177.345 ;
        RECT 67.645 176.605 67.975 177.130 ;
        RECT 68.145 176.735 68.315 177.345 ;
        RECT 68.485 176.690 68.815 177.125 ;
        RECT 68.485 176.605 68.865 176.690 ;
        RECT 69.035 176.620 69.325 177.345 ;
        RECT 67.775 176.435 67.975 176.605 ;
        RECT 68.640 176.565 68.865 176.605 ;
        RECT 66.730 176.105 67.605 176.435 ;
        RECT 67.775 176.105 68.525 176.435 ;
        RECT 65.540 174.965 65.790 175.295 ;
        RECT 66.730 175.265 66.900 176.105 ;
        RECT 67.775 175.900 67.965 176.105 ;
        RECT 68.695 175.985 68.865 176.565 ;
        RECT 68.650 175.935 68.865 175.985 ;
        RECT 67.070 175.525 67.965 175.900 ;
        RECT 68.475 175.855 68.865 175.935 ;
        RECT 66.015 175.095 66.900 175.265 ;
        RECT 67.080 174.795 67.395 175.295 ;
        RECT 67.625 174.965 67.965 175.525 ;
        RECT 68.135 174.795 68.305 175.805 ;
        RECT 68.475 175.010 68.805 175.855 ;
        RECT 69.035 174.795 69.325 175.960 ;
        RECT 69.505 174.975 69.765 177.165 ;
        RECT 70.025 176.975 70.695 177.345 ;
        RECT 70.875 176.795 71.185 177.165 ;
        RECT 69.955 176.595 71.185 176.795 ;
        RECT 69.955 175.925 70.245 176.595 ;
        RECT 71.365 176.415 71.595 177.055 ;
        RECT 71.775 176.615 72.065 177.345 ;
        RECT 72.345 176.795 72.515 177.085 ;
        RECT 72.685 176.965 73.015 177.345 ;
        RECT 72.345 176.625 73.010 176.795 ;
        RECT 70.425 176.105 70.890 176.415 ;
        RECT 71.070 176.105 71.595 176.415 ;
        RECT 71.775 176.105 72.075 176.435 ;
        RECT 69.955 175.705 70.725 175.925 ;
        RECT 69.935 174.795 70.275 175.525 ;
        RECT 70.455 174.975 70.725 175.705 ;
        RECT 70.905 175.685 72.065 175.925 ;
        RECT 72.260 175.805 72.610 176.455 ;
        RECT 70.905 174.975 71.135 175.685 ;
        RECT 71.305 174.795 71.635 175.505 ;
        RECT 71.805 174.975 72.065 175.685 ;
        RECT 72.780 175.635 73.010 176.625 ;
        RECT 72.345 175.465 73.010 175.635 ;
        RECT 72.345 174.965 72.515 175.465 ;
        RECT 72.685 174.795 73.015 175.295 ;
        RECT 73.185 174.965 73.370 177.085 ;
        RECT 73.625 176.885 73.875 177.345 ;
        RECT 74.045 176.895 74.380 177.065 ;
        RECT 74.575 176.895 75.250 177.065 ;
        RECT 74.045 176.755 74.215 176.895 ;
        RECT 73.540 175.765 73.820 176.715 ;
        RECT 73.990 176.625 74.215 176.755 ;
        RECT 73.990 175.520 74.160 176.625 ;
        RECT 74.385 176.475 74.910 176.695 ;
        RECT 74.330 175.710 74.570 176.305 ;
        RECT 74.740 175.775 74.910 176.475 ;
        RECT 75.080 176.115 75.250 176.895 ;
        RECT 75.570 176.845 75.940 177.345 ;
        RECT 76.120 176.895 76.525 177.065 ;
        RECT 76.695 176.895 77.480 177.065 ;
        RECT 76.120 176.665 76.290 176.895 ;
        RECT 75.460 176.365 76.290 176.665 ;
        RECT 76.675 176.395 77.140 176.725 ;
        RECT 75.460 176.335 75.660 176.365 ;
        RECT 75.780 176.115 75.950 176.185 ;
        RECT 75.080 175.945 75.950 176.115 ;
        RECT 75.440 175.855 75.950 175.945 ;
        RECT 73.990 175.390 74.295 175.520 ;
        RECT 74.740 175.410 75.270 175.775 ;
        RECT 73.610 174.795 73.875 175.255 ;
        RECT 74.045 174.965 74.295 175.390 ;
        RECT 75.440 175.240 75.610 175.855 ;
        RECT 74.505 175.070 75.610 175.240 ;
        RECT 75.780 174.795 75.950 175.595 ;
        RECT 76.120 175.295 76.290 176.365 ;
        RECT 76.460 175.465 76.650 176.185 ;
        RECT 76.820 175.435 77.140 176.395 ;
        RECT 77.310 176.435 77.480 176.895 ;
        RECT 77.755 176.815 77.965 177.345 ;
        RECT 78.225 176.605 78.555 177.130 ;
        RECT 78.725 176.735 78.895 177.345 ;
        RECT 79.065 176.690 79.395 177.125 ;
        RECT 79.665 176.690 79.995 177.125 ;
        RECT 80.165 176.735 80.335 177.345 ;
        RECT 79.065 176.605 79.445 176.690 ;
        RECT 78.355 176.435 78.555 176.605 ;
        RECT 79.220 176.565 79.445 176.605 ;
        RECT 77.310 176.105 78.185 176.435 ;
        RECT 78.355 176.105 79.105 176.435 ;
        RECT 76.120 174.965 76.370 175.295 ;
        RECT 77.310 175.265 77.480 176.105 ;
        RECT 78.355 175.900 78.545 176.105 ;
        RECT 79.275 175.985 79.445 176.565 ;
        RECT 79.230 175.935 79.445 175.985 ;
        RECT 77.650 175.525 78.545 175.900 ;
        RECT 79.055 175.855 79.445 175.935 ;
        RECT 79.615 176.605 79.995 176.690 ;
        RECT 80.505 176.605 80.835 177.130 ;
        RECT 81.095 176.815 81.305 177.345 ;
        RECT 81.580 176.895 82.365 177.065 ;
        RECT 82.535 176.895 82.940 177.065 ;
        RECT 79.615 176.565 79.840 176.605 ;
        RECT 79.615 175.985 79.785 176.565 ;
        RECT 80.505 176.435 80.705 176.605 ;
        RECT 81.580 176.435 81.750 176.895 ;
        RECT 79.955 176.105 80.705 176.435 ;
        RECT 80.875 176.105 81.750 176.435 ;
        RECT 79.615 175.935 79.830 175.985 ;
        RECT 79.615 175.855 80.005 175.935 ;
        RECT 76.595 175.095 77.480 175.265 ;
        RECT 77.660 174.795 77.975 175.295 ;
        RECT 78.205 174.965 78.545 175.525 ;
        RECT 78.715 174.795 78.885 175.805 ;
        RECT 79.055 175.010 79.385 175.855 ;
        RECT 79.675 175.010 80.005 175.855 ;
        RECT 80.515 175.900 80.705 176.105 ;
        RECT 80.175 174.795 80.345 175.805 ;
        RECT 80.515 175.525 81.410 175.900 ;
        RECT 80.515 174.965 80.855 175.525 ;
        RECT 81.085 174.795 81.400 175.295 ;
        RECT 81.580 175.265 81.750 176.105 ;
        RECT 81.920 176.395 82.385 176.725 ;
        RECT 82.770 176.665 82.940 176.895 ;
        RECT 83.120 176.845 83.490 177.345 ;
        RECT 83.810 176.895 84.485 177.065 ;
        RECT 84.680 176.895 85.015 177.065 ;
        RECT 81.920 175.435 82.240 176.395 ;
        RECT 82.770 176.365 83.600 176.665 ;
        RECT 82.410 175.465 82.600 176.185 ;
        RECT 82.770 175.295 82.940 176.365 ;
        RECT 83.400 176.335 83.600 176.365 ;
        RECT 83.110 176.115 83.280 176.185 ;
        RECT 83.810 176.115 83.980 176.895 ;
        RECT 84.845 176.755 85.015 176.895 ;
        RECT 85.185 176.885 85.435 177.345 ;
        RECT 83.110 175.945 83.980 176.115 ;
        RECT 84.150 176.475 84.675 176.695 ;
        RECT 84.845 176.625 85.070 176.755 ;
        RECT 83.110 175.855 83.620 175.945 ;
        RECT 81.580 175.095 82.465 175.265 ;
        RECT 82.690 174.965 82.940 175.295 ;
        RECT 83.110 174.795 83.280 175.595 ;
        RECT 83.450 175.240 83.620 175.855 ;
        RECT 84.150 175.775 84.320 176.475 ;
        RECT 83.790 175.410 84.320 175.775 ;
        RECT 84.490 175.710 84.730 176.305 ;
        RECT 84.900 175.520 85.070 176.625 ;
        RECT 85.240 175.765 85.520 176.715 ;
        RECT 84.765 175.390 85.070 175.520 ;
        RECT 83.450 175.070 84.555 175.240 ;
        RECT 84.765 174.965 85.015 175.390 ;
        RECT 85.185 174.795 85.450 175.255 ;
        RECT 85.690 174.965 85.875 177.085 ;
        RECT 86.045 176.965 86.375 177.345 ;
        RECT 86.545 176.795 86.715 177.085 ;
        RECT 86.050 176.625 86.715 176.795 ;
        RECT 86.050 175.635 86.280 176.625 ;
        RECT 86.975 176.605 87.360 177.175 ;
        RECT 87.530 176.885 87.855 177.345 ;
        RECT 88.375 176.715 88.655 177.175 ;
        RECT 86.450 175.805 86.800 176.455 ;
        RECT 86.975 175.935 87.255 176.605 ;
        RECT 87.530 176.545 88.655 176.715 ;
        RECT 87.530 176.435 87.980 176.545 ;
        RECT 87.425 176.105 87.980 176.435 ;
        RECT 88.845 176.375 89.245 177.175 ;
        RECT 89.645 176.885 89.915 177.345 ;
        RECT 90.085 176.715 90.370 177.175 ;
        RECT 86.050 175.465 86.715 175.635 ;
        RECT 86.045 174.795 86.375 175.295 ;
        RECT 86.545 174.965 86.715 175.465 ;
        RECT 86.975 174.965 87.360 175.935 ;
        RECT 87.530 175.645 87.980 176.105 ;
        RECT 88.150 175.815 89.245 176.375 ;
        RECT 87.530 175.425 88.655 175.645 ;
        RECT 87.530 174.795 87.855 175.255 ;
        RECT 88.375 174.965 88.655 175.425 ;
        RECT 88.845 174.965 89.245 175.815 ;
        RECT 89.415 176.545 90.370 176.715 ;
        RECT 90.655 176.575 94.165 177.345 ;
        RECT 94.795 176.620 95.085 177.345 ;
        RECT 95.255 176.800 100.600 177.345 ;
        RECT 100.775 176.800 106.120 177.345 ;
        RECT 89.415 175.645 89.625 176.545 ;
        RECT 89.795 175.815 90.485 176.375 ;
        RECT 90.655 176.055 92.305 176.575 ;
        RECT 92.475 175.885 94.165 176.405 ;
        RECT 96.840 175.970 97.180 176.800 ;
        RECT 89.415 175.425 90.370 175.645 ;
        RECT 89.645 174.795 89.915 175.255 ;
        RECT 90.085 174.965 90.370 175.425 ;
        RECT 90.655 174.795 94.165 175.885 ;
        RECT 94.795 174.795 95.085 175.960 ;
        RECT 98.660 175.230 99.010 176.480 ;
        RECT 102.360 175.970 102.700 176.800 ;
        RECT 106.295 176.575 109.805 177.345 ;
        RECT 110.435 176.605 110.925 177.175 ;
        RECT 111.095 176.775 111.325 177.175 ;
        RECT 111.495 176.945 111.915 177.345 ;
        RECT 112.085 176.775 112.255 177.175 ;
        RECT 111.095 176.605 112.255 176.775 ;
        RECT 112.425 176.605 112.875 177.345 ;
        RECT 113.045 176.605 113.485 177.165 ;
        RECT 113.675 176.835 113.915 177.345 ;
        RECT 114.085 176.835 114.375 177.175 ;
        RECT 114.605 176.835 114.920 177.345 ;
        RECT 104.180 175.230 104.530 176.480 ;
        RECT 106.295 176.055 107.945 176.575 ;
        RECT 108.115 175.885 109.805 176.405 ;
        RECT 95.255 174.795 100.600 175.230 ;
        RECT 100.775 174.795 106.120 175.230 ;
        RECT 106.295 174.795 109.805 175.885 ;
        RECT 110.435 175.935 110.605 176.605 ;
        RECT 110.775 176.105 111.180 176.435 ;
        RECT 110.435 175.765 111.205 175.935 ;
        RECT 110.445 174.795 110.775 175.595 ;
        RECT 110.955 175.135 111.205 175.765 ;
        RECT 111.395 175.305 111.645 176.435 ;
        RECT 111.845 176.105 112.090 176.435 ;
        RECT 112.275 176.155 112.665 176.435 ;
        RECT 111.845 175.305 112.045 176.105 ;
        RECT 112.835 175.985 113.005 176.435 ;
        RECT 112.215 175.815 113.005 175.985 ;
        RECT 112.215 175.135 112.385 175.815 ;
        RECT 110.955 174.965 112.385 175.135 ;
        RECT 112.555 174.795 112.870 175.645 ;
        RECT 113.175 175.595 113.485 176.605 ;
        RECT 113.715 176.495 113.915 176.665 ;
        RECT 113.720 176.105 113.915 176.495 ;
        RECT 114.085 175.935 114.265 176.835 ;
        RECT 115.090 176.775 115.260 177.045 ;
        RECT 115.430 176.945 115.760 177.345 ;
        RECT 115.960 176.815 116.250 177.165 ;
        RECT 116.445 176.985 116.775 177.345 ;
        RECT 116.945 176.815 117.175 177.120 ;
        RECT 114.435 176.105 114.845 176.665 ;
        RECT 115.090 176.605 115.785 176.775 ;
        RECT 115.960 176.645 117.175 176.815 ;
        RECT 115.015 175.935 115.185 176.435 ;
        RECT 113.045 174.965 113.485 175.595 ;
        RECT 113.725 175.765 115.185 175.935 ;
        RECT 113.725 175.590 114.085 175.765 ;
        RECT 115.355 175.595 115.785 176.605 ;
        RECT 117.365 176.475 117.535 177.040 ;
        RECT 117.820 176.945 118.150 177.345 ;
        RECT 118.320 176.775 118.490 177.045 ;
        RECT 118.660 176.835 118.975 177.345 ;
        RECT 119.205 176.835 119.495 177.175 ;
        RECT 119.665 176.835 119.905 177.345 ;
        RECT 116.020 176.325 116.280 176.435 ;
        RECT 116.015 176.155 116.280 176.325 ;
        RECT 116.020 176.105 116.280 176.155 ;
        RECT 116.460 176.105 116.845 176.435 ;
        RECT 117.015 176.305 117.535 176.475 ;
        RECT 117.795 176.605 118.490 176.775 ;
        RECT 114.670 174.795 114.840 175.595 ;
        RECT 115.010 175.425 115.785 175.595 ;
        RECT 115.010 174.965 115.340 175.425 ;
        RECT 115.510 174.795 115.680 175.255 ;
        RECT 115.960 174.795 116.280 175.935 ;
        RECT 116.460 175.055 116.655 176.105 ;
        RECT 117.015 175.925 117.185 176.305 ;
        RECT 116.835 175.645 117.185 175.925 ;
        RECT 117.375 175.775 117.620 176.135 ;
        RECT 116.835 174.965 117.165 175.645 ;
        RECT 117.795 175.595 118.225 176.605 ;
        RECT 118.395 175.935 118.565 176.435 ;
        RECT 118.735 176.105 119.145 176.665 ;
        RECT 119.315 175.935 119.495 176.835 ;
        RECT 119.665 176.495 119.865 176.665 ;
        RECT 120.555 176.620 120.845 177.345 ;
        RECT 121.220 176.565 121.720 177.175 ;
        RECT 119.665 176.105 119.860 176.495 ;
        RECT 121.015 176.105 121.365 176.355 ;
        RECT 118.395 175.765 119.855 175.935 ;
        RECT 117.365 174.795 117.620 175.595 ;
        RECT 117.795 175.425 118.570 175.595 ;
        RECT 117.900 174.795 118.070 175.255 ;
        RECT 118.240 174.965 118.570 175.425 ;
        RECT 118.740 174.795 118.910 175.595 ;
        RECT 119.495 175.590 119.855 175.765 ;
        RECT 120.555 174.795 120.845 175.960 ;
        RECT 121.550 175.935 121.720 176.565 ;
        RECT 122.350 176.695 122.680 177.175 ;
        RECT 122.850 176.885 123.075 177.345 ;
        RECT 123.245 176.695 123.575 177.175 ;
        RECT 122.350 176.525 123.575 176.695 ;
        RECT 123.765 176.545 124.015 177.345 ;
        RECT 124.185 176.545 124.525 177.175 ;
        RECT 121.890 176.155 122.220 176.355 ;
        RECT 122.390 176.155 122.720 176.355 ;
        RECT 122.890 176.155 123.310 176.355 ;
        RECT 123.485 176.185 124.180 176.355 ;
        RECT 123.485 175.935 123.655 176.185 ;
        RECT 124.350 175.935 124.525 176.545 ;
        RECT 124.700 176.525 124.975 177.345 ;
        RECT 125.145 176.705 125.475 177.175 ;
        RECT 125.645 176.875 125.815 177.345 ;
        RECT 125.985 176.705 126.315 177.175 ;
        RECT 126.485 176.875 126.775 177.345 ;
        RECT 125.145 176.695 126.315 176.705 ;
        RECT 125.145 176.525 126.745 176.695 ;
        RECT 124.700 176.155 125.420 176.355 ;
        RECT 125.590 176.155 126.360 176.355 ;
        RECT 126.530 175.985 126.745 176.525 ;
        RECT 126.995 176.575 128.665 177.345 ;
        RECT 129.385 176.795 129.555 177.175 ;
        RECT 129.735 176.965 130.065 177.345 ;
        RECT 129.385 176.625 130.050 176.795 ;
        RECT 130.245 176.670 130.505 177.175 ;
        RECT 126.995 176.055 127.745 176.575 ;
        RECT 121.220 175.765 123.655 175.935 ;
        RECT 121.220 174.965 121.550 175.765 ;
        RECT 121.720 174.795 122.050 175.595 ;
        RECT 122.350 174.965 122.680 175.765 ;
        RECT 123.325 174.795 123.575 175.595 ;
        RECT 123.845 174.795 124.015 175.935 ;
        RECT 124.185 174.965 124.525 175.935 ;
        RECT 124.700 175.765 125.815 175.975 ;
        RECT 124.700 174.965 124.975 175.765 ;
        RECT 125.145 174.795 125.475 175.595 ;
        RECT 125.645 175.135 125.815 175.765 ;
        RECT 125.985 175.815 126.765 175.985 ;
        RECT 127.915 175.885 128.665 176.405 ;
        RECT 129.315 176.075 129.645 176.445 ;
        RECT 129.880 176.370 130.050 176.625 ;
        RECT 129.880 176.040 130.165 176.370 ;
        RECT 129.880 175.895 130.050 176.040 ;
        RECT 125.985 175.765 126.745 175.815 ;
        RECT 125.985 175.305 126.315 175.765 ;
        RECT 126.485 175.135 126.785 175.595 ;
        RECT 125.645 174.965 126.785 175.135 ;
        RECT 126.995 174.795 128.665 175.885 ;
        RECT 129.385 175.725 130.050 175.895 ;
        RECT 130.335 175.870 130.505 176.670 ;
        RECT 130.765 176.795 130.935 177.085 ;
        RECT 131.105 176.965 131.435 177.345 ;
        RECT 130.765 176.625 131.430 176.795 ;
        RECT 129.385 174.965 129.555 175.725 ;
        RECT 129.735 174.795 130.065 175.555 ;
        RECT 130.235 174.965 130.505 175.870 ;
        RECT 130.680 175.805 131.030 176.455 ;
        RECT 131.200 175.635 131.430 176.625 ;
        RECT 130.765 175.465 131.430 175.635 ;
        RECT 130.765 174.965 130.935 175.465 ;
        RECT 131.105 174.795 131.435 175.295 ;
        RECT 131.605 174.965 131.790 177.085 ;
        RECT 132.045 176.885 132.295 177.345 ;
        RECT 132.465 176.895 132.800 177.065 ;
        RECT 132.995 176.895 133.670 177.065 ;
        RECT 132.465 176.755 132.635 176.895 ;
        RECT 131.960 175.765 132.240 176.715 ;
        RECT 132.410 176.625 132.635 176.755 ;
        RECT 132.410 175.520 132.580 176.625 ;
        RECT 132.805 176.475 133.330 176.695 ;
        RECT 132.750 175.710 132.990 176.305 ;
        RECT 133.160 175.775 133.330 176.475 ;
        RECT 133.500 176.115 133.670 176.895 ;
        RECT 133.990 176.845 134.360 177.345 ;
        RECT 134.540 176.895 134.945 177.065 ;
        RECT 135.115 176.895 135.900 177.065 ;
        RECT 134.540 176.665 134.710 176.895 ;
        RECT 133.880 176.365 134.710 176.665 ;
        RECT 135.095 176.395 135.560 176.725 ;
        RECT 133.880 176.335 134.080 176.365 ;
        RECT 134.200 176.115 134.370 176.185 ;
        RECT 133.500 175.945 134.370 176.115 ;
        RECT 133.860 175.855 134.370 175.945 ;
        RECT 132.410 175.390 132.715 175.520 ;
        RECT 133.160 175.410 133.690 175.775 ;
        RECT 132.030 174.795 132.295 175.255 ;
        RECT 132.465 174.965 132.715 175.390 ;
        RECT 133.860 175.240 134.030 175.855 ;
        RECT 132.925 175.070 134.030 175.240 ;
        RECT 134.200 174.795 134.370 175.595 ;
        RECT 134.540 175.295 134.710 176.365 ;
        RECT 134.880 175.465 135.070 176.185 ;
        RECT 135.240 175.435 135.560 176.395 ;
        RECT 135.730 176.435 135.900 176.895 ;
        RECT 136.175 176.815 136.385 177.345 ;
        RECT 136.645 176.605 136.975 177.130 ;
        RECT 137.145 176.735 137.315 177.345 ;
        RECT 137.485 176.690 137.815 177.125 ;
        RECT 137.485 176.605 137.865 176.690 ;
        RECT 136.775 176.435 136.975 176.605 ;
        RECT 137.640 176.565 137.865 176.605 ;
        RECT 135.730 176.105 136.605 176.435 ;
        RECT 136.775 176.105 137.525 176.435 ;
        RECT 134.540 174.965 134.790 175.295 ;
        RECT 135.730 175.265 135.900 176.105 ;
        RECT 136.775 175.900 136.965 176.105 ;
        RECT 137.695 175.985 137.865 176.565 ;
        RECT 137.650 175.935 137.865 175.985 ;
        RECT 136.070 175.525 136.965 175.900 ;
        RECT 137.475 175.855 137.865 175.935 ;
        RECT 138.035 176.605 138.420 177.175 ;
        RECT 138.590 176.885 138.915 177.345 ;
        RECT 139.435 176.715 139.715 177.175 ;
        RECT 138.035 175.935 138.315 176.605 ;
        RECT 138.590 176.545 139.715 176.715 ;
        RECT 138.590 176.435 139.040 176.545 ;
        RECT 138.485 176.105 139.040 176.435 ;
        RECT 139.905 176.375 140.305 177.175 ;
        RECT 140.705 176.885 140.975 177.345 ;
        RECT 141.145 176.715 141.430 177.175 ;
        RECT 135.015 175.095 135.900 175.265 ;
        RECT 136.080 174.795 136.395 175.295 ;
        RECT 136.625 174.965 136.965 175.525 ;
        RECT 137.135 174.795 137.305 175.805 ;
        RECT 137.475 175.010 137.805 175.855 ;
        RECT 138.035 174.965 138.420 175.935 ;
        RECT 138.590 175.645 139.040 176.105 ;
        RECT 139.210 175.815 140.305 176.375 ;
        RECT 138.590 175.425 139.715 175.645 ;
        RECT 138.590 174.795 138.915 175.255 ;
        RECT 139.435 174.965 139.715 175.425 ;
        RECT 139.905 174.965 140.305 175.815 ;
        RECT 140.475 176.545 141.430 176.715 ;
        RECT 141.715 176.595 142.925 177.345 ;
        RECT 140.475 175.645 140.685 176.545 ;
        RECT 140.855 175.815 141.545 176.375 ;
        RECT 141.715 175.885 142.235 176.425 ;
        RECT 142.405 176.055 142.925 176.595 ;
        RECT 140.475 175.425 141.430 175.645 ;
        RECT 140.705 174.795 140.975 175.255 ;
        RECT 141.145 174.965 141.430 175.425 ;
        RECT 141.715 174.795 142.925 175.885 ;
        RECT 17.430 174.625 143.010 174.795 ;
        RECT 17.515 173.535 18.725 174.625 ;
        RECT 18.895 173.535 20.565 174.625 ;
        RECT 21.285 173.955 21.455 174.455 ;
        RECT 21.625 174.125 21.955 174.625 ;
        RECT 21.285 173.785 21.950 173.955 ;
        RECT 17.515 172.825 18.035 173.365 ;
        RECT 18.205 172.995 18.725 173.535 ;
        RECT 18.895 172.845 19.645 173.365 ;
        RECT 19.815 173.015 20.565 173.535 ;
        RECT 21.200 172.965 21.550 173.615 ;
        RECT 17.515 172.075 18.725 172.825 ;
        RECT 18.895 172.075 20.565 172.845 ;
        RECT 21.720 172.795 21.950 173.785 ;
        RECT 21.285 172.625 21.950 172.795 ;
        RECT 21.285 172.335 21.455 172.625 ;
        RECT 21.625 172.075 21.955 172.455 ;
        RECT 22.125 172.335 22.310 174.455 ;
        RECT 22.550 174.165 22.815 174.625 ;
        RECT 22.985 174.030 23.235 174.455 ;
        RECT 23.445 174.180 24.550 174.350 ;
        RECT 22.930 173.900 23.235 174.030 ;
        RECT 22.480 172.705 22.760 173.655 ;
        RECT 22.930 172.795 23.100 173.900 ;
        RECT 23.270 173.115 23.510 173.710 ;
        RECT 23.680 173.645 24.210 174.010 ;
        RECT 23.680 172.945 23.850 173.645 ;
        RECT 24.380 173.565 24.550 174.180 ;
        RECT 24.720 173.825 24.890 174.625 ;
        RECT 25.060 174.125 25.310 174.455 ;
        RECT 25.535 174.155 26.420 174.325 ;
        RECT 24.380 173.475 24.890 173.565 ;
        RECT 22.930 172.665 23.155 172.795 ;
        RECT 23.325 172.725 23.850 172.945 ;
        RECT 24.020 173.305 24.890 173.475 ;
        RECT 22.565 172.075 22.815 172.535 ;
        RECT 22.985 172.525 23.155 172.665 ;
        RECT 24.020 172.525 24.190 173.305 ;
        RECT 24.720 173.235 24.890 173.305 ;
        RECT 24.400 173.055 24.600 173.085 ;
        RECT 25.060 173.055 25.230 174.125 ;
        RECT 25.400 173.235 25.590 173.955 ;
        RECT 24.400 172.755 25.230 173.055 ;
        RECT 25.760 173.025 26.080 173.985 ;
        RECT 22.985 172.355 23.320 172.525 ;
        RECT 23.515 172.355 24.190 172.525 ;
        RECT 24.510 172.075 24.880 172.575 ;
        RECT 25.060 172.525 25.230 172.755 ;
        RECT 25.615 172.695 26.080 173.025 ;
        RECT 26.250 173.315 26.420 174.155 ;
        RECT 26.600 174.125 26.915 174.625 ;
        RECT 27.145 173.895 27.485 174.455 ;
        RECT 26.590 173.520 27.485 173.895 ;
        RECT 27.655 173.615 27.825 174.625 ;
        RECT 27.295 173.315 27.485 173.520 ;
        RECT 27.995 173.565 28.325 174.410 ;
        RECT 28.565 173.655 28.895 174.440 ;
        RECT 27.995 173.485 28.385 173.565 ;
        RECT 28.565 173.485 29.245 173.655 ;
        RECT 29.425 173.485 29.755 174.625 ;
        RECT 28.170 173.435 28.385 173.485 ;
        RECT 26.250 172.985 27.125 173.315 ;
        RECT 27.295 172.985 28.045 173.315 ;
        RECT 26.250 172.525 26.420 172.985 ;
        RECT 27.295 172.815 27.495 172.985 ;
        RECT 28.215 172.855 28.385 173.435 ;
        RECT 28.555 173.065 28.905 173.315 ;
        RECT 29.075 172.885 29.245 173.485 ;
        RECT 30.395 173.460 30.685 174.625 ;
        RECT 30.855 173.535 32.525 174.625 ;
        RECT 29.415 173.065 29.765 173.315 ;
        RECT 28.160 172.815 28.385 172.855 ;
        RECT 25.060 172.355 25.465 172.525 ;
        RECT 25.635 172.355 26.420 172.525 ;
        RECT 26.695 172.075 26.905 172.605 ;
        RECT 27.165 172.290 27.495 172.815 ;
        RECT 28.005 172.730 28.385 172.815 ;
        RECT 27.665 172.075 27.835 172.685 ;
        RECT 28.005 172.295 28.335 172.730 ;
        RECT 28.575 172.075 28.815 172.885 ;
        RECT 28.985 172.245 29.315 172.885 ;
        RECT 29.485 172.075 29.755 172.885 ;
        RECT 30.855 172.845 31.605 173.365 ;
        RECT 31.775 173.015 32.525 173.535 ;
        RECT 33.245 173.695 33.415 174.455 ;
        RECT 33.630 173.865 33.960 174.625 ;
        RECT 33.245 173.525 33.960 173.695 ;
        RECT 34.130 173.550 34.385 174.455 ;
        RECT 33.155 172.975 33.510 173.345 ;
        RECT 33.790 173.315 33.960 173.525 ;
        RECT 33.790 172.985 34.045 173.315 ;
        RECT 30.395 172.075 30.685 172.800 ;
        RECT 30.855 172.075 32.525 172.845 ;
        RECT 33.790 172.795 33.960 172.985 ;
        RECT 34.215 172.820 34.385 173.550 ;
        RECT 34.560 173.475 34.820 174.625 ;
        RECT 35.495 174.165 35.710 174.625 ;
        RECT 35.880 173.995 36.210 174.455 ;
        RECT 35.040 173.825 36.210 173.995 ;
        RECT 36.380 173.825 36.630 174.625 ;
        RECT 37.305 173.905 37.635 174.625 ;
        RECT 33.245 172.625 33.960 172.795 ;
        RECT 33.245 172.245 33.415 172.625 ;
        RECT 33.630 172.075 33.960 172.455 ;
        RECT 34.130 172.245 34.385 172.820 ;
        RECT 34.560 172.075 34.820 172.915 ;
        RECT 35.040 172.535 35.410 173.825 ;
        RECT 36.840 173.655 37.120 173.815 ;
        RECT 35.785 173.485 37.120 173.655 ;
        RECT 35.785 173.315 35.955 173.485 ;
        RECT 35.580 173.065 35.955 173.315 ;
        RECT 36.125 173.065 36.600 173.305 ;
        RECT 36.770 173.065 37.120 173.305 ;
        RECT 37.295 173.265 37.525 173.605 ;
        RECT 37.815 173.265 38.030 174.380 ;
        RECT 38.225 173.680 38.555 174.455 ;
        RECT 38.725 173.850 39.435 174.625 ;
        RECT 38.225 173.465 39.375 173.680 ;
        RECT 37.295 173.065 37.625 173.265 ;
        RECT 37.815 173.085 38.265 173.265 ;
        RECT 37.935 173.065 38.265 173.085 ;
        RECT 38.435 173.065 38.905 173.295 ;
        RECT 35.785 172.895 35.955 173.065 ;
        RECT 39.090 172.895 39.375 173.465 ;
        RECT 39.605 173.020 39.885 174.455 ;
        RECT 35.785 172.725 37.120 172.895 ;
        RECT 35.040 172.245 35.790 172.535 ;
        RECT 36.300 172.075 36.630 172.535 ;
        RECT 36.850 172.515 37.120 172.725 ;
        RECT 37.295 172.705 38.475 172.895 ;
        RECT 37.295 172.245 37.635 172.705 ;
        RECT 38.145 172.625 38.475 172.705 ;
        RECT 38.665 172.705 39.375 172.895 ;
        RECT 38.665 172.565 38.965 172.705 ;
        RECT 38.650 172.555 38.965 172.565 ;
        RECT 38.640 172.545 38.965 172.555 ;
        RECT 38.630 172.540 38.965 172.545 ;
        RECT 37.805 172.075 37.975 172.535 ;
        RECT 38.625 172.530 38.965 172.540 ;
        RECT 38.620 172.525 38.965 172.530 ;
        RECT 38.615 172.515 38.965 172.525 ;
        RECT 38.610 172.510 38.965 172.515 ;
        RECT 38.605 172.245 38.965 172.510 ;
        RECT 39.205 172.075 39.375 172.535 ;
        RECT 39.545 172.245 39.885 173.020 ;
        RECT 40.055 172.355 40.335 174.455 ;
        RECT 40.525 173.865 41.310 174.625 ;
        RECT 41.705 173.795 42.090 174.455 ;
        RECT 41.705 173.695 42.115 173.795 ;
        RECT 40.505 173.485 42.115 173.695 ;
        RECT 42.415 173.605 42.615 174.395 ;
        RECT 40.505 172.885 40.780 173.485 ;
        RECT 42.285 173.435 42.615 173.605 ;
        RECT 42.785 173.445 43.105 174.625 ;
        RECT 43.330 173.755 43.615 174.625 ;
        RECT 43.785 173.995 44.045 174.455 ;
        RECT 44.220 174.165 44.475 174.625 ;
        RECT 44.645 173.995 44.905 174.455 ;
        RECT 43.785 173.825 44.905 173.995 ;
        RECT 45.075 173.825 45.385 174.625 ;
        RECT 43.785 173.575 44.045 173.825 ;
        RECT 45.555 173.655 45.865 174.455 ;
        RECT 42.285 173.315 42.465 173.435 ;
        RECT 40.950 173.065 41.305 173.315 ;
        RECT 41.500 173.265 41.965 173.315 ;
        RECT 41.495 173.095 41.965 173.265 ;
        RECT 41.500 173.065 41.965 173.095 ;
        RECT 42.135 173.065 42.465 173.315 ;
        RECT 43.290 173.405 44.045 173.575 ;
        RECT 44.835 173.485 45.865 173.655 ;
        RECT 42.640 173.065 43.105 173.265 ;
        RECT 43.290 172.895 43.695 173.405 ;
        RECT 44.835 173.235 45.005 173.485 ;
        RECT 43.865 173.065 45.005 173.235 ;
        RECT 40.505 172.705 41.755 172.885 ;
        RECT 41.390 172.635 41.755 172.705 ;
        RECT 41.925 172.685 43.105 172.855 ;
        RECT 43.290 172.725 44.940 172.895 ;
        RECT 45.175 172.745 45.525 173.315 ;
        RECT 40.565 172.075 40.735 172.535 ;
        RECT 41.925 172.465 42.255 172.685 ;
        RECT 41.005 172.285 42.255 172.465 ;
        RECT 42.425 172.075 42.595 172.515 ;
        RECT 42.765 172.270 43.105 172.685 ;
        RECT 43.335 172.075 43.615 172.555 ;
        RECT 43.785 172.335 44.045 172.725 ;
        RECT 44.220 172.075 44.475 172.555 ;
        RECT 44.645 172.335 44.940 172.725 ;
        RECT 45.695 172.575 45.865 173.485 ;
        RECT 45.120 172.075 45.395 172.555 ;
        RECT 45.565 172.245 45.865 172.575 ;
        RECT 46.035 173.905 46.495 174.455 ;
        RECT 46.685 173.905 47.015 174.625 ;
        RECT 46.035 172.535 46.285 173.905 ;
        RECT 47.215 173.735 47.515 174.285 ;
        RECT 47.685 173.955 47.965 174.625 ;
        RECT 46.575 173.565 47.515 173.735 ;
        RECT 46.575 173.315 46.745 173.565 ;
        RECT 47.885 173.315 48.150 173.675 ;
        RECT 48.855 173.565 49.185 174.410 ;
        RECT 49.355 173.615 49.525 174.625 ;
        RECT 49.695 173.895 50.035 174.455 ;
        RECT 50.265 174.125 50.580 174.625 ;
        RECT 50.760 174.155 51.645 174.325 ;
        RECT 46.455 172.985 46.745 173.315 ;
        RECT 46.915 173.065 47.255 173.315 ;
        RECT 47.475 173.065 48.150 173.315 ;
        RECT 48.795 173.485 49.185 173.565 ;
        RECT 49.695 173.520 50.590 173.895 ;
        RECT 48.795 173.435 49.010 173.485 ;
        RECT 46.575 172.895 46.745 172.985 ;
        RECT 46.575 172.705 47.965 172.895 ;
        RECT 48.795 172.855 48.965 173.435 ;
        RECT 49.695 173.315 49.885 173.520 ;
        RECT 50.760 173.315 50.930 174.155 ;
        RECT 51.870 174.125 52.120 174.455 ;
        RECT 49.135 172.985 49.885 173.315 ;
        RECT 50.055 172.985 50.930 173.315 ;
        RECT 48.795 172.815 49.020 172.855 ;
        RECT 49.685 172.815 49.885 172.985 ;
        RECT 48.795 172.730 49.175 172.815 ;
        RECT 46.035 172.245 46.595 172.535 ;
        RECT 46.765 172.075 47.015 172.535 ;
        RECT 47.635 172.345 47.965 172.705 ;
        RECT 48.845 172.295 49.175 172.730 ;
        RECT 49.345 172.075 49.515 172.685 ;
        RECT 49.685 172.290 50.015 172.815 ;
        RECT 50.275 172.075 50.485 172.605 ;
        RECT 50.760 172.525 50.930 172.985 ;
        RECT 51.100 173.025 51.420 173.985 ;
        RECT 51.590 173.235 51.780 173.955 ;
        RECT 51.950 173.055 52.120 174.125 ;
        RECT 52.290 173.825 52.460 174.625 ;
        RECT 52.630 174.180 53.735 174.350 ;
        RECT 52.630 173.565 52.800 174.180 ;
        RECT 53.945 174.030 54.195 174.455 ;
        RECT 54.365 174.165 54.630 174.625 ;
        RECT 52.970 173.645 53.500 174.010 ;
        RECT 53.945 173.900 54.250 174.030 ;
        RECT 52.290 173.475 52.800 173.565 ;
        RECT 52.290 173.305 53.160 173.475 ;
        RECT 52.290 173.235 52.460 173.305 ;
        RECT 52.580 173.055 52.780 173.085 ;
        RECT 51.100 172.695 51.565 173.025 ;
        RECT 51.950 172.755 52.780 173.055 ;
        RECT 51.950 172.525 52.120 172.755 ;
        RECT 50.760 172.355 51.545 172.525 ;
        RECT 51.715 172.355 52.120 172.525 ;
        RECT 52.300 172.075 52.670 172.575 ;
        RECT 52.990 172.525 53.160 173.305 ;
        RECT 53.330 172.945 53.500 173.645 ;
        RECT 53.670 173.115 53.910 173.710 ;
        RECT 53.330 172.725 53.855 172.945 ;
        RECT 54.080 172.795 54.250 173.900 ;
        RECT 54.025 172.665 54.250 172.795 ;
        RECT 54.420 172.705 54.700 173.655 ;
        RECT 54.025 172.525 54.195 172.665 ;
        RECT 52.990 172.355 53.665 172.525 ;
        RECT 53.860 172.355 54.195 172.525 ;
        RECT 54.365 172.075 54.615 172.535 ;
        RECT 54.870 172.335 55.055 174.455 ;
        RECT 55.225 174.125 55.555 174.625 ;
        RECT 55.725 173.955 55.895 174.455 ;
        RECT 55.230 173.785 55.895 173.955 ;
        RECT 55.230 172.795 55.460 173.785 ;
        RECT 55.630 172.965 55.980 173.615 ;
        RECT 56.155 173.460 56.445 174.625 ;
        RECT 56.615 174.195 56.955 174.455 ;
        RECT 55.230 172.625 55.895 172.795 ;
        RECT 55.225 172.075 55.555 172.455 ;
        RECT 55.725 172.335 55.895 172.625 ;
        RECT 56.155 172.075 56.445 172.800 ;
        RECT 56.615 172.795 56.875 174.195 ;
        RECT 57.125 173.825 57.455 174.625 ;
        RECT 57.920 173.655 58.170 174.455 ;
        RECT 58.355 173.905 58.685 174.625 ;
        RECT 58.905 173.655 59.155 174.455 ;
        RECT 59.325 174.245 59.660 174.625 ;
        RECT 57.065 173.485 59.255 173.655 ;
        RECT 57.065 173.315 57.380 173.485 ;
        RECT 57.050 173.065 57.380 173.315 ;
        RECT 56.615 172.285 56.955 172.795 ;
        RECT 57.125 172.075 57.395 172.875 ;
        RECT 57.575 172.345 57.855 173.315 ;
        RECT 58.035 172.345 58.335 173.315 ;
        RECT 58.515 172.350 58.865 173.315 ;
        RECT 59.085 172.575 59.255 173.485 ;
        RECT 59.425 172.755 59.665 174.065 ;
        RECT 59.835 173.535 61.045 174.625 ;
        RECT 61.305 173.955 61.475 174.455 ;
        RECT 61.645 174.125 61.975 174.625 ;
        RECT 61.305 173.785 61.970 173.955 ;
        RECT 59.835 172.825 60.355 173.365 ;
        RECT 60.525 172.995 61.045 173.535 ;
        RECT 61.220 172.965 61.570 173.615 ;
        RECT 59.085 172.245 59.580 172.575 ;
        RECT 59.835 172.075 61.045 172.825 ;
        RECT 61.740 172.795 61.970 173.785 ;
        RECT 61.305 172.625 61.970 172.795 ;
        RECT 61.305 172.335 61.475 172.625 ;
        RECT 61.645 172.075 61.975 172.455 ;
        RECT 62.145 172.335 62.330 174.455 ;
        RECT 62.570 174.165 62.835 174.625 ;
        RECT 63.005 174.030 63.255 174.455 ;
        RECT 63.465 174.180 64.570 174.350 ;
        RECT 62.950 173.900 63.255 174.030 ;
        RECT 62.500 172.705 62.780 173.655 ;
        RECT 62.950 172.795 63.120 173.900 ;
        RECT 63.290 173.115 63.530 173.710 ;
        RECT 63.700 173.645 64.230 174.010 ;
        RECT 63.700 172.945 63.870 173.645 ;
        RECT 64.400 173.565 64.570 174.180 ;
        RECT 64.740 173.825 64.910 174.625 ;
        RECT 65.080 174.125 65.330 174.455 ;
        RECT 65.555 174.155 66.440 174.325 ;
        RECT 64.400 173.475 64.910 173.565 ;
        RECT 62.950 172.665 63.175 172.795 ;
        RECT 63.345 172.725 63.870 172.945 ;
        RECT 64.040 173.305 64.910 173.475 ;
        RECT 62.585 172.075 62.835 172.535 ;
        RECT 63.005 172.525 63.175 172.665 ;
        RECT 64.040 172.525 64.210 173.305 ;
        RECT 64.740 173.235 64.910 173.305 ;
        RECT 64.420 173.055 64.620 173.085 ;
        RECT 65.080 173.055 65.250 174.125 ;
        RECT 65.420 173.235 65.610 173.955 ;
        RECT 64.420 172.755 65.250 173.055 ;
        RECT 65.780 173.025 66.100 173.985 ;
        RECT 63.005 172.355 63.340 172.525 ;
        RECT 63.535 172.355 64.210 172.525 ;
        RECT 64.530 172.075 64.900 172.575 ;
        RECT 65.080 172.525 65.250 172.755 ;
        RECT 65.635 172.695 66.100 173.025 ;
        RECT 66.270 173.315 66.440 174.155 ;
        RECT 66.620 174.125 66.935 174.625 ;
        RECT 67.165 173.895 67.505 174.455 ;
        RECT 66.610 173.520 67.505 173.895 ;
        RECT 67.675 173.615 67.845 174.625 ;
        RECT 67.315 173.315 67.505 173.520 ;
        RECT 68.015 173.565 68.345 174.410 ;
        RECT 68.015 173.485 68.405 173.565 ;
        RECT 68.575 173.485 68.855 174.625 ;
        RECT 68.190 173.435 68.405 173.485 ;
        RECT 69.025 173.475 69.355 174.455 ;
        RECT 69.525 173.485 69.785 174.625 ;
        RECT 69.955 173.535 71.165 174.625 ;
        RECT 66.270 172.985 67.145 173.315 ;
        RECT 67.315 172.985 68.065 173.315 ;
        RECT 66.270 172.525 66.440 172.985 ;
        RECT 67.315 172.815 67.515 172.985 ;
        RECT 68.235 172.855 68.405 173.435 ;
        RECT 68.585 173.045 68.920 173.315 ;
        RECT 69.090 172.875 69.260 173.475 ;
        RECT 69.430 173.065 69.765 173.315 ;
        RECT 68.180 172.815 68.405 172.855 ;
        RECT 65.080 172.355 65.485 172.525 ;
        RECT 65.655 172.355 66.440 172.525 ;
        RECT 66.715 172.075 66.925 172.605 ;
        RECT 67.185 172.290 67.515 172.815 ;
        RECT 68.025 172.730 68.405 172.815 ;
        RECT 67.685 172.075 67.855 172.685 ;
        RECT 68.025 172.295 68.355 172.730 ;
        RECT 68.575 172.075 68.885 172.875 ;
        RECT 69.090 172.245 69.785 172.875 ;
        RECT 69.955 172.825 70.475 173.365 ;
        RECT 70.645 172.995 71.165 173.535 ;
        RECT 71.335 173.485 71.720 174.455 ;
        RECT 71.890 174.165 72.215 174.625 ;
        RECT 72.735 173.995 73.015 174.455 ;
        RECT 71.890 173.775 73.015 173.995 ;
        RECT 69.955 172.075 71.165 172.825 ;
        RECT 71.335 172.815 71.615 173.485 ;
        RECT 71.890 173.315 72.340 173.775 ;
        RECT 73.205 173.605 73.605 174.455 ;
        RECT 74.005 174.165 74.275 174.625 ;
        RECT 74.445 173.995 74.730 174.455 ;
        RECT 71.785 172.985 72.340 173.315 ;
        RECT 72.510 173.045 73.605 173.605 ;
        RECT 71.890 172.875 72.340 172.985 ;
        RECT 71.335 172.245 71.720 172.815 ;
        RECT 71.890 172.705 73.015 172.875 ;
        RECT 71.890 172.075 72.215 172.535 ;
        RECT 72.735 172.245 73.015 172.705 ;
        RECT 73.205 172.245 73.605 173.045 ;
        RECT 73.775 173.775 74.730 173.995 ;
        RECT 73.775 172.875 73.985 173.775 ;
        RECT 74.155 173.045 74.845 173.605 ;
        RECT 75.015 173.485 75.400 174.445 ;
        RECT 75.615 173.825 75.905 174.625 ;
        RECT 76.075 174.285 77.440 174.455 ;
        RECT 76.075 173.655 76.245 174.285 ;
        RECT 75.570 173.485 76.245 173.655 ;
        RECT 73.775 172.705 74.730 172.875 ;
        RECT 74.005 172.075 74.275 172.535 ;
        RECT 74.445 172.245 74.730 172.705 ;
        RECT 75.015 172.815 75.190 173.485 ;
        RECT 75.570 173.315 75.740 173.485 ;
        RECT 76.415 173.315 76.740 174.115 ;
        RECT 77.110 174.075 77.440 174.285 ;
        RECT 77.110 173.825 78.065 174.075 ;
        RECT 75.375 173.065 75.740 173.315 ;
        RECT 75.935 173.065 76.185 173.315 ;
        RECT 75.375 172.985 75.565 173.065 ;
        RECT 75.935 172.985 76.105 173.065 ;
        RECT 76.395 172.985 76.740 173.315 ;
        RECT 76.910 172.985 77.185 173.650 ;
        RECT 77.370 172.985 77.725 173.650 ;
        RECT 77.895 172.815 78.065 173.825 ;
        RECT 78.235 173.485 78.525 174.625 ;
        RECT 78.695 173.485 78.970 174.455 ;
        RECT 79.180 173.825 79.460 174.625 ;
        RECT 79.630 174.115 81.245 174.445 ;
        RECT 79.630 173.775 80.805 173.945 ;
        RECT 79.630 173.655 79.800 173.775 ;
        RECT 79.140 173.485 79.800 173.655 ;
        RECT 78.250 172.985 78.525 173.315 ;
        RECT 75.015 172.245 75.525 172.815 ;
        RECT 76.070 172.645 77.470 172.815 ;
        RECT 75.695 172.075 75.865 172.635 ;
        RECT 76.070 172.245 76.400 172.645 ;
        RECT 76.575 172.075 76.905 172.475 ;
        RECT 77.140 172.455 77.470 172.645 ;
        RECT 77.640 172.625 78.065 172.815 ;
        RECT 78.695 172.750 78.865 173.485 ;
        RECT 79.140 173.315 79.310 173.485 ;
        RECT 80.060 173.315 80.305 173.605 ;
        RECT 80.475 173.485 80.805 173.775 ;
        RECT 81.065 173.315 81.235 173.875 ;
        RECT 81.485 173.485 81.745 174.625 ;
        RECT 81.915 173.460 82.205 174.625 ;
        RECT 82.835 173.865 83.350 174.275 ;
        RECT 83.585 173.865 83.755 174.625 ;
        RECT 83.925 174.285 85.955 174.455 ;
        RECT 79.035 172.985 79.310 173.315 ;
        RECT 79.480 172.985 80.305 173.315 ;
        RECT 80.520 172.985 81.235 173.315 ;
        RECT 81.405 173.065 81.740 173.315 ;
        RECT 79.140 172.815 79.310 172.985 ;
        RECT 80.985 172.895 81.235 172.985 ;
        RECT 82.835 173.055 83.175 173.865 ;
        RECT 83.925 173.620 84.095 174.285 ;
        RECT 84.490 173.945 85.615 174.115 ;
        RECT 83.345 173.430 84.095 173.620 ;
        RECT 84.265 173.605 85.275 173.775 ;
        RECT 78.235 172.455 78.525 172.725 ;
        RECT 77.140 172.245 78.525 172.455 ;
        RECT 78.695 172.405 78.970 172.750 ;
        RECT 79.140 172.645 80.805 172.815 ;
        RECT 79.160 172.075 79.535 172.475 ;
        RECT 79.705 172.295 79.875 172.645 ;
        RECT 80.045 172.075 80.375 172.475 ;
        RECT 80.545 172.245 80.805 172.645 ;
        RECT 80.985 172.475 81.315 172.895 ;
        RECT 81.485 172.075 81.745 172.895 ;
        RECT 82.835 172.885 84.065 173.055 ;
        RECT 81.915 172.075 82.205 172.800 ;
        RECT 83.110 172.280 83.355 172.885 ;
        RECT 83.575 172.075 84.085 172.610 ;
        RECT 84.265 172.245 84.455 173.605 ;
        RECT 84.625 172.925 84.900 173.405 ;
        RECT 84.625 172.755 84.905 172.925 ;
        RECT 85.105 172.805 85.275 173.605 ;
        RECT 85.445 172.815 85.615 173.945 ;
        RECT 85.785 173.315 85.955 174.285 ;
        RECT 86.125 173.485 86.295 174.625 ;
        RECT 86.465 173.485 86.800 174.455 ;
        RECT 86.985 173.655 87.315 174.440 ;
        RECT 86.985 173.485 87.665 173.655 ;
        RECT 87.845 173.485 88.175 174.625 ;
        RECT 88.355 174.190 93.700 174.625 ;
        RECT 85.785 172.985 85.980 173.315 ;
        RECT 86.205 172.985 86.460 173.315 ;
        RECT 86.205 172.815 86.375 172.985 ;
        RECT 86.630 172.815 86.800 173.485 ;
        RECT 86.975 173.065 87.325 173.315 ;
        RECT 87.495 172.885 87.665 173.485 ;
        RECT 87.835 173.065 88.185 173.315 ;
        RECT 84.625 172.245 84.900 172.755 ;
        RECT 85.445 172.645 86.375 172.815 ;
        RECT 85.445 172.610 85.620 172.645 ;
        RECT 85.090 172.245 85.620 172.610 ;
        RECT 86.045 172.075 86.375 172.475 ;
        RECT 86.545 172.245 86.800 172.815 ;
        RECT 86.995 172.075 87.235 172.885 ;
        RECT 87.405 172.245 87.735 172.885 ;
        RECT 87.905 172.075 88.175 172.885 ;
        RECT 89.940 172.620 90.280 173.450 ;
        RECT 91.760 172.940 92.110 174.190 ;
        RECT 93.875 173.535 95.085 174.625 ;
        RECT 93.875 172.825 94.395 173.365 ;
        RECT 94.565 172.995 95.085 173.535 ;
        RECT 95.260 173.485 95.595 174.455 ;
        RECT 95.765 173.485 95.935 174.625 ;
        RECT 96.105 174.285 98.135 174.455 ;
        RECT 88.355 172.075 93.700 172.620 ;
        RECT 93.875 172.075 95.085 172.825 ;
        RECT 95.260 172.815 95.430 173.485 ;
        RECT 96.105 173.315 96.275 174.285 ;
        RECT 95.600 172.985 95.855 173.315 ;
        RECT 96.080 172.985 96.275 173.315 ;
        RECT 96.445 173.945 97.570 174.115 ;
        RECT 95.685 172.815 95.855 172.985 ;
        RECT 96.445 172.815 96.615 173.945 ;
        RECT 95.260 172.245 95.515 172.815 ;
        RECT 95.685 172.645 96.615 172.815 ;
        RECT 96.785 173.605 97.795 173.775 ;
        RECT 96.785 172.805 96.955 173.605 ;
        RECT 97.160 173.265 97.435 173.405 ;
        RECT 97.155 173.095 97.435 173.265 ;
        RECT 96.440 172.610 96.615 172.645 ;
        RECT 95.685 172.075 96.015 172.475 ;
        RECT 96.440 172.245 96.970 172.610 ;
        RECT 97.160 172.245 97.435 173.095 ;
        RECT 97.605 172.245 97.795 173.605 ;
        RECT 97.965 173.620 98.135 174.285 ;
        RECT 98.305 173.865 98.475 174.625 ;
        RECT 98.710 173.865 99.225 174.275 ;
        RECT 97.965 173.430 98.715 173.620 ;
        RECT 98.885 173.055 99.225 173.865 ;
        RECT 97.995 172.885 99.225 173.055 ;
        RECT 99.395 173.485 99.780 174.455 ;
        RECT 99.950 174.165 100.275 174.625 ;
        RECT 100.795 173.995 101.075 174.455 ;
        RECT 99.950 173.775 101.075 173.995 ;
        RECT 97.975 172.075 98.485 172.610 ;
        RECT 98.705 172.280 98.950 172.885 ;
        RECT 99.395 172.815 99.675 173.485 ;
        RECT 99.950 173.315 100.400 173.775 ;
        RECT 101.265 173.605 101.665 174.455 ;
        RECT 102.065 174.165 102.335 174.625 ;
        RECT 102.505 173.995 102.790 174.455 ;
        RECT 99.845 172.985 100.400 173.315 ;
        RECT 100.570 173.045 101.665 173.605 ;
        RECT 99.950 172.875 100.400 172.985 ;
        RECT 99.395 172.245 99.780 172.815 ;
        RECT 99.950 172.705 101.075 172.875 ;
        RECT 99.950 172.075 100.275 172.535 ;
        RECT 100.795 172.245 101.075 172.705 ;
        RECT 101.265 172.245 101.665 173.045 ;
        RECT 101.835 173.775 102.790 173.995 ;
        RECT 103.190 173.995 103.475 174.455 ;
        RECT 103.645 174.165 103.915 174.625 ;
        RECT 103.190 173.775 104.145 173.995 ;
        RECT 101.835 172.875 102.045 173.775 ;
        RECT 102.215 173.045 102.905 173.605 ;
        RECT 103.075 173.045 103.765 173.605 ;
        RECT 103.935 172.875 104.145 173.775 ;
        RECT 101.835 172.705 102.790 172.875 ;
        RECT 102.065 172.075 102.335 172.535 ;
        RECT 102.505 172.245 102.790 172.705 ;
        RECT 103.190 172.705 104.145 172.875 ;
        RECT 104.315 173.605 104.715 174.455 ;
        RECT 104.905 173.995 105.185 174.455 ;
        RECT 105.705 174.165 106.030 174.625 ;
        RECT 104.905 173.775 106.030 173.995 ;
        RECT 104.315 173.045 105.410 173.605 ;
        RECT 105.580 173.315 106.030 173.775 ;
        RECT 106.200 173.485 106.585 174.455 ;
        RECT 103.190 172.245 103.475 172.705 ;
        RECT 103.645 172.075 103.915 172.535 ;
        RECT 104.315 172.245 104.715 173.045 ;
        RECT 105.580 172.985 106.135 173.315 ;
        RECT 105.580 172.875 106.030 172.985 ;
        RECT 104.905 172.705 106.030 172.875 ;
        RECT 106.305 172.815 106.585 173.485 ;
        RECT 107.675 173.460 107.965 174.625 ;
        RECT 108.175 174.285 109.315 174.455 ;
        RECT 108.175 173.825 108.475 174.285 ;
        RECT 108.645 173.655 108.975 174.115 ;
        RECT 104.905 172.245 105.185 172.705 ;
        RECT 105.705 172.075 106.030 172.535 ;
        RECT 106.200 172.245 106.585 172.815 ;
        RECT 108.215 173.435 108.975 173.655 ;
        RECT 109.145 173.655 109.315 174.285 ;
        RECT 109.485 173.825 109.815 174.625 ;
        RECT 109.985 173.655 110.260 174.455 ;
        RECT 109.145 173.445 110.260 173.655 ;
        RECT 110.445 173.655 110.775 174.440 ;
        RECT 110.445 173.485 111.125 173.655 ;
        RECT 111.305 173.485 111.635 174.625 ;
        RECT 111.815 173.485 112.075 174.625 ;
        RECT 108.215 172.895 108.430 173.435 ;
        RECT 108.600 173.065 109.370 173.265 ;
        RECT 109.540 173.065 110.260 173.265 ;
        RECT 110.435 173.065 110.785 173.315 ;
        RECT 107.675 172.075 107.965 172.800 ;
        RECT 108.215 172.725 109.815 172.895 ;
        RECT 108.645 172.715 109.815 172.725 ;
        RECT 108.185 172.075 108.475 172.545 ;
        RECT 108.645 172.245 108.975 172.715 ;
        RECT 109.145 172.075 109.315 172.545 ;
        RECT 109.485 172.245 109.815 172.715 ;
        RECT 109.985 172.075 110.260 172.895 ;
        RECT 110.955 172.885 111.125 173.485 ;
        RECT 112.245 173.475 112.575 174.455 ;
        RECT 112.745 173.485 113.025 174.625 ;
        RECT 113.655 174.115 114.845 174.405 ;
        RECT 113.675 173.775 114.845 173.945 ;
        RECT 115.015 173.825 115.295 174.625 ;
        RECT 113.675 173.485 114.000 173.775 ;
        RECT 114.675 173.655 114.845 173.775 ;
        RECT 111.295 173.065 111.645 173.315 ;
        RECT 111.835 173.065 112.170 173.315 ;
        RECT 110.455 172.075 110.695 172.885 ;
        RECT 110.865 172.245 111.195 172.885 ;
        RECT 111.365 172.075 111.635 172.885 ;
        RECT 112.340 172.875 112.510 173.475 ;
        RECT 114.170 173.315 114.365 173.605 ;
        RECT 114.675 173.485 115.335 173.655 ;
        RECT 115.505 173.485 115.780 174.455 ;
        RECT 115.165 173.315 115.335 173.485 ;
        RECT 112.680 173.045 113.015 173.315 ;
        RECT 113.655 172.985 114.000 173.315 ;
        RECT 114.170 172.985 114.995 173.315 ;
        RECT 115.165 172.985 115.440 173.315 ;
        RECT 111.815 172.245 112.510 172.875 ;
        RECT 112.715 172.075 113.025 172.875 ;
        RECT 115.165 172.815 115.335 172.985 ;
        RECT 113.670 172.645 115.335 172.815 ;
        RECT 115.610 172.750 115.780 173.485 ;
        RECT 116.110 173.615 116.410 174.455 ;
        RECT 116.605 173.785 116.855 174.625 ;
        RECT 117.445 174.035 118.250 174.455 ;
        RECT 117.025 173.865 118.590 174.035 ;
        RECT 117.025 173.615 117.195 173.865 ;
        RECT 116.110 173.445 117.195 173.615 ;
        RECT 115.955 172.985 116.285 173.275 ;
        RECT 116.455 172.815 116.625 173.445 ;
        RECT 117.365 173.315 117.685 173.695 ;
        RECT 117.875 173.605 118.250 173.695 ;
        RECT 117.855 173.435 118.250 173.605 ;
        RECT 118.420 173.615 118.590 173.865 ;
        RECT 118.760 173.785 119.090 174.625 ;
        RECT 119.260 173.865 119.925 174.455 ;
        RECT 120.095 174.115 121.285 174.405 ;
        RECT 118.420 173.445 119.340 173.615 ;
        RECT 116.795 173.065 117.125 173.275 ;
        RECT 117.305 173.065 117.685 173.315 ;
        RECT 117.875 173.275 118.250 173.435 ;
        RECT 119.170 173.275 119.340 173.445 ;
        RECT 117.875 173.065 118.360 173.275 ;
        RECT 118.550 173.065 119.000 173.275 ;
        RECT 119.170 173.065 119.505 173.275 ;
        RECT 119.675 172.895 119.925 173.865 ;
        RECT 120.115 173.775 121.285 173.945 ;
        RECT 121.455 173.825 121.735 174.625 ;
        RECT 120.115 173.485 120.440 173.775 ;
        RECT 121.115 173.655 121.285 173.775 ;
        RECT 120.610 173.315 120.805 173.605 ;
        RECT 121.115 173.485 121.775 173.655 ;
        RECT 121.945 173.485 122.220 174.455 ;
        RECT 122.580 173.655 122.970 173.830 ;
        RECT 123.455 173.825 123.785 174.625 ;
        RECT 123.955 173.835 124.490 174.455 ;
        RECT 122.580 173.485 124.005 173.655 ;
        RECT 121.605 173.315 121.775 173.485 ;
        RECT 120.095 172.985 120.440 173.315 ;
        RECT 120.610 172.985 121.435 173.315 ;
        RECT 121.605 172.985 121.880 173.315 ;
        RECT 113.670 172.295 113.925 172.645 ;
        RECT 114.095 172.075 114.425 172.475 ;
        RECT 114.595 172.295 114.765 172.645 ;
        RECT 114.935 172.075 115.315 172.475 ;
        RECT 115.505 172.405 115.780 172.750 ;
        RECT 116.115 172.635 116.625 172.815 ;
        RECT 117.030 172.725 118.730 172.895 ;
        RECT 117.030 172.635 117.415 172.725 ;
        RECT 116.115 172.245 116.445 172.635 ;
        RECT 116.615 172.295 117.800 172.465 ;
        RECT 118.060 172.075 118.230 172.545 ;
        RECT 118.400 172.260 118.730 172.725 ;
        RECT 118.900 172.075 119.070 172.895 ;
        RECT 119.240 172.255 119.925 172.895 ;
        RECT 121.605 172.815 121.775 172.985 ;
        RECT 120.110 172.645 121.775 172.815 ;
        RECT 122.050 172.750 122.220 173.485 ;
        RECT 122.455 172.755 122.810 173.315 ;
        RECT 120.110 172.295 120.365 172.645 ;
        RECT 120.535 172.075 120.865 172.475 ;
        RECT 121.035 172.295 121.205 172.645 ;
        RECT 121.375 172.075 121.755 172.475 ;
        RECT 121.945 172.405 122.220 172.750 ;
        RECT 122.980 172.585 123.150 173.485 ;
        RECT 123.320 172.755 123.585 173.315 ;
        RECT 123.835 172.985 124.005 173.485 ;
        RECT 124.175 172.815 124.490 173.835 ;
        RECT 124.695 173.535 125.905 174.625 ;
        RECT 122.560 172.075 122.800 172.585 ;
        RECT 122.980 172.255 123.260 172.585 ;
        RECT 123.490 172.075 123.705 172.585 ;
        RECT 123.875 172.245 124.490 172.815 ;
        RECT 124.695 172.825 125.215 173.365 ;
        RECT 125.385 172.995 125.905 173.535 ;
        RECT 126.080 174.235 126.415 174.455 ;
        RECT 127.420 174.245 127.775 174.625 ;
        RECT 126.080 173.615 126.335 174.235 ;
        RECT 126.585 174.075 126.815 174.115 ;
        RECT 127.945 174.075 128.195 174.455 ;
        RECT 126.585 173.875 128.195 174.075 ;
        RECT 126.585 173.785 126.770 173.875 ;
        RECT 127.360 173.865 128.195 173.875 ;
        RECT 128.445 173.845 128.695 174.625 ;
        RECT 128.865 173.775 129.125 174.455 ;
        RECT 126.925 173.675 127.255 173.705 ;
        RECT 126.925 173.615 128.725 173.675 ;
        RECT 126.080 173.505 128.785 173.615 ;
        RECT 126.080 173.445 127.255 173.505 ;
        RECT 128.585 173.470 128.785 173.505 ;
        RECT 126.075 173.065 126.565 173.265 ;
        RECT 126.755 173.065 127.230 173.275 ;
        RECT 124.695 172.075 125.905 172.825 ;
        RECT 126.080 172.075 126.535 172.840 ;
        RECT 127.010 172.665 127.230 173.065 ;
        RECT 127.475 173.065 127.805 173.275 ;
        RECT 127.475 172.665 127.685 173.065 ;
        RECT 127.975 173.030 128.385 173.335 ;
        RECT 128.615 172.895 128.785 173.470 ;
        RECT 128.515 172.775 128.785 172.895 ;
        RECT 127.940 172.730 128.785 172.775 ;
        RECT 127.940 172.605 128.695 172.730 ;
        RECT 127.940 172.455 128.110 172.605 ;
        RECT 128.955 172.575 129.125 173.775 ;
        RECT 129.295 173.865 129.810 174.275 ;
        RECT 130.045 173.865 130.215 174.625 ;
        RECT 130.385 174.285 132.415 174.455 ;
        RECT 129.295 173.055 129.635 173.865 ;
        RECT 130.385 173.620 130.555 174.285 ;
        RECT 130.950 173.945 132.075 174.115 ;
        RECT 129.805 173.430 130.555 173.620 ;
        RECT 130.725 173.605 131.735 173.775 ;
        RECT 129.295 172.885 130.525 173.055 ;
        RECT 126.810 172.245 128.110 172.455 ;
        RECT 128.365 172.075 128.695 172.435 ;
        RECT 128.865 172.245 129.125 172.575 ;
        RECT 129.570 172.280 129.815 172.885 ;
        RECT 130.035 172.075 130.545 172.610 ;
        RECT 130.725 172.245 130.915 173.605 ;
        RECT 131.085 173.265 131.360 173.405 ;
        RECT 131.085 173.095 131.365 173.265 ;
        RECT 131.085 172.245 131.360 173.095 ;
        RECT 131.565 172.805 131.735 173.605 ;
        RECT 131.905 172.815 132.075 173.945 ;
        RECT 132.245 173.315 132.415 174.285 ;
        RECT 132.585 173.485 132.755 174.625 ;
        RECT 132.925 173.485 133.260 174.455 ;
        RECT 132.245 172.985 132.440 173.315 ;
        RECT 132.665 172.985 132.920 173.315 ;
        RECT 132.665 172.815 132.835 172.985 ;
        RECT 133.090 172.815 133.260 173.485 ;
        RECT 133.435 173.460 133.725 174.625 ;
        RECT 133.985 173.955 134.155 174.455 ;
        RECT 134.325 174.125 134.655 174.625 ;
        RECT 133.985 173.785 134.650 173.955 ;
        RECT 133.900 172.965 134.250 173.615 ;
        RECT 131.905 172.645 132.835 172.815 ;
        RECT 131.905 172.610 132.080 172.645 ;
        RECT 131.550 172.245 132.080 172.610 ;
        RECT 132.505 172.075 132.835 172.475 ;
        RECT 133.005 172.245 133.260 172.815 ;
        RECT 133.435 172.075 133.725 172.800 ;
        RECT 134.420 172.795 134.650 173.785 ;
        RECT 133.985 172.625 134.650 172.795 ;
        RECT 133.985 172.335 134.155 172.625 ;
        RECT 134.325 172.075 134.655 172.455 ;
        RECT 134.825 172.335 135.010 174.455 ;
        RECT 135.250 174.165 135.515 174.625 ;
        RECT 135.685 174.030 135.935 174.455 ;
        RECT 136.145 174.180 137.250 174.350 ;
        RECT 135.630 173.900 135.935 174.030 ;
        RECT 135.180 172.705 135.460 173.655 ;
        RECT 135.630 172.795 135.800 173.900 ;
        RECT 135.970 173.115 136.210 173.710 ;
        RECT 136.380 173.645 136.910 174.010 ;
        RECT 136.380 172.945 136.550 173.645 ;
        RECT 137.080 173.565 137.250 174.180 ;
        RECT 137.420 173.825 137.590 174.625 ;
        RECT 137.760 174.125 138.010 174.455 ;
        RECT 138.235 174.155 139.120 174.325 ;
        RECT 137.080 173.475 137.590 173.565 ;
        RECT 135.630 172.665 135.855 172.795 ;
        RECT 136.025 172.725 136.550 172.945 ;
        RECT 136.720 173.305 137.590 173.475 ;
        RECT 135.265 172.075 135.515 172.535 ;
        RECT 135.685 172.525 135.855 172.665 ;
        RECT 136.720 172.525 136.890 173.305 ;
        RECT 137.420 173.235 137.590 173.305 ;
        RECT 137.100 173.055 137.300 173.085 ;
        RECT 137.760 173.055 137.930 174.125 ;
        RECT 138.100 173.235 138.290 173.955 ;
        RECT 137.100 172.755 137.930 173.055 ;
        RECT 138.460 173.025 138.780 173.985 ;
        RECT 135.685 172.355 136.020 172.525 ;
        RECT 136.215 172.355 136.890 172.525 ;
        RECT 137.210 172.075 137.580 172.575 ;
        RECT 137.760 172.525 137.930 172.755 ;
        RECT 138.315 172.695 138.780 173.025 ;
        RECT 138.950 173.315 139.120 174.155 ;
        RECT 139.300 174.125 139.615 174.625 ;
        RECT 139.845 173.895 140.185 174.455 ;
        RECT 139.290 173.520 140.185 173.895 ;
        RECT 140.355 173.615 140.525 174.625 ;
        RECT 139.995 173.315 140.185 173.520 ;
        RECT 140.695 173.565 141.025 174.410 ;
        RECT 140.695 173.485 141.085 173.565 ;
        RECT 140.870 173.435 141.085 173.485 ;
        RECT 138.950 172.985 139.825 173.315 ;
        RECT 139.995 172.985 140.745 173.315 ;
        RECT 138.950 172.525 139.120 172.985 ;
        RECT 139.995 172.815 140.195 172.985 ;
        RECT 140.915 172.855 141.085 173.435 ;
        RECT 141.715 173.535 142.925 174.625 ;
        RECT 141.715 172.995 142.235 173.535 ;
        RECT 140.860 172.815 141.085 172.855 ;
        RECT 142.405 172.825 142.925 173.365 ;
        RECT 137.760 172.355 138.165 172.525 ;
        RECT 138.335 172.355 139.120 172.525 ;
        RECT 139.395 172.075 139.605 172.605 ;
        RECT 139.865 172.290 140.195 172.815 ;
        RECT 140.705 172.730 141.085 172.815 ;
        RECT 140.365 172.075 140.535 172.685 ;
        RECT 140.705 172.295 141.035 172.730 ;
        RECT 141.715 172.075 142.925 172.825 ;
        RECT 17.430 171.905 143.010 172.075 ;
        RECT 17.515 171.155 18.725 171.905 ;
        RECT 17.515 170.615 18.035 171.155 ;
        RECT 18.895 171.135 20.565 171.905 ;
        RECT 18.205 170.445 18.725 170.985 ;
        RECT 18.895 170.615 19.645 171.135 ;
        RECT 20.745 171.095 21.015 171.905 ;
        RECT 21.185 171.095 21.515 171.735 ;
        RECT 21.685 171.095 21.925 171.905 ;
        RECT 22.120 171.650 22.455 171.695 ;
        RECT 22.115 171.185 22.455 171.650 ;
        RECT 22.625 171.525 22.955 171.905 ;
        RECT 23.415 171.565 23.685 171.570 ;
        RECT 23.415 171.395 23.725 171.565 ;
        RECT 19.815 170.445 20.565 170.965 ;
        RECT 20.735 170.665 21.085 170.915 ;
        RECT 21.255 170.495 21.425 171.095 ;
        RECT 21.595 170.665 21.945 170.915 ;
        RECT 22.115 170.495 22.285 171.185 ;
        RECT 22.455 170.665 22.715 170.995 ;
        RECT 17.515 169.355 18.725 170.445 ;
        RECT 18.895 169.355 20.565 170.445 ;
        RECT 20.745 169.355 21.075 170.495 ;
        RECT 21.255 170.325 21.935 170.495 ;
        RECT 21.605 169.540 21.935 170.325 ;
        RECT 22.115 169.525 22.375 170.495 ;
        RECT 22.545 170.115 22.715 170.665 ;
        RECT 22.885 170.295 23.225 171.325 ;
        RECT 23.415 170.295 23.685 171.395 ;
        RECT 23.910 170.295 24.190 171.570 ;
        RECT 24.390 171.405 24.620 171.735 ;
        RECT 24.865 171.525 25.195 171.905 ;
        RECT 24.390 170.115 24.560 171.405 ;
        RECT 25.365 171.335 25.540 171.735 ;
        RECT 24.910 171.165 25.540 171.335 ;
        RECT 25.795 171.255 26.055 171.735 ;
        RECT 26.225 171.365 26.475 171.905 ;
        RECT 24.910 170.995 25.080 171.165 ;
        RECT 24.730 170.665 25.080 170.995 ;
        RECT 22.545 169.945 24.560 170.115 ;
        RECT 24.910 170.145 25.080 170.665 ;
        RECT 25.260 170.315 25.625 170.995 ;
        RECT 25.795 170.225 25.965 171.255 ;
        RECT 26.645 171.225 26.865 171.685 ;
        RECT 26.615 171.200 26.865 171.225 ;
        RECT 26.135 170.605 26.365 171.000 ;
        RECT 26.535 170.775 26.865 171.200 ;
        RECT 27.035 171.525 27.925 171.695 ;
        RECT 27.035 170.800 27.205 171.525 ;
        RECT 28.180 171.405 28.675 171.735 ;
        RECT 27.375 170.970 27.925 171.355 ;
        RECT 27.035 170.730 27.925 170.800 ;
        RECT 27.030 170.705 27.925 170.730 ;
        RECT 27.020 170.690 27.925 170.705 ;
        RECT 27.015 170.675 27.925 170.690 ;
        RECT 27.005 170.670 27.925 170.675 ;
        RECT 27.000 170.660 27.925 170.670 ;
        RECT 26.995 170.650 27.925 170.660 ;
        RECT 26.985 170.645 27.925 170.650 ;
        RECT 26.975 170.635 27.925 170.645 ;
        RECT 26.965 170.630 27.925 170.635 ;
        RECT 26.965 170.625 27.300 170.630 ;
        RECT 26.950 170.620 27.300 170.625 ;
        RECT 26.935 170.610 27.300 170.620 ;
        RECT 26.910 170.605 27.300 170.610 ;
        RECT 26.135 170.600 27.300 170.605 ;
        RECT 26.135 170.565 27.270 170.600 ;
        RECT 26.135 170.540 27.235 170.565 ;
        RECT 26.135 170.510 27.205 170.540 ;
        RECT 26.135 170.480 27.185 170.510 ;
        RECT 26.135 170.450 27.165 170.480 ;
        RECT 26.135 170.440 27.095 170.450 ;
        RECT 26.135 170.430 27.070 170.440 ;
        RECT 26.135 170.415 27.050 170.430 ;
        RECT 26.135 170.400 27.030 170.415 ;
        RECT 26.240 170.390 27.025 170.400 ;
        RECT 26.240 170.355 27.010 170.390 ;
        RECT 24.910 169.975 25.540 170.145 ;
        RECT 22.570 169.355 22.900 169.765 ;
        RECT 23.100 169.525 23.270 169.945 ;
        RECT 23.485 169.355 24.155 169.765 ;
        RECT 24.390 169.525 24.560 169.945 ;
        RECT 24.865 169.355 25.195 169.795 ;
        RECT 25.365 169.525 25.540 169.975 ;
        RECT 25.795 169.525 26.070 170.225 ;
        RECT 26.240 170.105 26.995 170.355 ;
        RECT 27.165 170.035 27.495 170.280 ;
        RECT 27.665 170.180 27.925 170.630 ;
        RECT 27.310 170.010 27.495 170.035 ;
        RECT 27.310 169.910 27.925 170.010 ;
        RECT 28.095 169.915 28.335 171.225 ;
        RECT 28.505 170.495 28.675 171.405 ;
        RECT 28.895 170.665 29.245 171.630 ;
        RECT 29.425 170.665 29.725 171.635 ;
        RECT 29.905 170.665 30.185 171.635 ;
        RECT 30.365 171.105 30.635 171.905 ;
        RECT 30.805 171.185 31.145 171.695 ;
        RECT 30.380 170.665 30.710 170.915 ;
        RECT 30.380 170.495 30.695 170.665 ;
        RECT 28.505 170.325 30.695 170.495 ;
        RECT 26.240 169.355 26.495 169.900 ;
        RECT 26.665 169.525 27.145 169.865 ;
        RECT 27.320 169.355 27.925 169.910 ;
        RECT 28.100 169.355 28.435 169.735 ;
        RECT 28.605 169.525 28.855 170.325 ;
        RECT 29.075 169.355 29.405 170.075 ;
        RECT 29.590 169.525 29.840 170.325 ;
        RECT 30.305 169.355 30.635 170.155 ;
        RECT 30.885 169.785 31.145 171.185 ;
        RECT 31.315 171.135 33.905 171.905 ;
        RECT 31.315 170.615 32.525 171.135 ;
        RECT 34.280 171.125 34.780 171.735 ;
        RECT 32.695 170.445 33.905 170.965 ;
        RECT 34.075 170.665 34.425 170.915 ;
        RECT 34.610 170.495 34.780 171.125 ;
        RECT 35.410 171.255 35.740 171.735 ;
        RECT 35.910 171.445 36.135 171.905 ;
        RECT 36.305 171.255 36.635 171.735 ;
        RECT 35.410 171.085 36.635 171.255 ;
        RECT 36.825 171.105 37.075 171.905 ;
        RECT 37.245 171.105 37.585 171.735 ;
        RECT 38.460 171.425 38.760 171.905 ;
        RECT 38.930 171.255 39.190 171.710 ;
        RECT 39.360 171.425 39.620 171.905 ;
        RECT 39.790 171.255 40.050 171.710 ;
        RECT 40.220 171.425 40.480 171.905 ;
        RECT 40.650 171.255 40.910 171.710 ;
        RECT 41.080 171.425 41.340 171.905 ;
        RECT 41.510 171.255 41.770 171.710 ;
        RECT 41.940 171.380 42.200 171.905 ;
        RECT 34.950 170.715 35.280 170.915 ;
        RECT 35.450 170.715 35.780 170.915 ;
        RECT 35.950 170.715 36.370 170.915 ;
        RECT 36.545 170.745 37.240 170.915 ;
        RECT 36.545 170.495 36.715 170.745 ;
        RECT 37.410 170.495 37.585 171.105 ;
        RECT 30.805 169.525 31.145 169.785 ;
        RECT 31.315 169.355 33.905 170.445 ;
        RECT 34.280 170.325 36.715 170.495 ;
        RECT 34.280 169.525 34.610 170.325 ;
        RECT 34.780 169.355 35.110 170.155 ;
        RECT 35.410 169.525 35.740 170.325 ;
        RECT 36.385 169.355 36.635 170.155 ;
        RECT 36.905 169.355 37.075 170.495 ;
        RECT 37.245 169.525 37.585 170.495 ;
        RECT 38.460 171.085 41.770 171.255 ;
        RECT 38.460 170.495 39.430 171.085 ;
        RECT 42.370 170.915 42.620 171.725 ;
        RECT 42.800 171.445 43.045 171.905 ;
        RECT 39.600 170.665 42.620 170.915 ;
        RECT 42.790 170.665 43.105 171.275 ;
        RECT 43.275 171.180 43.565 171.905 ;
        RECT 43.745 171.255 44.075 171.730 ;
        RECT 44.245 171.425 44.415 171.905 ;
        RECT 44.585 171.255 44.915 171.730 ;
        RECT 45.085 171.425 45.255 171.905 ;
        RECT 45.425 171.255 45.755 171.730 ;
        RECT 45.925 171.425 46.095 171.905 ;
        RECT 46.265 171.255 46.595 171.730 ;
        RECT 46.765 171.425 46.935 171.905 ;
        RECT 47.105 171.255 47.435 171.730 ;
        RECT 47.605 171.425 47.775 171.905 ;
        RECT 47.945 171.730 48.195 171.735 ;
        RECT 47.945 171.255 48.275 171.730 ;
        RECT 48.445 171.425 48.615 171.905 ;
        RECT 48.865 171.730 49.035 171.735 ;
        RECT 48.785 171.255 49.115 171.730 ;
        RECT 49.285 171.425 49.455 171.905 ;
        RECT 49.705 171.730 49.875 171.735 ;
        RECT 49.625 171.255 49.955 171.730 ;
        RECT 50.125 171.425 50.295 171.905 ;
        RECT 50.465 171.255 50.795 171.730 ;
        RECT 50.965 171.425 51.135 171.905 ;
        RECT 51.305 171.255 51.635 171.730 ;
        RECT 51.805 171.425 51.975 171.905 ;
        RECT 52.145 171.255 52.475 171.730 ;
        RECT 52.645 171.425 52.815 171.905 ;
        RECT 52.985 171.255 53.315 171.730 ;
        RECT 53.485 171.425 53.655 171.905 ;
        RECT 53.825 171.255 54.155 171.730 ;
        RECT 54.325 171.425 54.495 171.905 ;
        RECT 55.020 171.425 55.320 171.905 ;
        RECT 55.490 171.255 55.750 171.710 ;
        RECT 55.920 171.425 56.180 171.905 ;
        RECT 56.350 171.255 56.610 171.710 ;
        RECT 56.780 171.425 57.040 171.905 ;
        RECT 57.210 171.255 57.470 171.710 ;
        RECT 57.640 171.425 57.900 171.905 ;
        RECT 58.070 171.255 58.330 171.710 ;
        RECT 58.500 171.380 58.760 171.905 ;
        RECT 43.745 171.085 45.255 171.255 ;
        RECT 45.425 171.085 47.775 171.255 ;
        RECT 47.945 171.085 54.605 171.255 ;
        RECT 45.085 170.915 45.255 171.085 ;
        RECT 47.600 170.915 47.775 171.085 ;
        RECT 43.740 170.715 44.915 170.915 ;
        RECT 45.085 170.715 47.395 170.915 ;
        RECT 47.600 170.715 54.160 170.915 ;
        RECT 38.460 170.255 41.770 170.495 ;
        RECT 38.465 169.355 38.760 170.085 ;
        RECT 38.930 169.530 39.190 170.255 ;
        RECT 39.360 169.355 39.620 170.085 ;
        RECT 39.790 169.530 40.050 170.255 ;
        RECT 40.220 169.355 40.480 170.085 ;
        RECT 40.650 169.530 40.910 170.255 ;
        RECT 41.080 169.355 41.340 170.085 ;
        RECT 41.510 169.530 41.770 170.255 ;
        RECT 41.940 169.355 42.200 170.465 ;
        RECT 42.370 169.530 42.620 170.665 ;
        RECT 45.085 170.545 45.255 170.715 ;
        RECT 47.600 170.545 47.775 170.715 ;
        RECT 54.330 170.545 54.605 171.085 ;
        RECT 42.800 169.355 43.095 170.465 ;
        RECT 43.275 169.355 43.565 170.520 ;
        RECT 43.745 170.375 45.255 170.545 ;
        RECT 45.425 170.375 47.775 170.545 ;
        RECT 47.945 170.375 54.605 170.545 ;
        RECT 55.020 171.085 58.330 171.255 ;
        RECT 55.020 170.495 55.990 171.085 ;
        RECT 58.930 170.915 59.180 171.725 ;
        RECT 59.360 171.445 59.605 171.905 ;
        RECT 56.160 170.665 59.180 170.915 ;
        RECT 59.350 170.665 59.665 171.275 ;
        RECT 59.855 171.095 60.095 171.905 ;
        RECT 60.265 171.095 60.595 171.735 ;
        RECT 60.765 171.095 61.035 171.905 ;
        RECT 61.215 171.360 66.560 171.905 ;
        RECT 59.835 170.665 60.185 170.915 ;
        RECT 43.745 169.525 44.075 170.375 ;
        RECT 44.245 169.355 44.415 170.205 ;
        RECT 44.585 169.525 44.915 170.375 ;
        RECT 45.085 169.355 45.255 170.205 ;
        RECT 45.425 169.525 45.755 170.375 ;
        RECT 45.925 169.355 46.095 170.155 ;
        RECT 46.265 169.525 46.595 170.375 ;
        RECT 46.765 169.355 46.935 170.155 ;
        RECT 47.105 169.525 47.435 170.375 ;
        RECT 47.605 169.355 47.775 170.155 ;
        RECT 47.945 169.525 48.275 170.375 ;
        RECT 48.445 169.355 48.615 170.155 ;
        RECT 48.785 169.525 49.115 170.375 ;
        RECT 49.285 169.355 49.455 170.155 ;
        RECT 49.625 169.525 49.955 170.375 ;
        RECT 50.125 169.355 50.295 170.155 ;
        RECT 50.465 169.525 50.795 170.375 ;
        RECT 50.965 169.355 51.135 170.155 ;
        RECT 51.305 169.525 51.635 170.375 ;
        RECT 51.805 169.355 51.975 170.155 ;
        RECT 52.145 169.525 52.475 170.375 ;
        RECT 52.645 169.355 52.815 170.155 ;
        RECT 52.985 169.525 53.315 170.375 ;
        RECT 53.485 169.355 53.655 170.155 ;
        RECT 53.825 169.525 54.155 170.375 ;
        RECT 55.020 170.255 58.330 170.495 ;
        RECT 54.325 169.355 54.495 170.155 ;
        RECT 55.025 169.355 55.320 170.085 ;
        RECT 55.490 169.530 55.750 170.255 ;
        RECT 55.920 169.355 56.180 170.085 ;
        RECT 56.350 169.530 56.610 170.255 ;
        RECT 56.780 169.355 57.040 170.085 ;
        RECT 57.210 169.530 57.470 170.255 ;
        RECT 57.640 169.355 57.900 170.085 ;
        RECT 58.070 169.530 58.330 170.255 ;
        RECT 58.500 169.355 58.760 170.465 ;
        RECT 58.930 169.530 59.180 170.665 ;
        RECT 60.355 170.495 60.525 171.095 ;
        RECT 60.695 170.665 61.045 170.915 ;
        RECT 62.800 170.530 63.140 171.360 ;
        RECT 66.735 171.135 68.405 171.905 ;
        RECT 69.035 171.180 69.325 171.905 ;
        RECT 69.545 171.250 69.875 171.685 ;
        RECT 70.045 171.295 70.215 171.905 ;
        RECT 69.495 171.165 69.875 171.250 ;
        RECT 70.385 171.165 70.715 171.690 ;
        RECT 70.975 171.375 71.185 171.905 ;
        RECT 71.460 171.455 72.245 171.625 ;
        RECT 72.415 171.455 72.820 171.625 ;
        RECT 59.360 169.355 59.655 170.465 ;
        RECT 59.845 170.325 60.525 170.495 ;
        RECT 59.845 169.540 60.175 170.325 ;
        RECT 60.705 169.355 61.035 170.495 ;
        RECT 64.620 169.790 64.970 171.040 ;
        RECT 66.735 170.615 67.485 171.135 ;
        RECT 69.495 171.125 69.720 171.165 ;
        RECT 67.655 170.445 68.405 170.965 ;
        RECT 69.495 170.545 69.665 171.125 ;
        RECT 70.385 170.995 70.585 171.165 ;
        RECT 71.460 170.995 71.630 171.455 ;
        RECT 69.835 170.665 70.585 170.995 ;
        RECT 70.755 170.665 71.630 170.995 ;
        RECT 61.215 169.355 66.560 169.790 ;
        RECT 66.735 169.355 68.405 170.445 ;
        RECT 69.035 169.355 69.325 170.520 ;
        RECT 69.495 170.495 69.710 170.545 ;
        RECT 69.495 170.415 69.885 170.495 ;
        RECT 69.555 169.570 69.885 170.415 ;
        RECT 70.395 170.460 70.585 170.665 ;
        RECT 70.055 169.355 70.225 170.365 ;
        RECT 70.395 170.085 71.290 170.460 ;
        RECT 70.395 169.525 70.735 170.085 ;
        RECT 70.965 169.355 71.280 169.855 ;
        RECT 71.460 169.825 71.630 170.665 ;
        RECT 71.800 170.955 72.265 171.285 ;
        RECT 72.650 171.225 72.820 171.455 ;
        RECT 73.000 171.405 73.370 171.905 ;
        RECT 73.690 171.455 74.365 171.625 ;
        RECT 74.560 171.455 74.895 171.625 ;
        RECT 71.800 169.995 72.120 170.955 ;
        RECT 72.650 170.925 73.480 171.225 ;
        RECT 72.290 170.025 72.480 170.745 ;
        RECT 72.650 169.855 72.820 170.925 ;
        RECT 73.280 170.895 73.480 170.925 ;
        RECT 72.990 170.675 73.160 170.745 ;
        RECT 73.690 170.675 73.860 171.455 ;
        RECT 74.725 171.315 74.895 171.455 ;
        RECT 75.065 171.445 75.315 171.905 ;
        RECT 72.990 170.505 73.860 170.675 ;
        RECT 74.030 171.035 74.555 171.255 ;
        RECT 74.725 171.185 74.950 171.315 ;
        RECT 72.990 170.415 73.500 170.505 ;
        RECT 71.460 169.655 72.345 169.825 ;
        RECT 72.570 169.525 72.820 169.855 ;
        RECT 72.990 169.355 73.160 170.155 ;
        RECT 73.330 169.800 73.500 170.415 ;
        RECT 74.030 170.335 74.200 171.035 ;
        RECT 73.670 169.970 74.200 170.335 ;
        RECT 74.370 170.270 74.610 170.865 ;
        RECT 74.780 170.080 74.950 171.185 ;
        RECT 75.120 170.325 75.400 171.275 ;
        RECT 74.645 169.950 74.950 170.080 ;
        RECT 73.330 169.630 74.435 169.800 ;
        RECT 74.645 169.525 74.895 169.950 ;
        RECT 75.065 169.355 75.330 169.815 ;
        RECT 75.570 169.525 75.755 171.645 ;
        RECT 75.925 171.525 76.255 171.905 ;
        RECT 76.425 171.355 76.595 171.645 ;
        RECT 75.930 171.185 76.595 171.355 ;
        RECT 75.930 170.195 76.160 171.185 ;
        RECT 76.330 170.365 76.680 171.015 ;
        RECT 75.930 170.025 76.595 170.195 ;
        RECT 75.925 169.355 76.255 169.855 ;
        RECT 76.425 169.525 76.595 170.025 ;
        RECT 76.865 169.535 77.125 171.725 ;
        RECT 77.385 171.535 78.055 171.905 ;
        RECT 78.235 171.355 78.545 171.725 ;
        RECT 77.315 171.155 78.545 171.355 ;
        RECT 77.315 170.485 77.605 171.155 ;
        RECT 78.725 170.975 78.955 171.615 ;
        RECT 79.135 171.175 79.425 171.905 ;
        RECT 79.650 171.165 80.265 171.735 ;
        RECT 80.435 171.395 80.650 171.905 ;
        RECT 80.880 171.395 81.160 171.725 ;
        RECT 81.340 171.395 81.580 171.905 ;
        RECT 81.915 171.445 82.475 171.735 ;
        RECT 82.645 171.445 82.895 171.905 ;
        RECT 77.785 170.665 78.250 170.975 ;
        RECT 78.430 170.665 78.955 170.975 ;
        RECT 79.135 170.665 79.435 170.995 ;
        RECT 77.315 170.265 78.085 170.485 ;
        RECT 77.295 169.355 77.635 170.085 ;
        RECT 77.815 169.535 78.085 170.265 ;
        RECT 78.265 170.245 79.425 170.485 ;
        RECT 78.265 169.535 78.495 170.245 ;
        RECT 78.665 169.355 78.995 170.065 ;
        RECT 79.165 169.535 79.425 170.245 ;
        RECT 79.650 170.145 79.965 171.165 ;
        RECT 80.135 170.495 80.305 170.995 ;
        RECT 80.555 170.665 80.820 171.225 ;
        RECT 80.990 170.495 81.160 171.395 ;
        RECT 81.330 170.665 81.685 171.225 ;
        RECT 80.135 170.325 81.560 170.495 ;
        RECT 79.650 169.525 80.185 170.145 ;
        RECT 80.355 169.355 80.685 170.155 ;
        RECT 81.170 170.150 81.560 170.325 ;
        RECT 81.915 170.075 82.165 171.445 ;
        RECT 83.515 171.275 83.845 171.635 ;
        RECT 82.455 171.085 83.845 171.275 ;
        RECT 84.330 171.275 84.615 171.735 ;
        RECT 84.785 171.445 85.055 171.905 ;
        RECT 84.330 171.105 85.285 171.275 ;
        RECT 82.455 170.995 82.625 171.085 ;
        RECT 82.335 170.665 82.625 170.995 ;
        RECT 82.795 170.665 83.135 170.915 ;
        RECT 83.355 170.665 84.030 170.915 ;
        RECT 82.455 170.415 82.625 170.665 ;
        RECT 82.455 170.245 83.395 170.415 ;
        RECT 83.765 170.305 84.030 170.665 ;
        RECT 84.215 170.375 84.905 170.935 ;
        RECT 81.915 169.525 82.375 170.075 ;
        RECT 82.565 169.355 82.895 170.075 ;
        RECT 83.095 169.695 83.395 170.245 ;
        RECT 85.075 170.205 85.285 171.105 ;
        RECT 83.565 169.355 83.845 170.025 ;
        RECT 84.330 169.985 85.285 170.205 ;
        RECT 85.455 170.935 85.855 171.735 ;
        RECT 86.045 171.275 86.325 171.735 ;
        RECT 86.845 171.445 87.170 171.905 ;
        RECT 86.045 171.105 87.170 171.275 ;
        RECT 87.340 171.165 87.725 171.735 ;
        RECT 86.720 170.995 87.170 171.105 ;
        RECT 85.455 170.375 86.550 170.935 ;
        RECT 86.720 170.665 87.275 170.995 ;
        RECT 84.330 169.525 84.615 169.985 ;
        RECT 84.785 169.355 85.055 169.815 ;
        RECT 85.455 169.525 85.855 170.375 ;
        RECT 86.720 170.205 87.170 170.665 ;
        RECT 87.445 170.495 87.725 171.165 ;
        RECT 86.045 169.985 87.170 170.205 ;
        RECT 86.045 169.525 86.325 169.985 ;
        RECT 86.845 169.355 87.170 169.815 ;
        RECT 87.340 169.525 87.725 170.495 ;
        RECT 87.900 171.165 88.155 171.735 ;
        RECT 88.325 171.505 88.655 171.905 ;
        RECT 89.080 171.370 89.610 171.735 ;
        RECT 89.080 171.335 89.255 171.370 ;
        RECT 88.325 171.165 89.255 171.335 ;
        RECT 87.900 170.495 88.070 171.165 ;
        RECT 88.325 170.995 88.495 171.165 ;
        RECT 88.240 170.665 88.495 170.995 ;
        RECT 88.720 170.665 88.915 170.995 ;
        RECT 87.900 169.525 88.235 170.495 ;
        RECT 88.405 169.355 88.575 170.495 ;
        RECT 88.745 169.695 88.915 170.665 ;
        RECT 89.085 170.035 89.255 171.165 ;
        RECT 89.425 170.375 89.595 171.175 ;
        RECT 89.800 170.885 90.075 171.735 ;
        RECT 89.795 170.715 90.075 170.885 ;
        RECT 89.800 170.575 90.075 170.715 ;
        RECT 90.245 170.375 90.435 171.735 ;
        RECT 90.615 171.370 91.125 171.905 ;
        RECT 91.345 171.095 91.590 171.700 ;
        RECT 92.035 171.135 94.625 171.905 ;
        RECT 94.795 171.180 95.085 171.905 ;
        RECT 95.305 171.250 95.635 171.685 ;
        RECT 95.805 171.295 95.975 171.905 ;
        RECT 95.255 171.165 95.635 171.250 ;
        RECT 96.145 171.165 96.475 171.690 ;
        RECT 96.735 171.375 96.945 171.905 ;
        RECT 97.220 171.455 98.005 171.625 ;
        RECT 98.175 171.455 98.580 171.625 ;
        RECT 90.635 170.925 91.865 171.095 ;
        RECT 89.425 170.205 90.435 170.375 ;
        RECT 90.605 170.360 91.355 170.550 ;
        RECT 89.085 169.865 90.210 170.035 ;
        RECT 90.605 169.695 90.775 170.360 ;
        RECT 91.525 170.115 91.865 170.925 ;
        RECT 92.035 170.615 93.245 171.135 ;
        RECT 95.255 171.125 95.480 171.165 ;
        RECT 93.415 170.445 94.625 170.965 ;
        RECT 95.255 170.545 95.425 171.125 ;
        RECT 96.145 170.995 96.345 171.165 ;
        RECT 97.220 170.995 97.390 171.455 ;
        RECT 95.595 170.665 96.345 170.995 ;
        RECT 96.515 170.665 97.390 170.995 ;
        RECT 88.745 169.525 90.775 169.695 ;
        RECT 90.945 169.355 91.115 170.115 ;
        RECT 91.350 169.705 91.865 170.115 ;
        RECT 92.035 169.355 94.625 170.445 ;
        RECT 94.795 169.355 95.085 170.520 ;
        RECT 95.255 170.495 95.470 170.545 ;
        RECT 95.255 170.415 95.645 170.495 ;
        RECT 95.315 169.570 95.645 170.415 ;
        RECT 96.155 170.460 96.345 170.665 ;
        RECT 95.815 169.355 95.985 170.365 ;
        RECT 96.155 170.085 97.050 170.460 ;
        RECT 96.155 169.525 96.495 170.085 ;
        RECT 96.725 169.355 97.040 169.855 ;
        RECT 97.220 169.825 97.390 170.665 ;
        RECT 97.560 170.955 98.025 171.285 ;
        RECT 98.410 171.225 98.580 171.455 ;
        RECT 98.760 171.405 99.130 171.905 ;
        RECT 99.450 171.455 100.125 171.625 ;
        RECT 100.320 171.455 100.655 171.625 ;
        RECT 97.560 169.995 97.880 170.955 ;
        RECT 98.410 170.925 99.240 171.225 ;
        RECT 98.050 170.025 98.240 170.745 ;
        RECT 98.410 169.855 98.580 170.925 ;
        RECT 99.040 170.895 99.240 170.925 ;
        RECT 98.750 170.675 98.920 170.745 ;
        RECT 99.450 170.675 99.620 171.455 ;
        RECT 100.485 171.315 100.655 171.455 ;
        RECT 100.825 171.445 101.075 171.905 ;
        RECT 98.750 170.505 99.620 170.675 ;
        RECT 99.790 171.035 100.315 171.255 ;
        RECT 100.485 171.185 100.710 171.315 ;
        RECT 98.750 170.415 99.260 170.505 ;
        RECT 97.220 169.655 98.105 169.825 ;
        RECT 98.330 169.525 98.580 169.855 ;
        RECT 98.750 169.355 98.920 170.155 ;
        RECT 99.090 169.800 99.260 170.415 ;
        RECT 99.790 170.335 99.960 171.035 ;
        RECT 99.430 169.970 99.960 170.335 ;
        RECT 100.130 170.270 100.370 170.865 ;
        RECT 100.540 170.080 100.710 171.185 ;
        RECT 100.880 170.325 101.160 171.275 ;
        RECT 100.405 169.950 100.710 170.080 ;
        RECT 99.090 169.630 100.195 169.800 ;
        RECT 100.405 169.525 100.655 169.950 ;
        RECT 100.825 169.355 101.090 169.815 ;
        RECT 101.330 169.525 101.515 171.645 ;
        RECT 101.685 171.525 102.015 171.905 ;
        RECT 102.185 171.355 102.355 171.645 ;
        RECT 101.690 171.185 102.355 171.355 ;
        RECT 102.615 171.405 102.875 171.735 ;
        RECT 103.045 171.545 103.375 171.905 ;
        RECT 103.630 171.525 104.930 171.735 ;
        RECT 102.615 171.395 102.845 171.405 ;
        RECT 101.690 170.195 101.920 171.185 ;
        RECT 102.090 170.365 102.440 171.015 ;
        RECT 102.615 170.205 102.785 171.395 ;
        RECT 103.630 171.375 103.800 171.525 ;
        RECT 103.045 171.250 103.800 171.375 ;
        RECT 102.955 171.205 103.800 171.250 ;
        RECT 102.955 171.085 103.225 171.205 ;
        RECT 102.955 170.510 103.125 171.085 ;
        RECT 103.355 170.645 103.765 170.950 ;
        RECT 104.055 170.915 104.265 171.315 ;
        RECT 103.935 170.705 104.265 170.915 ;
        RECT 104.510 170.915 104.730 171.315 ;
        RECT 105.205 171.140 105.660 171.905 ;
        RECT 104.510 170.705 104.985 170.915 ;
        RECT 105.175 170.715 105.665 170.915 ;
        RECT 102.955 170.475 103.155 170.510 ;
        RECT 104.485 170.475 105.660 170.535 ;
        RECT 102.955 170.365 105.660 170.475 ;
        RECT 103.015 170.305 104.815 170.365 ;
        RECT 104.485 170.275 104.815 170.305 ;
        RECT 101.690 170.025 102.355 170.195 ;
        RECT 101.685 169.355 102.015 169.855 ;
        RECT 102.185 169.525 102.355 170.025 ;
        RECT 102.615 169.525 102.875 170.205 ;
        RECT 103.045 169.355 103.295 170.135 ;
        RECT 103.545 170.105 104.380 170.115 ;
        RECT 104.970 170.105 105.155 170.195 ;
        RECT 103.545 169.905 105.155 170.105 ;
        RECT 103.545 169.525 103.795 169.905 ;
        RECT 104.925 169.865 105.155 169.905 ;
        RECT 105.405 169.745 105.660 170.365 ;
        RECT 103.965 169.355 104.320 169.735 ;
        RECT 105.325 169.525 105.660 169.745 ;
        RECT 105.840 170.305 106.175 171.725 ;
        RECT 106.355 171.535 107.100 171.905 ;
        RECT 107.665 171.365 107.920 171.725 ;
        RECT 108.100 171.535 108.430 171.905 ;
        RECT 108.610 171.365 108.835 171.725 ;
        RECT 106.350 171.175 108.835 171.365 ;
        RECT 106.350 170.485 106.575 171.175 ;
        RECT 109.055 171.135 112.565 171.905 ;
        RECT 106.775 170.665 107.055 170.995 ;
        RECT 107.235 170.665 107.810 170.995 ;
        RECT 107.990 170.665 108.425 170.995 ;
        RECT 108.605 170.665 108.875 170.995 ;
        RECT 109.055 170.615 110.705 171.135 ;
        RECT 106.350 170.305 108.845 170.485 ;
        RECT 110.875 170.445 112.565 170.965 ;
        RECT 105.840 169.535 106.105 170.305 ;
        RECT 106.275 169.355 106.605 170.075 ;
        RECT 106.795 169.895 107.985 170.125 ;
        RECT 106.795 169.535 107.055 169.895 ;
        RECT 107.225 169.355 107.555 169.725 ;
        RECT 107.725 169.535 107.985 169.895 ;
        RECT 108.555 169.535 108.845 170.305 ;
        RECT 109.055 169.355 112.565 170.445 ;
        RECT 113.655 169.525 113.935 171.625 ;
        RECT 114.165 171.445 114.335 171.905 ;
        RECT 114.605 171.515 115.855 171.695 ;
        RECT 114.990 171.275 115.355 171.345 ;
        RECT 114.105 171.095 115.355 171.275 ;
        RECT 115.525 171.295 115.855 171.515 ;
        RECT 116.025 171.465 116.195 171.905 ;
        RECT 116.365 171.295 116.705 171.710 ;
        RECT 115.525 171.125 116.705 171.295 ;
        RECT 114.105 170.495 114.380 171.095 ;
        RECT 114.550 170.665 114.905 170.915 ;
        RECT 115.100 170.885 115.565 170.915 ;
        RECT 115.095 170.715 115.565 170.885 ;
        RECT 115.100 170.665 115.565 170.715 ;
        RECT 115.735 170.665 116.065 170.915 ;
        RECT 116.240 170.715 116.705 170.915 ;
        RECT 115.885 170.545 116.065 170.665 ;
        RECT 114.105 170.285 115.715 170.495 ;
        RECT 115.885 170.375 116.215 170.545 ;
        RECT 115.305 170.185 115.715 170.285 ;
        RECT 114.125 169.355 114.910 170.115 ;
        RECT 115.305 169.525 115.690 170.185 ;
        RECT 116.015 169.585 116.215 170.375 ;
        RECT 116.385 169.355 116.705 170.535 ;
        RECT 116.885 169.535 117.145 171.725 ;
        RECT 117.405 171.535 118.075 171.905 ;
        RECT 118.255 171.355 118.565 171.725 ;
        RECT 117.335 171.155 118.565 171.355 ;
        RECT 117.335 170.485 117.625 171.155 ;
        RECT 118.745 170.975 118.975 171.615 ;
        RECT 119.155 171.175 119.445 171.905 ;
        RECT 120.555 171.180 120.845 171.905 ;
        RECT 121.175 171.345 121.505 171.735 ;
        RECT 121.675 171.515 122.860 171.685 ;
        RECT 123.120 171.435 123.290 171.905 ;
        RECT 121.175 171.165 121.685 171.345 ;
        RECT 117.805 170.665 118.270 170.975 ;
        RECT 118.450 170.665 118.975 170.975 ;
        RECT 119.155 170.665 119.455 170.995 ;
        RECT 121.015 170.705 121.345 170.995 ;
        RECT 121.515 170.535 121.685 171.165 ;
        RECT 122.090 171.255 122.475 171.345 ;
        RECT 123.460 171.255 123.790 171.720 ;
        RECT 122.090 171.085 123.790 171.255 ;
        RECT 123.960 171.085 124.130 171.905 ;
        RECT 124.300 171.085 124.985 171.725 ;
        RECT 125.160 171.140 125.615 171.905 ;
        RECT 125.890 171.525 127.190 171.735 ;
        RECT 127.445 171.545 127.775 171.905 ;
        RECT 127.020 171.375 127.190 171.525 ;
        RECT 127.945 171.405 128.205 171.735 ;
        RECT 121.855 170.705 122.185 170.915 ;
        RECT 122.365 170.665 122.745 170.915 ;
        RECT 117.335 170.265 118.105 170.485 ;
        RECT 117.315 169.355 117.655 170.085 ;
        RECT 117.835 169.535 118.105 170.265 ;
        RECT 118.285 170.245 119.445 170.485 ;
        RECT 118.285 169.535 118.515 170.245 ;
        RECT 118.685 169.355 119.015 170.065 ;
        RECT 119.185 169.535 119.445 170.245 ;
        RECT 120.555 169.355 120.845 170.520 ;
        RECT 121.170 170.365 122.255 170.535 ;
        RECT 121.170 169.525 121.470 170.365 ;
        RECT 121.665 169.355 121.915 170.195 ;
        RECT 122.085 170.115 122.255 170.365 ;
        RECT 122.425 170.285 122.745 170.665 ;
        RECT 122.935 170.705 123.420 170.915 ;
        RECT 123.610 170.705 124.060 170.915 ;
        RECT 124.230 170.705 124.565 170.915 ;
        RECT 122.935 170.545 123.310 170.705 ;
        RECT 122.915 170.375 123.310 170.545 ;
        RECT 124.230 170.535 124.400 170.705 ;
        RECT 122.935 170.285 123.310 170.375 ;
        RECT 123.480 170.365 124.400 170.535 ;
        RECT 123.480 170.115 123.650 170.365 ;
        RECT 122.085 169.945 123.650 170.115 ;
        RECT 122.505 169.525 123.310 169.945 ;
        RECT 123.820 169.355 124.150 170.195 ;
        RECT 124.735 170.115 124.985 171.085 ;
        RECT 126.090 170.915 126.310 171.315 ;
        RECT 125.155 170.715 125.645 170.915 ;
        RECT 125.835 170.705 126.310 170.915 ;
        RECT 126.555 170.915 126.765 171.315 ;
        RECT 127.020 171.250 127.775 171.375 ;
        RECT 127.020 171.205 127.865 171.250 ;
        RECT 127.595 171.085 127.865 171.205 ;
        RECT 126.555 170.705 126.885 170.915 ;
        RECT 127.055 170.645 127.465 170.950 ;
        RECT 124.320 169.525 124.985 170.115 ;
        RECT 125.160 170.475 126.335 170.535 ;
        RECT 127.695 170.510 127.865 171.085 ;
        RECT 127.665 170.475 127.865 170.510 ;
        RECT 125.160 170.365 127.865 170.475 ;
        RECT 125.160 169.745 125.415 170.365 ;
        RECT 126.005 170.305 127.805 170.365 ;
        RECT 126.005 170.275 126.335 170.305 ;
        RECT 128.035 170.205 128.205 171.405 ;
        RECT 128.380 171.140 128.835 171.905 ;
        RECT 129.110 171.525 130.410 171.735 ;
        RECT 130.665 171.545 130.995 171.905 ;
        RECT 130.240 171.375 130.410 171.525 ;
        RECT 131.165 171.405 131.425 171.735 ;
        RECT 131.195 171.395 131.425 171.405 ;
        RECT 129.310 170.915 129.530 171.315 ;
        RECT 128.375 170.715 128.865 170.915 ;
        RECT 129.055 170.705 129.530 170.915 ;
        RECT 129.775 170.915 129.985 171.315 ;
        RECT 130.240 171.250 130.995 171.375 ;
        RECT 130.240 171.205 131.085 171.250 ;
        RECT 130.815 171.085 131.085 171.205 ;
        RECT 129.775 170.705 130.105 170.915 ;
        RECT 130.275 170.645 130.685 170.950 ;
        RECT 125.665 170.105 125.850 170.195 ;
        RECT 126.440 170.105 127.275 170.115 ;
        RECT 125.665 169.905 127.275 170.105 ;
        RECT 125.665 169.865 125.895 169.905 ;
        RECT 125.160 169.525 125.495 169.745 ;
        RECT 126.500 169.355 126.855 169.735 ;
        RECT 127.025 169.525 127.275 169.905 ;
        RECT 127.525 169.355 127.775 170.135 ;
        RECT 127.945 169.525 128.205 170.205 ;
        RECT 128.380 170.475 129.555 170.535 ;
        RECT 130.915 170.510 131.085 171.085 ;
        RECT 130.885 170.475 131.085 170.510 ;
        RECT 128.380 170.365 131.085 170.475 ;
        RECT 128.380 169.745 128.635 170.365 ;
        RECT 129.225 170.305 131.025 170.365 ;
        RECT 129.225 170.275 129.555 170.305 ;
        RECT 131.255 170.205 131.425 171.395 ;
        RECT 131.870 171.095 132.115 171.700 ;
        RECT 132.335 171.370 132.845 171.905 ;
        RECT 128.885 170.105 129.070 170.195 ;
        RECT 129.660 170.105 130.495 170.115 ;
        RECT 128.885 169.905 130.495 170.105 ;
        RECT 128.885 169.865 129.115 169.905 ;
        RECT 128.380 169.525 128.715 169.745 ;
        RECT 129.720 169.355 130.075 169.735 ;
        RECT 130.245 169.525 130.495 169.905 ;
        RECT 130.745 169.355 130.995 170.135 ;
        RECT 131.165 169.525 131.425 170.205 ;
        RECT 131.595 170.925 132.825 171.095 ;
        RECT 131.595 170.115 131.935 170.925 ;
        RECT 132.105 170.360 132.855 170.550 ;
        RECT 131.595 169.705 132.110 170.115 ;
        RECT 132.345 169.355 132.515 170.115 ;
        RECT 132.685 169.695 132.855 170.360 ;
        RECT 133.025 170.375 133.215 171.735 ;
        RECT 133.385 171.225 133.660 171.735 ;
        RECT 133.850 171.370 134.380 171.735 ;
        RECT 134.805 171.505 135.135 171.905 ;
        RECT 134.205 171.335 134.380 171.370 ;
        RECT 133.385 171.055 133.665 171.225 ;
        RECT 133.385 170.575 133.660 171.055 ;
        RECT 133.865 170.375 134.035 171.175 ;
        RECT 133.025 170.205 134.035 170.375 ;
        RECT 134.205 171.165 135.135 171.335 ;
        RECT 135.305 171.165 135.560 171.735 ;
        RECT 135.825 171.355 135.995 171.735 ;
        RECT 136.175 171.525 136.505 171.905 ;
        RECT 135.825 171.185 136.490 171.355 ;
        RECT 136.685 171.230 136.945 171.735 ;
        RECT 134.205 170.035 134.375 171.165 ;
        RECT 134.965 170.995 135.135 171.165 ;
        RECT 133.250 169.865 134.375 170.035 ;
        RECT 134.545 170.665 134.740 170.995 ;
        RECT 134.965 170.665 135.220 170.995 ;
        RECT 134.545 169.695 134.715 170.665 ;
        RECT 135.390 170.495 135.560 171.165 ;
        RECT 135.755 170.635 136.085 171.005 ;
        RECT 136.320 170.930 136.490 171.185 ;
        RECT 132.685 169.525 134.715 169.695 ;
        RECT 134.885 169.355 135.055 170.495 ;
        RECT 135.225 169.525 135.560 170.495 ;
        RECT 136.320 170.600 136.605 170.930 ;
        RECT 136.320 170.455 136.490 170.600 ;
        RECT 135.825 170.285 136.490 170.455 ;
        RECT 136.775 170.430 136.945 171.230 ;
        RECT 135.825 169.525 135.995 170.285 ;
        RECT 136.175 169.355 136.505 170.115 ;
        RECT 136.675 169.525 136.945 170.430 ;
        RECT 137.115 171.165 137.500 171.735 ;
        RECT 137.670 171.445 137.995 171.905 ;
        RECT 138.515 171.275 138.795 171.735 ;
        RECT 137.115 170.495 137.395 171.165 ;
        RECT 137.670 171.105 138.795 171.275 ;
        RECT 137.670 170.995 138.120 171.105 ;
        RECT 137.565 170.665 138.120 170.995 ;
        RECT 138.985 170.935 139.385 171.735 ;
        RECT 139.785 171.445 140.055 171.905 ;
        RECT 140.225 171.275 140.510 171.735 ;
        RECT 137.115 169.525 137.500 170.495 ;
        RECT 137.670 170.205 138.120 170.665 ;
        RECT 138.290 170.375 139.385 170.935 ;
        RECT 137.670 169.985 138.795 170.205 ;
        RECT 137.670 169.355 137.995 169.815 ;
        RECT 138.515 169.525 138.795 169.985 ;
        RECT 138.985 169.525 139.385 170.375 ;
        RECT 139.555 171.105 140.510 171.275 ;
        RECT 141.715 171.155 142.925 171.905 ;
        RECT 139.555 170.205 139.765 171.105 ;
        RECT 139.935 170.375 140.625 170.935 ;
        RECT 141.715 170.445 142.235 170.985 ;
        RECT 142.405 170.615 142.925 171.155 ;
        RECT 139.555 169.985 140.510 170.205 ;
        RECT 139.785 169.355 140.055 169.815 ;
        RECT 140.225 169.525 140.510 169.985 ;
        RECT 141.715 169.355 142.925 170.445 ;
        RECT 17.430 169.185 143.010 169.355 ;
        RECT 17.515 168.095 18.725 169.185 ;
        RECT 18.895 168.750 24.240 169.185 ;
        RECT 17.515 167.385 18.035 167.925 ;
        RECT 18.205 167.555 18.725 168.095 ;
        RECT 17.515 166.635 18.725 167.385 ;
        RECT 20.480 167.180 20.820 168.010 ;
        RECT 22.300 167.500 22.650 168.750 ;
        RECT 25.345 168.575 25.675 169.005 ;
        RECT 25.855 168.745 26.050 169.185 ;
        RECT 26.220 168.575 26.550 169.005 ;
        RECT 25.345 168.405 26.550 168.575 ;
        RECT 25.345 168.075 26.240 168.405 ;
        RECT 26.720 168.235 26.995 169.005 ;
        RECT 26.410 168.045 26.995 168.235 ;
        RECT 27.175 168.095 29.765 169.185 ;
        RECT 25.350 167.545 25.645 167.875 ;
        RECT 25.825 167.545 26.240 167.875 ;
        RECT 18.895 166.635 24.240 167.180 ;
        RECT 25.345 166.635 25.645 167.365 ;
        RECT 25.825 166.925 26.055 167.545 ;
        RECT 26.410 167.375 26.585 168.045 ;
        RECT 26.255 167.195 26.585 167.375 ;
        RECT 26.755 167.225 26.995 167.875 ;
        RECT 27.175 167.405 28.385 167.925 ;
        RECT 28.555 167.575 29.765 168.095 ;
        RECT 30.395 168.020 30.685 169.185 ;
        RECT 30.855 168.095 32.525 169.185 ;
        RECT 33.155 168.675 34.345 168.965 ;
        RECT 30.855 167.405 31.605 167.925 ;
        RECT 31.775 167.575 32.525 168.095 ;
        RECT 33.175 168.335 34.345 168.505 ;
        RECT 34.515 168.385 34.795 169.185 ;
        RECT 33.175 168.045 33.500 168.335 ;
        RECT 34.175 168.215 34.345 168.335 ;
        RECT 33.670 167.875 33.865 168.165 ;
        RECT 34.175 168.045 34.835 168.215 ;
        RECT 35.005 168.045 35.280 169.015 ;
        RECT 36.375 168.045 36.655 169.185 ;
        RECT 34.665 167.875 34.835 168.045 ;
        RECT 33.155 167.545 33.500 167.875 ;
        RECT 33.670 167.545 34.495 167.875 ;
        RECT 34.665 167.545 34.940 167.875 ;
        RECT 26.255 166.815 26.480 167.195 ;
        RECT 26.650 166.635 26.980 167.025 ;
        RECT 27.175 166.635 29.765 167.405 ;
        RECT 30.395 166.635 30.685 167.360 ;
        RECT 30.855 166.635 32.525 167.405 ;
        RECT 34.665 167.375 34.835 167.545 ;
        RECT 33.170 167.205 34.835 167.375 ;
        RECT 35.110 167.310 35.280 168.045 ;
        RECT 36.825 168.035 37.155 169.015 ;
        RECT 37.325 168.045 37.585 169.185 ;
        RECT 37.960 168.215 38.290 169.015 ;
        RECT 38.460 168.385 38.790 169.185 ;
        RECT 39.090 168.215 39.420 169.015 ;
        RECT 40.065 168.385 40.315 169.185 ;
        RECT 37.960 168.045 40.395 168.215 ;
        RECT 40.585 168.045 40.755 169.185 ;
        RECT 40.925 168.045 41.265 169.015 ;
        RECT 36.385 167.605 36.720 167.875 ;
        RECT 36.890 167.435 37.060 168.035 ;
        RECT 37.230 167.625 37.565 167.875 ;
        RECT 37.755 167.625 38.105 167.875 ;
        RECT 33.170 166.855 33.425 167.205 ;
        RECT 33.595 166.635 33.925 167.035 ;
        RECT 34.095 166.855 34.265 167.205 ;
        RECT 34.435 166.635 34.815 167.035 ;
        RECT 35.005 166.965 35.280 167.310 ;
        RECT 36.375 166.635 36.685 167.435 ;
        RECT 36.890 166.805 37.585 167.435 ;
        RECT 38.290 167.415 38.460 168.045 ;
        RECT 38.630 167.625 38.960 167.825 ;
        RECT 39.130 167.625 39.460 167.825 ;
        RECT 39.630 167.625 40.050 167.825 ;
        RECT 40.225 167.795 40.395 168.045 ;
        RECT 40.225 167.625 40.920 167.795 ;
        RECT 37.960 166.805 38.460 167.415 ;
        RECT 39.090 167.285 40.315 167.455 ;
        RECT 41.090 167.435 41.265 168.045 ;
        RECT 39.090 166.805 39.420 167.285 ;
        RECT 39.590 166.635 39.815 167.095 ;
        RECT 39.985 166.805 40.315 167.285 ;
        RECT 40.505 166.635 40.755 167.435 ;
        RECT 40.925 166.805 41.265 167.435 ;
        RECT 41.435 168.045 41.710 169.015 ;
        RECT 41.920 168.385 42.200 169.185 ;
        RECT 42.370 168.675 43.985 169.005 ;
        RECT 42.370 168.335 43.545 168.505 ;
        RECT 42.370 168.215 42.540 168.335 ;
        RECT 41.880 168.045 42.540 168.215 ;
        RECT 41.435 167.310 41.605 168.045 ;
        RECT 41.880 167.875 42.050 168.045 ;
        RECT 42.800 167.875 43.045 168.165 ;
        RECT 43.215 168.045 43.545 168.335 ;
        RECT 43.805 167.875 43.975 168.435 ;
        RECT 44.225 168.045 44.485 169.185 ;
        RECT 44.840 168.215 45.230 168.390 ;
        RECT 45.715 168.385 46.045 169.185 ;
        RECT 46.215 168.395 46.750 169.015 ;
        RECT 44.840 168.045 46.265 168.215 ;
        RECT 41.775 167.545 42.050 167.875 ;
        RECT 42.220 167.545 43.045 167.875 ;
        RECT 43.260 167.545 43.975 167.875 ;
        RECT 44.145 167.625 44.480 167.875 ;
        RECT 41.880 167.375 42.050 167.545 ;
        RECT 43.725 167.455 43.975 167.545 ;
        RECT 41.435 166.965 41.710 167.310 ;
        RECT 41.880 167.205 43.545 167.375 ;
        RECT 41.900 166.635 42.275 167.035 ;
        RECT 42.445 166.855 42.615 167.205 ;
        RECT 42.785 166.635 43.115 167.035 ;
        RECT 43.285 166.805 43.545 167.205 ;
        RECT 43.725 167.035 44.055 167.455 ;
        RECT 44.225 166.635 44.485 167.455 ;
        RECT 44.715 167.315 45.070 167.875 ;
        RECT 45.240 167.145 45.410 168.045 ;
        RECT 45.580 167.315 45.845 167.875 ;
        RECT 46.095 167.545 46.265 168.045 ;
        RECT 46.435 167.375 46.750 168.395 ;
        RECT 46.955 168.095 50.465 169.185 ;
        RECT 50.720 168.565 50.895 169.015 ;
        RECT 51.065 168.745 51.395 169.185 ;
        RECT 51.700 168.595 51.870 169.015 ;
        RECT 52.105 168.775 52.775 169.185 ;
        RECT 52.990 168.595 53.160 169.015 ;
        RECT 53.360 168.775 53.690 169.185 ;
        RECT 50.720 168.395 51.350 168.565 ;
        RECT 44.820 166.635 45.060 167.145 ;
        RECT 45.240 166.815 45.520 167.145 ;
        RECT 45.750 166.635 45.965 167.145 ;
        RECT 46.135 166.805 46.750 167.375 ;
        RECT 46.955 167.405 48.605 167.925 ;
        RECT 48.775 167.575 50.465 168.095 ;
        RECT 50.635 167.545 51.000 168.225 ;
        RECT 51.180 167.875 51.350 168.395 ;
        RECT 51.700 168.425 53.715 168.595 ;
        RECT 51.180 167.545 51.530 167.875 ;
        RECT 46.955 166.635 50.465 167.405 ;
        RECT 51.180 167.375 51.350 167.545 ;
        RECT 50.720 167.205 51.350 167.375 ;
        RECT 50.720 166.805 50.895 167.205 ;
        RECT 51.700 167.135 51.870 168.425 ;
        RECT 51.065 166.635 51.395 167.015 ;
        RECT 51.640 166.805 51.870 167.135 ;
        RECT 52.070 166.970 52.350 168.245 ;
        RECT 52.575 168.165 52.845 168.245 ;
        RECT 52.535 167.995 52.845 168.165 ;
        RECT 52.575 166.970 52.845 167.995 ;
        RECT 53.035 167.215 53.375 168.245 ;
        RECT 53.545 167.875 53.715 168.425 ;
        RECT 53.885 168.045 54.145 169.015 ;
        RECT 54.325 168.045 54.655 169.185 ;
        RECT 55.185 168.215 55.515 169.000 ;
        RECT 54.835 168.045 55.515 168.215 ;
        RECT 53.545 167.545 53.805 167.875 ;
        RECT 53.975 167.355 54.145 168.045 ;
        RECT 54.315 167.625 54.665 167.875 ;
        RECT 54.835 167.445 55.005 168.045 ;
        RECT 56.155 168.020 56.445 169.185 ;
        RECT 56.615 168.350 57.000 169.185 ;
        RECT 57.170 168.180 57.430 168.985 ;
        RECT 57.600 168.350 57.860 169.185 ;
        RECT 58.030 168.180 58.285 168.985 ;
        RECT 58.460 168.350 58.720 169.185 ;
        RECT 58.890 168.180 59.145 168.985 ;
        RECT 59.320 168.350 59.665 169.185 ;
        RECT 56.615 168.010 59.645 168.180 ;
        RECT 59.835 168.095 63.345 169.185 ;
        RECT 55.175 167.625 55.525 167.875 ;
        RECT 56.615 167.445 56.915 168.010 ;
        RECT 57.090 167.615 59.305 167.840 ;
        RECT 59.475 167.445 59.645 168.010 ;
        RECT 53.305 166.635 53.635 167.015 ;
        RECT 53.805 166.890 54.145 167.355 ;
        RECT 53.805 166.845 54.140 166.890 ;
        RECT 54.325 166.635 54.595 167.445 ;
        RECT 54.765 166.805 55.095 167.445 ;
        RECT 55.265 166.635 55.505 167.445 ;
        RECT 56.155 166.635 56.445 167.360 ;
        RECT 56.615 167.275 59.645 167.445 ;
        RECT 59.835 167.405 61.485 167.925 ;
        RECT 61.655 167.575 63.345 168.095 ;
        RECT 64.445 168.075 64.740 169.185 ;
        RECT 64.920 167.875 65.170 169.010 ;
        RECT 65.340 168.075 65.600 169.185 ;
        RECT 65.770 168.285 66.030 169.010 ;
        RECT 66.200 168.455 66.460 169.185 ;
        RECT 66.630 168.285 66.890 169.010 ;
        RECT 67.060 168.455 67.320 169.185 ;
        RECT 67.490 168.285 67.750 169.010 ;
        RECT 67.920 168.455 68.180 169.185 ;
        RECT 68.350 168.285 68.610 169.010 ;
        RECT 68.780 168.455 69.075 169.185 ;
        RECT 65.770 168.045 69.080 168.285 ;
        RECT 57.135 166.635 57.435 167.105 ;
        RECT 57.605 166.830 57.860 167.275 ;
        RECT 58.030 166.635 58.290 167.105 ;
        RECT 58.460 166.830 58.720 167.275 ;
        RECT 58.890 166.635 59.185 167.105 ;
        RECT 59.835 166.635 63.345 167.405 ;
        RECT 64.435 167.265 64.750 167.875 ;
        RECT 64.920 167.625 67.940 167.875 ;
        RECT 64.495 166.635 64.740 167.095 ;
        RECT 64.920 166.815 65.170 167.625 ;
        RECT 68.110 167.455 69.080 168.045 ;
        RECT 69.505 168.165 69.835 169.015 ;
        RECT 70.005 168.335 70.175 169.185 ;
        RECT 70.345 168.165 70.675 169.015 ;
        RECT 70.845 168.335 71.015 169.185 ;
        RECT 71.185 168.165 71.515 169.015 ;
        RECT 71.685 168.385 71.855 169.185 ;
        RECT 72.025 168.165 72.355 169.015 ;
        RECT 72.525 168.385 72.695 169.185 ;
        RECT 72.865 168.165 73.195 169.015 ;
        RECT 73.365 168.385 73.535 169.185 ;
        RECT 73.705 168.165 74.035 169.015 ;
        RECT 74.205 168.385 74.375 169.185 ;
        RECT 74.545 168.165 74.875 169.015 ;
        RECT 75.045 168.385 75.215 169.185 ;
        RECT 75.385 168.165 75.715 169.015 ;
        RECT 75.885 168.385 76.055 169.185 ;
        RECT 76.225 168.165 76.555 169.015 ;
        RECT 76.725 168.385 76.895 169.185 ;
        RECT 77.065 168.165 77.395 169.015 ;
        RECT 77.565 168.385 77.735 169.185 ;
        RECT 77.905 168.165 78.235 169.015 ;
        RECT 78.405 168.385 78.575 169.185 ;
        RECT 78.745 168.165 79.075 169.015 ;
        RECT 79.245 168.385 79.415 169.185 ;
        RECT 79.585 168.165 79.915 169.015 ;
        RECT 80.085 168.385 80.255 169.185 ;
        RECT 69.505 167.995 71.015 168.165 ;
        RECT 71.185 167.995 73.535 168.165 ;
        RECT 73.705 167.995 80.365 168.165 ;
        RECT 80.535 168.045 80.795 169.185 ;
        RECT 80.965 168.035 81.295 169.015 ;
        RECT 81.465 168.045 81.745 169.185 ;
        RECT 70.845 167.825 71.015 167.995 ;
        RECT 73.360 167.825 73.535 167.995 ;
        RECT 69.500 167.625 70.675 167.825 ;
        RECT 70.845 167.625 73.155 167.825 ;
        RECT 73.360 167.625 79.920 167.825 ;
        RECT 70.845 167.455 71.015 167.625 ;
        RECT 73.360 167.455 73.535 167.625 ;
        RECT 80.090 167.455 80.365 167.995 ;
        RECT 80.555 167.625 80.890 167.875 ;
        RECT 65.770 167.285 69.080 167.455 ;
        RECT 69.505 167.285 71.015 167.455 ;
        RECT 71.185 167.285 73.535 167.455 ;
        RECT 73.705 167.285 80.365 167.455 ;
        RECT 81.060 167.435 81.230 168.035 ;
        RECT 81.915 168.020 82.205 169.185 ;
        RECT 82.895 168.125 83.225 168.970 ;
        RECT 83.395 168.175 83.565 169.185 ;
        RECT 83.735 168.455 84.075 169.015 ;
        RECT 84.305 168.685 84.620 169.185 ;
        RECT 84.800 168.715 85.685 168.885 ;
        RECT 82.835 168.045 83.225 168.125 ;
        RECT 83.735 168.080 84.630 168.455 ;
        RECT 82.835 167.995 83.050 168.045 ;
        RECT 81.400 167.605 81.735 167.875 ;
        RECT 65.340 166.635 65.600 167.160 ;
        RECT 65.770 166.830 66.030 167.285 ;
        RECT 66.200 166.635 66.460 167.115 ;
        RECT 66.630 166.830 66.890 167.285 ;
        RECT 67.060 166.635 67.320 167.115 ;
        RECT 67.490 166.830 67.750 167.285 ;
        RECT 67.920 166.635 68.180 167.115 ;
        RECT 68.350 166.830 68.610 167.285 ;
        RECT 68.780 166.635 69.080 167.115 ;
        RECT 69.505 166.810 69.835 167.285 ;
        RECT 70.005 166.635 70.175 167.115 ;
        RECT 70.345 166.810 70.675 167.285 ;
        RECT 70.845 166.635 71.015 167.115 ;
        RECT 71.185 166.810 71.515 167.285 ;
        RECT 71.685 166.635 71.855 167.115 ;
        RECT 72.025 166.810 72.355 167.285 ;
        RECT 72.525 166.635 72.695 167.115 ;
        RECT 72.865 166.810 73.195 167.285 ;
        RECT 73.365 166.635 73.535 167.115 ;
        RECT 73.705 166.810 74.035 167.285 ;
        RECT 73.705 166.805 73.955 166.810 ;
        RECT 74.205 166.635 74.375 167.115 ;
        RECT 74.545 166.810 74.875 167.285 ;
        RECT 74.625 166.805 74.795 166.810 ;
        RECT 75.045 166.635 75.215 167.115 ;
        RECT 75.385 166.810 75.715 167.285 ;
        RECT 75.465 166.805 75.635 166.810 ;
        RECT 75.885 166.635 76.055 167.115 ;
        RECT 76.225 166.810 76.555 167.285 ;
        RECT 76.725 166.635 76.895 167.115 ;
        RECT 77.065 166.810 77.395 167.285 ;
        RECT 77.565 166.635 77.735 167.115 ;
        RECT 77.905 166.810 78.235 167.285 ;
        RECT 78.405 166.635 78.575 167.115 ;
        RECT 78.745 166.810 79.075 167.285 ;
        RECT 79.245 166.635 79.415 167.115 ;
        RECT 79.585 166.810 79.915 167.285 ;
        RECT 80.085 166.635 80.255 167.115 ;
        RECT 80.535 166.805 81.230 167.435 ;
        RECT 81.435 166.635 81.745 167.435 ;
        RECT 82.835 167.415 83.005 167.995 ;
        RECT 83.735 167.875 83.925 168.080 ;
        RECT 84.800 167.875 84.970 168.715 ;
        RECT 85.910 168.685 86.160 169.015 ;
        RECT 83.175 167.545 83.925 167.875 ;
        RECT 84.095 167.545 84.970 167.875 ;
        RECT 82.835 167.375 83.060 167.415 ;
        RECT 83.725 167.375 83.925 167.545 ;
        RECT 81.915 166.635 82.205 167.360 ;
        RECT 82.835 167.290 83.215 167.375 ;
        RECT 82.885 166.855 83.215 167.290 ;
        RECT 83.385 166.635 83.555 167.245 ;
        RECT 83.725 166.850 84.055 167.375 ;
        RECT 84.315 166.635 84.525 167.165 ;
        RECT 84.800 167.085 84.970 167.545 ;
        RECT 85.140 167.585 85.460 168.545 ;
        RECT 85.630 167.795 85.820 168.515 ;
        RECT 85.990 167.615 86.160 168.685 ;
        RECT 86.330 168.385 86.500 169.185 ;
        RECT 86.670 168.740 87.775 168.910 ;
        RECT 86.670 168.125 86.840 168.740 ;
        RECT 87.985 168.590 88.235 169.015 ;
        RECT 88.405 168.725 88.670 169.185 ;
        RECT 87.010 168.205 87.540 168.570 ;
        RECT 87.985 168.460 88.290 168.590 ;
        RECT 86.330 168.035 86.840 168.125 ;
        RECT 86.330 167.865 87.200 168.035 ;
        RECT 86.330 167.795 86.500 167.865 ;
        RECT 86.620 167.615 86.820 167.645 ;
        RECT 85.140 167.255 85.605 167.585 ;
        RECT 85.990 167.315 86.820 167.615 ;
        RECT 85.990 167.085 86.160 167.315 ;
        RECT 84.800 166.915 85.585 167.085 ;
        RECT 85.755 166.915 86.160 167.085 ;
        RECT 86.340 166.635 86.710 167.135 ;
        RECT 87.030 167.085 87.200 167.865 ;
        RECT 87.370 167.505 87.540 168.205 ;
        RECT 87.710 167.675 87.950 168.270 ;
        RECT 87.370 167.285 87.895 167.505 ;
        RECT 88.120 167.355 88.290 168.460 ;
        RECT 88.065 167.225 88.290 167.355 ;
        RECT 88.460 167.265 88.740 168.215 ;
        RECT 88.065 167.085 88.235 167.225 ;
        RECT 87.030 166.915 87.705 167.085 ;
        RECT 87.900 166.915 88.235 167.085 ;
        RECT 88.405 166.635 88.655 167.095 ;
        RECT 88.910 166.895 89.095 169.015 ;
        RECT 89.265 168.685 89.595 169.185 ;
        RECT 89.765 168.515 89.935 169.015 ;
        RECT 89.270 168.345 89.935 168.515 ;
        RECT 90.285 168.515 90.455 169.015 ;
        RECT 90.625 168.685 90.955 169.185 ;
        RECT 90.285 168.345 90.950 168.515 ;
        RECT 89.270 167.355 89.500 168.345 ;
        RECT 89.670 167.525 90.020 168.175 ;
        RECT 90.200 167.525 90.550 168.175 ;
        RECT 90.720 167.355 90.950 168.345 ;
        RECT 89.270 167.185 89.935 167.355 ;
        RECT 89.265 166.635 89.595 167.015 ;
        RECT 89.765 166.895 89.935 167.185 ;
        RECT 90.285 167.185 90.950 167.355 ;
        RECT 90.285 166.895 90.455 167.185 ;
        RECT 90.625 166.635 90.955 167.015 ;
        RECT 91.125 166.895 91.310 169.015 ;
        RECT 91.550 168.725 91.815 169.185 ;
        RECT 91.985 168.590 92.235 169.015 ;
        RECT 92.445 168.740 93.550 168.910 ;
        RECT 91.930 168.460 92.235 168.590 ;
        RECT 91.480 167.265 91.760 168.215 ;
        RECT 91.930 167.355 92.100 168.460 ;
        RECT 92.270 167.675 92.510 168.270 ;
        RECT 92.680 168.205 93.210 168.570 ;
        RECT 92.680 167.505 92.850 168.205 ;
        RECT 93.380 168.125 93.550 168.740 ;
        RECT 93.720 168.385 93.890 169.185 ;
        RECT 94.060 168.685 94.310 169.015 ;
        RECT 94.535 168.715 95.420 168.885 ;
        RECT 93.380 168.035 93.890 168.125 ;
        RECT 91.930 167.225 92.155 167.355 ;
        RECT 92.325 167.285 92.850 167.505 ;
        RECT 93.020 167.865 93.890 168.035 ;
        RECT 91.565 166.635 91.815 167.095 ;
        RECT 91.985 167.085 92.155 167.225 ;
        RECT 93.020 167.085 93.190 167.865 ;
        RECT 93.720 167.795 93.890 167.865 ;
        RECT 93.400 167.615 93.600 167.645 ;
        RECT 94.060 167.615 94.230 168.685 ;
        RECT 94.400 167.795 94.590 168.515 ;
        RECT 93.400 167.315 94.230 167.615 ;
        RECT 94.760 167.585 95.080 168.545 ;
        RECT 91.985 166.915 92.320 167.085 ;
        RECT 92.515 166.915 93.190 167.085 ;
        RECT 93.510 166.635 93.880 167.135 ;
        RECT 94.060 167.085 94.230 167.315 ;
        RECT 94.615 167.255 95.080 167.585 ;
        RECT 95.250 167.875 95.420 168.715 ;
        RECT 95.600 168.685 95.915 169.185 ;
        RECT 96.145 168.455 96.485 169.015 ;
        RECT 95.590 168.080 96.485 168.455 ;
        RECT 96.655 168.175 96.825 169.185 ;
        RECT 96.295 167.875 96.485 168.080 ;
        RECT 96.995 168.125 97.325 168.970 ;
        RECT 96.995 168.045 97.385 168.125 ;
        RECT 97.555 168.095 99.225 169.185 ;
        RECT 99.455 168.125 99.785 168.970 ;
        RECT 99.955 168.175 100.125 169.185 ;
        RECT 100.295 168.455 100.635 169.015 ;
        RECT 100.865 168.685 101.180 169.185 ;
        RECT 101.360 168.715 102.245 168.885 ;
        RECT 97.170 167.995 97.385 168.045 ;
        RECT 95.250 167.545 96.125 167.875 ;
        RECT 96.295 167.545 97.045 167.875 ;
        RECT 95.250 167.085 95.420 167.545 ;
        RECT 96.295 167.375 96.495 167.545 ;
        RECT 97.215 167.415 97.385 167.995 ;
        RECT 97.160 167.375 97.385 167.415 ;
        RECT 94.060 166.915 94.465 167.085 ;
        RECT 94.635 166.915 95.420 167.085 ;
        RECT 95.695 166.635 95.905 167.165 ;
        RECT 96.165 166.850 96.495 167.375 ;
        RECT 97.005 167.290 97.385 167.375 ;
        RECT 97.555 167.405 98.305 167.925 ;
        RECT 98.475 167.575 99.225 168.095 ;
        RECT 99.395 168.045 99.785 168.125 ;
        RECT 100.295 168.080 101.190 168.455 ;
        RECT 99.395 167.995 99.610 168.045 ;
        RECT 99.395 167.415 99.565 167.995 ;
        RECT 100.295 167.875 100.485 168.080 ;
        RECT 101.360 167.875 101.530 168.715 ;
        RECT 102.470 168.685 102.720 169.015 ;
        RECT 99.735 167.545 100.485 167.875 ;
        RECT 100.655 167.545 101.530 167.875 ;
        RECT 96.665 166.635 96.835 167.245 ;
        RECT 97.005 166.855 97.335 167.290 ;
        RECT 97.555 166.635 99.225 167.405 ;
        RECT 99.395 167.375 99.620 167.415 ;
        RECT 100.285 167.375 100.485 167.545 ;
        RECT 99.395 167.290 99.775 167.375 ;
        RECT 99.445 166.855 99.775 167.290 ;
        RECT 99.945 166.635 100.115 167.245 ;
        RECT 100.285 166.850 100.615 167.375 ;
        RECT 100.875 166.635 101.085 167.165 ;
        RECT 101.360 167.085 101.530 167.545 ;
        RECT 101.700 167.585 102.020 168.545 ;
        RECT 102.190 167.795 102.380 168.515 ;
        RECT 102.550 167.615 102.720 168.685 ;
        RECT 102.890 168.385 103.060 169.185 ;
        RECT 103.230 168.740 104.335 168.910 ;
        RECT 103.230 168.125 103.400 168.740 ;
        RECT 104.545 168.590 104.795 169.015 ;
        RECT 104.965 168.725 105.230 169.185 ;
        RECT 103.570 168.205 104.100 168.570 ;
        RECT 104.545 168.460 104.850 168.590 ;
        RECT 102.890 168.035 103.400 168.125 ;
        RECT 102.890 167.865 103.760 168.035 ;
        RECT 102.890 167.795 103.060 167.865 ;
        RECT 103.180 167.615 103.380 167.645 ;
        RECT 101.700 167.255 102.165 167.585 ;
        RECT 102.550 167.315 103.380 167.615 ;
        RECT 102.550 167.085 102.720 167.315 ;
        RECT 101.360 166.915 102.145 167.085 ;
        RECT 102.315 166.915 102.720 167.085 ;
        RECT 102.900 166.635 103.270 167.135 ;
        RECT 103.590 167.085 103.760 167.865 ;
        RECT 103.930 167.505 104.100 168.205 ;
        RECT 104.270 167.675 104.510 168.270 ;
        RECT 103.930 167.285 104.455 167.505 ;
        RECT 104.680 167.355 104.850 168.460 ;
        RECT 104.625 167.225 104.850 167.355 ;
        RECT 105.020 167.265 105.300 168.215 ;
        RECT 104.625 167.085 104.795 167.225 ;
        RECT 103.590 166.915 104.265 167.085 ;
        RECT 104.460 166.915 104.795 167.085 ;
        RECT 104.965 166.635 105.215 167.095 ;
        RECT 105.470 166.895 105.655 169.015 ;
        RECT 105.825 168.685 106.155 169.185 ;
        RECT 106.325 168.515 106.495 169.015 ;
        RECT 105.830 168.345 106.495 168.515 ;
        RECT 105.830 167.355 106.060 168.345 ;
        RECT 106.230 167.525 106.580 168.175 ;
        RECT 107.675 168.020 107.965 169.185 ;
        RECT 108.250 168.555 108.535 169.015 ;
        RECT 108.705 168.725 108.975 169.185 ;
        RECT 108.250 168.335 109.205 168.555 ;
        RECT 108.135 167.605 108.825 168.165 ;
        RECT 108.995 167.435 109.205 168.335 ;
        RECT 105.830 167.185 106.495 167.355 ;
        RECT 105.825 166.635 106.155 167.015 ;
        RECT 106.325 166.895 106.495 167.185 ;
        RECT 107.675 166.635 107.965 167.360 ;
        RECT 108.250 167.265 109.205 167.435 ;
        RECT 109.375 168.165 109.775 169.015 ;
        RECT 109.965 168.555 110.245 169.015 ;
        RECT 110.765 168.725 111.090 169.185 ;
        RECT 109.965 168.335 111.090 168.555 ;
        RECT 109.375 167.605 110.470 168.165 ;
        RECT 110.640 167.875 111.090 168.335 ;
        RECT 111.260 168.045 111.645 169.015 ;
        RECT 108.250 166.805 108.535 167.265 ;
        RECT 108.705 166.635 108.975 167.095 ;
        RECT 109.375 166.805 109.775 167.605 ;
        RECT 110.640 167.545 111.195 167.875 ;
        RECT 110.640 167.435 111.090 167.545 ;
        RECT 109.965 167.265 111.090 167.435 ;
        RECT 111.365 167.375 111.645 168.045 ;
        RECT 109.965 166.805 110.245 167.265 ;
        RECT 110.765 166.635 111.090 167.095 ;
        RECT 111.260 166.805 111.645 167.375 ;
        RECT 111.815 168.385 112.255 169.015 ;
        RECT 111.815 167.375 112.125 168.385 ;
        RECT 112.430 168.335 112.745 169.185 ;
        RECT 112.915 168.845 114.345 169.015 ;
        RECT 112.915 168.165 113.085 168.845 ;
        RECT 112.295 167.995 113.085 168.165 ;
        RECT 112.295 167.545 112.465 167.995 ;
        RECT 113.255 167.875 113.455 168.675 ;
        RECT 112.635 167.545 113.025 167.825 ;
        RECT 113.210 167.545 113.455 167.875 ;
        RECT 113.655 167.545 113.905 168.675 ;
        RECT 114.095 168.215 114.345 168.845 ;
        RECT 114.525 168.385 114.855 169.185 ;
        RECT 114.095 168.045 114.865 168.215 ;
        RECT 114.120 167.545 114.525 167.875 ;
        RECT 114.695 167.375 114.865 168.045 ;
        RECT 111.815 166.815 112.255 167.375 ;
        RECT 112.425 166.635 112.875 167.375 ;
        RECT 113.045 167.205 114.205 167.375 ;
        RECT 113.045 166.805 113.215 167.205 ;
        RECT 113.385 166.635 113.805 167.035 ;
        RECT 113.975 166.805 114.205 167.205 ;
        RECT 114.375 166.805 114.865 167.375 ;
        RECT 115.045 168.125 115.375 168.975 ;
        RECT 115.045 167.995 115.265 168.125 ;
        RECT 115.545 168.045 115.795 169.185 ;
        RECT 115.985 168.545 116.235 168.965 ;
        RECT 116.465 168.715 116.795 169.185 ;
        RECT 117.025 168.545 117.275 168.965 ;
        RECT 115.985 168.375 117.275 168.545 ;
        RECT 117.455 168.545 117.785 168.975 ;
        RECT 117.455 168.375 117.910 168.545 ;
        RECT 115.045 167.360 115.235 167.995 ;
        RECT 115.975 167.875 116.190 168.205 ;
        RECT 115.405 167.545 115.715 167.875 ;
        RECT 115.885 167.545 116.190 167.875 ;
        RECT 116.365 167.545 116.650 168.205 ;
        RECT 116.845 167.545 117.110 168.205 ;
        RECT 117.325 167.545 117.570 168.205 ;
        RECT 115.545 167.375 115.715 167.545 ;
        RECT 117.740 167.375 117.910 168.375 ;
        RECT 118.255 168.095 119.925 169.185 ;
        RECT 115.045 166.850 115.375 167.360 ;
        RECT 115.545 167.205 117.910 167.375 ;
        RECT 118.255 167.405 119.005 167.925 ;
        RECT 119.175 167.575 119.925 168.095 ;
        RECT 120.115 168.295 120.375 169.005 ;
        RECT 120.545 168.475 120.875 169.185 ;
        RECT 121.045 168.295 121.275 169.005 ;
        RECT 120.115 168.055 121.275 168.295 ;
        RECT 121.455 168.275 121.725 169.005 ;
        RECT 121.905 168.455 122.245 169.185 ;
        RECT 121.455 168.055 122.225 168.275 ;
        RECT 120.105 167.545 120.405 167.875 ;
        RECT 120.585 167.565 121.110 167.875 ;
        RECT 121.290 167.565 121.755 167.875 ;
        RECT 115.545 166.635 115.875 167.035 ;
        RECT 116.925 166.865 117.255 167.205 ;
        RECT 117.425 166.635 117.755 167.035 ;
        RECT 118.255 166.635 119.925 167.405 ;
        RECT 120.115 166.635 120.405 167.365 ;
        RECT 120.585 166.925 120.815 167.565 ;
        RECT 121.935 167.385 122.225 168.055 ;
        RECT 120.995 167.185 122.225 167.385 ;
        RECT 120.995 166.815 121.305 167.185 ;
        RECT 121.485 166.635 122.155 167.005 ;
        RECT 122.415 166.815 122.675 169.005 ;
        RECT 122.890 168.395 123.425 169.015 ;
        RECT 122.890 167.375 123.205 168.395 ;
        RECT 123.595 168.385 123.925 169.185 ;
        RECT 125.155 168.750 130.500 169.185 ;
        RECT 124.410 168.215 124.800 168.390 ;
        RECT 123.375 168.045 124.800 168.215 ;
        RECT 123.375 167.545 123.545 168.045 ;
        RECT 122.890 166.805 123.505 167.375 ;
        RECT 123.795 167.315 124.060 167.875 ;
        RECT 124.230 167.145 124.400 168.045 ;
        RECT 124.570 167.315 124.925 167.875 ;
        RECT 126.740 167.180 127.080 168.010 ;
        RECT 128.560 167.500 128.910 168.750 ;
        RECT 131.685 168.255 131.855 169.015 ;
        RECT 132.070 168.425 132.400 169.185 ;
        RECT 131.685 168.085 132.400 168.255 ;
        RECT 132.570 168.110 132.825 169.015 ;
        RECT 131.595 167.535 131.950 167.905 ;
        RECT 132.230 167.875 132.400 168.085 ;
        RECT 132.230 167.545 132.485 167.875 ;
        RECT 132.230 167.355 132.400 167.545 ;
        RECT 132.655 167.380 132.825 168.110 ;
        RECT 133.000 168.035 133.260 169.185 ;
        RECT 133.435 168.020 133.725 169.185 ;
        RECT 133.900 168.045 134.235 169.015 ;
        RECT 134.405 168.045 134.575 169.185 ;
        RECT 134.745 168.845 136.775 169.015 ;
        RECT 131.685 167.185 132.400 167.355 ;
        RECT 123.675 166.635 123.890 167.145 ;
        RECT 124.120 166.815 124.400 167.145 ;
        RECT 124.580 166.635 124.820 167.145 ;
        RECT 125.155 166.635 130.500 167.180 ;
        RECT 131.685 166.805 131.855 167.185 ;
        RECT 132.070 166.635 132.400 167.015 ;
        RECT 132.570 166.805 132.825 167.380 ;
        RECT 133.000 166.635 133.260 167.475 ;
        RECT 133.900 167.375 134.070 168.045 ;
        RECT 134.745 167.875 134.915 168.845 ;
        RECT 134.240 167.545 134.495 167.875 ;
        RECT 134.720 167.545 134.915 167.875 ;
        RECT 135.085 168.505 136.210 168.675 ;
        RECT 134.325 167.375 134.495 167.545 ;
        RECT 135.085 167.375 135.255 168.505 ;
        RECT 133.435 166.635 133.725 167.360 ;
        RECT 133.900 166.805 134.155 167.375 ;
        RECT 134.325 167.205 135.255 167.375 ;
        RECT 135.425 168.165 136.435 168.335 ;
        RECT 135.425 167.365 135.595 168.165 ;
        RECT 135.800 167.485 136.075 167.965 ;
        RECT 135.795 167.315 136.075 167.485 ;
        RECT 135.080 167.170 135.255 167.205 ;
        RECT 134.325 166.635 134.655 167.035 ;
        RECT 135.080 166.805 135.610 167.170 ;
        RECT 135.800 166.805 136.075 167.315 ;
        RECT 136.245 166.805 136.435 168.165 ;
        RECT 136.605 168.180 136.775 168.845 ;
        RECT 136.945 168.425 137.115 169.185 ;
        RECT 137.350 168.425 137.865 168.835 ;
        RECT 136.605 167.990 137.355 168.180 ;
        RECT 137.525 167.615 137.865 168.425 ;
        RECT 136.635 167.445 137.865 167.615 ;
        RECT 138.035 168.045 138.420 169.015 ;
        RECT 138.590 168.725 138.915 169.185 ;
        RECT 139.435 168.555 139.715 169.015 ;
        RECT 138.590 168.335 139.715 168.555 ;
        RECT 136.615 166.635 137.125 167.170 ;
        RECT 137.345 166.840 137.590 167.445 ;
        RECT 138.035 167.375 138.315 168.045 ;
        RECT 138.590 167.875 139.040 168.335 ;
        RECT 139.905 168.165 140.305 169.015 ;
        RECT 140.705 168.725 140.975 169.185 ;
        RECT 141.145 168.555 141.430 169.015 ;
        RECT 138.485 167.545 139.040 167.875 ;
        RECT 139.210 167.605 140.305 168.165 ;
        RECT 138.590 167.435 139.040 167.545 ;
        RECT 138.035 166.805 138.420 167.375 ;
        RECT 138.590 167.265 139.715 167.435 ;
        RECT 138.590 166.635 138.915 167.095 ;
        RECT 139.435 166.805 139.715 167.265 ;
        RECT 139.905 166.805 140.305 167.605 ;
        RECT 140.475 168.335 141.430 168.555 ;
        RECT 140.475 167.435 140.685 168.335 ;
        RECT 140.855 167.605 141.545 168.165 ;
        RECT 141.715 168.095 142.925 169.185 ;
        RECT 141.715 167.555 142.235 168.095 ;
        RECT 140.475 167.265 141.430 167.435 ;
        RECT 142.405 167.385 142.925 167.925 ;
        RECT 140.705 166.635 140.975 167.095 ;
        RECT 141.145 166.805 141.430 167.265 ;
        RECT 141.715 166.635 142.925 167.385 ;
        RECT 17.430 166.465 143.010 166.635 ;
        RECT 17.515 165.715 18.725 166.465 ;
        RECT 17.515 165.175 18.035 165.715 ;
        RECT 18.895 165.695 21.485 166.465 ;
        RECT 22.165 166.075 22.495 166.465 ;
        RECT 22.665 165.895 22.835 166.215 ;
        RECT 23.005 166.075 23.335 166.465 ;
        RECT 23.750 166.065 24.705 166.235 ;
        RECT 22.115 165.725 24.365 165.895 ;
        RECT 18.205 165.005 18.725 165.545 ;
        RECT 18.895 165.175 20.105 165.695 ;
        RECT 20.275 165.005 21.485 165.525 ;
        RECT 17.515 163.915 18.725 165.005 ;
        RECT 18.895 163.915 21.485 165.005 ;
        RECT 22.115 164.765 22.285 165.725 ;
        RECT 22.455 165.105 22.700 165.555 ;
        RECT 22.870 165.275 23.420 165.475 ;
        RECT 23.590 165.305 23.965 165.475 ;
        RECT 23.590 165.105 23.760 165.305 ;
        RECT 24.135 165.225 24.365 165.725 ;
        RECT 22.455 164.935 23.760 165.105 ;
        RECT 24.535 165.185 24.705 166.065 ;
        RECT 24.875 165.630 25.165 166.465 ;
        RECT 25.340 166.065 25.675 166.465 ;
        RECT 25.845 165.895 26.050 166.295 ;
        RECT 26.260 165.985 26.535 166.465 ;
        RECT 26.745 165.965 27.005 166.295 ;
        RECT 25.365 165.725 26.050 165.895 ;
        RECT 24.535 165.015 25.165 165.185 ;
        RECT 22.115 164.085 22.495 164.765 ;
        RECT 23.085 163.915 23.255 164.765 ;
        RECT 23.425 164.595 24.665 164.765 ;
        RECT 23.425 164.085 23.755 164.595 ;
        RECT 23.925 163.915 24.095 164.425 ;
        RECT 24.265 164.085 24.665 164.595 ;
        RECT 24.845 164.085 25.165 165.015 ;
        RECT 25.365 164.695 25.705 165.725 ;
        RECT 25.875 165.055 26.125 165.555 ;
        RECT 26.305 165.225 26.665 165.805 ;
        RECT 26.835 165.055 27.005 165.965 ;
        RECT 27.175 165.695 29.765 166.465 ;
        RECT 29.935 165.725 30.400 166.270 ;
        RECT 27.175 165.175 28.385 165.695 ;
        RECT 25.875 164.885 27.005 165.055 ;
        RECT 28.555 165.005 29.765 165.525 ;
        RECT 25.365 164.520 26.030 164.695 ;
        RECT 25.340 163.915 25.675 164.340 ;
        RECT 25.845 164.115 26.030 164.520 ;
        RECT 26.235 163.915 26.565 164.695 ;
        RECT 26.735 164.115 27.005 164.885 ;
        RECT 27.175 163.915 29.765 165.005 ;
        RECT 29.935 164.765 30.105 165.725 ;
        RECT 30.905 165.645 31.075 166.465 ;
        RECT 31.245 165.815 31.575 166.295 ;
        RECT 31.745 166.075 32.095 166.465 ;
        RECT 32.265 165.895 32.495 166.295 ;
        RECT 31.985 165.815 32.495 165.895 ;
        RECT 31.245 165.725 32.495 165.815 ;
        RECT 32.665 165.725 32.985 166.205 ;
        RECT 31.245 165.645 32.155 165.725 ;
        RECT 30.275 165.105 30.520 165.555 ;
        RECT 30.780 165.275 31.475 165.475 ;
        RECT 31.645 165.305 32.245 165.475 ;
        RECT 31.645 165.105 31.815 165.305 ;
        RECT 32.475 165.135 32.645 165.555 ;
        RECT 30.275 164.935 31.815 165.105 ;
        RECT 31.985 164.965 32.645 165.135 ;
        RECT 31.985 164.765 32.155 164.965 ;
        RECT 32.815 164.795 32.985 165.725 ;
        RECT 29.935 164.595 32.155 164.765 ;
        RECT 32.325 164.595 32.985 164.795 ;
        RECT 33.155 165.725 33.620 166.270 ;
        RECT 33.155 164.765 33.325 165.725 ;
        RECT 34.125 165.645 34.295 166.465 ;
        RECT 34.465 165.815 34.795 166.295 ;
        RECT 34.965 166.075 35.315 166.465 ;
        RECT 35.485 165.895 35.715 166.295 ;
        RECT 35.205 165.815 35.715 165.895 ;
        RECT 34.465 165.725 35.715 165.815 ;
        RECT 35.885 165.725 36.205 166.205 ;
        RECT 34.465 165.645 35.375 165.725 ;
        RECT 33.495 165.105 33.740 165.555 ;
        RECT 34.000 165.275 34.695 165.475 ;
        RECT 34.865 165.305 35.465 165.475 ;
        RECT 34.865 165.105 35.035 165.305 ;
        RECT 35.695 165.135 35.865 165.555 ;
        RECT 33.495 164.935 35.035 165.105 ;
        RECT 35.205 164.965 35.865 165.135 ;
        RECT 35.205 164.765 35.375 164.965 ;
        RECT 36.035 164.795 36.205 165.725 ;
        RECT 36.375 165.695 38.965 166.465 ;
        RECT 39.610 165.895 39.865 166.245 ;
        RECT 40.035 166.065 40.365 166.465 ;
        RECT 40.535 165.895 40.705 166.245 ;
        RECT 40.875 166.065 41.255 166.465 ;
        RECT 39.610 165.725 41.275 165.895 ;
        RECT 41.445 165.790 41.720 166.135 ;
        RECT 36.375 165.175 37.585 165.695 ;
        RECT 41.105 165.555 41.275 165.725 ;
        RECT 37.755 165.005 38.965 165.525 ;
        RECT 39.595 165.225 39.940 165.555 ;
        RECT 40.110 165.225 40.935 165.555 ;
        RECT 41.105 165.225 41.380 165.555 ;
        RECT 33.155 164.595 35.375 164.765 ;
        RECT 35.545 164.595 36.205 164.795 ;
        RECT 29.935 163.915 30.235 164.425 ;
        RECT 30.405 164.085 30.735 164.595 ;
        RECT 32.325 164.425 32.495 164.595 ;
        RECT 30.905 163.915 31.535 164.425 ;
        RECT 32.115 164.255 32.495 164.425 ;
        RECT 32.665 163.915 32.965 164.425 ;
        RECT 33.155 163.915 33.455 164.425 ;
        RECT 33.625 164.085 33.955 164.595 ;
        RECT 35.545 164.425 35.715 164.595 ;
        RECT 34.125 163.915 34.755 164.425 ;
        RECT 35.335 164.255 35.715 164.425 ;
        RECT 35.885 163.915 36.185 164.425 ;
        RECT 36.375 163.915 38.965 165.005 ;
        RECT 39.615 164.765 39.940 165.055 ;
        RECT 40.110 164.935 40.305 165.225 ;
        RECT 41.105 165.055 41.275 165.225 ;
        RECT 41.550 165.055 41.720 165.790 ;
        RECT 41.895 165.715 43.105 166.465 ;
        RECT 43.275 165.740 43.565 166.465 ;
        RECT 43.825 165.815 43.995 166.295 ;
        RECT 44.165 165.985 44.495 166.465 ;
        RECT 44.720 166.045 46.255 166.295 ;
        RECT 44.720 165.815 44.890 166.045 ;
        RECT 41.895 165.175 42.415 165.715 ;
        RECT 43.825 165.645 44.890 165.815 ;
        RECT 40.615 164.885 41.275 165.055 ;
        RECT 40.615 164.765 40.785 164.885 ;
        RECT 39.615 164.595 40.785 164.765 ;
        RECT 39.595 164.135 40.785 164.425 ;
        RECT 40.955 163.915 41.235 164.715 ;
        RECT 41.445 164.085 41.720 165.055 ;
        RECT 42.585 165.005 43.105 165.545 ;
        RECT 45.070 165.475 45.350 165.875 ;
        RECT 43.740 165.265 44.090 165.475 ;
        RECT 44.260 165.275 44.705 165.475 ;
        RECT 44.875 165.275 45.350 165.475 ;
        RECT 45.620 165.475 45.905 165.875 ;
        RECT 46.085 165.815 46.255 166.045 ;
        RECT 46.425 165.985 46.755 166.465 ;
        RECT 46.970 165.965 47.225 166.295 ;
        RECT 47.040 165.885 47.225 165.965 ;
        RECT 47.415 165.920 52.760 166.465 ;
        RECT 52.985 166.075 53.315 166.465 ;
        RECT 46.085 165.645 46.885 165.815 ;
        RECT 45.620 165.275 45.950 165.475 ;
        RECT 46.120 165.445 46.485 165.475 ;
        RECT 46.120 165.275 46.495 165.445 ;
        RECT 46.715 165.095 46.885 165.645 ;
        RECT 41.895 163.915 43.105 165.005 ;
        RECT 43.275 163.915 43.565 165.080 ;
        RECT 43.825 164.925 46.885 165.095 ;
        RECT 43.825 164.085 43.995 164.925 ;
        RECT 47.055 164.755 47.225 165.885 ;
        RECT 49.000 165.090 49.340 165.920 ;
        RECT 53.485 165.895 53.655 166.215 ;
        RECT 53.825 166.075 54.155 166.465 ;
        RECT 54.570 166.065 55.525 166.235 ;
        RECT 52.935 165.725 55.185 165.895 ;
        RECT 44.165 164.255 44.495 164.755 ;
        RECT 44.665 164.515 46.300 164.755 ;
        RECT 44.665 164.425 44.895 164.515 ;
        RECT 45.005 164.255 45.335 164.295 ;
        RECT 44.165 164.085 45.335 164.255 ;
        RECT 45.525 163.915 45.880 164.335 ;
        RECT 46.050 164.085 46.300 164.515 ;
        RECT 46.470 163.915 46.800 164.675 ;
        RECT 46.970 164.085 47.225 164.755 ;
        RECT 50.820 164.350 51.170 165.600 ;
        RECT 52.935 164.765 53.105 165.725 ;
        RECT 53.275 165.105 53.520 165.555 ;
        RECT 53.690 165.275 54.240 165.475 ;
        RECT 54.410 165.305 54.785 165.475 ;
        RECT 54.410 165.105 54.580 165.305 ;
        RECT 54.955 165.225 55.185 165.725 ;
        RECT 53.275 164.935 54.580 165.105 ;
        RECT 55.355 165.185 55.525 166.065 ;
        RECT 55.695 165.630 55.985 166.465 ;
        RECT 56.160 166.065 56.495 166.465 ;
        RECT 56.665 165.895 56.870 166.295 ;
        RECT 57.080 165.985 57.355 166.465 ;
        RECT 57.565 165.965 57.825 166.295 ;
        RECT 56.185 165.725 56.870 165.895 ;
        RECT 55.355 165.015 55.985 165.185 ;
        RECT 47.415 163.915 52.760 164.350 ;
        RECT 52.935 164.085 53.315 164.765 ;
        RECT 53.905 163.915 54.075 164.765 ;
        RECT 54.245 164.595 55.485 164.765 ;
        RECT 54.245 164.085 54.575 164.595 ;
        RECT 54.745 163.915 54.915 164.425 ;
        RECT 55.085 164.085 55.485 164.595 ;
        RECT 55.665 164.085 55.985 165.015 ;
        RECT 56.185 164.695 56.525 165.725 ;
        RECT 56.695 165.055 56.945 165.555 ;
        RECT 57.125 165.225 57.485 165.805 ;
        RECT 57.655 165.055 57.825 165.965 ;
        RECT 57.995 165.920 63.340 166.465 ;
        RECT 59.580 165.090 59.920 165.920 ;
        RECT 63.515 165.695 65.185 166.465 ;
        RECT 65.360 165.935 65.650 166.285 ;
        RECT 65.845 166.105 66.175 166.465 ;
        RECT 66.345 165.935 66.575 166.240 ;
        RECT 65.360 165.765 66.575 165.935 ;
        RECT 66.765 165.785 66.935 166.160 ;
        RECT 56.695 164.885 57.825 165.055 ;
        RECT 56.185 164.520 56.850 164.695 ;
        RECT 56.160 163.915 56.495 164.340 ;
        RECT 56.665 164.115 56.850 164.520 ;
        RECT 57.055 163.915 57.385 164.695 ;
        RECT 57.555 164.115 57.825 164.885 ;
        RECT 61.400 164.350 61.750 165.600 ;
        RECT 63.515 165.175 64.265 165.695 ;
        RECT 66.765 165.615 66.965 165.785 ;
        RECT 67.195 165.695 68.865 166.465 ;
        RECT 69.035 165.740 69.325 166.465 ;
        RECT 69.585 165.915 69.755 166.205 ;
        RECT 69.925 166.085 70.255 166.465 ;
        RECT 69.585 165.745 70.250 165.915 ;
        RECT 66.765 165.595 66.935 165.615 ;
        RECT 64.435 165.005 65.185 165.525 ;
        RECT 65.420 165.445 65.680 165.555 ;
        RECT 65.415 165.275 65.680 165.445 ;
        RECT 65.420 165.225 65.680 165.275 ;
        RECT 65.860 165.225 66.245 165.555 ;
        RECT 66.415 165.425 66.935 165.595 ;
        RECT 57.995 163.915 63.340 164.350 ;
        RECT 63.515 163.915 65.185 165.005 ;
        RECT 65.360 163.915 65.680 165.055 ;
        RECT 65.860 164.175 66.055 165.225 ;
        RECT 66.415 165.045 66.585 165.425 ;
        RECT 66.235 164.765 66.585 165.045 ;
        RECT 66.775 164.895 67.020 165.255 ;
        RECT 67.195 165.175 67.945 165.695 ;
        RECT 68.115 165.005 68.865 165.525 ;
        RECT 66.235 164.085 66.565 164.765 ;
        RECT 66.765 163.915 67.020 164.715 ;
        RECT 67.195 163.915 68.865 165.005 ;
        RECT 69.035 163.915 69.325 165.080 ;
        RECT 69.500 164.925 69.850 165.575 ;
        RECT 70.020 164.755 70.250 165.745 ;
        RECT 69.585 164.585 70.250 164.755 ;
        RECT 69.585 164.085 69.755 164.585 ;
        RECT 69.925 163.915 70.255 164.415 ;
        RECT 70.425 164.085 70.610 166.205 ;
        RECT 70.865 166.005 71.115 166.465 ;
        RECT 71.285 166.015 71.620 166.185 ;
        RECT 71.815 166.015 72.490 166.185 ;
        RECT 71.285 165.875 71.455 166.015 ;
        RECT 70.780 164.885 71.060 165.835 ;
        RECT 71.230 165.745 71.455 165.875 ;
        RECT 71.230 164.640 71.400 165.745 ;
        RECT 71.625 165.595 72.150 165.815 ;
        RECT 71.570 164.830 71.810 165.425 ;
        RECT 71.980 164.895 72.150 165.595 ;
        RECT 72.320 165.235 72.490 166.015 ;
        RECT 72.810 165.965 73.180 166.465 ;
        RECT 73.360 166.015 73.765 166.185 ;
        RECT 73.935 166.015 74.720 166.185 ;
        RECT 73.360 165.785 73.530 166.015 ;
        RECT 72.700 165.485 73.530 165.785 ;
        RECT 73.915 165.515 74.380 165.845 ;
        RECT 72.700 165.455 72.900 165.485 ;
        RECT 73.020 165.235 73.190 165.305 ;
        RECT 72.320 165.065 73.190 165.235 ;
        RECT 72.680 164.975 73.190 165.065 ;
        RECT 71.230 164.510 71.535 164.640 ;
        RECT 71.980 164.530 72.510 164.895 ;
        RECT 70.850 163.915 71.115 164.375 ;
        RECT 71.285 164.085 71.535 164.510 ;
        RECT 72.680 164.360 72.850 164.975 ;
        RECT 71.745 164.190 72.850 164.360 ;
        RECT 73.020 163.915 73.190 164.715 ;
        RECT 73.360 164.415 73.530 165.485 ;
        RECT 73.700 164.585 73.890 165.305 ;
        RECT 74.060 164.555 74.380 165.515 ;
        RECT 74.550 165.555 74.720 166.015 ;
        RECT 74.995 165.935 75.205 166.465 ;
        RECT 75.465 165.725 75.795 166.250 ;
        RECT 75.965 165.855 76.135 166.465 ;
        RECT 76.305 165.810 76.635 166.245 ;
        RECT 76.305 165.725 76.685 165.810 ;
        RECT 75.595 165.555 75.795 165.725 ;
        RECT 76.460 165.685 76.685 165.725 ;
        RECT 74.550 165.225 75.425 165.555 ;
        RECT 75.595 165.225 76.345 165.555 ;
        RECT 73.360 164.085 73.610 164.415 ;
        RECT 74.550 164.385 74.720 165.225 ;
        RECT 75.595 165.020 75.785 165.225 ;
        RECT 76.515 165.105 76.685 165.685 ;
        RECT 76.855 165.715 78.065 166.465 ;
        RECT 78.350 165.835 78.635 166.295 ;
        RECT 78.805 166.005 79.075 166.465 ;
        RECT 76.855 165.175 77.375 165.715 ;
        RECT 78.350 165.665 79.305 165.835 ;
        RECT 76.470 165.055 76.685 165.105 ;
        RECT 74.890 164.645 75.785 165.020 ;
        RECT 76.295 164.975 76.685 165.055 ;
        RECT 77.545 165.005 78.065 165.545 ;
        RECT 73.835 164.215 74.720 164.385 ;
        RECT 74.900 163.915 75.215 164.415 ;
        RECT 75.445 164.085 75.785 164.645 ;
        RECT 75.955 163.915 76.125 164.925 ;
        RECT 76.295 164.130 76.625 164.975 ;
        RECT 76.855 163.915 78.065 165.005 ;
        RECT 78.235 164.935 78.925 165.495 ;
        RECT 79.095 164.765 79.305 165.665 ;
        RECT 78.350 164.545 79.305 164.765 ;
        RECT 79.475 165.495 79.875 166.295 ;
        RECT 80.065 165.835 80.345 166.295 ;
        RECT 80.865 166.005 81.190 166.465 ;
        RECT 80.065 165.665 81.190 165.835 ;
        RECT 81.360 165.725 81.745 166.295 ;
        RECT 80.740 165.555 81.190 165.665 ;
        RECT 79.475 164.935 80.570 165.495 ;
        RECT 80.740 165.225 81.295 165.555 ;
        RECT 78.350 164.085 78.635 164.545 ;
        RECT 78.805 163.915 79.075 164.375 ;
        RECT 79.475 164.085 79.875 164.935 ;
        RECT 80.740 164.765 81.190 165.225 ;
        RECT 81.465 165.055 81.745 165.725 ;
        RECT 80.065 164.545 81.190 164.765 ;
        RECT 80.065 164.085 80.345 164.545 ;
        RECT 80.865 163.915 81.190 164.375 ;
        RECT 81.360 164.085 81.745 165.055 ;
        RECT 81.920 165.725 82.175 166.295 ;
        RECT 82.345 166.065 82.675 166.465 ;
        RECT 83.100 165.930 83.630 166.295 ;
        RECT 83.820 166.125 84.095 166.295 ;
        RECT 83.815 165.955 84.095 166.125 ;
        RECT 83.100 165.895 83.275 165.930 ;
        RECT 82.345 165.725 83.275 165.895 ;
        RECT 81.920 165.055 82.090 165.725 ;
        RECT 82.345 165.555 82.515 165.725 ;
        RECT 82.260 165.225 82.515 165.555 ;
        RECT 82.740 165.225 82.935 165.555 ;
        RECT 81.920 164.085 82.255 165.055 ;
        RECT 82.425 163.915 82.595 165.055 ;
        RECT 82.765 164.255 82.935 165.225 ;
        RECT 83.105 164.595 83.275 165.725 ;
        RECT 83.445 164.935 83.615 165.735 ;
        RECT 83.820 165.135 84.095 165.955 ;
        RECT 84.265 164.935 84.455 166.295 ;
        RECT 84.635 165.930 85.145 166.465 ;
        RECT 85.365 165.655 85.610 166.260 ;
        RECT 86.060 165.725 86.315 166.295 ;
        RECT 86.485 166.065 86.815 166.465 ;
        RECT 87.240 165.930 87.770 166.295 ;
        RECT 87.240 165.895 87.415 165.930 ;
        RECT 86.485 165.725 87.415 165.895 ;
        RECT 84.655 165.485 85.885 165.655 ;
        RECT 83.445 164.765 84.455 164.935 ;
        RECT 84.625 164.920 85.375 165.110 ;
        RECT 83.105 164.425 84.230 164.595 ;
        RECT 84.625 164.255 84.795 164.920 ;
        RECT 85.545 164.675 85.885 165.485 ;
        RECT 82.765 164.085 84.795 164.255 ;
        RECT 84.965 163.915 85.135 164.675 ;
        RECT 85.370 164.265 85.885 164.675 ;
        RECT 86.060 165.055 86.230 165.725 ;
        RECT 86.485 165.555 86.655 165.725 ;
        RECT 86.400 165.225 86.655 165.555 ;
        RECT 86.880 165.225 87.075 165.555 ;
        RECT 86.060 164.085 86.395 165.055 ;
        RECT 86.565 163.915 86.735 165.055 ;
        RECT 86.905 164.255 87.075 165.225 ;
        RECT 87.245 164.595 87.415 165.725 ;
        RECT 87.585 164.935 87.755 165.735 ;
        RECT 87.960 165.445 88.235 166.295 ;
        RECT 87.955 165.275 88.235 165.445 ;
        RECT 87.960 165.135 88.235 165.275 ;
        RECT 88.405 164.935 88.595 166.295 ;
        RECT 88.775 165.930 89.285 166.465 ;
        RECT 89.505 165.655 89.750 166.260 ;
        RECT 90.195 165.695 93.705 166.465 ;
        RECT 94.795 165.740 95.085 166.465 ;
        RECT 95.255 165.695 97.845 166.465 ;
        RECT 98.075 166.005 98.320 166.465 ;
        RECT 88.795 165.485 90.025 165.655 ;
        RECT 87.585 164.765 88.595 164.935 ;
        RECT 88.765 164.920 89.515 165.110 ;
        RECT 87.245 164.425 88.370 164.595 ;
        RECT 88.765 164.255 88.935 164.920 ;
        RECT 89.685 164.675 90.025 165.485 ;
        RECT 90.195 165.175 91.845 165.695 ;
        RECT 92.015 165.005 93.705 165.525 ;
        RECT 95.255 165.175 96.465 165.695 ;
        RECT 86.905 164.085 88.935 164.255 ;
        RECT 89.105 163.915 89.275 164.675 ;
        RECT 89.510 164.265 90.025 164.675 ;
        RECT 90.195 163.915 93.705 165.005 ;
        RECT 94.795 163.915 95.085 165.080 ;
        RECT 96.635 165.005 97.845 165.525 ;
        RECT 98.015 165.225 98.330 165.835 ;
        RECT 98.500 165.475 98.750 166.285 ;
        RECT 98.920 165.940 99.180 166.465 ;
        RECT 99.350 165.815 99.610 166.270 ;
        RECT 99.780 165.985 100.040 166.465 ;
        RECT 100.210 165.815 100.470 166.270 ;
        RECT 100.640 165.985 100.900 166.465 ;
        RECT 101.070 165.815 101.330 166.270 ;
        RECT 101.500 165.985 101.760 166.465 ;
        RECT 101.930 165.815 102.190 166.270 ;
        RECT 102.360 165.985 102.660 166.465 ;
        RECT 99.350 165.645 102.660 165.815 ;
        RECT 98.500 165.225 101.520 165.475 ;
        RECT 95.255 163.915 97.845 165.005 ;
        RECT 98.025 163.915 98.320 165.025 ;
        RECT 98.500 164.090 98.750 165.225 ;
        RECT 101.690 165.055 102.660 165.645 ;
        RECT 103.075 165.695 105.665 166.465 ;
        RECT 103.075 165.175 104.285 165.695 ;
        RECT 106.295 165.665 106.605 166.465 ;
        RECT 106.810 165.665 107.505 166.295 ;
        RECT 107.675 165.920 113.020 166.465 ;
        RECT 98.920 163.915 99.180 165.025 ;
        RECT 99.350 164.815 102.660 165.055 ;
        RECT 104.455 165.005 105.665 165.525 ;
        RECT 106.305 165.225 106.640 165.495 ;
        RECT 106.810 165.065 106.980 165.665 ;
        RECT 107.150 165.225 107.485 165.475 ;
        RECT 109.260 165.090 109.600 165.920 ;
        RECT 113.195 165.695 116.705 166.465 ;
        RECT 117.335 165.815 117.595 166.295 ;
        RECT 117.765 165.925 118.015 166.465 ;
        RECT 99.350 164.090 99.610 164.815 ;
        RECT 99.780 163.915 100.040 164.645 ;
        RECT 100.210 164.090 100.470 164.815 ;
        RECT 100.640 163.915 100.900 164.645 ;
        RECT 101.070 164.090 101.330 164.815 ;
        RECT 101.500 163.915 101.760 164.645 ;
        RECT 101.930 164.090 102.190 164.815 ;
        RECT 102.360 163.915 102.655 164.645 ;
        RECT 103.075 163.915 105.665 165.005 ;
        RECT 106.295 163.915 106.575 165.055 ;
        RECT 106.745 164.085 107.075 165.065 ;
        RECT 107.245 163.915 107.505 165.055 ;
        RECT 111.080 164.350 111.430 165.600 ;
        RECT 113.195 165.175 114.845 165.695 ;
        RECT 115.015 165.005 116.705 165.525 ;
        RECT 107.675 163.915 113.020 164.350 ;
        RECT 113.195 163.915 116.705 165.005 ;
        RECT 117.335 164.785 117.505 165.815 ;
        RECT 118.185 165.760 118.405 166.245 ;
        RECT 117.675 165.165 117.905 165.560 ;
        RECT 118.075 165.335 118.405 165.760 ;
        RECT 118.575 166.085 119.465 166.255 ;
        RECT 118.575 165.360 118.745 166.085 ;
        RECT 118.915 165.530 119.465 165.915 ;
        RECT 120.555 165.740 120.845 166.465 ;
        RECT 121.220 165.685 121.720 166.295 ;
        RECT 118.575 165.290 119.465 165.360 ;
        RECT 118.570 165.265 119.465 165.290 ;
        RECT 118.560 165.250 119.465 165.265 ;
        RECT 118.555 165.235 119.465 165.250 ;
        RECT 118.545 165.230 119.465 165.235 ;
        RECT 118.540 165.220 119.465 165.230 ;
        RECT 121.015 165.225 121.365 165.475 ;
        RECT 118.535 165.210 119.465 165.220 ;
        RECT 118.525 165.205 119.465 165.210 ;
        RECT 118.515 165.195 119.465 165.205 ;
        RECT 118.505 165.190 119.465 165.195 ;
        RECT 118.505 165.185 118.840 165.190 ;
        RECT 118.490 165.180 118.840 165.185 ;
        RECT 118.475 165.170 118.840 165.180 ;
        RECT 118.450 165.165 118.840 165.170 ;
        RECT 117.675 165.160 118.840 165.165 ;
        RECT 117.675 165.125 118.810 165.160 ;
        RECT 117.675 165.100 118.775 165.125 ;
        RECT 117.675 165.070 118.745 165.100 ;
        RECT 117.675 165.040 118.725 165.070 ;
        RECT 117.675 165.010 118.705 165.040 ;
        RECT 117.675 165.000 118.635 165.010 ;
        RECT 117.675 164.990 118.610 165.000 ;
        RECT 117.675 164.975 118.590 164.990 ;
        RECT 117.675 164.960 118.570 164.975 ;
        RECT 117.780 164.950 118.565 164.960 ;
        RECT 117.780 164.915 118.550 164.950 ;
        RECT 117.335 164.085 117.610 164.785 ;
        RECT 117.780 164.665 118.535 164.915 ;
        RECT 118.705 164.595 119.035 164.840 ;
        RECT 119.205 164.740 119.465 165.190 ;
        RECT 118.850 164.570 119.035 164.595 ;
        RECT 118.850 164.470 119.465 164.570 ;
        RECT 117.780 163.915 118.035 164.460 ;
        RECT 118.205 164.085 118.685 164.425 ;
        RECT 118.860 163.915 119.465 164.470 ;
        RECT 120.555 163.915 120.845 165.080 ;
        RECT 121.550 165.055 121.720 165.685 ;
        RECT 122.350 165.815 122.680 166.295 ;
        RECT 122.850 166.005 123.075 166.465 ;
        RECT 123.245 165.815 123.575 166.295 ;
        RECT 122.350 165.645 123.575 165.815 ;
        RECT 123.765 165.665 124.015 166.465 ;
        RECT 124.185 165.665 124.525 166.295 ;
        RECT 121.890 165.275 122.220 165.475 ;
        RECT 122.390 165.275 122.720 165.475 ;
        RECT 122.890 165.275 123.310 165.475 ;
        RECT 123.485 165.305 124.180 165.475 ;
        RECT 123.485 165.055 123.655 165.305 ;
        RECT 124.350 165.055 124.525 165.665 ;
        RECT 124.695 165.695 128.205 166.465 ;
        RECT 128.375 165.715 129.585 166.465 ;
        RECT 129.845 165.915 130.015 166.295 ;
        RECT 130.195 166.085 130.525 166.465 ;
        RECT 129.845 165.745 130.510 165.915 ;
        RECT 130.705 165.790 130.965 166.295 ;
        RECT 124.695 165.175 126.345 165.695 ;
        RECT 121.220 164.885 123.655 165.055 ;
        RECT 121.220 164.085 121.550 164.885 ;
        RECT 121.720 163.915 122.050 164.715 ;
        RECT 122.350 164.085 122.680 164.885 ;
        RECT 123.325 163.915 123.575 164.715 ;
        RECT 123.845 163.915 124.015 165.055 ;
        RECT 124.185 164.085 124.525 165.055 ;
        RECT 126.515 165.005 128.205 165.525 ;
        RECT 128.375 165.175 128.895 165.715 ;
        RECT 129.065 165.005 129.585 165.545 ;
        RECT 129.775 165.195 130.105 165.565 ;
        RECT 130.340 165.490 130.510 165.745 ;
        RECT 130.340 165.160 130.625 165.490 ;
        RECT 130.340 165.015 130.510 165.160 ;
        RECT 124.695 163.915 128.205 165.005 ;
        RECT 128.375 163.915 129.585 165.005 ;
        RECT 129.845 164.845 130.510 165.015 ;
        RECT 130.795 164.990 130.965 165.790 ;
        RECT 131.225 165.915 131.395 166.205 ;
        RECT 131.565 166.085 131.895 166.465 ;
        RECT 131.225 165.745 131.890 165.915 ;
        RECT 129.845 164.085 130.015 164.845 ;
        RECT 130.195 163.915 130.525 164.675 ;
        RECT 130.695 164.085 130.965 164.990 ;
        RECT 131.140 164.925 131.490 165.575 ;
        RECT 131.660 164.755 131.890 165.745 ;
        RECT 131.225 164.585 131.890 164.755 ;
        RECT 131.225 164.085 131.395 164.585 ;
        RECT 131.565 163.915 131.895 164.415 ;
        RECT 132.065 164.085 132.250 166.205 ;
        RECT 132.505 166.005 132.755 166.465 ;
        RECT 132.925 166.015 133.260 166.185 ;
        RECT 133.455 166.015 134.130 166.185 ;
        RECT 132.925 165.875 133.095 166.015 ;
        RECT 132.420 164.885 132.700 165.835 ;
        RECT 132.870 165.745 133.095 165.875 ;
        RECT 132.870 164.640 133.040 165.745 ;
        RECT 133.265 165.595 133.790 165.815 ;
        RECT 133.210 164.830 133.450 165.425 ;
        RECT 133.620 164.895 133.790 165.595 ;
        RECT 133.960 165.235 134.130 166.015 ;
        RECT 134.450 165.965 134.820 166.465 ;
        RECT 135.000 166.015 135.405 166.185 ;
        RECT 135.575 166.015 136.360 166.185 ;
        RECT 135.000 165.785 135.170 166.015 ;
        RECT 134.340 165.485 135.170 165.785 ;
        RECT 135.555 165.515 136.020 165.845 ;
        RECT 134.340 165.455 134.540 165.485 ;
        RECT 134.660 165.235 134.830 165.305 ;
        RECT 133.960 165.065 134.830 165.235 ;
        RECT 134.320 164.975 134.830 165.065 ;
        RECT 132.870 164.510 133.175 164.640 ;
        RECT 133.620 164.530 134.150 164.895 ;
        RECT 132.490 163.915 132.755 164.375 ;
        RECT 132.925 164.085 133.175 164.510 ;
        RECT 134.320 164.360 134.490 164.975 ;
        RECT 133.385 164.190 134.490 164.360 ;
        RECT 134.660 163.915 134.830 164.715 ;
        RECT 135.000 164.415 135.170 165.485 ;
        RECT 135.340 164.585 135.530 165.305 ;
        RECT 135.700 164.555 136.020 165.515 ;
        RECT 136.190 165.555 136.360 166.015 ;
        RECT 136.635 165.935 136.845 166.465 ;
        RECT 137.105 165.725 137.435 166.250 ;
        RECT 137.605 165.855 137.775 166.465 ;
        RECT 137.945 165.810 138.275 166.245 ;
        RECT 137.945 165.725 138.325 165.810 ;
        RECT 137.235 165.555 137.435 165.725 ;
        RECT 138.100 165.685 138.325 165.725 ;
        RECT 136.190 165.225 137.065 165.555 ;
        RECT 137.235 165.225 137.985 165.555 ;
        RECT 135.000 164.085 135.250 164.415 ;
        RECT 136.190 164.385 136.360 165.225 ;
        RECT 137.235 165.020 137.425 165.225 ;
        RECT 138.155 165.105 138.325 165.685 ;
        RECT 138.110 165.055 138.325 165.105 ;
        RECT 136.530 164.645 137.425 165.020 ;
        RECT 137.935 164.975 138.325 165.055 ;
        RECT 138.495 165.790 138.755 166.295 ;
        RECT 138.935 166.085 139.265 166.465 ;
        RECT 139.445 165.915 139.615 166.295 ;
        RECT 138.495 164.990 138.665 165.790 ;
        RECT 138.950 165.745 139.615 165.915 ;
        RECT 139.965 165.915 140.135 166.295 ;
        RECT 140.350 166.085 140.680 166.465 ;
        RECT 139.965 165.745 140.680 165.915 ;
        RECT 138.950 165.490 139.120 165.745 ;
        RECT 138.835 165.160 139.120 165.490 ;
        RECT 139.355 165.195 139.685 165.565 ;
        RECT 139.875 165.195 140.230 165.565 ;
        RECT 140.510 165.555 140.680 165.745 ;
        RECT 140.850 165.720 141.105 166.295 ;
        RECT 140.510 165.225 140.765 165.555 ;
        RECT 138.950 165.015 139.120 165.160 ;
        RECT 140.510 165.015 140.680 165.225 ;
        RECT 135.475 164.215 136.360 164.385 ;
        RECT 136.540 163.915 136.855 164.415 ;
        RECT 137.085 164.085 137.425 164.645 ;
        RECT 137.595 163.915 137.765 164.925 ;
        RECT 137.935 164.130 138.265 164.975 ;
        RECT 138.495 164.085 138.765 164.990 ;
        RECT 138.950 164.845 139.615 165.015 ;
        RECT 138.935 163.915 139.265 164.675 ;
        RECT 139.445 164.085 139.615 164.845 ;
        RECT 139.965 164.845 140.680 165.015 ;
        RECT 140.935 164.990 141.105 165.720 ;
        RECT 141.280 165.625 141.540 166.465 ;
        RECT 141.715 165.715 142.925 166.465 ;
        RECT 139.965 164.085 140.135 164.845 ;
        RECT 140.350 163.915 140.680 164.675 ;
        RECT 140.850 164.085 141.105 164.990 ;
        RECT 141.280 163.915 141.540 165.065 ;
        RECT 141.715 165.005 142.235 165.545 ;
        RECT 142.405 165.175 142.925 165.715 ;
        RECT 141.715 163.915 142.925 165.005 ;
        RECT 17.430 163.745 143.010 163.915 ;
        RECT 17.515 162.655 18.725 163.745 ;
        RECT 17.515 161.945 18.035 162.485 ;
        RECT 18.205 162.115 18.725 162.655 ;
        RECT 18.975 162.815 19.155 163.575 ;
        RECT 19.335 162.985 19.665 163.745 ;
        RECT 18.975 162.645 19.650 162.815 ;
        RECT 19.835 162.670 20.105 163.575 ;
        RECT 19.480 162.500 19.650 162.645 ;
        RECT 18.915 162.095 19.255 162.465 ;
        RECT 19.480 162.170 19.755 162.500 ;
        RECT 17.515 161.195 18.725 161.945 ;
        RECT 19.480 161.915 19.650 162.170 ;
        RECT 18.985 161.745 19.650 161.915 ;
        RECT 19.925 161.870 20.105 162.670 ;
        RECT 20.275 162.655 21.485 163.745 ;
        RECT 18.985 161.365 19.155 161.745 ;
        RECT 19.335 161.195 19.665 161.575 ;
        RECT 19.845 161.365 20.105 161.870 ;
        RECT 20.275 161.945 20.795 162.485 ;
        RECT 20.965 162.115 21.485 162.655 ;
        RECT 20.275 161.195 21.485 161.945 ;
        RECT 21.655 161.365 21.915 163.575 ;
        RECT 22.085 163.365 22.415 163.745 ;
        RECT 22.840 163.195 23.010 163.575 ;
        RECT 23.270 163.365 23.600 163.745 ;
        RECT 23.795 163.195 23.965 163.575 ;
        RECT 24.175 163.365 24.505 163.745 ;
        RECT 24.755 163.195 24.945 163.575 ;
        RECT 25.185 163.365 25.515 163.745 ;
        RECT 25.825 163.245 26.085 163.575 ;
        RECT 22.085 163.025 24.035 163.195 ;
        RECT 22.085 162.105 22.255 163.025 ;
        RECT 22.625 162.435 22.820 162.745 ;
        RECT 23.090 162.435 23.275 162.745 ;
        RECT 22.565 162.105 22.820 162.435 ;
        RECT 23.045 162.105 23.275 162.435 ;
        RECT 22.085 161.195 22.415 161.575 ;
        RECT 22.625 161.530 22.820 162.105 ;
        RECT 23.090 161.525 23.275 162.105 ;
        RECT 23.525 161.535 23.695 162.435 ;
        RECT 23.865 162.035 24.035 163.025 ;
        RECT 24.205 163.025 24.945 163.195 ;
        RECT 24.205 162.515 24.375 163.025 ;
        RECT 24.545 162.685 25.125 162.855 ;
        RECT 25.395 162.735 25.745 163.065 ;
        RECT 24.955 162.565 25.125 162.685 ;
        RECT 25.915 162.565 26.085 163.245 ;
        RECT 24.205 162.345 24.775 162.515 ;
        RECT 24.955 162.395 26.085 162.565 ;
        RECT 23.865 161.705 24.415 162.035 ;
        RECT 24.605 161.865 24.775 162.345 ;
        RECT 24.945 162.055 25.565 162.225 ;
        RECT 25.355 161.875 25.565 162.055 ;
        RECT 24.605 161.535 25.005 161.865 ;
        RECT 25.915 161.695 26.085 162.395 ;
        RECT 23.525 161.365 25.005 161.535 ;
        RECT 25.185 161.195 25.515 161.575 ;
        RECT 25.825 161.365 26.085 161.695 ;
        RECT 26.255 162.605 26.515 163.575 ;
        RECT 26.710 163.335 27.040 163.745 ;
        RECT 27.240 163.155 27.410 163.575 ;
        RECT 27.625 163.335 28.295 163.745 ;
        RECT 28.530 163.155 28.700 163.575 ;
        RECT 29.005 163.305 29.335 163.745 ;
        RECT 26.685 162.985 28.700 163.155 ;
        RECT 29.505 163.125 29.680 163.575 ;
        RECT 26.255 161.915 26.425 162.605 ;
        RECT 26.685 162.435 26.855 162.985 ;
        RECT 26.595 162.105 26.855 162.435 ;
        RECT 26.255 161.450 26.595 161.915 ;
        RECT 27.025 161.775 27.365 162.805 ;
        RECT 27.555 162.725 27.825 162.805 ;
        RECT 27.555 162.555 27.865 162.725 ;
        RECT 26.260 161.405 26.595 161.450 ;
        RECT 26.765 161.195 27.095 161.575 ;
        RECT 27.555 161.530 27.825 162.555 ;
        RECT 28.050 161.530 28.330 162.805 ;
        RECT 28.530 161.695 28.700 162.985 ;
        RECT 29.050 162.955 29.680 163.125 ;
        RECT 29.050 162.435 29.220 162.955 ;
        RECT 28.870 162.105 29.220 162.435 ;
        RECT 29.400 162.105 29.765 162.785 ;
        RECT 30.395 162.580 30.685 163.745 ;
        RECT 31.325 162.605 31.655 163.745 ;
        RECT 32.185 162.775 32.515 163.560 ;
        RECT 31.835 162.605 32.515 162.775 ;
        RECT 32.695 162.655 35.285 163.745 ;
        RECT 31.315 162.185 31.665 162.435 ;
        RECT 29.050 161.935 29.220 162.105 ;
        RECT 31.835 162.005 32.005 162.605 ;
        RECT 32.175 162.185 32.525 162.435 ;
        RECT 29.050 161.765 29.680 161.935 ;
        RECT 28.530 161.365 28.760 161.695 ;
        RECT 29.005 161.195 29.335 161.575 ;
        RECT 29.505 161.365 29.680 161.765 ;
        RECT 30.395 161.195 30.685 161.920 ;
        RECT 31.325 161.195 31.595 162.005 ;
        RECT 31.765 161.365 32.095 162.005 ;
        RECT 32.265 161.195 32.505 162.005 ;
        RECT 32.695 161.965 33.905 162.485 ;
        RECT 34.075 162.135 35.285 162.655 ;
        RECT 35.495 162.795 35.785 163.565 ;
        RECT 36.355 163.205 36.615 163.565 ;
        RECT 36.785 163.375 37.115 163.745 ;
        RECT 37.285 163.205 37.545 163.565 ;
        RECT 36.355 162.975 37.545 163.205 ;
        RECT 37.735 163.025 38.065 163.745 ;
        RECT 38.235 162.795 38.500 163.565 ;
        RECT 35.495 162.615 37.990 162.795 ;
        RECT 35.465 162.105 35.735 162.435 ;
        RECT 35.915 162.105 36.350 162.435 ;
        RECT 36.530 162.105 37.105 162.435 ;
        RECT 37.285 162.105 37.565 162.435 ;
        RECT 32.695 161.195 35.285 161.965 ;
        RECT 37.765 161.925 37.990 162.615 ;
        RECT 35.505 161.735 37.990 161.925 ;
        RECT 35.505 161.375 35.730 161.735 ;
        RECT 35.910 161.195 36.240 161.565 ;
        RECT 36.420 161.375 36.675 161.735 ;
        RECT 37.240 161.195 37.985 161.565 ;
        RECT 38.165 161.375 38.500 162.795 ;
        RECT 38.675 162.670 39.015 163.745 ;
        RECT 39.200 163.405 41.250 163.525 ;
        RECT 39.195 163.235 41.250 163.405 ;
        RECT 39.185 162.435 39.425 163.030 ;
        RECT 39.620 162.895 41.250 163.065 ;
        RECT 41.420 162.945 41.700 163.745 ;
        RECT 39.620 162.605 39.940 162.895 ;
        RECT 41.080 162.775 41.250 162.895 ;
        RECT 38.675 161.865 39.015 162.435 ;
        RECT 39.185 162.105 39.840 162.435 ;
        RECT 40.110 162.105 40.850 162.725 ;
        RECT 41.080 162.605 41.740 162.775 ;
        RECT 41.910 162.605 42.185 163.575 ;
        RECT 41.570 162.435 41.740 162.605 ;
        RECT 41.020 162.105 41.400 162.435 ;
        RECT 41.570 162.105 41.845 162.435 ;
        RECT 38.675 161.195 39.015 161.695 ;
        RECT 39.185 161.415 39.430 162.105 ;
        RECT 41.570 161.935 41.740 162.105 ;
        RECT 40.155 161.765 41.740 161.935 ;
        RECT 42.015 161.870 42.185 162.605 ;
        RECT 39.625 161.195 39.955 161.695 ;
        RECT 40.155 161.415 40.325 161.765 ;
        RECT 40.500 161.195 40.830 161.595 ;
        RECT 41.000 161.415 41.170 161.765 ;
        RECT 41.340 161.195 41.720 161.595 ;
        RECT 41.910 161.525 42.185 161.870 ;
        RECT 43.310 162.955 43.845 163.575 ;
        RECT 43.310 161.935 43.625 162.955 ;
        RECT 44.015 162.945 44.345 163.745 ;
        RECT 44.830 162.775 45.220 162.950 ;
        RECT 43.795 162.605 45.220 162.775 ;
        RECT 45.575 162.655 49.085 163.745 ;
        RECT 43.795 162.105 43.965 162.605 ;
        RECT 43.310 161.365 43.925 161.935 ;
        RECT 44.215 161.875 44.480 162.435 ;
        RECT 44.650 161.705 44.820 162.605 ;
        RECT 44.990 161.875 45.345 162.435 ;
        RECT 45.575 161.965 47.225 162.485 ;
        RECT 47.395 162.135 49.085 162.655 ;
        RECT 44.095 161.195 44.310 161.705 ;
        RECT 44.540 161.375 44.820 161.705 ;
        RECT 45.000 161.195 45.240 161.705 ;
        RECT 45.575 161.195 49.085 161.965 ;
        RECT 49.725 161.375 49.985 163.565 ;
        RECT 50.155 163.015 50.495 163.745 ;
        RECT 50.675 162.835 50.945 163.565 ;
        RECT 50.175 162.615 50.945 162.835 ;
        RECT 51.125 162.855 51.355 163.565 ;
        RECT 51.525 163.035 51.855 163.745 ;
        RECT 52.025 162.855 52.285 163.565 ;
        RECT 53.235 163.105 53.565 163.535 ;
        RECT 51.125 162.615 52.285 162.855 ;
        RECT 53.110 162.935 53.565 163.105 ;
        RECT 53.745 163.105 53.995 163.525 ;
        RECT 54.225 163.275 54.555 163.745 ;
        RECT 54.785 163.105 55.035 163.525 ;
        RECT 53.745 162.935 55.035 163.105 ;
        RECT 50.175 161.945 50.465 162.615 ;
        RECT 50.645 162.125 51.110 162.435 ;
        RECT 51.290 162.125 51.815 162.435 ;
        RECT 50.175 161.745 51.405 161.945 ;
        RECT 50.245 161.195 50.915 161.565 ;
        RECT 51.095 161.375 51.405 161.745 ;
        RECT 51.585 161.485 51.815 162.125 ;
        RECT 51.995 162.105 52.295 162.435 ;
        RECT 53.110 161.935 53.280 162.935 ;
        RECT 53.450 162.105 53.695 162.765 ;
        RECT 53.910 162.105 54.175 162.765 ;
        RECT 54.370 162.105 54.655 162.765 ;
        RECT 54.830 162.435 55.045 162.765 ;
        RECT 55.225 162.605 55.475 163.745 ;
        RECT 55.645 162.685 55.975 163.535 ;
        RECT 54.830 162.105 55.135 162.435 ;
        RECT 55.305 162.105 55.615 162.435 ;
        RECT 55.305 161.935 55.475 162.105 ;
        RECT 51.995 161.195 52.285 161.925 ;
        RECT 53.110 161.765 55.475 161.935 ;
        RECT 55.785 161.920 55.975 162.685 ;
        RECT 56.155 162.580 56.445 163.745 ;
        RECT 56.675 162.685 57.005 163.530 ;
        RECT 57.175 162.735 57.345 163.745 ;
        RECT 57.515 163.015 57.855 163.575 ;
        RECT 58.085 163.245 58.400 163.745 ;
        RECT 58.580 163.275 59.465 163.445 ;
        RECT 56.615 162.605 57.005 162.685 ;
        RECT 57.515 162.640 58.410 163.015 ;
        RECT 56.615 162.555 56.830 162.605 ;
        RECT 56.615 161.975 56.785 162.555 ;
        RECT 57.515 162.435 57.705 162.640 ;
        RECT 58.580 162.435 58.750 163.275 ;
        RECT 59.690 163.245 59.940 163.575 ;
        RECT 56.955 162.105 57.705 162.435 ;
        RECT 57.875 162.105 58.750 162.435 ;
        RECT 56.615 161.935 56.840 161.975 ;
        RECT 57.505 161.935 57.705 162.105 ;
        RECT 53.265 161.195 53.595 161.595 ;
        RECT 53.765 161.425 54.095 161.765 ;
        RECT 55.145 161.195 55.475 161.595 ;
        RECT 55.645 161.410 55.975 161.920 ;
        RECT 56.155 161.195 56.445 161.920 ;
        RECT 56.615 161.850 56.995 161.935 ;
        RECT 56.665 161.415 56.995 161.850 ;
        RECT 57.165 161.195 57.335 161.805 ;
        RECT 57.505 161.410 57.835 161.935 ;
        RECT 58.095 161.195 58.305 161.725 ;
        RECT 58.580 161.645 58.750 162.105 ;
        RECT 58.920 162.145 59.240 163.105 ;
        RECT 59.410 162.355 59.600 163.075 ;
        RECT 59.770 162.175 59.940 163.245 ;
        RECT 60.110 162.945 60.280 163.745 ;
        RECT 60.450 163.300 61.555 163.470 ;
        RECT 60.450 162.685 60.620 163.300 ;
        RECT 61.765 163.150 62.015 163.575 ;
        RECT 62.185 163.285 62.450 163.745 ;
        RECT 60.790 162.765 61.320 163.130 ;
        RECT 61.765 163.020 62.070 163.150 ;
        RECT 60.110 162.595 60.620 162.685 ;
        RECT 60.110 162.425 60.980 162.595 ;
        RECT 60.110 162.355 60.280 162.425 ;
        RECT 60.400 162.175 60.600 162.205 ;
        RECT 58.920 161.815 59.385 162.145 ;
        RECT 59.770 161.875 60.600 162.175 ;
        RECT 59.770 161.645 59.940 161.875 ;
        RECT 58.580 161.475 59.365 161.645 ;
        RECT 59.535 161.475 59.940 161.645 ;
        RECT 60.120 161.195 60.490 161.695 ;
        RECT 60.810 161.645 60.980 162.425 ;
        RECT 61.150 162.065 61.320 162.765 ;
        RECT 61.490 162.235 61.730 162.830 ;
        RECT 61.150 161.845 61.675 162.065 ;
        RECT 61.900 161.915 62.070 163.020 ;
        RECT 61.845 161.785 62.070 161.915 ;
        RECT 62.240 161.825 62.520 162.775 ;
        RECT 61.845 161.645 62.015 161.785 ;
        RECT 60.810 161.475 61.485 161.645 ;
        RECT 61.680 161.475 62.015 161.645 ;
        RECT 62.185 161.195 62.435 161.655 ;
        RECT 62.690 161.455 62.875 163.575 ;
        RECT 63.045 163.245 63.375 163.745 ;
        RECT 63.545 163.075 63.715 163.575 ;
        RECT 63.975 163.310 69.320 163.745 ;
        RECT 63.050 162.905 63.715 163.075 ;
        RECT 63.050 161.915 63.280 162.905 ;
        RECT 63.450 162.085 63.800 162.735 ;
        RECT 63.050 161.745 63.715 161.915 ;
        RECT 63.045 161.195 63.375 161.575 ;
        RECT 63.545 161.455 63.715 161.745 ;
        RECT 65.560 161.740 65.900 162.570 ;
        RECT 67.380 162.060 67.730 163.310 ;
        RECT 69.495 163.190 70.100 163.745 ;
        RECT 70.275 163.235 70.755 163.575 ;
        RECT 70.925 163.200 71.180 163.745 ;
        RECT 69.495 163.090 70.110 163.190 ;
        RECT 69.925 163.065 70.110 163.090 ;
        RECT 69.495 162.470 69.755 162.920 ;
        RECT 69.925 162.820 70.255 163.065 ;
        RECT 70.425 162.745 71.180 162.995 ;
        RECT 71.350 162.875 71.625 163.575 ;
        RECT 72.255 163.190 72.860 163.745 ;
        RECT 73.035 163.235 73.515 163.575 ;
        RECT 73.685 163.200 73.940 163.745 ;
        RECT 72.255 163.090 72.870 163.190 ;
        RECT 72.685 163.065 72.870 163.090 ;
        RECT 70.410 162.710 71.180 162.745 ;
        RECT 70.395 162.700 71.180 162.710 ;
        RECT 70.390 162.685 71.285 162.700 ;
        RECT 70.370 162.670 71.285 162.685 ;
        RECT 70.350 162.660 71.285 162.670 ;
        RECT 70.325 162.650 71.285 162.660 ;
        RECT 70.255 162.620 71.285 162.650 ;
        RECT 70.235 162.590 71.285 162.620 ;
        RECT 70.215 162.560 71.285 162.590 ;
        RECT 70.185 162.535 71.285 162.560 ;
        RECT 70.150 162.500 71.285 162.535 ;
        RECT 70.120 162.495 71.285 162.500 ;
        RECT 70.120 162.490 70.510 162.495 ;
        RECT 70.120 162.480 70.485 162.490 ;
        RECT 70.120 162.475 70.470 162.480 ;
        RECT 70.120 162.470 70.455 162.475 ;
        RECT 69.495 162.465 70.455 162.470 ;
        RECT 69.495 162.455 70.445 162.465 ;
        RECT 69.495 162.450 70.435 162.455 ;
        RECT 69.495 162.440 70.425 162.450 ;
        RECT 69.495 162.430 70.420 162.440 ;
        RECT 69.495 162.425 70.415 162.430 ;
        RECT 69.495 162.410 70.405 162.425 ;
        RECT 69.495 162.395 70.400 162.410 ;
        RECT 69.495 162.370 70.390 162.395 ;
        RECT 69.495 162.300 70.385 162.370 ;
        RECT 69.495 161.745 70.045 162.130 ;
        RECT 63.975 161.195 69.320 161.740 ;
        RECT 70.215 161.575 70.385 162.300 ;
        RECT 69.495 161.405 70.385 161.575 ;
        RECT 70.555 161.900 70.885 162.325 ;
        RECT 71.055 162.100 71.285 162.495 ;
        RECT 70.555 161.415 70.775 161.900 ;
        RECT 71.455 161.845 71.625 162.875 ;
        RECT 72.255 162.470 72.515 162.920 ;
        RECT 72.685 162.820 73.015 163.065 ;
        RECT 73.185 162.745 73.940 162.995 ;
        RECT 74.110 162.875 74.385 163.575 ;
        RECT 73.170 162.710 73.940 162.745 ;
        RECT 73.155 162.700 73.940 162.710 ;
        RECT 73.150 162.685 74.045 162.700 ;
        RECT 73.130 162.670 74.045 162.685 ;
        RECT 73.110 162.660 74.045 162.670 ;
        RECT 73.085 162.650 74.045 162.660 ;
        RECT 73.015 162.620 74.045 162.650 ;
        RECT 72.995 162.590 74.045 162.620 ;
        RECT 72.975 162.560 74.045 162.590 ;
        RECT 72.945 162.535 74.045 162.560 ;
        RECT 72.910 162.500 74.045 162.535 ;
        RECT 72.880 162.495 74.045 162.500 ;
        RECT 72.880 162.490 73.270 162.495 ;
        RECT 72.880 162.480 73.245 162.490 ;
        RECT 72.880 162.475 73.230 162.480 ;
        RECT 72.880 162.470 73.215 162.475 ;
        RECT 72.255 162.465 73.215 162.470 ;
        RECT 72.255 162.455 73.205 162.465 ;
        RECT 72.255 162.450 73.195 162.455 ;
        RECT 72.255 162.440 73.185 162.450 ;
        RECT 72.255 162.430 73.180 162.440 ;
        RECT 72.255 162.425 73.175 162.430 ;
        RECT 72.255 162.410 73.165 162.425 ;
        RECT 72.255 162.395 73.160 162.410 ;
        RECT 72.255 162.370 73.150 162.395 ;
        RECT 72.255 162.300 73.145 162.370 ;
        RECT 70.945 161.195 71.195 161.735 ;
        RECT 71.365 161.365 71.625 161.845 ;
        RECT 72.255 161.745 72.805 162.130 ;
        RECT 72.975 161.575 73.145 162.300 ;
        RECT 72.255 161.405 73.145 161.575 ;
        RECT 73.315 161.900 73.645 162.325 ;
        RECT 73.815 162.100 74.045 162.495 ;
        RECT 73.315 161.415 73.535 161.900 ;
        RECT 74.215 161.845 74.385 162.875 ;
        RECT 73.705 161.195 73.955 161.735 ;
        RECT 74.125 161.365 74.385 161.845 ;
        RECT 74.555 162.605 74.895 163.575 ;
        RECT 75.065 162.605 75.235 163.745 ;
        RECT 75.505 162.945 75.755 163.745 ;
        RECT 76.400 162.775 76.730 163.575 ;
        RECT 77.030 162.945 77.360 163.745 ;
        RECT 77.530 162.775 77.860 163.575 ;
        RECT 75.425 162.605 77.860 162.775 ;
        RECT 78.235 162.605 78.510 163.575 ;
        RECT 78.720 162.945 79.000 163.745 ;
        RECT 79.170 163.405 81.220 163.525 ;
        RECT 79.170 163.235 81.225 163.405 ;
        RECT 79.170 162.895 80.800 163.065 ;
        RECT 79.170 162.775 79.340 162.895 ;
        RECT 78.680 162.605 79.340 162.775 ;
        RECT 74.555 161.995 74.730 162.605 ;
        RECT 75.425 162.355 75.595 162.605 ;
        RECT 74.900 162.185 75.595 162.355 ;
        RECT 75.770 162.185 76.190 162.385 ;
        RECT 76.360 162.185 76.690 162.385 ;
        RECT 76.860 162.185 77.190 162.385 ;
        RECT 74.555 161.365 74.895 161.995 ;
        RECT 75.065 161.195 75.315 161.995 ;
        RECT 75.505 161.845 76.730 162.015 ;
        RECT 75.505 161.365 75.835 161.845 ;
        RECT 76.005 161.195 76.230 161.655 ;
        RECT 76.400 161.365 76.730 161.845 ;
        RECT 77.360 161.975 77.530 162.605 ;
        RECT 77.715 162.185 78.065 162.435 ;
        RECT 77.360 161.365 77.860 161.975 ;
        RECT 78.235 161.870 78.405 162.605 ;
        RECT 78.680 162.435 78.850 162.605 ;
        RECT 78.575 162.105 78.850 162.435 ;
        RECT 79.020 162.105 79.400 162.435 ;
        RECT 79.570 162.105 80.310 162.725 ;
        RECT 80.480 162.605 80.800 162.895 ;
        RECT 80.995 162.435 81.235 163.030 ;
        RECT 81.405 162.670 81.745 163.745 ;
        RECT 81.915 162.580 82.205 163.745 ;
        RECT 83.410 163.115 83.695 163.575 ;
        RECT 83.865 163.285 84.135 163.745 ;
        RECT 83.410 162.895 84.365 163.115 ;
        RECT 80.580 162.105 81.235 162.435 ;
        RECT 78.680 161.935 78.850 162.105 ;
        RECT 78.235 161.525 78.510 161.870 ;
        RECT 78.680 161.765 80.265 161.935 ;
        RECT 78.700 161.195 79.080 161.595 ;
        RECT 79.250 161.415 79.420 161.765 ;
        RECT 79.590 161.195 79.920 161.595 ;
        RECT 80.095 161.415 80.265 161.765 ;
        RECT 80.465 161.195 80.795 161.695 ;
        RECT 80.990 161.415 81.235 162.105 ;
        RECT 81.405 161.865 81.745 162.435 ;
        RECT 83.295 162.165 83.985 162.725 ;
        RECT 84.155 161.995 84.365 162.895 ;
        RECT 81.405 161.195 81.745 161.695 ;
        RECT 81.915 161.195 82.205 161.920 ;
        RECT 83.410 161.825 84.365 161.995 ;
        RECT 84.535 162.725 84.935 163.575 ;
        RECT 85.125 163.115 85.405 163.575 ;
        RECT 85.925 163.285 86.250 163.745 ;
        RECT 85.125 162.895 86.250 163.115 ;
        RECT 84.535 162.165 85.630 162.725 ;
        RECT 85.800 162.435 86.250 162.895 ;
        RECT 86.420 162.605 86.805 163.575 ;
        RECT 83.410 161.365 83.695 161.825 ;
        RECT 83.865 161.195 84.135 161.655 ;
        RECT 84.535 161.365 84.935 162.165 ;
        RECT 85.800 162.105 86.355 162.435 ;
        RECT 85.800 161.995 86.250 162.105 ;
        RECT 85.125 161.825 86.250 161.995 ;
        RECT 86.525 161.935 86.805 162.605 ;
        RECT 86.975 162.985 87.490 163.395 ;
        RECT 87.725 162.985 87.895 163.745 ;
        RECT 88.065 163.405 90.095 163.575 ;
        RECT 86.975 162.175 87.315 162.985 ;
        RECT 88.065 162.740 88.235 163.405 ;
        RECT 88.630 163.065 89.755 163.235 ;
        RECT 87.485 162.550 88.235 162.740 ;
        RECT 88.405 162.725 89.415 162.895 ;
        RECT 86.975 162.005 88.205 162.175 ;
        RECT 85.125 161.365 85.405 161.825 ;
        RECT 85.925 161.195 86.250 161.655 ;
        RECT 86.420 161.365 86.805 161.935 ;
        RECT 87.250 161.400 87.495 162.005 ;
        RECT 87.715 161.195 88.225 161.730 ;
        RECT 88.405 161.365 88.595 162.725 ;
        RECT 88.765 162.045 89.040 162.525 ;
        RECT 88.765 161.875 89.045 162.045 ;
        RECT 89.245 161.925 89.415 162.725 ;
        RECT 89.585 161.935 89.755 163.065 ;
        RECT 89.925 162.435 90.095 163.405 ;
        RECT 90.265 162.605 90.435 163.745 ;
        RECT 90.605 162.605 90.940 163.575 ;
        RECT 91.230 163.115 91.515 163.575 ;
        RECT 91.685 163.285 91.955 163.745 ;
        RECT 91.230 162.895 92.185 163.115 ;
        RECT 89.925 162.105 90.120 162.435 ;
        RECT 90.345 162.105 90.600 162.435 ;
        RECT 90.345 161.935 90.515 162.105 ;
        RECT 90.770 161.935 90.940 162.605 ;
        RECT 91.115 162.165 91.805 162.725 ;
        RECT 91.975 161.995 92.185 162.895 ;
        RECT 88.765 161.365 89.040 161.875 ;
        RECT 89.585 161.765 90.515 161.935 ;
        RECT 89.585 161.730 89.760 161.765 ;
        RECT 89.230 161.365 89.760 161.730 ;
        RECT 90.185 161.195 90.515 161.595 ;
        RECT 90.685 161.365 90.940 161.935 ;
        RECT 91.230 161.825 92.185 161.995 ;
        RECT 92.355 162.725 92.755 163.575 ;
        RECT 92.945 163.115 93.225 163.575 ;
        RECT 93.745 163.285 94.070 163.745 ;
        RECT 92.945 162.895 94.070 163.115 ;
        RECT 92.355 162.165 93.450 162.725 ;
        RECT 93.620 162.435 94.070 162.895 ;
        RECT 94.240 162.605 94.625 163.575 ;
        RECT 91.230 161.365 91.515 161.825 ;
        RECT 91.685 161.195 91.955 161.655 ;
        RECT 92.355 161.365 92.755 162.165 ;
        RECT 93.620 162.105 94.175 162.435 ;
        RECT 93.620 161.995 94.070 162.105 ;
        RECT 92.945 161.825 94.070 161.995 ;
        RECT 94.345 161.935 94.625 162.605 ;
        RECT 92.945 161.365 93.225 161.825 ;
        RECT 93.745 161.195 94.070 161.655 ;
        RECT 94.240 161.365 94.625 161.935 ;
        RECT 95.260 162.605 95.595 163.575 ;
        RECT 95.765 162.605 95.935 163.745 ;
        RECT 96.105 163.405 98.135 163.575 ;
        RECT 95.260 161.935 95.430 162.605 ;
        RECT 96.105 162.435 96.275 163.405 ;
        RECT 95.600 162.105 95.855 162.435 ;
        RECT 96.080 162.105 96.275 162.435 ;
        RECT 96.445 163.065 97.570 163.235 ;
        RECT 95.685 161.935 95.855 162.105 ;
        RECT 96.445 161.935 96.615 163.065 ;
        RECT 95.260 161.365 95.515 161.935 ;
        RECT 95.685 161.765 96.615 161.935 ;
        RECT 96.785 162.725 97.795 162.895 ;
        RECT 96.785 161.925 96.955 162.725 ;
        RECT 96.440 161.730 96.615 161.765 ;
        RECT 95.685 161.195 96.015 161.595 ;
        RECT 96.440 161.365 96.970 161.730 ;
        RECT 97.160 161.705 97.435 162.525 ;
        RECT 97.155 161.535 97.435 161.705 ;
        RECT 97.160 161.365 97.435 161.535 ;
        RECT 97.605 161.365 97.795 162.725 ;
        RECT 97.965 162.740 98.135 163.405 ;
        RECT 98.305 162.985 98.475 163.745 ;
        RECT 98.710 162.985 99.225 163.395 ;
        RECT 97.965 162.550 98.715 162.740 ;
        RECT 98.885 162.175 99.225 162.985 ;
        RECT 99.395 162.655 100.605 163.745 ;
        RECT 100.890 163.115 101.175 163.575 ;
        RECT 101.345 163.285 101.615 163.745 ;
        RECT 100.890 162.895 101.845 163.115 ;
        RECT 97.995 162.005 99.225 162.175 ;
        RECT 97.975 161.195 98.485 161.730 ;
        RECT 98.705 161.400 98.950 162.005 ;
        RECT 99.395 161.945 99.915 162.485 ;
        RECT 100.085 162.115 100.605 162.655 ;
        RECT 100.775 162.165 101.465 162.725 ;
        RECT 101.635 161.995 101.845 162.895 ;
        RECT 99.395 161.195 100.605 161.945 ;
        RECT 100.890 161.825 101.845 161.995 ;
        RECT 102.015 162.725 102.415 163.575 ;
        RECT 102.605 163.115 102.885 163.575 ;
        RECT 103.405 163.285 103.730 163.745 ;
        RECT 102.605 162.895 103.730 163.115 ;
        RECT 102.015 162.165 103.110 162.725 ;
        RECT 103.280 162.435 103.730 162.895 ;
        RECT 103.900 162.605 104.285 163.575 ;
        RECT 104.455 162.655 107.045 163.745 ;
        RECT 100.890 161.365 101.175 161.825 ;
        RECT 101.345 161.195 101.615 161.655 ;
        RECT 102.015 161.365 102.415 162.165 ;
        RECT 103.280 162.105 103.835 162.435 ;
        RECT 103.280 161.995 103.730 162.105 ;
        RECT 102.605 161.825 103.730 161.995 ;
        RECT 104.005 161.935 104.285 162.605 ;
        RECT 102.605 161.365 102.885 161.825 ;
        RECT 103.405 161.195 103.730 161.655 ;
        RECT 103.900 161.365 104.285 161.935 ;
        RECT 104.455 161.965 105.665 162.485 ;
        RECT 105.835 162.135 107.045 162.655 ;
        RECT 107.675 162.580 107.965 163.745 ;
        RECT 108.135 163.310 113.480 163.745 ;
        RECT 104.455 161.195 107.045 161.965 ;
        RECT 107.675 161.195 107.965 161.920 ;
        RECT 109.720 161.740 110.060 162.570 ;
        RECT 111.540 162.060 111.890 163.310 ;
        RECT 113.655 162.655 117.165 163.745 ;
        RECT 117.995 163.075 118.275 163.745 ;
        RECT 118.445 162.855 118.745 163.405 ;
        RECT 118.945 163.025 119.275 163.745 ;
        RECT 119.465 163.025 119.925 163.575 ;
        RECT 113.655 161.965 115.305 162.485 ;
        RECT 115.475 162.135 117.165 162.655 ;
        RECT 117.810 162.435 118.075 162.795 ;
        RECT 118.445 162.685 119.385 162.855 ;
        RECT 119.215 162.435 119.385 162.685 ;
        RECT 117.810 162.185 118.485 162.435 ;
        RECT 118.705 162.185 119.045 162.435 ;
        RECT 119.215 162.105 119.505 162.435 ;
        RECT 119.215 162.015 119.385 162.105 ;
        RECT 108.135 161.195 113.480 161.740 ;
        RECT 113.655 161.195 117.165 161.965 ;
        RECT 117.995 161.825 119.385 162.015 ;
        RECT 117.995 161.465 118.325 161.825 ;
        RECT 119.675 161.655 119.925 163.025 ;
        RECT 118.945 161.195 119.195 161.655 ;
        RECT 119.365 161.365 119.925 161.655 ;
        RECT 120.095 162.635 120.355 163.575 ;
        RECT 120.525 163.345 120.855 163.745 ;
        RECT 122.000 163.480 122.255 163.575 ;
        RECT 121.115 163.310 122.255 163.480 ;
        RECT 122.425 163.365 122.755 163.535 ;
        RECT 121.115 163.085 121.285 163.310 ;
        RECT 120.525 162.915 121.285 163.085 ;
        RECT 122.000 163.175 122.255 163.310 ;
        RECT 120.095 161.920 120.270 162.635 ;
        RECT 120.525 162.435 120.695 162.915 ;
        RECT 121.550 162.825 121.720 163.015 ;
        RECT 122.000 163.005 122.410 163.175 ;
        RECT 120.440 162.105 120.695 162.435 ;
        RECT 120.920 162.105 121.250 162.725 ;
        RECT 121.550 162.655 122.070 162.825 ;
        RECT 121.420 162.105 121.710 162.485 ;
        RECT 121.900 161.935 122.070 162.655 ;
        RECT 120.095 161.365 120.355 161.920 ;
        RECT 121.190 161.765 122.070 161.935 ;
        RECT 122.240 161.980 122.410 163.005 ;
        RECT 122.585 163.115 122.755 163.365 ;
        RECT 122.925 163.285 123.175 163.745 ;
        RECT 123.345 163.115 123.525 163.575 ;
        RECT 122.585 162.945 123.525 163.115 ;
        RECT 123.980 162.775 124.310 163.575 ;
        RECT 124.480 162.945 124.810 163.745 ;
        RECT 125.110 162.775 125.440 163.575 ;
        RECT 126.085 162.945 126.335 163.745 ;
        RECT 122.610 162.465 123.090 162.765 ;
        RECT 122.240 161.810 122.590 161.980 ;
        RECT 122.830 161.875 123.090 162.465 ;
        RECT 123.290 161.875 123.550 162.765 ;
        RECT 123.980 162.605 126.415 162.775 ;
        RECT 126.605 162.605 126.775 163.745 ;
        RECT 126.945 162.605 127.285 163.575 ;
        RECT 123.775 162.185 124.125 162.435 ;
        RECT 124.310 161.975 124.480 162.605 ;
        RECT 124.650 162.185 124.980 162.385 ;
        RECT 125.150 162.185 125.480 162.385 ;
        RECT 125.650 162.185 126.070 162.385 ;
        RECT 126.245 162.355 126.415 162.605 ;
        RECT 126.245 162.185 126.940 162.355 ;
        RECT 120.525 161.195 120.955 161.640 ;
        RECT 121.190 161.365 121.360 161.765 ;
        RECT 121.530 161.195 122.250 161.595 ;
        RECT 122.420 161.365 122.590 161.810 ;
        RECT 123.165 161.195 123.565 161.705 ;
        RECT 123.980 161.365 124.480 161.975 ;
        RECT 125.110 161.845 126.335 162.015 ;
        RECT 127.110 161.995 127.285 162.605 ;
        RECT 127.460 163.355 127.795 163.575 ;
        RECT 128.800 163.365 129.155 163.745 ;
        RECT 127.460 162.735 127.715 163.355 ;
        RECT 127.965 163.195 128.195 163.235 ;
        RECT 129.325 163.195 129.575 163.575 ;
        RECT 127.965 162.995 129.575 163.195 ;
        RECT 127.965 162.905 128.150 162.995 ;
        RECT 128.740 162.985 129.575 162.995 ;
        RECT 129.825 162.965 130.075 163.745 ;
        RECT 130.245 162.895 130.505 163.575 ;
        RECT 128.305 162.795 128.635 162.825 ;
        RECT 128.305 162.735 130.105 162.795 ;
        RECT 127.460 162.625 130.165 162.735 ;
        RECT 127.460 162.565 128.635 162.625 ;
        RECT 129.965 162.590 130.165 162.625 ;
        RECT 127.455 162.185 127.945 162.385 ;
        RECT 128.135 162.185 128.610 162.395 ;
        RECT 125.110 161.365 125.440 161.845 ;
        RECT 125.610 161.195 125.835 161.655 ;
        RECT 126.005 161.365 126.335 161.845 ;
        RECT 126.525 161.195 126.775 161.995 ;
        RECT 126.945 161.365 127.285 161.995 ;
        RECT 127.460 161.195 127.915 161.960 ;
        RECT 128.390 161.785 128.610 162.185 ;
        RECT 128.855 162.185 129.185 162.395 ;
        RECT 128.855 161.785 129.065 162.185 ;
        RECT 129.355 162.150 129.765 162.455 ;
        RECT 129.995 162.015 130.165 162.590 ;
        RECT 129.895 161.895 130.165 162.015 ;
        RECT 129.320 161.850 130.165 161.895 ;
        RECT 129.320 161.725 130.075 161.850 ;
        RECT 129.320 161.575 129.490 161.725 ;
        RECT 130.335 161.695 130.505 162.895 ;
        RECT 130.675 162.655 133.265 163.745 ;
        RECT 128.190 161.365 129.490 161.575 ;
        RECT 129.745 161.195 130.075 161.555 ;
        RECT 130.245 161.365 130.505 161.695 ;
        RECT 130.675 161.965 131.885 162.485 ;
        RECT 132.055 162.135 133.265 162.655 ;
        RECT 133.435 162.580 133.725 163.745 ;
        RECT 133.900 162.605 134.235 163.575 ;
        RECT 134.405 162.605 134.575 163.745 ;
        RECT 134.745 163.405 136.775 163.575 ;
        RECT 130.675 161.195 133.265 161.965 ;
        RECT 133.900 161.935 134.070 162.605 ;
        RECT 134.745 162.435 134.915 163.405 ;
        RECT 134.240 162.105 134.495 162.435 ;
        RECT 134.720 162.105 134.915 162.435 ;
        RECT 135.085 163.065 136.210 163.235 ;
        RECT 134.325 161.935 134.495 162.105 ;
        RECT 135.085 161.935 135.255 163.065 ;
        RECT 133.435 161.195 133.725 161.920 ;
        RECT 133.900 161.365 134.155 161.935 ;
        RECT 134.325 161.765 135.255 161.935 ;
        RECT 135.425 162.725 136.435 162.895 ;
        RECT 135.425 161.925 135.595 162.725 ;
        RECT 135.800 162.045 136.075 162.525 ;
        RECT 135.795 161.875 136.075 162.045 ;
        RECT 135.080 161.730 135.255 161.765 ;
        RECT 134.325 161.195 134.655 161.595 ;
        RECT 135.080 161.365 135.610 161.730 ;
        RECT 135.800 161.365 136.075 161.875 ;
        RECT 136.245 161.365 136.435 162.725 ;
        RECT 136.605 162.740 136.775 163.405 ;
        RECT 136.945 162.985 137.115 163.745 ;
        RECT 137.350 162.985 137.865 163.395 ;
        RECT 136.605 162.550 137.355 162.740 ;
        RECT 137.525 162.175 137.865 162.985 ;
        RECT 136.635 162.005 137.865 162.175 ;
        RECT 138.035 162.605 138.420 163.575 ;
        RECT 138.590 163.285 138.915 163.745 ;
        RECT 139.435 163.115 139.715 163.575 ;
        RECT 138.590 162.895 139.715 163.115 ;
        RECT 136.615 161.195 137.125 161.730 ;
        RECT 137.345 161.400 137.590 162.005 ;
        RECT 138.035 161.935 138.315 162.605 ;
        RECT 138.590 162.435 139.040 162.895 ;
        RECT 139.905 162.725 140.305 163.575 ;
        RECT 140.705 163.285 140.975 163.745 ;
        RECT 141.145 163.115 141.430 163.575 ;
        RECT 138.485 162.105 139.040 162.435 ;
        RECT 139.210 162.165 140.305 162.725 ;
        RECT 138.590 161.995 139.040 162.105 ;
        RECT 138.035 161.365 138.420 161.935 ;
        RECT 138.590 161.825 139.715 161.995 ;
        RECT 138.590 161.195 138.915 161.655 ;
        RECT 139.435 161.365 139.715 161.825 ;
        RECT 139.905 161.365 140.305 162.165 ;
        RECT 140.475 162.895 141.430 163.115 ;
        RECT 140.475 161.995 140.685 162.895 ;
        RECT 140.855 162.165 141.545 162.725 ;
        RECT 141.715 162.655 142.925 163.745 ;
        RECT 141.715 162.115 142.235 162.655 ;
        RECT 140.475 161.825 141.430 161.995 ;
        RECT 142.405 161.945 142.925 162.485 ;
        RECT 140.705 161.195 140.975 161.655 ;
        RECT 141.145 161.365 141.430 161.825 ;
        RECT 141.715 161.195 142.925 161.945 ;
        RECT 17.430 161.025 143.010 161.195 ;
        RECT 17.515 160.275 18.725 161.025 ;
        RECT 17.515 159.735 18.035 160.275 ;
        RECT 18.895 160.255 20.565 161.025 ;
        RECT 21.245 160.370 21.575 160.805 ;
        RECT 21.745 160.415 21.915 161.025 ;
        RECT 21.195 160.285 21.575 160.370 ;
        RECT 22.085 160.285 22.415 160.810 ;
        RECT 22.675 160.495 22.885 161.025 ;
        RECT 23.160 160.575 23.945 160.745 ;
        RECT 24.115 160.575 24.520 160.745 ;
        RECT 18.205 159.565 18.725 160.105 ;
        RECT 18.895 159.735 19.645 160.255 ;
        RECT 21.195 160.245 21.420 160.285 ;
        RECT 19.815 159.565 20.565 160.085 ;
        RECT 17.515 158.475 18.725 159.565 ;
        RECT 18.895 158.475 20.565 159.565 ;
        RECT 21.195 159.665 21.365 160.245 ;
        RECT 22.085 160.115 22.285 160.285 ;
        RECT 23.160 160.115 23.330 160.575 ;
        RECT 21.535 159.785 22.285 160.115 ;
        RECT 22.455 159.785 23.330 160.115 ;
        RECT 21.195 159.615 21.410 159.665 ;
        RECT 21.195 159.535 21.585 159.615 ;
        RECT 21.255 158.690 21.585 159.535 ;
        RECT 22.095 159.580 22.285 159.785 ;
        RECT 21.755 158.475 21.925 159.485 ;
        RECT 22.095 159.205 22.990 159.580 ;
        RECT 22.095 158.645 22.435 159.205 ;
        RECT 22.665 158.475 22.980 158.975 ;
        RECT 23.160 158.945 23.330 159.785 ;
        RECT 23.500 160.075 23.965 160.405 ;
        RECT 24.350 160.345 24.520 160.575 ;
        RECT 24.700 160.525 25.070 161.025 ;
        RECT 25.390 160.575 26.065 160.745 ;
        RECT 26.260 160.575 26.595 160.745 ;
        RECT 23.500 159.115 23.820 160.075 ;
        RECT 24.350 160.045 25.180 160.345 ;
        RECT 23.990 159.145 24.180 159.865 ;
        RECT 24.350 158.975 24.520 160.045 ;
        RECT 24.980 160.015 25.180 160.045 ;
        RECT 24.690 159.795 24.860 159.865 ;
        RECT 25.390 159.795 25.560 160.575 ;
        RECT 26.425 160.435 26.595 160.575 ;
        RECT 26.765 160.565 27.015 161.025 ;
        RECT 24.690 159.625 25.560 159.795 ;
        RECT 25.730 160.155 26.255 160.375 ;
        RECT 26.425 160.305 26.650 160.435 ;
        RECT 24.690 159.535 25.200 159.625 ;
        RECT 23.160 158.775 24.045 158.945 ;
        RECT 24.270 158.645 24.520 158.975 ;
        RECT 24.690 158.475 24.860 159.275 ;
        RECT 25.030 158.920 25.200 159.535 ;
        RECT 25.730 159.455 25.900 160.155 ;
        RECT 25.370 159.090 25.900 159.455 ;
        RECT 26.070 159.390 26.310 159.985 ;
        RECT 26.480 159.200 26.650 160.305 ;
        RECT 26.820 159.445 27.100 160.395 ;
        RECT 26.345 159.070 26.650 159.200 ;
        RECT 25.030 158.750 26.135 158.920 ;
        RECT 26.345 158.645 26.595 159.070 ;
        RECT 26.765 158.475 27.030 158.935 ;
        RECT 27.270 158.645 27.455 160.765 ;
        RECT 27.625 160.645 27.955 161.025 ;
        RECT 28.125 160.475 28.295 160.765 ;
        RECT 27.630 160.305 28.295 160.475 ;
        RECT 27.630 159.315 27.860 160.305 ;
        RECT 28.555 160.255 31.145 161.025 ;
        RECT 31.780 160.375 32.050 160.585 ;
        RECT 32.270 160.565 32.600 161.025 ;
        RECT 33.110 160.565 33.860 160.855 ;
        RECT 28.030 159.485 28.380 160.135 ;
        RECT 28.555 159.735 29.765 160.255 ;
        RECT 31.780 160.205 33.115 160.375 ;
        RECT 29.935 159.565 31.145 160.085 ;
        RECT 32.945 160.035 33.115 160.205 ;
        RECT 31.780 159.795 32.130 160.035 ;
        RECT 32.300 159.795 32.775 160.035 ;
        RECT 32.945 159.785 33.320 160.035 ;
        RECT 32.945 159.615 33.115 159.785 ;
        RECT 27.630 159.145 28.295 159.315 ;
        RECT 27.625 158.475 27.955 158.975 ;
        RECT 28.125 158.645 28.295 159.145 ;
        RECT 28.555 158.475 31.145 159.565 ;
        RECT 31.780 159.445 33.115 159.615 ;
        RECT 31.780 159.285 32.060 159.445 ;
        RECT 33.490 159.275 33.860 160.565 ;
        RECT 34.080 160.260 34.535 161.025 ;
        RECT 34.810 160.645 36.110 160.855 ;
        RECT 36.365 160.665 36.695 161.025 ;
        RECT 35.940 160.495 36.110 160.645 ;
        RECT 36.865 160.525 37.125 160.855 ;
        RECT 36.895 160.515 37.125 160.525 ;
        RECT 35.010 160.035 35.230 160.435 ;
        RECT 34.075 159.835 34.565 160.035 ;
        RECT 34.755 159.825 35.230 160.035 ;
        RECT 35.475 160.035 35.685 160.435 ;
        RECT 35.940 160.370 36.695 160.495 ;
        RECT 35.940 160.325 36.785 160.370 ;
        RECT 36.515 160.205 36.785 160.325 ;
        RECT 35.475 159.825 35.805 160.035 ;
        RECT 35.975 159.765 36.385 160.070 ;
        RECT 32.270 158.475 32.520 159.275 ;
        RECT 32.690 159.105 33.860 159.275 ;
        RECT 34.080 159.595 35.255 159.655 ;
        RECT 36.615 159.630 36.785 160.205 ;
        RECT 36.585 159.595 36.785 159.630 ;
        RECT 34.080 159.485 36.785 159.595 ;
        RECT 32.690 158.645 33.020 159.105 ;
        RECT 33.190 158.475 33.405 158.935 ;
        RECT 34.080 158.865 34.335 159.485 ;
        RECT 34.925 159.425 36.725 159.485 ;
        RECT 34.925 159.395 35.255 159.425 ;
        RECT 36.955 159.325 37.125 160.515 ;
        RECT 37.295 160.275 38.505 161.025 ;
        RECT 38.675 160.285 39.015 160.855 ;
        RECT 39.210 160.360 39.380 161.025 ;
        RECT 39.660 160.685 39.880 160.730 ;
        RECT 39.655 160.515 39.880 160.685 ;
        RECT 40.050 160.545 40.495 160.715 ;
        RECT 39.660 160.375 39.880 160.515 ;
        RECT 37.295 159.735 37.815 160.275 ;
        RECT 37.985 159.565 38.505 160.105 ;
        RECT 34.585 159.225 34.770 159.315 ;
        RECT 35.360 159.225 36.195 159.235 ;
        RECT 34.585 159.025 36.195 159.225 ;
        RECT 34.585 158.985 34.815 159.025 ;
        RECT 34.080 158.645 34.415 158.865 ;
        RECT 35.420 158.475 35.775 158.855 ;
        RECT 35.945 158.645 36.195 159.025 ;
        RECT 36.445 158.475 36.695 159.255 ;
        RECT 36.865 158.645 37.125 159.325 ;
        RECT 37.295 158.475 38.505 159.565 ;
        RECT 38.675 159.315 38.850 160.285 ;
        RECT 39.660 160.205 40.155 160.375 ;
        RECT 39.020 159.665 39.190 160.115 ;
        RECT 39.360 159.835 39.810 160.035 ;
        RECT 39.980 160.010 40.155 160.205 ;
        RECT 40.325 159.755 40.495 160.545 ;
        RECT 40.665 160.420 40.915 160.790 ;
        RECT 40.745 160.035 40.915 160.420 ;
        RECT 41.085 160.385 41.335 160.790 ;
        RECT 41.505 160.555 41.675 161.025 ;
        RECT 41.845 160.385 42.185 160.790 ;
        RECT 41.085 160.205 42.185 160.385 ;
        RECT 43.275 160.300 43.565 161.025 ;
        RECT 43.735 160.255 45.405 161.025 ;
        RECT 45.585 160.665 47.655 160.855 ;
        RECT 47.885 160.665 48.215 161.025 ;
        RECT 48.745 160.665 49.075 161.025 ;
        RECT 49.605 160.665 49.935 161.025 ;
        RECT 46.535 160.645 47.655 160.665 ;
        RECT 40.745 159.865 40.940 160.035 ;
        RECT 39.020 159.495 39.415 159.665 ;
        RECT 40.325 159.615 40.600 159.755 ;
        RECT 38.675 158.645 38.935 159.315 ;
        RECT 39.245 159.225 39.415 159.495 ;
        RECT 39.585 159.395 40.600 159.615 ;
        RECT 40.770 159.615 40.940 159.865 ;
        RECT 41.110 159.785 41.670 160.035 ;
        RECT 40.770 159.225 41.325 159.615 ;
        RECT 39.245 159.055 41.325 159.225 ;
        RECT 39.105 158.475 39.435 158.875 ;
        RECT 40.305 158.475 40.705 158.875 ;
        RECT 40.995 158.820 41.325 159.055 ;
        RECT 41.495 158.685 41.670 159.785 ;
        RECT 41.840 159.465 42.185 160.035 ;
        RECT 43.735 159.735 44.485 160.255 ;
        RECT 41.840 158.475 42.185 159.295 ;
        RECT 43.275 158.475 43.565 159.640 ;
        RECT 44.655 159.565 45.405 160.085 ;
        RECT 43.735 158.475 45.405 159.565 ;
        RECT 45.575 159.140 45.865 160.115 ;
        RECT 46.035 159.570 46.365 160.440 ;
        RECT 46.535 160.220 46.725 160.645 ;
        RECT 49.245 160.475 49.435 160.595 ;
        RECT 46.895 160.265 49.435 160.475 ;
        RECT 49.605 160.035 49.945 160.345 ;
        RECT 50.175 160.225 50.870 160.855 ;
        RECT 51.075 160.225 51.385 161.025 ;
        RECT 51.640 160.455 51.815 160.855 ;
        RECT 51.985 160.645 52.315 161.025 ;
        RECT 52.560 160.525 52.790 160.855 ;
        RECT 51.640 160.285 52.270 160.455 ;
        RECT 46.535 159.745 47.395 160.035 ;
        RECT 47.855 159.755 48.825 160.035 ;
        RECT 48.995 159.865 49.945 160.035 ;
        RECT 49.050 159.815 49.945 159.865 ;
        RECT 50.195 159.785 50.530 160.035 ;
        RECT 50.700 159.625 50.870 160.225 ;
        RECT 52.100 160.115 52.270 160.285 ;
        RECT 51.040 159.785 51.375 160.055 ;
        RECT 46.035 159.400 48.645 159.570 ;
        RECT 45.605 158.475 45.865 158.935 ;
        RECT 46.035 158.645 46.295 159.400 ;
        RECT 46.465 158.475 46.795 159.195 ;
        RECT 46.965 158.645 47.155 159.400 ;
        RECT 47.325 158.475 47.655 159.195 ;
        RECT 47.885 158.815 48.145 159.010 ;
        RECT 48.315 158.985 48.645 159.400 ;
        RECT 48.815 159.415 49.935 159.585 ;
        RECT 48.815 158.815 49.005 159.415 ;
        RECT 47.885 158.645 49.005 158.815 ;
        RECT 49.175 158.475 49.505 159.245 ;
        RECT 49.675 158.645 49.935 159.415 ;
        RECT 50.175 158.475 50.435 159.615 ;
        RECT 50.605 158.645 50.935 159.625 ;
        RECT 51.105 158.475 51.385 159.615 ;
        RECT 51.555 159.435 51.920 160.115 ;
        RECT 52.100 159.785 52.450 160.115 ;
        RECT 52.100 159.265 52.270 159.785 ;
        RECT 51.640 159.095 52.270 159.265 ;
        RECT 52.620 159.235 52.790 160.525 ;
        RECT 52.990 159.415 53.270 160.690 ;
        RECT 53.495 160.685 53.765 160.690 ;
        RECT 53.455 160.515 53.765 160.685 ;
        RECT 54.225 160.645 54.555 161.025 ;
        RECT 54.725 160.770 55.060 160.815 ;
        RECT 53.495 159.415 53.765 160.515 ;
        RECT 53.955 159.415 54.295 160.445 ;
        RECT 54.725 160.305 55.065 160.770 ;
        RECT 55.285 160.370 55.615 160.805 ;
        RECT 55.785 160.415 55.955 161.025 ;
        RECT 54.465 159.785 54.725 160.115 ;
        RECT 54.465 159.235 54.635 159.785 ;
        RECT 54.895 159.615 55.065 160.305 ;
        RECT 51.640 158.645 51.815 159.095 ;
        RECT 52.620 159.065 54.635 159.235 ;
        RECT 51.985 158.475 52.315 158.915 ;
        RECT 52.620 158.645 52.790 159.065 ;
        RECT 53.025 158.475 53.695 158.885 ;
        RECT 53.910 158.645 54.080 159.065 ;
        RECT 54.280 158.475 54.610 158.885 ;
        RECT 54.805 158.645 55.065 159.615 ;
        RECT 55.235 160.285 55.615 160.370 ;
        RECT 56.125 160.285 56.455 160.810 ;
        RECT 56.715 160.495 56.925 161.025 ;
        RECT 57.200 160.575 57.985 160.745 ;
        RECT 58.155 160.575 58.560 160.745 ;
        RECT 55.235 160.245 55.460 160.285 ;
        RECT 55.235 159.665 55.405 160.245 ;
        RECT 56.125 160.115 56.325 160.285 ;
        RECT 57.200 160.115 57.370 160.575 ;
        RECT 55.575 159.785 56.325 160.115 ;
        RECT 56.495 159.785 57.370 160.115 ;
        RECT 55.235 159.615 55.450 159.665 ;
        RECT 55.235 159.535 55.625 159.615 ;
        RECT 55.295 158.690 55.625 159.535 ;
        RECT 56.135 159.580 56.325 159.785 ;
        RECT 55.795 158.475 55.965 159.485 ;
        RECT 56.135 159.205 57.030 159.580 ;
        RECT 56.135 158.645 56.475 159.205 ;
        RECT 56.705 158.475 57.020 158.975 ;
        RECT 57.200 158.945 57.370 159.785 ;
        RECT 57.540 160.075 58.005 160.405 ;
        RECT 58.390 160.345 58.560 160.575 ;
        RECT 58.740 160.525 59.110 161.025 ;
        RECT 59.430 160.575 60.105 160.745 ;
        RECT 60.300 160.575 60.635 160.745 ;
        RECT 57.540 159.115 57.860 160.075 ;
        RECT 58.390 160.045 59.220 160.345 ;
        RECT 58.030 159.145 58.220 159.865 ;
        RECT 58.390 158.975 58.560 160.045 ;
        RECT 59.020 160.015 59.220 160.045 ;
        RECT 58.730 159.795 58.900 159.865 ;
        RECT 59.430 159.795 59.600 160.575 ;
        RECT 60.465 160.435 60.635 160.575 ;
        RECT 60.805 160.565 61.055 161.025 ;
        RECT 58.730 159.625 59.600 159.795 ;
        RECT 59.770 160.155 60.295 160.375 ;
        RECT 60.465 160.305 60.690 160.435 ;
        RECT 58.730 159.535 59.240 159.625 ;
        RECT 57.200 158.775 58.085 158.945 ;
        RECT 58.310 158.645 58.560 158.975 ;
        RECT 58.730 158.475 58.900 159.275 ;
        RECT 59.070 158.920 59.240 159.535 ;
        RECT 59.770 159.455 59.940 160.155 ;
        RECT 59.410 159.090 59.940 159.455 ;
        RECT 60.110 159.390 60.350 159.985 ;
        RECT 60.520 159.200 60.690 160.305 ;
        RECT 60.860 159.445 61.140 160.395 ;
        RECT 60.385 159.070 60.690 159.200 ;
        RECT 59.070 158.750 60.175 158.920 ;
        RECT 60.385 158.645 60.635 159.070 ;
        RECT 60.805 158.475 61.070 158.935 ;
        RECT 61.310 158.645 61.495 160.765 ;
        RECT 61.665 160.645 61.995 161.025 ;
        RECT 62.600 160.770 62.935 160.815 ;
        RECT 62.165 160.475 62.335 160.765 ;
        RECT 61.670 160.305 62.335 160.475 ;
        RECT 62.595 160.305 62.935 160.770 ;
        RECT 63.105 160.645 63.435 161.025 ;
        RECT 61.670 159.315 61.900 160.305 ;
        RECT 62.070 159.485 62.420 160.135 ;
        RECT 62.595 159.615 62.765 160.305 ;
        RECT 62.935 159.785 63.195 160.115 ;
        RECT 61.670 159.145 62.335 159.315 ;
        RECT 61.665 158.475 61.995 158.975 ;
        RECT 62.165 158.645 62.335 159.145 ;
        RECT 62.595 158.645 62.855 159.615 ;
        RECT 63.025 159.235 63.195 159.785 ;
        RECT 63.365 159.415 63.705 160.445 ;
        RECT 63.895 160.345 64.165 160.690 ;
        RECT 63.895 160.175 64.205 160.345 ;
        RECT 63.895 159.415 64.165 160.175 ;
        RECT 64.390 159.415 64.670 160.690 ;
        RECT 64.870 160.525 65.100 160.855 ;
        RECT 65.345 160.645 65.675 161.025 ;
        RECT 64.870 159.235 65.040 160.525 ;
        RECT 65.845 160.455 66.020 160.855 ;
        RECT 65.390 160.285 66.020 160.455 ;
        RECT 65.390 160.115 65.560 160.285 ;
        RECT 66.275 160.255 68.865 161.025 ;
        RECT 69.035 160.300 69.325 161.025 ;
        RECT 69.495 160.255 71.165 161.025 ;
        RECT 71.340 160.520 71.675 161.025 ;
        RECT 71.845 160.455 72.085 160.830 ;
        RECT 72.365 160.695 72.535 160.840 ;
        RECT 72.365 160.500 72.740 160.695 ;
        RECT 73.100 160.530 73.495 161.025 ;
        RECT 65.210 159.785 65.560 160.115 ;
        RECT 63.025 159.065 65.040 159.235 ;
        RECT 65.390 159.265 65.560 159.785 ;
        RECT 65.740 159.435 66.105 160.115 ;
        RECT 66.275 159.735 67.485 160.255 ;
        RECT 67.655 159.565 68.865 160.085 ;
        RECT 69.495 159.735 70.245 160.255 ;
        RECT 65.390 159.095 66.020 159.265 ;
        RECT 63.050 158.475 63.380 158.885 ;
        RECT 63.580 158.645 63.750 159.065 ;
        RECT 63.965 158.475 64.635 158.885 ;
        RECT 64.870 158.645 65.040 159.065 ;
        RECT 65.345 158.475 65.675 158.915 ;
        RECT 65.845 158.645 66.020 159.095 ;
        RECT 66.275 158.475 68.865 159.565 ;
        RECT 69.035 158.475 69.325 159.640 ;
        RECT 70.415 159.565 71.165 160.085 ;
        RECT 69.495 158.475 71.165 159.565 ;
        RECT 71.395 159.495 71.695 160.345 ;
        RECT 71.865 160.305 72.085 160.455 ;
        RECT 71.865 159.975 72.400 160.305 ;
        RECT 72.570 160.165 72.740 160.500 ;
        RECT 73.665 160.335 73.905 160.855 ;
        RECT 74.105 160.525 74.435 161.025 ;
        RECT 74.635 160.455 74.805 160.805 ;
        RECT 75.005 160.625 75.335 161.025 ;
        RECT 75.505 160.455 75.675 160.805 ;
        RECT 75.845 160.625 76.225 161.025 ;
        RECT 71.865 159.325 72.100 159.975 ;
        RECT 72.570 159.805 73.555 160.165 ;
        RECT 71.425 159.095 72.100 159.325 ;
        RECT 72.270 159.785 73.555 159.805 ;
        RECT 72.270 159.635 73.130 159.785 ;
        RECT 71.425 158.665 71.595 159.095 ;
        RECT 71.765 158.475 72.095 158.925 ;
        RECT 72.270 158.690 72.555 159.635 ;
        RECT 73.730 159.530 73.905 160.335 ;
        RECT 74.100 159.785 74.450 160.355 ;
        RECT 74.635 160.285 76.245 160.455 ;
        RECT 76.415 160.350 76.685 160.695 ;
        RECT 76.075 160.115 76.245 160.285 ;
        RECT 72.730 159.155 73.425 159.465 ;
        RECT 72.735 158.475 73.420 158.945 ;
        RECT 73.600 158.745 73.905 159.530 ;
        RECT 74.100 159.325 74.420 159.615 ;
        RECT 74.620 159.495 75.330 160.115 ;
        RECT 75.500 159.785 75.905 160.115 ;
        RECT 76.075 159.785 76.345 160.115 ;
        RECT 76.075 159.615 76.245 159.785 ;
        RECT 76.515 159.615 76.685 160.350 ;
        RECT 76.905 160.485 77.130 160.845 ;
        RECT 77.310 160.655 77.640 161.025 ;
        RECT 77.820 160.485 78.075 160.845 ;
        RECT 78.640 160.655 79.385 161.025 ;
        RECT 76.905 160.295 79.390 160.485 ;
        RECT 76.865 159.785 77.135 160.115 ;
        RECT 77.315 159.785 77.750 160.115 ;
        RECT 77.930 159.785 78.505 160.115 ;
        RECT 78.685 159.785 78.965 160.115 ;
        RECT 75.520 159.445 76.245 159.615 ;
        RECT 75.520 159.325 75.690 159.445 ;
        RECT 74.100 159.155 75.690 159.325 ;
        RECT 74.100 158.695 75.755 158.985 ;
        RECT 75.925 158.475 76.205 159.275 ;
        RECT 76.415 158.645 76.685 159.615 ;
        RECT 79.165 159.605 79.390 160.295 ;
        RECT 76.895 159.425 79.390 159.605 ;
        RECT 79.565 159.425 79.900 160.845 ;
        RECT 76.895 158.655 77.185 159.425 ;
        RECT 77.755 159.015 78.945 159.245 ;
        RECT 77.755 158.655 78.015 159.015 ;
        RECT 78.185 158.475 78.515 158.845 ;
        RECT 78.685 158.655 78.945 159.015 ;
        RECT 79.135 158.475 79.465 159.195 ;
        RECT 79.635 158.655 79.900 159.425 ;
        RECT 80.995 160.375 81.255 160.855 ;
        RECT 81.425 160.565 81.755 161.025 ;
        RECT 81.945 160.385 82.145 160.805 ;
        RECT 80.995 159.345 81.165 160.375 ;
        RECT 81.335 159.685 81.565 160.115 ;
        RECT 81.735 159.865 82.145 160.385 ;
        RECT 82.315 160.540 83.105 160.805 ;
        RECT 82.315 159.685 82.570 160.540 ;
        RECT 83.285 160.205 83.615 160.625 ;
        RECT 83.785 160.205 84.045 161.025 ;
        RECT 84.265 160.370 84.595 160.805 ;
        RECT 84.765 160.415 84.935 161.025 ;
        RECT 84.215 160.285 84.595 160.370 ;
        RECT 85.105 160.285 85.435 160.810 ;
        RECT 85.695 160.495 85.905 161.025 ;
        RECT 86.180 160.575 86.965 160.745 ;
        RECT 87.135 160.575 87.540 160.745 ;
        RECT 84.215 160.245 84.440 160.285 ;
        RECT 83.285 160.115 83.535 160.205 ;
        RECT 82.740 159.865 83.535 160.115 ;
        RECT 81.335 159.515 83.125 159.685 ;
        RECT 80.995 158.645 81.270 159.345 ;
        RECT 81.440 159.220 82.155 159.515 ;
        RECT 82.375 159.155 82.705 159.345 ;
        RECT 81.480 158.475 81.695 159.020 ;
        RECT 81.865 158.645 82.340 158.985 ;
        RECT 82.510 158.980 82.705 159.155 ;
        RECT 82.875 159.150 83.125 159.515 ;
        RECT 82.510 158.475 83.125 158.980 ;
        RECT 83.365 158.645 83.535 159.865 ;
        RECT 83.705 159.155 84.045 160.035 ;
        RECT 84.215 159.665 84.385 160.245 ;
        RECT 85.105 160.115 85.305 160.285 ;
        RECT 86.180 160.115 86.350 160.575 ;
        RECT 84.555 159.785 85.305 160.115 ;
        RECT 85.475 159.785 86.350 160.115 ;
        RECT 84.215 159.615 84.430 159.665 ;
        RECT 84.215 159.535 84.605 159.615 ;
        RECT 83.785 158.475 84.045 158.985 ;
        RECT 84.275 158.690 84.605 159.535 ;
        RECT 85.115 159.580 85.305 159.785 ;
        RECT 84.775 158.475 84.945 159.485 ;
        RECT 85.115 159.205 86.010 159.580 ;
        RECT 85.115 158.645 85.455 159.205 ;
        RECT 85.685 158.475 86.000 158.975 ;
        RECT 86.180 158.945 86.350 159.785 ;
        RECT 86.520 160.075 86.985 160.405 ;
        RECT 87.370 160.345 87.540 160.575 ;
        RECT 87.720 160.525 88.090 161.025 ;
        RECT 88.410 160.575 89.085 160.745 ;
        RECT 89.280 160.575 89.615 160.745 ;
        RECT 86.520 159.115 86.840 160.075 ;
        RECT 87.370 160.045 88.200 160.345 ;
        RECT 87.010 159.145 87.200 159.865 ;
        RECT 87.370 158.975 87.540 160.045 ;
        RECT 88.000 160.015 88.200 160.045 ;
        RECT 87.710 159.795 87.880 159.865 ;
        RECT 88.410 159.795 88.580 160.575 ;
        RECT 89.445 160.435 89.615 160.575 ;
        RECT 89.785 160.565 90.035 161.025 ;
        RECT 87.710 159.625 88.580 159.795 ;
        RECT 88.750 160.155 89.275 160.375 ;
        RECT 89.445 160.305 89.670 160.435 ;
        RECT 87.710 159.535 88.220 159.625 ;
        RECT 86.180 158.775 87.065 158.945 ;
        RECT 87.290 158.645 87.540 158.975 ;
        RECT 87.710 158.475 87.880 159.275 ;
        RECT 88.050 158.920 88.220 159.535 ;
        RECT 88.750 159.455 88.920 160.155 ;
        RECT 88.390 159.090 88.920 159.455 ;
        RECT 89.090 159.390 89.330 159.985 ;
        RECT 89.500 159.200 89.670 160.305 ;
        RECT 89.840 159.445 90.120 160.395 ;
        RECT 89.365 159.070 89.670 159.200 ;
        RECT 88.050 158.750 89.155 158.920 ;
        RECT 89.365 158.645 89.615 159.070 ;
        RECT 89.785 158.475 90.050 158.935 ;
        RECT 90.290 158.645 90.475 160.765 ;
        RECT 90.645 160.645 90.975 161.025 ;
        RECT 91.145 160.475 91.315 160.765 ;
        RECT 90.650 160.305 91.315 160.475 ;
        RECT 90.650 159.315 90.880 160.305 ;
        RECT 91.575 160.255 94.165 161.025 ;
        RECT 94.795 160.300 95.085 161.025 ;
        RECT 96.225 160.370 96.555 160.805 ;
        RECT 96.725 160.415 96.895 161.025 ;
        RECT 96.175 160.285 96.555 160.370 ;
        RECT 97.065 160.285 97.395 160.810 ;
        RECT 97.655 160.495 97.865 161.025 ;
        RECT 98.140 160.575 98.925 160.745 ;
        RECT 99.095 160.575 99.500 160.745 ;
        RECT 91.050 159.485 91.400 160.135 ;
        RECT 91.575 159.735 92.785 160.255 ;
        RECT 96.175 160.245 96.400 160.285 ;
        RECT 92.955 159.565 94.165 160.085 ;
        RECT 96.175 159.665 96.345 160.245 ;
        RECT 97.065 160.115 97.265 160.285 ;
        RECT 98.140 160.115 98.310 160.575 ;
        RECT 96.515 159.785 97.265 160.115 ;
        RECT 97.435 159.785 98.310 160.115 ;
        RECT 90.650 159.145 91.315 159.315 ;
        RECT 90.645 158.475 90.975 158.975 ;
        RECT 91.145 158.645 91.315 159.145 ;
        RECT 91.575 158.475 94.165 159.565 ;
        RECT 94.795 158.475 95.085 159.640 ;
        RECT 96.175 159.615 96.390 159.665 ;
        RECT 96.175 159.535 96.565 159.615 ;
        RECT 96.235 158.690 96.565 159.535 ;
        RECT 97.075 159.580 97.265 159.785 ;
        RECT 96.735 158.475 96.905 159.485 ;
        RECT 97.075 159.205 97.970 159.580 ;
        RECT 97.075 158.645 97.415 159.205 ;
        RECT 97.645 158.475 97.960 158.975 ;
        RECT 98.140 158.945 98.310 159.785 ;
        RECT 98.480 160.075 98.945 160.405 ;
        RECT 99.330 160.345 99.500 160.575 ;
        RECT 99.680 160.525 100.050 161.025 ;
        RECT 100.370 160.575 101.045 160.745 ;
        RECT 101.240 160.575 101.575 160.745 ;
        RECT 98.480 159.115 98.800 160.075 ;
        RECT 99.330 160.045 100.160 160.345 ;
        RECT 98.970 159.145 99.160 159.865 ;
        RECT 99.330 158.975 99.500 160.045 ;
        RECT 99.960 160.015 100.160 160.045 ;
        RECT 99.670 159.795 99.840 159.865 ;
        RECT 100.370 159.795 100.540 160.575 ;
        RECT 101.405 160.435 101.575 160.575 ;
        RECT 101.745 160.565 101.995 161.025 ;
        RECT 99.670 159.625 100.540 159.795 ;
        RECT 100.710 160.155 101.235 160.375 ;
        RECT 101.405 160.305 101.630 160.435 ;
        RECT 99.670 159.535 100.180 159.625 ;
        RECT 98.140 158.775 99.025 158.945 ;
        RECT 99.250 158.645 99.500 158.975 ;
        RECT 99.670 158.475 99.840 159.275 ;
        RECT 100.010 158.920 100.180 159.535 ;
        RECT 100.710 159.455 100.880 160.155 ;
        RECT 100.350 159.090 100.880 159.455 ;
        RECT 101.050 159.390 101.290 159.985 ;
        RECT 101.460 159.200 101.630 160.305 ;
        RECT 101.800 159.445 102.080 160.395 ;
        RECT 101.325 159.070 101.630 159.200 ;
        RECT 100.010 158.750 101.115 158.920 ;
        RECT 101.325 158.645 101.575 159.070 ;
        RECT 101.745 158.475 102.010 158.935 ;
        RECT 102.250 158.645 102.435 160.765 ;
        RECT 102.605 160.645 102.935 161.025 ;
        RECT 103.105 160.475 103.275 160.765 ;
        RECT 102.610 160.305 103.275 160.475 ;
        RECT 102.610 159.315 102.840 160.305 ;
        RECT 103.010 159.485 103.360 160.135 ;
        RECT 102.610 159.145 103.275 159.315 ;
        RECT 102.605 158.475 102.935 158.975 ;
        RECT 103.105 158.645 103.275 159.145 ;
        RECT 103.535 158.645 103.815 160.745 ;
        RECT 104.045 160.565 104.215 161.025 ;
        RECT 104.485 160.635 105.735 160.815 ;
        RECT 104.870 160.395 105.235 160.465 ;
        RECT 103.985 160.215 105.235 160.395 ;
        RECT 105.405 160.415 105.735 160.635 ;
        RECT 105.905 160.585 106.075 161.025 ;
        RECT 106.245 160.415 106.585 160.830 ;
        RECT 105.405 160.245 106.585 160.415 ;
        RECT 106.755 160.255 108.425 161.025 ;
        RECT 109.255 160.395 109.585 160.755 ;
        RECT 110.205 160.565 110.455 161.025 ;
        RECT 110.625 160.565 111.185 160.855 ;
        RECT 103.985 159.615 104.260 160.215 ;
        RECT 104.430 159.785 104.785 160.035 ;
        RECT 104.980 160.005 105.445 160.035 ;
        RECT 104.975 159.835 105.445 160.005 ;
        RECT 104.980 159.785 105.445 159.835 ;
        RECT 105.615 159.785 105.945 160.035 ;
        RECT 106.120 159.835 106.585 160.035 ;
        RECT 105.765 159.665 105.945 159.785 ;
        RECT 106.755 159.735 107.505 160.255 ;
        RECT 109.255 160.205 110.645 160.395 ;
        RECT 110.475 160.115 110.645 160.205 ;
        RECT 103.985 159.405 105.595 159.615 ;
        RECT 105.765 159.495 106.095 159.665 ;
        RECT 105.185 159.305 105.595 159.405 ;
        RECT 104.005 158.475 104.790 159.235 ;
        RECT 105.185 158.645 105.570 159.305 ;
        RECT 105.895 158.705 106.095 159.495 ;
        RECT 106.265 158.475 106.585 159.655 ;
        RECT 107.675 159.565 108.425 160.085 ;
        RECT 106.755 158.475 108.425 159.565 ;
        RECT 109.070 159.785 109.745 160.035 ;
        RECT 109.965 159.785 110.305 160.035 ;
        RECT 110.475 159.785 110.765 160.115 ;
        RECT 109.070 159.425 109.335 159.785 ;
        RECT 110.475 159.535 110.645 159.785 ;
        RECT 109.705 159.365 110.645 159.535 ;
        RECT 109.255 158.475 109.535 159.145 ;
        RECT 109.705 158.815 110.005 159.365 ;
        RECT 110.935 159.195 111.185 160.565 ;
        RECT 111.415 160.205 111.625 161.025 ;
        RECT 111.795 160.225 112.125 160.855 ;
        RECT 111.795 159.625 112.045 160.225 ;
        RECT 112.295 160.205 112.525 161.025 ;
        RECT 112.735 160.225 113.430 160.855 ;
        RECT 113.635 160.225 113.945 161.025 ;
        RECT 113.255 160.175 113.430 160.225 ;
        RECT 114.125 160.215 114.395 161.025 ;
        RECT 114.565 160.215 114.895 160.855 ;
        RECT 115.065 160.215 115.305 161.025 ;
        RECT 115.495 160.225 116.190 160.855 ;
        RECT 116.395 160.225 116.705 161.025 ;
        RECT 118.075 160.395 118.455 160.845 ;
        RECT 112.215 159.785 112.545 160.035 ;
        RECT 112.755 159.785 113.090 160.035 ;
        RECT 113.260 159.625 113.430 160.175 ;
        RECT 113.600 159.785 113.935 160.055 ;
        RECT 114.115 159.785 114.465 160.035 ;
        RECT 110.205 158.475 110.535 159.195 ;
        RECT 110.725 158.645 111.185 159.195 ;
        RECT 111.415 158.475 111.625 159.615 ;
        RECT 111.795 158.645 112.125 159.625 ;
        RECT 112.295 158.475 112.525 159.615 ;
        RECT 112.735 158.475 112.995 159.615 ;
        RECT 113.165 158.645 113.495 159.625 ;
        RECT 114.635 159.615 114.805 160.215 ;
        RECT 114.975 159.785 115.325 160.035 ;
        RECT 115.515 159.785 115.850 160.035 ;
        RECT 116.020 159.665 116.190 160.225 ;
        RECT 116.360 159.785 116.695 160.055 ;
        RECT 116.015 159.625 116.190 159.665 ;
        RECT 113.665 158.475 113.945 159.615 ;
        RECT 114.125 158.475 114.455 159.615 ;
        RECT 114.635 159.445 115.315 159.615 ;
        RECT 114.985 158.660 115.315 159.445 ;
        RECT 115.495 158.475 115.755 159.615 ;
        RECT 115.925 158.645 116.255 159.625 ;
        RECT 116.425 158.475 116.705 159.615 ;
        RECT 117.815 159.445 118.045 160.135 ;
        RECT 118.225 159.945 118.455 160.395 ;
        RECT 118.635 160.245 118.865 161.025 ;
        RECT 119.045 160.315 119.475 160.845 ;
        RECT 119.045 160.065 119.290 160.315 ;
        RECT 119.655 160.115 119.865 160.735 ;
        RECT 120.035 160.295 120.365 161.025 ;
        RECT 120.555 160.300 120.845 161.025 ;
        RECT 121.030 160.455 121.285 160.805 ;
        RECT 121.455 160.625 121.785 161.025 ;
        RECT 121.955 160.455 122.125 160.805 ;
        RECT 122.295 160.625 122.675 161.025 ;
        RECT 121.030 160.285 122.695 160.455 ;
        RECT 122.865 160.350 123.140 160.695 ;
        RECT 123.375 160.565 123.620 161.025 ;
        RECT 122.525 160.115 122.695 160.285 ;
        RECT 118.225 159.265 118.565 159.945 ;
        RECT 117.805 159.065 118.565 159.265 ;
        RECT 118.755 159.765 119.290 160.065 ;
        RECT 119.470 159.765 119.865 160.115 ;
        RECT 120.060 159.765 120.350 160.115 ;
        RECT 121.015 159.785 121.360 160.115 ;
        RECT 121.530 159.785 122.355 160.115 ;
        RECT 122.525 159.785 122.800 160.115 ;
        RECT 117.805 158.675 118.065 159.065 ;
        RECT 118.235 158.475 118.565 158.885 ;
        RECT 118.755 158.655 119.085 159.765 ;
        RECT 119.255 159.385 120.295 159.585 ;
        RECT 119.255 158.655 119.445 159.385 ;
        RECT 119.615 158.475 119.945 159.205 ;
        RECT 120.125 158.655 120.295 159.385 ;
        RECT 120.555 158.475 120.845 159.640 ;
        RECT 121.035 159.325 121.360 159.615 ;
        RECT 121.530 159.495 121.725 159.785 ;
        RECT 122.525 159.615 122.695 159.785 ;
        RECT 122.970 159.615 123.140 160.350 ;
        RECT 123.315 159.785 123.630 160.395 ;
        RECT 123.800 160.035 124.050 160.845 ;
        RECT 124.220 160.500 124.480 161.025 ;
        RECT 124.650 160.375 124.910 160.830 ;
        RECT 125.080 160.545 125.340 161.025 ;
        RECT 125.510 160.375 125.770 160.830 ;
        RECT 125.940 160.545 126.200 161.025 ;
        RECT 126.370 160.375 126.630 160.830 ;
        RECT 126.800 160.545 127.060 161.025 ;
        RECT 127.230 160.375 127.490 160.830 ;
        RECT 127.660 160.545 127.960 161.025 ;
        RECT 124.650 160.205 127.960 160.375 ;
        RECT 128.375 160.225 129.070 160.855 ;
        RECT 129.275 160.225 129.585 161.025 ;
        RECT 130.765 160.475 130.935 160.765 ;
        RECT 131.105 160.645 131.435 161.025 ;
        RECT 130.765 160.305 131.430 160.475 ;
        RECT 123.800 159.785 126.820 160.035 ;
        RECT 122.035 159.445 122.695 159.615 ;
        RECT 122.035 159.325 122.205 159.445 ;
        RECT 121.035 159.155 122.205 159.325 ;
        RECT 121.015 158.695 122.205 158.985 ;
        RECT 122.375 158.475 122.655 159.275 ;
        RECT 122.865 158.645 123.140 159.615 ;
        RECT 123.325 158.475 123.620 159.585 ;
        RECT 123.800 158.650 124.050 159.785 ;
        RECT 126.990 159.615 127.960 160.205 ;
        RECT 128.395 159.785 128.730 160.035 ;
        RECT 128.900 159.625 129.070 160.225 ;
        RECT 129.240 159.785 129.575 160.055 ;
        RECT 124.220 158.475 124.480 159.585 ;
        RECT 124.650 159.375 127.960 159.615 ;
        RECT 124.650 158.650 124.910 159.375 ;
        RECT 125.080 158.475 125.340 159.205 ;
        RECT 125.510 158.650 125.770 159.375 ;
        RECT 125.940 158.475 126.200 159.205 ;
        RECT 126.370 158.650 126.630 159.375 ;
        RECT 126.800 158.475 127.060 159.205 ;
        RECT 127.230 158.650 127.490 159.375 ;
        RECT 127.660 158.475 127.955 159.205 ;
        RECT 128.375 158.475 128.635 159.615 ;
        RECT 128.805 158.645 129.135 159.625 ;
        RECT 129.305 158.475 129.585 159.615 ;
        RECT 130.680 159.485 131.030 160.135 ;
        RECT 131.200 159.315 131.430 160.305 ;
        RECT 130.765 159.145 131.430 159.315 ;
        RECT 130.765 158.645 130.935 159.145 ;
        RECT 131.105 158.475 131.435 158.975 ;
        RECT 131.605 158.645 131.790 160.765 ;
        RECT 132.045 160.565 132.295 161.025 ;
        RECT 132.465 160.575 132.800 160.745 ;
        RECT 132.995 160.575 133.670 160.745 ;
        RECT 132.465 160.435 132.635 160.575 ;
        RECT 131.960 159.445 132.240 160.395 ;
        RECT 132.410 160.305 132.635 160.435 ;
        RECT 132.410 159.200 132.580 160.305 ;
        RECT 132.805 160.155 133.330 160.375 ;
        RECT 132.750 159.390 132.990 159.985 ;
        RECT 133.160 159.455 133.330 160.155 ;
        RECT 133.500 159.795 133.670 160.575 ;
        RECT 133.990 160.525 134.360 161.025 ;
        RECT 134.540 160.575 134.945 160.745 ;
        RECT 135.115 160.575 135.900 160.745 ;
        RECT 134.540 160.345 134.710 160.575 ;
        RECT 133.880 160.045 134.710 160.345 ;
        RECT 135.095 160.075 135.560 160.405 ;
        RECT 133.880 160.015 134.080 160.045 ;
        RECT 134.200 159.795 134.370 159.865 ;
        RECT 133.500 159.625 134.370 159.795 ;
        RECT 133.860 159.535 134.370 159.625 ;
        RECT 132.410 159.070 132.715 159.200 ;
        RECT 133.160 159.090 133.690 159.455 ;
        RECT 132.030 158.475 132.295 158.935 ;
        RECT 132.465 158.645 132.715 159.070 ;
        RECT 133.860 158.920 134.030 159.535 ;
        RECT 132.925 158.750 134.030 158.920 ;
        RECT 134.200 158.475 134.370 159.275 ;
        RECT 134.540 158.975 134.710 160.045 ;
        RECT 134.880 159.145 135.070 159.865 ;
        RECT 135.240 159.115 135.560 160.075 ;
        RECT 135.730 160.115 135.900 160.575 ;
        RECT 136.175 160.495 136.385 161.025 ;
        RECT 136.645 160.285 136.975 160.810 ;
        RECT 137.145 160.415 137.315 161.025 ;
        RECT 137.485 160.370 137.815 160.805 ;
        RECT 138.125 160.475 138.295 160.855 ;
        RECT 138.510 160.645 138.840 161.025 ;
        RECT 137.485 160.285 137.865 160.370 ;
        RECT 138.125 160.305 138.840 160.475 ;
        RECT 136.775 160.115 136.975 160.285 ;
        RECT 137.640 160.245 137.865 160.285 ;
        RECT 135.730 159.785 136.605 160.115 ;
        RECT 136.775 159.785 137.525 160.115 ;
        RECT 134.540 158.645 134.790 158.975 ;
        RECT 135.730 158.945 135.900 159.785 ;
        RECT 136.775 159.580 136.965 159.785 ;
        RECT 137.695 159.665 137.865 160.245 ;
        RECT 138.035 159.755 138.390 160.125 ;
        RECT 138.670 160.115 138.840 160.305 ;
        RECT 139.010 160.280 139.265 160.855 ;
        RECT 138.670 159.785 138.925 160.115 ;
        RECT 137.650 159.615 137.865 159.665 ;
        RECT 136.070 159.205 136.965 159.580 ;
        RECT 137.475 159.535 137.865 159.615 ;
        RECT 138.670 159.575 138.840 159.785 ;
        RECT 135.015 158.775 135.900 158.945 ;
        RECT 136.080 158.475 136.395 158.975 ;
        RECT 136.625 158.645 136.965 159.205 ;
        RECT 137.135 158.475 137.305 159.485 ;
        RECT 137.475 158.690 137.805 159.535 ;
        RECT 138.125 159.405 138.840 159.575 ;
        RECT 139.095 159.550 139.265 160.280 ;
        RECT 139.440 160.185 139.700 161.025 ;
        RECT 139.965 160.475 140.135 160.855 ;
        RECT 140.350 160.645 140.680 161.025 ;
        RECT 139.965 160.305 140.680 160.475 ;
        RECT 139.875 159.755 140.230 160.125 ;
        RECT 140.510 160.115 140.680 160.305 ;
        RECT 140.850 160.280 141.105 160.855 ;
        RECT 140.510 159.785 140.765 160.115 ;
        RECT 138.125 158.645 138.295 159.405 ;
        RECT 138.510 158.475 138.840 159.235 ;
        RECT 139.010 158.645 139.265 159.550 ;
        RECT 139.440 158.475 139.700 159.625 ;
        RECT 140.510 159.575 140.680 159.785 ;
        RECT 139.965 159.405 140.680 159.575 ;
        RECT 140.935 159.550 141.105 160.280 ;
        RECT 141.280 160.185 141.540 161.025 ;
        RECT 141.715 160.275 142.925 161.025 ;
        RECT 139.965 158.645 140.135 159.405 ;
        RECT 140.350 158.475 140.680 159.235 ;
        RECT 140.850 158.645 141.105 159.550 ;
        RECT 141.280 158.475 141.540 159.625 ;
        RECT 141.715 159.565 142.235 160.105 ;
        RECT 142.405 159.735 142.925 160.275 ;
        RECT 141.715 158.475 142.925 159.565 ;
        RECT 17.430 158.305 143.010 158.475 ;
        RECT 17.515 157.215 18.725 158.305 ;
        RECT 19.905 157.635 20.075 158.135 ;
        RECT 20.245 157.805 20.575 158.305 ;
        RECT 19.905 157.465 20.570 157.635 ;
        RECT 17.515 156.505 18.035 157.045 ;
        RECT 18.205 156.675 18.725 157.215 ;
        RECT 19.820 156.645 20.170 157.295 ;
        RECT 17.515 155.755 18.725 156.505 ;
        RECT 20.340 156.475 20.570 157.465 ;
        RECT 19.905 156.305 20.570 156.475 ;
        RECT 19.905 156.015 20.075 156.305 ;
        RECT 20.245 155.755 20.575 156.135 ;
        RECT 20.745 156.015 20.930 158.135 ;
        RECT 21.170 157.845 21.435 158.305 ;
        RECT 21.605 157.710 21.855 158.135 ;
        RECT 22.065 157.860 23.170 158.030 ;
        RECT 21.550 157.580 21.855 157.710 ;
        RECT 21.100 156.385 21.380 157.335 ;
        RECT 21.550 156.475 21.720 157.580 ;
        RECT 21.890 156.795 22.130 157.390 ;
        RECT 22.300 157.325 22.830 157.690 ;
        RECT 22.300 156.625 22.470 157.325 ;
        RECT 23.000 157.245 23.170 157.860 ;
        RECT 23.340 157.505 23.510 158.305 ;
        RECT 23.680 157.805 23.930 158.135 ;
        RECT 24.155 157.835 25.040 158.005 ;
        RECT 23.000 157.155 23.510 157.245 ;
        RECT 21.550 156.345 21.775 156.475 ;
        RECT 21.945 156.405 22.470 156.625 ;
        RECT 22.640 156.985 23.510 157.155 ;
        RECT 21.185 155.755 21.435 156.215 ;
        RECT 21.605 156.205 21.775 156.345 ;
        RECT 22.640 156.205 22.810 156.985 ;
        RECT 23.340 156.915 23.510 156.985 ;
        RECT 23.020 156.735 23.220 156.765 ;
        RECT 23.680 156.735 23.850 157.805 ;
        RECT 24.020 156.915 24.210 157.635 ;
        RECT 23.020 156.435 23.850 156.735 ;
        RECT 24.380 156.705 24.700 157.665 ;
        RECT 21.605 156.035 21.940 156.205 ;
        RECT 22.135 156.035 22.810 156.205 ;
        RECT 23.130 155.755 23.500 156.255 ;
        RECT 23.680 156.205 23.850 156.435 ;
        RECT 24.235 156.375 24.700 156.705 ;
        RECT 24.870 156.995 25.040 157.835 ;
        RECT 25.220 157.805 25.535 158.305 ;
        RECT 25.765 157.575 26.105 158.135 ;
        RECT 25.210 157.200 26.105 157.575 ;
        RECT 26.275 157.295 26.445 158.305 ;
        RECT 25.915 156.995 26.105 157.200 ;
        RECT 26.615 157.245 26.945 158.090 ;
        RECT 26.615 157.165 27.005 157.245 ;
        RECT 27.175 157.215 29.765 158.305 ;
        RECT 26.790 157.115 27.005 157.165 ;
        RECT 24.870 156.665 25.745 156.995 ;
        RECT 25.915 156.665 26.665 156.995 ;
        RECT 24.870 156.205 25.040 156.665 ;
        RECT 25.915 156.495 26.115 156.665 ;
        RECT 26.835 156.535 27.005 157.115 ;
        RECT 26.780 156.495 27.005 156.535 ;
        RECT 23.680 156.035 24.085 156.205 ;
        RECT 24.255 156.035 25.040 156.205 ;
        RECT 25.315 155.755 25.525 156.285 ;
        RECT 25.785 155.970 26.115 156.495 ;
        RECT 26.625 156.410 27.005 156.495 ;
        RECT 27.175 156.525 28.385 157.045 ;
        RECT 28.555 156.695 29.765 157.215 ;
        RECT 30.395 157.140 30.685 158.305 ;
        RECT 30.910 157.435 31.195 158.305 ;
        RECT 31.365 157.675 31.625 158.135 ;
        RECT 31.800 157.845 32.055 158.305 ;
        RECT 32.225 157.675 32.485 158.135 ;
        RECT 31.365 157.505 32.485 157.675 ;
        RECT 32.655 157.505 32.965 158.305 ;
        RECT 31.365 157.255 31.625 157.505 ;
        RECT 33.135 157.335 33.445 158.135 ;
        RECT 33.615 157.870 38.960 158.305 ;
        RECT 30.870 157.085 31.625 157.255 ;
        RECT 32.415 157.165 33.445 157.335 ;
        RECT 30.870 156.575 31.275 157.085 ;
        RECT 32.415 156.915 32.585 157.165 ;
        RECT 31.445 156.745 32.585 156.915 ;
        RECT 26.285 155.755 26.455 156.365 ;
        RECT 26.625 155.975 26.955 156.410 ;
        RECT 27.175 155.755 29.765 156.525 ;
        RECT 30.395 155.755 30.685 156.480 ;
        RECT 30.870 156.405 32.520 156.575 ;
        RECT 32.755 156.425 33.105 156.995 ;
        RECT 30.915 155.755 31.195 156.235 ;
        RECT 31.365 156.015 31.625 156.405 ;
        RECT 31.800 155.755 32.055 156.235 ;
        RECT 32.225 156.015 32.520 156.405 ;
        RECT 33.275 156.255 33.445 157.165 ;
        RECT 35.200 156.300 35.540 157.130 ;
        RECT 37.020 156.620 37.370 157.870 ;
        RECT 39.135 156.700 39.415 158.135 ;
        RECT 39.585 157.530 40.295 158.305 ;
        RECT 40.465 157.360 40.795 158.135 ;
        RECT 39.645 157.145 40.795 157.360 ;
        RECT 32.700 155.755 32.975 156.235 ;
        RECT 33.145 155.925 33.445 156.255 ;
        RECT 33.615 155.755 38.960 156.300 ;
        RECT 39.135 155.925 39.475 156.700 ;
        RECT 39.645 156.575 39.930 157.145 ;
        RECT 40.115 156.745 40.585 156.975 ;
        RECT 40.990 156.945 41.205 158.060 ;
        RECT 41.385 157.585 41.715 158.305 ;
        RECT 41.495 156.945 41.725 157.285 ;
        RECT 41.895 157.215 43.565 158.305 ;
        RECT 40.755 156.765 41.205 156.945 ;
        RECT 40.755 156.745 41.085 156.765 ;
        RECT 41.395 156.745 41.725 156.945 ;
        RECT 39.645 156.385 40.355 156.575 ;
        RECT 40.055 156.245 40.355 156.385 ;
        RECT 40.545 156.385 41.725 156.575 ;
        RECT 40.545 156.305 40.875 156.385 ;
        RECT 40.055 156.235 40.370 156.245 ;
        RECT 40.055 156.225 40.380 156.235 ;
        RECT 40.055 156.220 40.390 156.225 ;
        RECT 39.645 155.755 39.815 156.215 ;
        RECT 40.055 156.210 40.395 156.220 ;
        RECT 40.055 156.205 40.400 156.210 ;
        RECT 40.055 156.195 40.405 156.205 ;
        RECT 40.055 156.190 40.410 156.195 ;
        RECT 40.055 155.925 40.415 156.190 ;
        RECT 41.045 155.755 41.215 156.215 ;
        RECT 41.385 155.925 41.725 156.385 ;
        RECT 41.895 156.525 42.645 157.045 ;
        RECT 42.815 156.695 43.565 157.215 ;
        RECT 43.735 157.165 44.005 158.135 ;
        RECT 44.215 157.505 44.495 158.305 ;
        RECT 44.665 157.795 46.320 158.085 ;
        RECT 44.730 157.455 46.320 157.625 ;
        RECT 46.505 157.505 46.835 158.305 ;
        RECT 47.015 157.965 48.445 158.135 ;
        RECT 44.730 157.335 44.900 157.455 ;
        RECT 44.175 157.165 44.900 157.335 ;
        RECT 41.895 155.755 43.565 156.525 ;
        RECT 43.735 156.430 43.905 157.165 ;
        RECT 44.175 156.995 44.345 157.165 ;
        RECT 44.075 156.665 44.345 156.995 ;
        RECT 44.515 156.665 44.920 156.995 ;
        RECT 45.090 156.665 45.800 157.285 ;
        RECT 46.000 157.165 46.320 157.455 ;
        RECT 47.015 157.335 47.265 157.965 ;
        RECT 46.495 157.165 47.265 157.335 ;
        RECT 44.175 156.495 44.345 156.665 ;
        RECT 43.735 156.085 44.005 156.430 ;
        RECT 44.175 156.325 45.785 156.495 ;
        RECT 45.970 156.425 46.320 156.995 ;
        RECT 46.495 156.495 46.665 157.165 ;
        RECT 46.835 156.665 47.240 156.995 ;
        RECT 47.455 156.665 47.705 157.795 ;
        RECT 47.905 156.995 48.105 157.795 ;
        RECT 48.275 157.285 48.445 157.965 ;
        RECT 48.615 157.455 48.930 158.305 ;
        RECT 49.105 157.505 49.545 158.135 ;
        RECT 48.275 157.115 49.065 157.285 ;
        RECT 47.905 156.665 48.150 156.995 ;
        RECT 48.335 156.665 48.725 156.945 ;
        RECT 48.895 156.665 49.065 157.115 ;
        RECT 49.235 156.495 49.545 157.505 ;
        RECT 49.725 157.335 50.055 158.120 ;
        RECT 49.725 157.165 50.405 157.335 ;
        RECT 50.585 157.165 50.915 158.305 ;
        RECT 52.100 157.685 52.275 158.135 ;
        RECT 52.445 157.865 52.775 158.305 ;
        RECT 53.080 157.715 53.250 158.135 ;
        RECT 53.485 157.895 54.155 158.305 ;
        RECT 54.370 157.715 54.540 158.135 ;
        RECT 54.740 157.895 55.070 158.305 ;
        RECT 52.100 157.515 52.730 157.685 ;
        RECT 49.715 156.745 50.065 156.995 ;
        RECT 50.235 156.565 50.405 157.165 ;
        RECT 50.575 156.745 50.925 156.995 ;
        RECT 52.015 156.665 52.380 157.345 ;
        RECT 52.560 156.995 52.730 157.515 ;
        RECT 53.080 157.545 55.095 157.715 ;
        RECT 52.560 156.665 52.910 156.995 ;
        RECT 44.195 155.755 44.575 156.155 ;
        RECT 44.745 155.975 44.915 156.325 ;
        RECT 45.085 155.755 45.415 156.155 ;
        RECT 45.615 155.975 45.785 156.325 ;
        RECT 45.985 155.755 46.315 156.255 ;
        RECT 46.495 155.925 46.985 156.495 ;
        RECT 47.155 156.325 48.315 156.495 ;
        RECT 47.155 155.925 47.385 156.325 ;
        RECT 47.555 155.755 47.975 156.155 ;
        RECT 48.145 155.925 48.315 156.325 ;
        RECT 48.485 155.755 48.935 156.495 ;
        RECT 49.105 155.935 49.545 156.495 ;
        RECT 49.735 155.755 49.975 156.565 ;
        RECT 50.145 155.925 50.475 156.565 ;
        RECT 50.645 155.755 50.915 156.565 ;
        RECT 52.560 156.495 52.730 156.665 ;
        RECT 52.100 156.325 52.730 156.495 ;
        RECT 52.100 155.925 52.275 156.325 ;
        RECT 53.080 156.255 53.250 157.545 ;
        RECT 52.445 155.755 52.775 156.135 ;
        RECT 53.020 155.925 53.250 156.255 ;
        RECT 53.450 156.090 53.730 157.365 ;
        RECT 53.955 157.285 54.225 157.365 ;
        RECT 53.915 157.115 54.225 157.285 ;
        RECT 53.955 156.090 54.225 157.115 ;
        RECT 54.415 156.335 54.755 157.365 ;
        RECT 54.925 156.995 55.095 157.545 ;
        RECT 55.265 157.165 55.525 158.135 ;
        RECT 54.925 156.665 55.185 156.995 ;
        RECT 55.355 156.475 55.525 157.165 ;
        RECT 56.155 157.140 56.445 158.305 ;
        RECT 56.675 157.245 57.005 158.090 ;
        RECT 57.175 157.295 57.345 158.305 ;
        RECT 57.515 157.575 57.855 158.135 ;
        RECT 58.085 157.805 58.400 158.305 ;
        RECT 58.580 157.835 59.465 158.005 ;
        RECT 56.615 157.165 57.005 157.245 ;
        RECT 57.515 157.200 58.410 157.575 ;
        RECT 56.615 157.115 56.830 157.165 ;
        RECT 56.615 156.535 56.785 157.115 ;
        RECT 57.515 156.995 57.705 157.200 ;
        RECT 58.580 156.995 58.750 157.835 ;
        RECT 59.690 157.805 59.940 158.135 ;
        RECT 56.955 156.665 57.705 156.995 ;
        RECT 57.875 156.665 58.750 156.995 ;
        RECT 56.615 156.495 56.840 156.535 ;
        RECT 57.505 156.495 57.705 156.665 ;
        RECT 54.685 155.755 55.015 156.135 ;
        RECT 55.185 156.010 55.525 156.475 ;
        RECT 55.185 155.965 55.520 156.010 ;
        RECT 56.155 155.755 56.445 156.480 ;
        RECT 56.615 156.410 56.995 156.495 ;
        RECT 56.665 155.975 56.995 156.410 ;
        RECT 57.165 155.755 57.335 156.365 ;
        RECT 57.505 155.970 57.835 156.495 ;
        RECT 58.095 155.755 58.305 156.285 ;
        RECT 58.580 156.205 58.750 156.665 ;
        RECT 58.920 156.705 59.240 157.665 ;
        RECT 59.410 156.915 59.600 157.635 ;
        RECT 59.770 156.735 59.940 157.805 ;
        RECT 60.110 157.505 60.280 158.305 ;
        RECT 60.450 157.860 61.555 158.030 ;
        RECT 60.450 157.245 60.620 157.860 ;
        RECT 61.765 157.710 62.015 158.135 ;
        RECT 62.185 157.845 62.450 158.305 ;
        RECT 60.790 157.325 61.320 157.690 ;
        RECT 61.765 157.580 62.070 157.710 ;
        RECT 60.110 157.155 60.620 157.245 ;
        RECT 60.110 156.985 60.980 157.155 ;
        RECT 60.110 156.915 60.280 156.985 ;
        RECT 60.400 156.735 60.600 156.765 ;
        RECT 58.920 156.375 59.385 156.705 ;
        RECT 59.770 156.435 60.600 156.735 ;
        RECT 59.770 156.205 59.940 156.435 ;
        RECT 58.580 156.035 59.365 156.205 ;
        RECT 59.535 156.035 59.940 156.205 ;
        RECT 60.120 155.755 60.490 156.255 ;
        RECT 60.810 156.205 60.980 156.985 ;
        RECT 61.150 156.625 61.320 157.325 ;
        RECT 61.490 156.795 61.730 157.390 ;
        RECT 61.150 156.405 61.675 156.625 ;
        RECT 61.900 156.475 62.070 157.580 ;
        RECT 61.845 156.345 62.070 156.475 ;
        RECT 62.240 156.385 62.520 157.335 ;
        RECT 61.845 156.205 62.015 156.345 ;
        RECT 60.810 156.035 61.485 156.205 ;
        RECT 61.680 156.035 62.015 156.205 ;
        RECT 62.185 155.755 62.435 156.215 ;
        RECT 62.690 156.015 62.875 158.135 ;
        RECT 63.045 157.805 63.375 158.305 ;
        RECT 63.545 157.635 63.715 158.135 ;
        RECT 63.050 157.465 63.715 157.635 ;
        RECT 63.050 156.475 63.280 157.465 ;
        RECT 64.435 157.335 64.745 158.135 ;
        RECT 64.915 157.505 65.225 158.305 ;
        RECT 65.395 157.675 65.655 158.135 ;
        RECT 65.825 157.845 66.080 158.305 ;
        RECT 66.255 157.675 66.515 158.135 ;
        RECT 65.395 157.505 66.515 157.675 ;
        RECT 63.450 156.645 63.800 157.295 ;
        RECT 64.435 157.165 65.465 157.335 ;
        RECT 63.050 156.305 63.715 156.475 ;
        RECT 63.045 155.755 63.375 156.135 ;
        RECT 63.545 156.015 63.715 156.305 ;
        RECT 64.435 156.255 64.605 157.165 ;
        RECT 64.775 156.425 65.125 156.995 ;
        RECT 65.295 156.915 65.465 157.165 ;
        RECT 66.255 157.255 66.515 157.505 ;
        RECT 66.685 157.435 66.970 158.305 ;
        RECT 66.255 157.085 67.010 157.255 ;
        RECT 67.205 157.195 67.500 158.305 ;
        RECT 65.295 156.745 66.435 156.915 ;
        RECT 66.605 156.575 67.010 157.085 ;
        RECT 67.680 156.995 67.930 158.130 ;
        RECT 68.100 157.195 68.360 158.305 ;
        RECT 68.530 157.405 68.790 158.130 ;
        RECT 68.960 157.575 69.220 158.305 ;
        RECT 69.390 157.405 69.650 158.130 ;
        RECT 69.820 157.575 70.080 158.305 ;
        RECT 70.250 157.405 70.510 158.130 ;
        RECT 70.680 157.575 70.940 158.305 ;
        RECT 71.110 157.405 71.370 158.130 ;
        RECT 71.540 157.575 71.835 158.305 ;
        RECT 72.255 157.795 72.515 158.305 ;
        RECT 68.530 157.165 71.840 157.405 ;
        RECT 65.360 156.405 67.010 156.575 ;
        RECT 64.435 155.925 64.735 156.255 ;
        RECT 64.905 155.755 65.180 156.235 ;
        RECT 65.360 156.015 65.655 156.405 ;
        RECT 65.825 155.755 66.080 156.235 ;
        RECT 66.255 156.015 66.515 156.405 ;
        RECT 67.195 156.385 67.510 156.995 ;
        RECT 67.680 156.745 70.700 156.995 ;
        RECT 66.685 155.755 66.965 156.235 ;
        RECT 67.255 155.755 67.500 156.215 ;
        RECT 67.680 155.935 67.930 156.745 ;
        RECT 70.870 156.575 71.840 157.165 ;
        RECT 72.255 156.745 72.595 157.625 ;
        RECT 72.765 156.915 72.935 158.135 ;
        RECT 73.175 157.800 73.790 158.305 ;
        RECT 73.175 157.265 73.425 157.630 ;
        RECT 73.595 157.625 73.790 157.800 ;
        RECT 73.960 157.795 74.435 158.135 ;
        RECT 74.605 157.760 74.820 158.305 ;
        RECT 73.595 157.435 73.925 157.625 ;
        RECT 74.145 157.265 74.860 157.560 ;
        RECT 75.030 157.435 75.305 158.135 ;
        RECT 75.565 157.685 75.735 158.115 ;
        RECT 75.905 157.855 76.235 158.305 ;
        RECT 75.565 157.455 76.240 157.685 ;
        RECT 73.175 157.095 74.965 157.265 ;
        RECT 72.765 156.665 73.560 156.915 ;
        RECT 72.765 156.575 73.015 156.665 ;
        RECT 68.530 156.405 71.840 156.575 ;
        RECT 68.100 155.755 68.360 156.280 ;
        RECT 68.530 155.950 68.790 156.405 ;
        RECT 68.960 155.755 69.220 156.235 ;
        RECT 69.390 155.950 69.650 156.405 ;
        RECT 69.820 155.755 70.080 156.235 ;
        RECT 70.250 155.950 70.510 156.405 ;
        RECT 70.680 155.755 70.940 156.235 ;
        RECT 71.110 155.950 71.370 156.405 ;
        RECT 71.540 155.755 71.840 156.235 ;
        RECT 72.255 155.755 72.515 156.575 ;
        RECT 72.685 156.155 73.015 156.575 ;
        RECT 73.730 156.240 73.985 157.095 ;
        RECT 73.195 155.975 73.985 156.240 ;
        RECT 74.155 156.395 74.565 156.915 ;
        RECT 74.735 156.665 74.965 157.095 ;
        RECT 75.135 156.405 75.305 157.435 ;
        RECT 75.535 156.435 75.835 157.285 ;
        RECT 76.005 156.805 76.240 157.455 ;
        RECT 76.410 157.145 76.695 158.090 ;
        RECT 76.875 157.835 77.560 158.305 ;
        RECT 76.870 157.315 77.565 157.625 ;
        RECT 77.740 157.250 78.045 158.035 ;
        RECT 78.350 157.675 78.635 158.135 ;
        RECT 78.805 157.845 79.075 158.305 ;
        RECT 78.350 157.455 79.305 157.675 ;
        RECT 76.410 156.995 77.270 157.145 ;
        RECT 76.410 156.975 77.695 156.995 ;
        RECT 76.005 156.475 76.540 156.805 ;
        RECT 76.710 156.615 77.695 156.975 ;
        RECT 74.155 155.975 74.355 156.395 ;
        RECT 74.545 155.755 74.875 156.215 ;
        RECT 75.045 155.925 75.305 156.405 ;
        RECT 76.005 156.325 76.225 156.475 ;
        RECT 75.480 155.755 75.815 156.260 ;
        RECT 75.985 155.950 76.225 156.325 ;
        RECT 76.710 156.280 76.880 156.615 ;
        RECT 77.870 156.445 78.045 157.250 ;
        RECT 78.235 156.725 78.925 157.285 ;
        RECT 79.095 156.555 79.305 157.455 ;
        RECT 76.505 156.085 76.880 156.280 ;
        RECT 76.505 155.940 76.675 156.085 ;
        RECT 77.240 155.755 77.635 156.250 ;
        RECT 77.805 155.925 78.045 156.445 ;
        RECT 78.350 156.385 79.305 156.555 ;
        RECT 79.475 157.285 79.875 158.135 ;
        RECT 80.065 157.675 80.345 158.135 ;
        RECT 80.865 157.845 81.190 158.305 ;
        RECT 80.065 157.455 81.190 157.675 ;
        RECT 79.475 156.725 80.570 157.285 ;
        RECT 80.740 156.995 81.190 157.455 ;
        RECT 81.360 157.165 81.745 158.135 ;
        RECT 78.350 155.925 78.635 156.385 ;
        RECT 78.805 155.755 79.075 156.215 ;
        RECT 79.475 155.925 79.875 156.725 ;
        RECT 80.740 156.665 81.295 156.995 ;
        RECT 80.740 156.555 81.190 156.665 ;
        RECT 80.065 156.385 81.190 156.555 ;
        RECT 81.465 156.495 81.745 157.165 ;
        RECT 81.915 157.140 82.205 158.305 ;
        RECT 82.435 157.245 82.765 158.090 ;
        RECT 82.935 157.295 83.105 158.305 ;
        RECT 83.275 157.575 83.615 158.135 ;
        RECT 83.845 157.805 84.160 158.305 ;
        RECT 84.340 157.835 85.225 158.005 ;
        RECT 82.375 157.165 82.765 157.245 ;
        RECT 83.275 157.200 84.170 157.575 ;
        RECT 80.065 155.925 80.345 156.385 ;
        RECT 80.865 155.755 81.190 156.215 ;
        RECT 81.360 155.925 81.745 156.495 ;
        RECT 82.375 157.115 82.590 157.165 ;
        RECT 82.375 156.535 82.545 157.115 ;
        RECT 83.275 156.995 83.465 157.200 ;
        RECT 84.340 156.995 84.510 157.835 ;
        RECT 85.450 157.805 85.700 158.135 ;
        RECT 82.715 156.665 83.465 156.995 ;
        RECT 83.635 156.665 84.510 156.995 ;
        RECT 82.375 156.495 82.600 156.535 ;
        RECT 83.265 156.495 83.465 156.665 ;
        RECT 81.915 155.755 82.205 156.480 ;
        RECT 82.375 156.410 82.755 156.495 ;
        RECT 82.425 155.975 82.755 156.410 ;
        RECT 82.925 155.755 83.095 156.365 ;
        RECT 83.265 155.970 83.595 156.495 ;
        RECT 83.855 155.755 84.065 156.285 ;
        RECT 84.340 156.205 84.510 156.665 ;
        RECT 84.680 156.705 85.000 157.665 ;
        RECT 85.170 156.915 85.360 157.635 ;
        RECT 85.530 156.735 85.700 157.805 ;
        RECT 85.870 157.505 86.040 158.305 ;
        RECT 86.210 157.860 87.315 158.030 ;
        RECT 86.210 157.245 86.380 157.860 ;
        RECT 87.525 157.710 87.775 158.135 ;
        RECT 87.945 157.845 88.210 158.305 ;
        RECT 86.550 157.325 87.080 157.690 ;
        RECT 87.525 157.580 87.830 157.710 ;
        RECT 85.870 157.155 86.380 157.245 ;
        RECT 85.870 156.985 86.740 157.155 ;
        RECT 85.870 156.915 86.040 156.985 ;
        RECT 86.160 156.735 86.360 156.765 ;
        RECT 84.680 156.375 85.145 156.705 ;
        RECT 85.530 156.435 86.360 156.735 ;
        RECT 85.530 156.205 85.700 156.435 ;
        RECT 84.340 156.035 85.125 156.205 ;
        RECT 85.295 156.035 85.700 156.205 ;
        RECT 85.880 155.755 86.250 156.255 ;
        RECT 86.570 156.205 86.740 156.985 ;
        RECT 86.910 156.625 87.080 157.325 ;
        RECT 87.250 156.795 87.490 157.390 ;
        RECT 86.910 156.405 87.435 156.625 ;
        RECT 87.660 156.475 87.830 157.580 ;
        RECT 87.605 156.345 87.830 156.475 ;
        RECT 88.000 156.385 88.280 157.335 ;
        RECT 87.605 156.205 87.775 156.345 ;
        RECT 86.570 156.035 87.245 156.205 ;
        RECT 87.440 156.035 87.775 156.205 ;
        RECT 87.945 155.755 88.195 156.215 ;
        RECT 88.450 156.015 88.635 158.135 ;
        RECT 88.805 157.805 89.135 158.305 ;
        RECT 89.305 157.635 89.475 158.135 ;
        RECT 88.810 157.465 89.475 157.635 ;
        RECT 88.810 156.475 89.040 157.465 ;
        RECT 89.210 156.645 89.560 157.295 ;
        RECT 89.740 157.165 90.075 158.135 ;
        RECT 90.245 157.165 90.415 158.305 ;
        RECT 90.585 157.965 92.615 158.135 ;
        RECT 89.740 156.495 89.910 157.165 ;
        RECT 90.585 156.995 90.755 157.965 ;
        RECT 90.080 156.665 90.335 156.995 ;
        RECT 90.560 156.665 90.755 156.995 ;
        RECT 90.925 157.625 92.050 157.795 ;
        RECT 90.165 156.495 90.335 156.665 ;
        RECT 90.925 156.495 91.095 157.625 ;
        RECT 88.810 156.305 89.475 156.475 ;
        RECT 88.805 155.755 89.135 156.135 ;
        RECT 89.305 156.015 89.475 156.305 ;
        RECT 89.740 155.925 89.995 156.495 ;
        RECT 90.165 156.325 91.095 156.495 ;
        RECT 91.265 157.285 92.275 157.455 ;
        RECT 91.265 156.485 91.435 157.285 ;
        RECT 90.920 156.290 91.095 156.325 ;
        RECT 90.165 155.755 90.495 156.155 ;
        RECT 90.920 155.925 91.450 156.290 ;
        RECT 91.640 156.265 91.915 157.085 ;
        RECT 91.635 156.095 91.915 156.265 ;
        RECT 91.640 155.925 91.915 156.095 ;
        RECT 92.085 155.925 92.275 157.285 ;
        RECT 92.445 157.300 92.615 157.965 ;
        RECT 92.785 157.545 92.955 158.305 ;
        RECT 93.190 157.545 93.705 157.955 ;
        RECT 92.445 157.110 93.195 157.300 ;
        RECT 93.365 156.735 93.705 157.545 ;
        RECT 93.875 157.215 95.545 158.305 ;
        RECT 92.475 156.565 93.705 156.735 ;
        RECT 92.455 155.755 92.965 156.290 ;
        RECT 93.185 155.960 93.430 156.565 ;
        RECT 93.875 156.525 94.625 157.045 ;
        RECT 94.795 156.695 95.545 157.215 ;
        RECT 96.185 157.195 96.480 158.305 ;
        RECT 96.660 156.995 96.910 158.130 ;
        RECT 97.080 157.195 97.340 158.305 ;
        RECT 97.510 157.405 97.770 158.130 ;
        RECT 97.940 157.575 98.200 158.305 ;
        RECT 98.370 157.405 98.630 158.130 ;
        RECT 98.800 157.575 99.060 158.305 ;
        RECT 99.230 157.405 99.490 158.130 ;
        RECT 99.660 157.575 99.920 158.305 ;
        RECT 100.090 157.405 100.350 158.130 ;
        RECT 100.520 157.575 100.815 158.305 ;
        RECT 97.510 157.165 100.820 157.405 ;
        RECT 93.875 155.755 95.545 156.525 ;
        RECT 96.175 156.385 96.490 156.995 ;
        RECT 96.660 156.745 99.680 156.995 ;
        RECT 96.235 155.755 96.480 156.215 ;
        RECT 96.660 155.935 96.910 156.745 ;
        RECT 99.850 156.575 100.820 157.165 ;
        RECT 97.510 156.405 100.820 156.575 ;
        RECT 101.240 157.165 101.575 158.135 ;
        RECT 101.745 157.165 101.915 158.305 ;
        RECT 102.085 157.965 104.115 158.135 ;
        RECT 101.240 156.495 101.410 157.165 ;
        RECT 102.085 156.995 102.255 157.965 ;
        RECT 101.580 156.665 101.835 156.995 ;
        RECT 102.060 156.665 102.255 156.995 ;
        RECT 102.425 157.625 103.550 157.795 ;
        RECT 101.665 156.495 101.835 156.665 ;
        RECT 102.425 156.495 102.595 157.625 ;
        RECT 97.080 155.755 97.340 156.280 ;
        RECT 97.510 155.950 97.770 156.405 ;
        RECT 97.940 155.755 98.200 156.235 ;
        RECT 98.370 155.950 98.630 156.405 ;
        RECT 98.800 155.755 99.060 156.235 ;
        RECT 99.230 155.950 99.490 156.405 ;
        RECT 99.660 155.755 99.920 156.235 ;
        RECT 100.090 155.950 100.350 156.405 ;
        RECT 100.520 155.755 100.820 156.235 ;
        RECT 101.240 155.925 101.495 156.495 ;
        RECT 101.665 156.325 102.595 156.495 ;
        RECT 102.765 157.285 103.775 157.455 ;
        RECT 102.765 156.485 102.935 157.285 ;
        RECT 102.420 156.290 102.595 156.325 ;
        RECT 101.665 155.755 101.995 156.155 ;
        RECT 102.420 155.925 102.950 156.290 ;
        RECT 103.140 156.265 103.415 157.085 ;
        RECT 103.135 156.095 103.415 156.265 ;
        RECT 103.140 155.925 103.415 156.095 ;
        RECT 103.585 155.925 103.775 157.285 ;
        RECT 103.945 157.300 104.115 157.965 ;
        RECT 104.285 157.545 104.455 158.305 ;
        RECT 104.690 157.545 105.205 157.955 ;
        RECT 103.945 157.110 104.695 157.300 ;
        RECT 104.865 156.735 105.205 157.545 ;
        RECT 105.375 157.215 107.045 158.305 ;
        RECT 103.975 156.565 105.205 156.735 ;
        RECT 103.955 155.755 104.465 156.290 ;
        RECT 104.685 155.960 104.930 156.565 ;
        RECT 105.375 156.525 106.125 157.045 ;
        RECT 106.295 156.695 107.045 157.215 ;
        RECT 107.675 157.140 107.965 158.305 ;
        RECT 108.140 157.165 108.460 158.305 ;
        RECT 108.640 156.995 108.835 158.045 ;
        RECT 109.015 157.455 109.345 158.135 ;
        RECT 109.545 157.505 109.800 158.305 ;
        RECT 109.015 157.175 109.365 157.455 ;
        RECT 108.200 156.945 108.460 156.995 ;
        RECT 108.195 156.775 108.460 156.945 ;
        RECT 108.200 156.665 108.460 156.775 ;
        RECT 108.640 156.665 109.025 156.995 ;
        RECT 109.195 156.795 109.365 157.175 ;
        RECT 109.555 156.965 109.800 157.325 ;
        RECT 110.475 157.165 110.705 158.305 ;
        RECT 110.875 157.155 111.205 158.135 ;
        RECT 111.375 157.165 111.585 158.305 ;
        RECT 111.815 157.215 115.325 158.305 ;
        RECT 109.195 156.625 109.715 156.795 ;
        RECT 110.455 156.745 110.785 156.995 ;
        RECT 105.375 155.755 107.045 156.525 ;
        RECT 107.675 155.755 107.965 156.480 ;
        RECT 108.140 156.285 109.355 156.455 ;
        RECT 108.140 155.935 108.430 156.285 ;
        RECT 108.625 155.755 108.955 156.115 ;
        RECT 109.125 155.980 109.355 156.285 ;
        RECT 109.545 156.265 109.715 156.625 ;
        RECT 109.545 156.095 109.745 156.265 ;
        RECT 109.545 156.060 109.715 156.095 ;
        RECT 110.475 155.755 110.705 156.575 ;
        RECT 110.955 156.555 111.205 157.155 ;
        RECT 110.875 155.925 111.205 156.555 ;
        RECT 111.375 155.755 111.585 156.575 ;
        RECT 111.815 156.525 113.465 157.045 ;
        RECT 113.635 156.695 115.325 157.215 ;
        RECT 116.110 157.295 116.410 158.135 ;
        RECT 116.605 157.465 116.855 158.305 ;
        RECT 117.445 157.715 118.250 158.135 ;
        RECT 117.025 157.545 118.590 157.715 ;
        RECT 117.025 157.295 117.195 157.545 ;
        RECT 116.110 157.125 117.195 157.295 ;
        RECT 115.955 156.665 116.285 156.955 ;
        RECT 111.815 155.755 115.325 156.525 ;
        RECT 116.455 156.495 116.625 157.125 ;
        RECT 117.365 156.995 117.685 157.375 ;
        RECT 117.875 157.285 118.250 157.375 ;
        RECT 117.855 157.115 118.250 157.285 ;
        RECT 118.420 157.295 118.590 157.545 ;
        RECT 118.760 157.465 119.090 158.305 ;
        RECT 119.260 157.545 119.925 158.135 ;
        RECT 118.420 157.125 119.340 157.295 ;
        RECT 116.795 156.745 117.125 156.955 ;
        RECT 117.305 156.745 117.685 156.995 ;
        RECT 117.875 156.955 118.250 157.115 ;
        RECT 119.170 156.955 119.340 157.125 ;
        RECT 117.875 156.745 118.360 156.955 ;
        RECT 118.550 156.745 119.000 156.955 ;
        RECT 119.170 156.745 119.505 156.955 ;
        RECT 119.675 156.575 119.925 157.545 ;
        RECT 120.100 157.165 120.355 158.305 ;
        RECT 120.525 157.335 120.855 158.135 ;
        RECT 121.025 157.505 121.255 158.305 ;
        RECT 121.425 157.335 121.755 158.135 ;
        RECT 120.525 157.165 121.755 157.335 ;
        RECT 122.405 157.285 122.735 158.135 ;
        RECT 122.905 157.455 123.075 158.305 ;
        RECT 123.245 157.285 123.575 158.135 ;
        RECT 123.745 157.455 123.915 158.305 ;
        RECT 124.085 157.285 124.415 158.135 ;
        RECT 124.585 157.505 124.755 158.305 ;
        RECT 124.925 157.285 125.255 158.135 ;
        RECT 125.425 157.505 125.595 158.305 ;
        RECT 125.765 157.285 126.095 158.135 ;
        RECT 126.265 157.505 126.435 158.305 ;
        RECT 126.605 157.285 126.935 158.135 ;
        RECT 127.105 157.505 127.275 158.305 ;
        RECT 127.445 157.285 127.775 158.135 ;
        RECT 127.945 157.505 128.115 158.305 ;
        RECT 128.285 157.285 128.615 158.135 ;
        RECT 128.785 157.505 128.955 158.305 ;
        RECT 129.125 157.285 129.455 158.135 ;
        RECT 129.625 157.505 129.795 158.305 ;
        RECT 129.965 157.285 130.295 158.135 ;
        RECT 130.465 157.505 130.635 158.305 ;
        RECT 130.805 157.285 131.135 158.135 ;
        RECT 131.305 157.505 131.475 158.305 ;
        RECT 131.645 157.285 131.975 158.135 ;
        RECT 132.145 157.505 132.315 158.305 ;
        RECT 132.485 157.285 132.815 158.135 ;
        RECT 132.985 157.505 133.155 158.305 ;
        RECT 116.115 156.315 116.625 156.495 ;
        RECT 117.030 156.405 118.730 156.575 ;
        RECT 117.030 156.315 117.415 156.405 ;
        RECT 116.115 155.925 116.445 156.315 ;
        RECT 116.615 155.975 117.800 156.145 ;
        RECT 118.060 155.755 118.230 156.225 ;
        RECT 118.400 155.940 118.730 156.405 ;
        RECT 118.900 155.755 119.070 156.575 ;
        RECT 119.240 155.935 119.925 156.575 ;
        RECT 120.120 156.415 120.340 156.995 ;
        RECT 120.525 156.265 120.705 157.165 ;
        RECT 122.405 157.115 123.915 157.285 ;
        RECT 124.085 157.115 126.435 157.285 ;
        RECT 126.605 157.115 133.265 157.285 ;
        RECT 133.435 157.140 133.725 158.305 ;
        RECT 133.900 157.165 134.235 158.135 ;
        RECT 134.405 157.165 134.575 158.305 ;
        RECT 134.745 157.965 136.775 158.135 ;
        RECT 120.875 156.435 121.250 156.995 ;
        RECT 121.455 156.665 121.765 156.995 ;
        RECT 123.745 156.945 123.915 157.115 ;
        RECT 126.260 156.945 126.435 157.115 ;
        RECT 122.400 156.745 123.575 156.945 ;
        RECT 123.745 156.745 126.055 156.945 ;
        RECT 126.260 156.745 132.820 156.945 ;
        RECT 123.745 156.575 123.915 156.745 ;
        RECT 126.260 156.575 126.435 156.745 ;
        RECT 132.990 156.575 133.265 157.115 ;
        RECT 121.425 156.265 121.755 156.495 ;
        RECT 120.100 155.755 120.355 156.245 ;
        RECT 120.525 155.925 121.755 156.265 ;
        RECT 122.405 156.405 123.915 156.575 ;
        RECT 124.085 156.405 126.435 156.575 ;
        RECT 126.605 156.405 133.265 156.575 ;
        RECT 133.900 156.495 134.070 157.165 ;
        RECT 134.745 156.995 134.915 157.965 ;
        RECT 134.240 156.665 134.495 156.995 ;
        RECT 134.720 156.665 134.915 156.995 ;
        RECT 135.085 157.625 136.210 157.795 ;
        RECT 134.325 156.495 134.495 156.665 ;
        RECT 135.085 156.495 135.255 157.625 ;
        RECT 122.405 155.930 122.735 156.405 ;
        RECT 122.905 155.755 123.075 156.235 ;
        RECT 123.245 155.930 123.575 156.405 ;
        RECT 123.745 155.755 123.915 156.235 ;
        RECT 124.085 155.930 124.415 156.405 ;
        RECT 124.585 155.755 124.755 156.235 ;
        RECT 124.925 155.930 125.255 156.405 ;
        RECT 125.425 155.755 125.595 156.235 ;
        RECT 125.765 155.930 126.095 156.405 ;
        RECT 126.265 155.755 126.435 156.235 ;
        RECT 126.605 155.930 126.935 156.405 ;
        RECT 126.605 155.925 126.855 155.930 ;
        RECT 127.105 155.755 127.275 156.235 ;
        RECT 127.445 155.930 127.775 156.405 ;
        RECT 127.525 155.925 127.695 155.930 ;
        RECT 127.945 155.755 128.115 156.235 ;
        RECT 128.285 155.930 128.615 156.405 ;
        RECT 128.365 155.925 128.535 155.930 ;
        RECT 128.785 155.755 128.955 156.235 ;
        RECT 129.125 155.930 129.455 156.405 ;
        RECT 129.625 155.755 129.795 156.235 ;
        RECT 129.965 155.930 130.295 156.405 ;
        RECT 130.465 155.755 130.635 156.235 ;
        RECT 130.805 155.930 131.135 156.405 ;
        RECT 131.305 155.755 131.475 156.235 ;
        RECT 131.645 155.930 131.975 156.405 ;
        RECT 132.145 155.755 132.315 156.235 ;
        RECT 132.485 155.930 132.815 156.405 ;
        RECT 132.985 155.755 133.155 156.235 ;
        RECT 133.435 155.755 133.725 156.480 ;
        RECT 133.900 155.925 134.155 156.495 ;
        RECT 134.325 156.325 135.255 156.495 ;
        RECT 135.425 157.285 136.435 157.455 ;
        RECT 135.425 156.485 135.595 157.285 ;
        RECT 135.800 156.605 136.075 157.085 ;
        RECT 135.795 156.435 136.075 156.605 ;
        RECT 135.080 156.290 135.255 156.325 ;
        RECT 134.325 155.755 134.655 156.155 ;
        RECT 135.080 155.925 135.610 156.290 ;
        RECT 135.800 155.925 136.075 156.435 ;
        RECT 136.245 155.925 136.435 157.285 ;
        RECT 136.605 157.300 136.775 157.965 ;
        RECT 136.945 157.545 137.115 158.305 ;
        RECT 137.350 157.545 137.865 157.955 ;
        RECT 136.605 157.110 137.355 157.300 ;
        RECT 137.525 156.735 137.865 157.545 ;
        RECT 136.635 156.565 137.865 156.735 ;
        RECT 138.035 157.165 138.420 158.135 ;
        RECT 138.590 157.845 138.915 158.305 ;
        RECT 139.435 157.675 139.715 158.135 ;
        RECT 138.590 157.455 139.715 157.675 ;
        RECT 136.615 155.755 137.125 156.290 ;
        RECT 137.345 155.960 137.590 156.565 ;
        RECT 138.035 156.495 138.315 157.165 ;
        RECT 138.590 156.995 139.040 157.455 ;
        RECT 139.905 157.285 140.305 158.135 ;
        RECT 140.705 157.845 140.975 158.305 ;
        RECT 141.145 157.675 141.430 158.135 ;
        RECT 138.485 156.665 139.040 156.995 ;
        RECT 139.210 156.725 140.305 157.285 ;
        RECT 138.590 156.555 139.040 156.665 ;
        RECT 138.035 155.925 138.420 156.495 ;
        RECT 138.590 156.385 139.715 156.555 ;
        RECT 138.590 155.755 138.915 156.215 ;
        RECT 139.435 155.925 139.715 156.385 ;
        RECT 139.905 155.925 140.305 156.725 ;
        RECT 140.475 157.455 141.430 157.675 ;
        RECT 140.475 156.555 140.685 157.455 ;
        RECT 140.855 156.725 141.545 157.285 ;
        RECT 141.715 157.215 142.925 158.305 ;
        RECT 141.715 156.675 142.235 157.215 ;
        RECT 140.475 156.385 141.430 156.555 ;
        RECT 142.405 156.505 142.925 157.045 ;
        RECT 140.705 155.755 140.975 156.215 ;
        RECT 141.145 155.925 141.430 156.385 ;
        RECT 141.715 155.755 142.925 156.505 ;
        RECT 17.430 155.585 143.010 155.755 ;
        RECT 17.515 154.835 18.725 155.585 ;
        RECT 18.895 155.040 24.240 155.585 ;
        RECT 17.515 154.295 18.035 154.835 ;
        RECT 18.205 154.125 18.725 154.665 ;
        RECT 20.480 154.210 20.820 155.040 ;
        RECT 24.415 154.815 26.085 155.585 ;
        RECT 26.765 155.195 27.095 155.585 ;
        RECT 27.265 155.015 27.435 155.335 ;
        RECT 27.605 155.195 27.935 155.585 ;
        RECT 28.350 155.185 29.305 155.355 ;
        RECT 26.715 154.845 28.965 155.015 ;
        RECT 17.515 153.035 18.725 154.125 ;
        RECT 22.300 153.470 22.650 154.720 ;
        RECT 24.415 154.295 25.165 154.815 ;
        RECT 25.335 154.125 26.085 154.645 ;
        RECT 18.895 153.035 24.240 153.470 ;
        RECT 24.415 153.035 26.085 154.125 ;
        RECT 26.715 153.885 26.885 154.845 ;
        RECT 27.055 154.225 27.300 154.675 ;
        RECT 27.470 154.395 28.020 154.595 ;
        RECT 28.190 154.425 28.565 154.595 ;
        RECT 28.190 154.225 28.360 154.425 ;
        RECT 28.735 154.345 28.965 154.845 ;
        RECT 27.055 154.055 28.360 154.225 ;
        RECT 29.135 154.305 29.305 155.185 ;
        RECT 29.475 154.750 29.765 155.585 ;
        RECT 29.935 154.815 32.525 155.585 ;
        RECT 33.160 154.935 33.430 155.145 ;
        RECT 33.650 155.125 33.980 155.585 ;
        RECT 34.490 155.125 35.240 155.415 ;
        RECT 29.135 154.135 29.765 154.305 ;
        RECT 29.935 154.295 31.145 154.815 ;
        RECT 33.160 154.765 34.495 154.935 ;
        RECT 26.715 153.205 27.095 153.885 ;
        RECT 27.685 153.035 27.855 153.885 ;
        RECT 28.025 153.715 29.265 153.885 ;
        RECT 28.025 153.205 28.355 153.715 ;
        RECT 28.525 153.035 28.695 153.545 ;
        RECT 28.865 153.205 29.265 153.715 ;
        RECT 29.445 153.205 29.765 154.135 ;
        RECT 31.315 154.125 32.525 154.645 ;
        RECT 34.325 154.595 34.495 154.765 ;
        RECT 33.160 154.355 33.510 154.595 ;
        RECT 33.680 154.355 34.155 154.595 ;
        RECT 34.325 154.345 34.700 154.595 ;
        RECT 34.325 154.175 34.495 154.345 ;
        RECT 29.935 153.035 32.525 154.125 ;
        RECT 33.160 154.005 34.495 154.175 ;
        RECT 33.160 153.845 33.440 154.005 ;
        RECT 34.870 153.835 35.240 155.125 ;
        RECT 35.455 155.040 40.800 155.585 ;
        RECT 37.040 154.210 37.380 155.040 ;
        RECT 40.975 154.815 42.645 155.585 ;
        RECT 43.275 154.860 43.565 155.585 ;
        RECT 33.650 153.035 33.900 153.835 ;
        RECT 34.070 153.665 35.240 153.835 ;
        RECT 34.070 153.205 34.400 153.665 ;
        RECT 34.570 153.035 34.785 153.495 ;
        RECT 38.860 153.470 39.210 154.720 ;
        RECT 40.975 154.295 41.725 154.815 ;
        RECT 43.775 154.765 44.005 155.585 ;
        RECT 44.175 154.785 44.505 155.415 ;
        RECT 41.895 154.125 42.645 154.645 ;
        RECT 43.755 154.345 44.085 154.595 ;
        RECT 35.455 153.035 40.800 153.470 ;
        RECT 40.975 153.035 42.645 154.125 ;
        RECT 43.275 153.035 43.565 154.200 ;
        RECT 44.255 154.185 44.505 154.785 ;
        RECT 44.675 154.765 44.885 155.585 ;
        RECT 45.575 154.845 46.040 155.390 ;
        RECT 43.775 153.035 44.005 154.175 ;
        RECT 44.175 153.205 44.505 154.185 ;
        RECT 44.675 153.035 44.885 154.175 ;
        RECT 45.575 153.885 45.745 154.845 ;
        RECT 46.545 154.765 46.715 155.585 ;
        RECT 46.885 154.935 47.215 155.415 ;
        RECT 47.385 155.195 47.735 155.585 ;
        RECT 47.905 155.015 48.135 155.415 ;
        RECT 47.625 154.935 48.135 155.015 ;
        RECT 46.885 154.845 48.135 154.935 ;
        RECT 48.305 154.845 48.625 155.325 ;
        RECT 48.805 155.085 49.135 155.585 ;
        RECT 49.335 155.015 49.505 155.365 ;
        RECT 49.705 155.185 50.035 155.585 ;
        RECT 50.205 155.015 50.375 155.365 ;
        RECT 50.545 155.185 50.925 155.585 ;
        RECT 46.885 154.765 47.795 154.845 ;
        RECT 45.915 154.225 46.160 154.675 ;
        RECT 46.420 154.395 47.115 154.595 ;
        RECT 47.285 154.425 47.885 154.595 ;
        RECT 47.285 154.225 47.455 154.425 ;
        RECT 48.115 154.255 48.285 154.675 ;
        RECT 45.915 154.055 47.455 154.225 ;
        RECT 47.625 154.085 48.285 154.255 ;
        RECT 47.625 153.885 47.795 154.085 ;
        RECT 48.455 153.915 48.625 154.845 ;
        RECT 48.800 154.345 49.150 154.915 ;
        RECT 49.335 154.845 50.945 155.015 ;
        RECT 51.115 154.910 51.385 155.255 ;
        RECT 50.775 154.675 50.945 154.845 ;
        RECT 45.575 153.715 47.795 153.885 ;
        RECT 47.965 153.715 48.625 153.915 ;
        RECT 48.800 153.885 49.120 154.175 ;
        RECT 49.320 154.055 50.030 154.675 ;
        RECT 50.200 154.345 50.605 154.675 ;
        RECT 50.775 154.345 51.045 154.675 ;
        RECT 50.775 154.175 50.945 154.345 ;
        RECT 51.215 154.175 51.385 154.910 ;
        RECT 51.555 154.815 53.225 155.585 ;
        RECT 53.395 154.845 53.715 155.325 ;
        RECT 53.885 155.015 54.115 155.415 ;
        RECT 54.285 155.195 54.635 155.585 ;
        RECT 53.885 154.935 54.395 155.015 ;
        RECT 54.805 154.935 55.135 155.415 ;
        RECT 53.885 154.845 55.135 154.935 ;
        RECT 51.555 154.295 52.305 154.815 ;
        RECT 50.220 154.005 50.945 154.175 ;
        RECT 50.220 153.885 50.390 154.005 ;
        RECT 48.800 153.715 50.390 153.885 ;
        RECT 45.575 153.035 45.875 153.545 ;
        RECT 46.045 153.205 46.375 153.715 ;
        RECT 47.965 153.545 48.135 153.715 ;
        RECT 46.545 153.035 47.175 153.545 ;
        RECT 47.755 153.375 48.135 153.545 ;
        RECT 48.305 153.035 48.605 153.545 ;
        RECT 48.800 153.255 50.455 153.545 ;
        RECT 50.625 153.035 50.905 153.835 ;
        RECT 51.115 153.205 51.385 154.175 ;
        RECT 52.475 154.125 53.225 154.645 ;
        RECT 51.555 153.035 53.225 154.125 ;
        RECT 53.395 153.915 53.565 154.845 ;
        RECT 54.225 154.765 55.135 154.845 ;
        RECT 55.305 154.765 55.475 155.585 ;
        RECT 55.980 154.845 56.445 155.390 ;
        RECT 56.615 155.040 61.960 155.585 ;
        RECT 62.135 155.040 67.480 155.585 ;
        RECT 53.735 154.255 53.905 154.675 ;
        RECT 54.135 154.425 54.735 154.595 ;
        RECT 53.735 154.085 54.395 154.255 ;
        RECT 53.395 153.715 54.055 153.915 ;
        RECT 54.225 153.885 54.395 154.085 ;
        RECT 54.565 154.225 54.735 154.425 ;
        RECT 54.905 154.395 55.600 154.595 ;
        RECT 55.860 154.225 56.105 154.675 ;
        RECT 54.565 154.055 56.105 154.225 ;
        RECT 56.275 153.885 56.445 154.845 ;
        RECT 58.200 154.210 58.540 155.040 ;
        RECT 54.225 153.715 56.445 153.885 ;
        RECT 53.885 153.545 54.055 153.715 ;
        RECT 53.415 153.035 53.715 153.545 ;
        RECT 53.885 153.375 54.265 153.545 ;
        RECT 54.845 153.035 55.475 153.545 ;
        RECT 55.645 153.205 55.975 153.715 ;
        RECT 56.145 153.035 56.445 153.545 ;
        RECT 60.020 153.470 60.370 154.720 ;
        RECT 63.720 154.210 64.060 155.040 ;
        RECT 67.655 154.835 68.865 155.585 ;
        RECT 69.035 154.860 69.325 155.585 ;
        RECT 69.585 155.035 69.755 155.325 ;
        RECT 69.925 155.205 70.255 155.585 ;
        RECT 69.585 154.865 70.250 155.035 ;
        RECT 65.540 153.470 65.890 154.720 ;
        RECT 67.655 154.295 68.175 154.835 ;
        RECT 68.345 154.125 68.865 154.665 ;
        RECT 56.615 153.035 61.960 153.470 ;
        RECT 62.135 153.035 67.480 153.470 ;
        RECT 67.655 153.035 68.865 154.125 ;
        RECT 69.035 153.035 69.325 154.200 ;
        RECT 69.500 154.045 69.850 154.695 ;
        RECT 70.020 153.875 70.250 154.865 ;
        RECT 69.585 153.705 70.250 153.875 ;
        RECT 69.585 153.205 69.755 153.705 ;
        RECT 69.925 153.035 70.255 153.535 ;
        RECT 70.425 153.205 70.610 155.325 ;
        RECT 70.865 155.125 71.115 155.585 ;
        RECT 71.285 155.135 71.620 155.305 ;
        RECT 71.815 155.135 72.490 155.305 ;
        RECT 71.285 154.995 71.455 155.135 ;
        RECT 70.780 154.005 71.060 154.955 ;
        RECT 71.230 154.865 71.455 154.995 ;
        RECT 71.230 153.760 71.400 154.865 ;
        RECT 71.625 154.715 72.150 154.935 ;
        RECT 71.570 153.950 71.810 154.545 ;
        RECT 71.980 154.015 72.150 154.715 ;
        RECT 72.320 154.355 72.490 155.135 ;
        RECT 72.810 155.085 73.180 155.585 ;
        RECT 73.360 155.135 73.765 155.305 ;
        RECT 73.935 155.135 74.720 155.305 ;
        RECT 73.360 154.905 73.530 155.135 ;
        RECT 72.700 154.605 73.530 154.905 ;
        RECT 73.915 154.635 74.380 154.965 ;
        RECT 72.700 154.575 72.900 154.605 ;
        RECT 73.020 154.355 73.190 154.425 ;
        RECT 72.320 154.185 73.190 154.355 ;
        RECT 72.680 154.095 73.190 154.185 ;
        RECT 71.230 153.630 71.535 153.760 ;
        RECT 71.980 153.650 72.510 154.015 ;
        RECT 70.850 153.035 71.115 153.495 ;
        RECT 71.285 153.205 71.535 153.630 ;
        RECT 72.680 153.480 72.850 154.095 ;
        RECT 71.745 153.310 72.850 153.480 ;
        RECT 73.020 153.035 73.190 153.835 ;
        RECT 73.360 153.535 73.530 154.605 ;
        RECT 73.700 153.705 73.890 154.425 ;
        RECT 74.060 153.675 74.380 154.635 ;
        RECT 74.550 154.675 74.720 155.135 ;
        RECT 74.995 155.055 75.205 155.585 ;
        RECT 75.465 154.845 75.795 155.370 ;
        RECT 75.965 154.975 76.135 155.585 ;
        RECT 76.305 154.930 76.635 155.365 ;
        RECT 76.305 154.845 76.685 154.930 ;
        RECT 75.595 154.675 75.795 154.845 ;
        RECT 76.460 154.805 76.685 154.845 ;
        RECT 74.550 154.345 75.425 154.675 ;
        RECT 75.595 154.345 76.345 154.675 ;
        RECT 73.360 153.205 73.610 153.535 ;
        RECT 74.550 153.505 74.720 154.345 ;
        RECT 75.595 154.140 75.785 154.345 ;
        RECT 76.515 154.225 76.685 154.805 ;
        RECT 76.470 154.175 76.685 154.225 ;
        RECT 74.890 153.765 75.785 154.140 ;
        RECT 76.295 154.095 76.685 154.175 ;
        RECT 76.855 154.845 77.240 155.415 ;
        RECT 77.410 155.125 77.735 155.585 ;
        RECT 78.255 154.955 78.535 155.415 ;
        RECT 76.855 154.175 77.135 154.845 ;
        RECT 77.410 154.785 78.535 154.955 ;
        RECT 77.410 154.675 77.860 154.785 ;
        RECT 77.305 154.345 77.860 154.675 ;
        RECT 78.725 154.615 79.125 155.415 ;
        RECT 79.525 155.125 79.795 155.585 ;
        RECT 79.965 154.955 80.250 155.415 ;
        RECT 73.835 153.335 74.720 153.505 ;
        RECT 74.900 153.035 75.215 153.535 ;
        RECT 75.445 153.205 75.785 153.765 ;
        RECT 75.955 153.035 76.125 154.045 ;
        RECT 76.295 153.250 76.625 154.095 ;
        RECT 76.855 153.205 77.240 154.175 ;
        RECT 77.410 153.885 77.860 154.345 ;
        RECT 78.030 154.055 79.125 154.615 ;
        RECT 77.410 153.665 78.535 153.885 ;
        RECT 77.410 153.035 77.735 153.495 ;
        RECT 78.255 153.205 78.535 153.665 ;
        RECT 78.725 153.205 79.125 154.055 ;
        RECT 79.295 154.785 80.250 154.955 ;
        RECT 80.535 154.815 82.205 155.585 ;
        RECT 82.425 154.930 82.755 155.365 ;
        RECT 82.925 154.975 83.095 155.585 ;
        RECT 82.375 154.845 82.755 154.930 ;
        RECT 83.265 154.845 83.595 155.370 ;
        RECT 83.855 155.055 84.065 155.585 ;
        RECT 84.340 155.135 85.125 155.305 ;
        RECT 85.295 155.135 85.700 155.305 ;
        RECT 79.295 153.885 79.505 154.785 ;
        RECT 79.675 154.055 80.365 154.615 ;
        RECT 80.535 154.295 81.285 154.815 ;
        RECT 82.375 154.805 82.600 154.845 ;
        RECT 81.455 154.125 82.205 154.645 ;
        RECT 79.295 153.665 80.250 153.885 ;
        RECT 79.525 153.035 79.795 153.495 ;
        RECT 79.965 153.205 80.250 153.665 ;
        RECT 80.535 153.035 82.205 154.125 ;
        RECT 82.375 154.225 82.545 154.805 ;
        RECT 83.265 154.675 83.465 154.845 ;
        RECT 84.340 154.675 84.510 155.135 ;
        RECT 82.715 154.345 83.465 154.675 ;
        RECT 83.635 154.345 84.510 154.675 ;
        RECT 82.375 154.175 82.590 154.225 ;
        RECT 82.375 154.095 82.765 154.175 ;
        RECT 82.435 153.250 82.765 154.095 ;
        RECT 83.275 154.140 83.465 154.345 ;
        RECT 82.935 153.035 83.105 154.045 ;
        RECT 83.275 153.765 84.170 154.140 ;
        RECT 83.275 153.205 83.615 153.765 ;
        RECT 83.845 153.035 84.160 153.535 ;
        RECT 84.340 153.505 84.510 154.345 ;
        RECT 84.680 154.635 85.145 154.965 ;
        RECT 85.530 154.905 85.700 155.135 ;
        RECT 85.880 155.085 86.250 155.585 ;
        RECT 86.570 155.135 87.245 155.305 ;
        RECT 87.440 155.135 87.775 155.305 ;
        RECT 84.680 153.675 85.000 154.635 ;
        RECT 85.530 154.605 86.360 154.905 ;
        RECT 85.170 153.705 85.360 154.425 ;
        RECT 85.530 153.535 85.700 154.605 ;
        RECT 86.160 154.575 86.360 154.605 ;
        RECT 85.870 154.355 86.040 154.425 ;
        RECT 86.570 154.355 86.740 155.135 ;
        RECT 87.605 154.995 87.775 155.135 ;
        RECT 87.945 155.125 88.195 155.585 ;
        RECT 85.870 154.185 86.740 154.355 ;
        RECT 86.910 154.715 87.435 154.935 ;
        RECT 87.605 154.865 87.830 154.995 ;
        RECT 85.870 154.095 86.380 154.185 ;
        RECT 84.340 153.335 85.225 153.505 ;
        RECT 85.450 153.205 85.700 153.535 ;
        RECT 85.870 153.035 86.040 153.835 ;
        RECT 86.210 153.480 86.380 154.095 ;
        RECT 86.910 154.015 87.080 154.715 ;
        RECT 86.550 153.650 87.080 154.015 ;
        RECT 87.250 153.950 87.490 154.545 ;
        RECT 87.660 153.760 87.830 154.865 ;
        RECT 88.000 154.005 88.280 154.955 ;
        RECT 87.525 153.630 87.830 153.760 ;
        RECT 86.210 153.310 87.315 153.480 ;
        RECT 87.525 153.205 87.775 153.630 ;
        RECT 87.945 153.035 88.210 153.495 ;
        RECT 88.450 153.205 88.635 155.325 ;
        RECT 88.805 155.205 89.135 155.585 ;
        RECT 89.305 155.035 89.475 155.325 ;
        RECT 88.810 154.865 89.475 155.035 ;
        RECT 88.810 153.875 89.040 154.865 ;
        RECT 89.740 154.845 89.995 155.415 ;
        RECT 90.165 155.185 90.495 155.585 ;
        RECT 90.920 155.050 91.450 155.415 ;
        RECT 90.920 155.015 91.095 155.050 ;
        RECT 90.165 154.845 91.095 155.015 ;
        RECT 89.210 154.045 89.560 154.695 ;
        RECT 89.740 154.175 89.910 154.845 ;
        RECT 90.165 154.675 90.335 154.845 ;
        RECT 90.080 154.345 90.335 154.675 ;
        RECT 90.560 154.345 90.755 154.675 ;
        RECT 88.810 153.705 89.475 153.875 ;
        RECT 88.805 153.035 89.135 153.535 ;
        RECT 89.305 153.205 89.475 153.705 ;
        RECT 89.740 153.205 90.075 154.175 ;
        RECT 90.245 153.035 90.415 154.175 ;
        RECT 90.585 153.375 90.755 154.345 ;
        RECT 90.925 153.715 91.095 154.845 ;
        RECT 91.265 154.055 91.435 154.855 ;
        RECT 91.640 154.565 91.915 155.415 ;
        RECT 91.635 154.395 91.915 154.565 ;
        RECT 91.640 154.255 91.915 154.395 ;
        RECT 92.085 154.055 92.275 155.415 ;
        RECT 92.455 155.050 92.965 155.585 ;
        RECT 93.185 154.775 93.430 155.380 ;
        RECT 94.795 154.860 95.085 155.585 ;
        RECT 96.235 155.125 96.480 155.585 ;
        RECT 92.475 154.605 93.705 154.775 ;
        RECT 91.265 153.885 92.275 154.055 ;
        RECT 92.445 154.040 93.195 154.230 ;
        RECT 90.925 153.545 92.050 153.715 ;
        RECT 92.445 153.375 92.615 154.040 ;
        RECT 93.365 153.795 93.705 154.605 ;
        RECT 96.175 154.345 96.490 154.955 ;
        RECT 96.660 154.595 96.910 155.405 ;
        RECT 97.080 155.060 97.340 155.585 ;
        RECT 97.510 154.935 97.770 155.390 ;
        RECT 97.940 155.105 98.200 155.585 ;
        RECT 98.370 154.935 98.630 155.390 ;
        RECT 98.800 155.105 99.060 155.585 ;
        RECT 99.230 154.935 99.490 155.390 ;
        RECT 99.660 155.105 99.920 155.585 ;
        RECT 100.090 154.935 100.350 155.390 ;
        RECT 100.520 155.105 100.820 155.585 ;
        RECT 97.510 154.765 100.820 154.935 ;
        RECT 96.660 154.345 99.680 154.595 ;
        RECT 90.585 153.205 92.615 153.375 ;
        RECT 92.785 153.035 92.955 153.795 ;
        RECT 93.190 153.385 93.705 153.795 ;
        RECT 94.795 153.035 95.085 154.200 ;
        RECT 96.185 153.035 96.480 154.145 ;
        RECT 96.660 153.210 96.910 154.345 ;
        RECT 99.850 154.175 100.820 154.765 ;
        RECT 97.080 153.035 97.340 154.145 ;
        RECT 97.510 153.935 100.820 154.175 ;
        RECT 101.240 154.845 101.495 155.415 ;
        RECT 101.665 155.185 101.995 155.585 ;
        RECT 102.420 155.050 102.950 155.415 ;
        RECT 102.420 155.015 102.595 155.050 ;
        RECT 101.665 154.845 102.595 155.015 ;
        RECT 103.140 154.905 103.415 155.415 ;
        RECT 101.240 154.175 101.410 154.845 ;
        RECT 101.665 154.675 101.835 154.845 ;
        RECT 101.580 154.345 101.835 154.675 ;
        RECT 102.060 154.345 102.255 154.675 ;
        RECT 97.510 153.210 97.770 153.935 ;
        RECT 97.940 153.035 98.200 153.765 ;
        RECT 98.370 153.210 98.630 153.935 ;
        RECT 98.800 153.035 99.060 153.765 ;
        RECT 99.230 153.210 99.490 153.935 ;
        RECT 99.660 153.035 99.920 153.765 ;
        RECT 100.090 153.210 100.350 153.935 ;
        RECT 100.520 153.035 100.815 153.765 ;
        RECT 101.240 153.205 101.575 154.175 ;
        RECT 101.745 153.035 101.915 154.175 ;
        RECT 102.085 153.375 102.255 154.345 ;
        RECT 102.425 153.715 102.595 154.845 ;
        RECT 102.765 154.055 102.935 154.855 ;
        RECT 103.135 154.735 103.415 154.905 ;
        RECT 103.140 154.255 103.415 154.735 ;
        RECT 103.585 154.055 103.775 155.415 ;
        RECT 103.955 155.050 104.465 155.585 ;
        RECT 104.685 154.775 104.930 155.380 ;
        RECT 105.380 154.845 105.635 155.415 ;
        RECT 105.805 155.185 106.135 155.585 ;
        RECT 106.560 155.050 107.090 155.415 ;
        RECT 106.560 155.015 106.735 155.050 ;
        RECT 105.805 154.845 106.735 155.015 ;
        RECT 103.975 154.605 105.205 154.775 ;
        RECT 102.765 153.885 103.775 154.055 ;
        RECT 103.945 154.040 104.695 154.230 ;
        RECT 102.425 153.545 103.550 153.715 ;
        RECT 103.945 153.375 104.115 154.040 ;
        RECT 104.865 153.795 105.205 154.605 ;
        RECT 102.085 153.205 104.115 153.375 ;
        RECT 104.285 153.035 104.455 153.795 ;
        RECT 104.690 153.385 105.205 153.795 ;
        RECT 105.380 154.175 105.550 154.845 ;
        RECT 105.805 154.675 105.975 154.845 ;
        RECT 105.720 154.345 105.975 154.675 ;
        RECT 106.200 154.345 106.395 154.675 ;
        RECT 105.380 153.205 105.715 154.175 ;
        RECT 105.885 153.035 106.055 154.175 ;
        RECT 106.225 153.375 106.395 154.345 ;
        RECT 106.565 153.715 106.735 154.845 ;
        RECT 106.905 154.055 107.075 154.855 ;
        RECT 107.280 154.565 107.555 155.415 ;
        RECT 107.275 154.395 107.555 154.565 ;
        RECT 107.280 154.255 107.555 154.395 ;
        RECT 107.725 154.055 107.915 155.415 ;
        RECT 108.095 155.050 108.605 155.585 ;
        RECT 108.825 154.775 109.070 155.380 ;
        RECT 109.515 154.845 109.900 155.415 ;
        RECT 110.070 155.125 110.395 155.585 ;
        RECT 110.915 154.955 111.195 155.415 ;
        RECT 108.115 154.605 109.345 154.775 ;
        RECT 106.905 153.885 107.915 154.055 ;
        RECT 108.085 154.040 108.835 154.230 ;
        RECT 106.565 153.545 107.690 153.715 ;
        RECT 108.085 153.375 108.255 154.040 ;
        RECT 109.005 153.795 109.345 154.605 ;
        RECT 106.225 153.205 108.255 153.375 ;
        RECT 108.425 153.035 108.595 153.795 ;
        RECT 108.830 153.385 109.345 153.795 ;
        RECT 109.515 154.175 109.795 154.845 ;
        RECT 110.070 154.785 111.195 154.955 ;
        RECT 110.070 154.675 110.520 154.785 ;
        RECT 109.965 154.345 110.520 154.675 ;
        RECT 111.385 154.615 111.785 155.415 ;
        RECT 112.185 155.125 112.455 155.585 ;
        RECT 112.625 154.955 112.910 155.415 ;
        RECT 109.515 153.205 109.900 154.175 ;
        RECT 110.070 153.885 110.520 154.345 ;
        RECT 110.690 154.055 111.785 154.615 ;
        RECT 110.070 153.665 111.195 153.885 ;
        RECT 110.070 153.035 110.395 153.495 ;
        RECT 110.915 153.205 111.195 153.665 ;
        RECT 111.385 153.205 111.785 154.055 ;
        RECT 111.955 154.785 112.910 154.955 ;
        RECT 113.200 154.820 113.655 155.585 ;
        RECT 113.930 155.205 115.230 155.415 ;
        RECT 115.485 155.225 115.815 155.585 ;
        RECT 115.060 155.055 115.230 155.205 ;
        RECT 115.985 155.085 116.245 155.415 ;
        RECT 111.955 153.885 112.165 154.785 ;
        RECT 112.335 154.055 113.025 154.615 ;
        RECT 114.130 154.595 114.350 154.995 ;
        RECT 113.195 154.395 113.685 154.595 ;
        RECT 113.875 154.385 114.350 154.595 ;
        RECT 114.595 154.595 114.805 154.995 ;
        RECT 115.060 154.930 115.815 155.055 ;
        RECT 115.060 154.885 115.905 154.930 ;
        RECT 115.635 154.765 115.905 154.885 ;
        RECT 114.595 154.385 114.925 154.595 ;
        RECT 115.095 154.325 115.505 154.630 ;
        RECT 113.200 154.155 114.375 154.215 ;
        RECT 115.735 154.190 115.905 154.765 ;
        RECT 115.705 154.155 115.905 154.190 ;
        RECT 113.200 154.045 115.905 154.155 ;
        RECT 111.955 153.665 112.910 153.885 ;
        RECT 112.185 153.035 112.455 153.495 ;
        RECT 112.625 153.205 112.910 153.665 ;
        RECT 113.200 153.425 113.455 154.045 ;
        RECT 114.045 153.985 115.845 154.045 ;
        RECT 114.045 153.955 114.375 153.985 ;
        RECT 116.075 153.885 116.245 155.085 ;
        RECT 113.705 153.785 113.890 153.875 ;
        RECT 114.480 153.785 115.315 153.795 ;
        RECT 113.705 153.585 115.315 153.785 ;
        RECT 113.705 153.545 113.935 153.585 ;
        RECT 113.200 153.205 113.535 153.425 ;
        RECT 114.540 153.035 114.895 153.415 ;
        RECT 115.065 153.205 115.315 153.585 ;
        RECT 115.565 153.035 115.815 153.815 ;
        RECT 115.985 153.205 116.245 153.885 ;
        RECT 116.425 154.860 116.755 155.370 ;
        RECT 116.925 155.185 117.255 155.585 ;
        RECT 118.305 155.015 118.635 155.355 ;
        RECT 118.805 155.185 119.135 155.585 ;
        RECT 116.425 154.095 116.615 154.860 ;
        RECT 116.925 154.845 119.290 155.015 ;
        RECT 120.555 154.860 120.845 155.585 ;
        RECT 121.030 155.015 121.285 155.365 ;
        RECT 121.455 155.185 121.785 155.585 ;
        RECT 121.955 155.015 122.125 155.365 ;
        RECT 122.295 155.185 122.675 155.585 ;
        RECT 121.030 154.845 122.695 155.015 ;
        RECT 122.865 154.910 123.140 155.255 ;
        RECT 123.375 155.125 123.620 155.585 ;
        RECT 116.925 154.675 117.095 154.845 ;
        RECT 116.785 154.345 117.095 154.675 ;
        RECT 117.265 154.345 117.570 154.675 ;
        RECT 116.425 153.245 116.755 154.095 ;
        RECT 116.925 153.035 117.175 154.175 ;
        RECT 117.355 154.015 117.570 154.345 ;
        RECT 117.745 154.015 118.030 154.675 ;
        RECT 118.225 154.015 118.490 154.675 ;
        RECT 118.705 154.015 118.950 154.675 ;
        RECT 119.120 153.845 119.290 154.845 ;
        RECT 122.525 154.675 122.695 154.845 ;
        RECT 121.015 154.345 121.360 154.675 ;
        RECT 121.530 154.345 122.355 154.675 ;
        RECT 122.525 154.345 122.800 154.675 ;
        RECT 117.365 153.675 118.655 153.845 ;
        RECT 117.365 153.255 117.615 153.675 ;
        RECT 117.845 153.035 118.175 153.505 ;
        RECT 118.405 153.255 118.655 153.675 ;
        RECT 118.835 153.675 119.290 153.845 ;
        RECT 118.835 153.245 119.165 153.675 ;
        RECT 120.555 153.035 120.845 154.200 ;
        RECT 121.035 153.885 121.360 154.175 ;
        RECT 121.530 154.055 121.725 154.345 ;
        RECT 122.525 154.175 122.695 154.345 ;
        RECT 122.970 154.175 123.140 154.910 ;
        RECT 123.315 154.345 123.630 154.955 ;
        RECT 123.800 154.595 124.050 155.405 ;
        RECT 124.220 155.060 124.480 155.585 ;
        RECT 124.650 154.935 124.910 155.390 ;
        RECT 125.080 155.105 125.340 155.585 ;
        RECT 125.510 154.935 125.770 155.390 ;
        RECT 125.940 155.105 126.200 155.585 ;
        RECT 126.370 154.935 126.630 155.390 ;
        RECT 126.800 155.105 127.060 155.585 ;
        RECT 127.230 154.935 127.490 155.390 ;
        RECT 127.660 155.105 127.960 155.585 ;
        RECT 128.540 155.075 128.780 155.585 ;
        RECT 128.960 155.075 129.240 155.405 ;
        RECT 129.470 155.075 129.685 155.585 ;
        RECT 124.650 154.765 127.960 154.935 ;
        RECT 123.800 154.345 126.820 154.595 ;
        RECT 122.035 154.005 122.695 154.175 ;
        RECT 122.035 153.885 122.205 154.005 ;
        RECT 121.035 153.715 122.205 153.885 ;
        RECT 121.015 153.255 122.205 153.545 ;
        RECT 122.375 153.035 122.655 153.835 ;
        RECT 122.865 153.205 123.140 154.175 ;
        RECT 123.325 153.035 123.620 154.145 ;
        RECT 123.800 153.210 124.050 154.345 ;
        RECT 126.990 154.175 127.960 154.765 ;
        RECT 128.435 154.345 128.790 154.905 ;
        RECT 128.960 154.175 129.130 155.075 ;
        RECT 129.300 154.345 129.565 154.905 ;
        RECT 129.855 154.845 130.470 155.415 ;
        RECT 130.765 155.035 130.935 155.325 ;
        RECT 131.105 155.205 131.435 155.585 ;
        RECT 130.765 154.865 131.430 155.035 ;
        RECT 129.815 154.175 129.985 154.675 ;
        RECT 124.220 153.035 124.480 154.145 ;
        RECT 124.650 153.935 127.960 154.175 ;
        RECT 128.560 154.005 129.985 154.175 ;
        RECT 124.650 153.210 124.910 153.935 ;
        RECT 125.080 153.035 125.340 153.765 ;
        RECT 125.510 153.210 125.770 153.935 ;
        RECT 125.940 153.035 126.200 153.765 ;
        RECT 126.370 153.210 126.630 153.935 ;
        RECT 126.800 153.035 127.060 153.765 ;
        RECT 127.230 153.210 127.490 153.935 ;
        RECT 128.560 153.830 128.950 154.005 ;
        RECT 127.660 153.035 127.955 153.765 ;
        RECT 129.435 153.035 129.765 153.835 ;
        RECT 130.155 153.825 130.470 154.845 ;
        RECT 130.680 154.045 131.030 154.695 ;
        RECT 131.200 153.875 131.430 154.865 ;
        RECT 129.935 153.205 130.470 153.825 ;
        RECT 130.765 153.705 131.430 153.875 ;
        RECT 130.765 153.205 130.935 153.705 ;
        RECT 131.105 153.035 131.435 153.535 ;
        RECT 131.605 153.205 131.790 155.325 ;
        RECT 132.045 155.125 132.295 155.585 ;
        RECT 132.465 155.135 132.800 155.305 ;
        RECT 132.995 155.135 133.670 155.305 ;
        RECT 132.465 154.995 132.635 155.135 ;
        RECT 131.960 154.005 132.240 154.955 ;
        RECT 132.410 154.865 132.635 154.995 ;
        RECT 132.410 153.760 132.580 154.865 ;
        RECT 132.805 154.715 133.330 154.935 ;
        RECT 132.750 153.950 132.990 154.545 ;
        RECT 133.160 154.015 133.330 154.715 ;
        RECT 133.500 154.355 133.670 155.135 ;
        RECT 133.990 155.085 134.360 155.585 ;
        RECT 134.540 155.135 134.945 155.305 ;
        RECT 135.115 155.135 135.900 155.305 ;
        RECT 134.540 154.905 134.710 155.135 ;
        RECT 133.880 154.605 134.710 154.905 ;
        RECT 135.095 154.635 135.560 154.965 ;
        RECT 133.880 154.575 134.080 154.605 ;
        RECT 134.200 154.355 134.370 154.425 ;
        RECT 133.500 154.185 134.370 154.355 ;
        RECT 133.860 154.095 134.370 154.185 ;
        RECT 132.410 153.630 132.715 153.760 ;
        RECT 133.160 153.650 133.690 154.015 ;
        RECT 132.030 153.035 132.295 153.495 ;
        RECT 132.465 153.205 132.715 153.630 ;
        RECT 133.860 153.480 134.030 154.095 ;
        RECT 132.925 153.310 134.030 153.480 ;
        RECT 134.200 153.035 134.370 153.835 ;
        RECT 134.540 153.535 134.710 154.605 ;
        RECT 134.880 153.705 135.070 154.425 ;
        RECT 135.240 153.675 135.560 154.635 ;
        RECT 135.730 154.675 135.900 155.135 ;
        RECT 136.175 155.055 136.385 155.585 ;
        RECT 136.645 154.845 136.975 155.370 ;
        RECT 137.145 154.975 137.315 155.585 ;
        RECT 137.485 154.930 137.815 155.365 ;
        RECT 138.125 155.035 138.295 155.415 ;
        RECT 138.475 155.205 138.805 155.585 ;
        RECT 137.485 154.845 137.865 154.930 ;
        RECT 138.125 154.865 138.790 155.035 ;
        RECT 138.985 154.910 139.245 155.415 ;
        RECT 136.775 154.675 136.975 154.845 ;
        RECT 137.640 154.805 137.865 154.845 ;
        RECT 135.730 154.345 136.605 154.675 ;
        RECT 136.775 154.345 137.525 154.675 ;
        RECT 134.540 153.205 134.790 153.535 ;
        RECT 135.730 153.505 135.900 154.345 ;
        RECT 136.775 154.140 136.965 154.345 ;
        RECT 137.695 154.225 137.865 154.805 ;
        RECT 138.055 154.315 138.385 154.685 ;
        RECT 138.620 154.610 138.790 154.865 ;
        RECT 137.650 154.175 137.865 154.225 ;
        RECT 136.070 153.765 136.965 154.140 ;
        RECT 137.475 154.095 137.865 154.175 ;
        RECT 138.620 154.280 138.905 154.610 ;
        RECT 138.620 154.135 138.790 154.280 ;
        RECT 135.015 153.335 135.900 153.505 ;
        RECT 136.080 153.035 136.395 153.535 ;
        RECT 136.625 153.205 136.965 153.765 ;
        RECT 137.135 153.035 137.305 154.045 ;
        RECT 137.475 153.250 137.805 154.095 ;
        RECT 138.125 153.965 138.790 154.135 ;
        RECT 139.075 154.110 139.245 154.910 ;
        RECT 139.965 155.035 140.135 155.415 ;
        RECT 140.350 155.205 140.680 155.585 ;
        RECT 139.965 154.865 140.680 155.035 ;
        RECT 139.875 154.315 140.230 154.685 ;
        RECT 140.510 154.675 140.680 154.865 ;
        RECT 140.850 154.840 141.105 155.415 ;
        RECT 140.510 154.345 140.765 154.675 ;
        RECT 140.510 154.135 140.680 154.345 ;
        RECT 138.125 153.205 138.295 153.965 ;
        RECT 138.475 153.035 138.805 153.795 ;
        RECT 138.975 153.205 139.245 154.110 ;
        RECT 139.965 153.965 140.680 154.135 ;
        RECT 140.935 154.110 141.105 154.840 ;
        RECT 141.280 154.745 141.540 155.585 ;
        RECT 141.715 154.835 142.925 155.585 ;
        RECT 139.965 153.205 140.135 153.965 ;
        RECT 140.350 153.035 140.680 153.795 ;
        RECT 140.850 153.205 141.105 154.110 ;
        RECT 141.280 153.035 141.540 154.185 ;
        RECT 141.715 154.125 142.235 154.665 ;
        RECT 142.405 154.295 142.925 154.835 ;
        RECT 141.715 153.035 142.925 154.125 ;
        RECT 17.430 152.865 143.010 153.035 ;
        RECT 17.515 151.775 18.725 152.865 ;
        RECT 18.895 152.430 24.240 152.865 ;
        RECT 24.415 152.430 29.760 152.865 ;
        RECT 17.515 151.065 18.035 151.605 ;
        RECT 18.205 151.235 18.725 151.775 ;
        RECT 17.515 150.315 18.725 151.065 ;
        RECT 20.480 150.860 20.820 151.690 ;
        RECT 22.300 151.180 22.650 152.430 ;
        RECT 26.000 150.860 26.340 151.690 ;
        RECT 27.820 151.180 28.170 152.430 ;
        RECT 30.395 151.700 30.685 152.865 ;
        RECT 30.855 152.430 36.200 152.865 ;
        RECT 18.895 150.315 24.240 150.860 ;
        RECT 24.415 150.315 29.760 150.860 ;
        RECT 30.395 150.315 30.685 151.040 ;
        RECT 32.440 150.860 32.780 151.690 ;
        RECT 34.260 151.180 34.610 152.430 ;
        RECT 36.375 151.775 38.045 152.865 ;
        RECT 36.375 151.085 37.125 151.605 ;
        RECT 37.295 151.255 38.045 151.775 ;
        RECT 38.215 151.845 38.590 152.695 ;
        RECT 38.760 152.065 39.010 152.865 ;
        RECT 39.180 152.235 39.430 152.695 ;
        RECT 39.600 152.405 39.850 152.865 ;
        RECT 40.020 152.235 40.270 152.695 ;
        RECT 40.440 152.405 40.690 152.865 ;
        RECT 40.860 152.235 41.110 152.695 ;
        RECT 41.280 152.405 41.530 152.865 ;
        RECT 41.700 152.235 41.950 152.695 ;
        RECT 39.180 152.015 41.950 152.235 ;
        RECT 42.165 152.235 42.480 152.695 ;
        RECT 42.650 152.405 42.900 152.865 ;
        RECT 43.070 152.235 43.320 152.695 ;
        RECT 43.490 152.405 43.740 152.865 ;
        RECT 43.910 152.445 45.880 152.695 ;
        RECT 43.910 152.235 44.120 152.445 ;
        RECT 46.090 152.275 46.380 152.695 ;
        RECT 42.165 152.015 44.120 152.235 ;
        RECT 44.290 152.015 46.380 152.275 ;
        RECT 46.550 152.065 46.800 152.865 ;
        RECT 39.180 151.845 39.430 152.015 ;
        RECT 46.090 151.895 46.380 152.015 ;
        RECT 46.970 151.895 47.220 152.695 ;
        RECT 47.390 152.065 47.640 152.865 ;
        RECT 47.810 151.895 48.165 152.695 ;
        RECT 48.335 152.430 53.680 152.865 ;
        RECT 38.215 151.675 39.430 151.845 ;
        RECT 39.815 151.675 43.860 151.845 ;
        RECT 44.030 151.675 45.900 151.845 ;
        RECT 46.090 151.675 48.165 151.895 ;
        RECT 38.215 151.135 38.450 151.675 ;
        RECT 39.815 151.505 39.985 151.675 ;
        RECT 43.690 151.505 43.860 151.675 ;
        RECT 45.730 151.505 45.900 151.675 ;
        RECT 38.620 151.305 39.985 151.505 ;
        RECT 40.305 151.305 43.520 151.505 ;
        RECT 43.690 151.305 45.560 151.505 ;
        RECT 45.730 151.305 47.775 151.505 ;
        RECT 47.945 151.135 48.165 151.675 ;
        RECT 30.855 150.315 36.200 150.860 ;
        RECT 36.375 150.315 38.045 151.085 ;
        RECT 38.215 150.875 39.890 151.135 ;
        RECT 40.060 150.955 41.990 151.135 ;
        RECT 40.060 150.705 40.310 150.955 ;
        RECT 38.300 150.485 40.310 150.705 ;
        RECT 40.480 150.315 40.650 150.785 ;
        RECT 40.820 150.485 41.150 150.955 ;
        RECT 41.320 150.315 41.490 150.785 ;
        RECT 41.660 150.485 41.990 150.955 ;
        RECT 42.165 150.315 42.440 151.135 ;
        RECT 42.610 150.965 46.340 151.135 ;
        RECT 42.610 150.955 45.560 150.965 ;
        RECT 42.610 150.485 42.940 150.955 ;
        RECT 43.110 150.315 43.280 150.785 ;
        RECT 43.450 150.485 43.780 150.955 ;
        RECT 43.950 150.315 44.120 150.785 ;
        RECT 44.290 150.485 44.620 150.955 ;
        RECT 44.790 150.315 44.960 150.785 ;
        RECT 45.130 150.485 45.460 150.955 ;
        RECT 45.630 150.315 45.900 150.785 ;
        RECT 46.090 150.705 46.340 150.965 ;
        RECT 46.510 150.875 48.165 151.135 ;
        RECT 49.920 150.860 50.260 151.690 ;
        RECT 51.740 151.180 52.090 152.430 ;
        RECT 53.855 151.775 55.525 152.865 ;
        RECT 53.855 151.085 54.605 151.605 ;
        RECT 54.775 151.255 55.525 151.775 ;
        RECT 56.155 151.700 56.445 152.865 ;
        RECT 56.615 152.430 61.960 152.865 ;
        RECT 62.135 152.430 67.480 152.865 ;
        RECT 46.090 150.535 48.100 150.705 ;
        RECT 48.335 150.315 53.680 150.860 ;
        RECT 53.855 150.315 55.525 151.085 ;
        RECT 56.155 150.315 56.445 151.040 ;
        RECT 58.200 150.860 58.540 151.690 ;
        RECT 60.020 151.180 60.370 152.430 ;
        RECT 63.720 150.860 64.060 151.690 ;
        RECT 65.540 151.180 65.890 152.430 ;
        RECT 67.655 151.775 70.245 152.865 ;
        RECT 67.655 151.085 68.865 151.605 ;
        RECT 69.035 151.255 70.245 151.775 ;
        RECT 70.880 151.725 71.215 152.695 ;
        RECT 71.385 151.725 71.555 152.865 ;
        RECT 71.725 152.525 73.755 152.695 ;
        RECT 56.615 150.315 61.960 150.860 ;
        RECT 62.135 150.315 67.480 150.860 ;
        RECT 67.655 150.315 70.245 151.085 ;
        RECT 70.880 151.055 71.050 151.725 ;
        RECT 71.725 151.555 71.895 152.525 ;
        RECT 71.220 151.225 71.475 151.555 ;
        RECT 71.700 151.225 71.895 151.555 ;
        RECT 72.065 152.185 73.190 152.355 ;
        RECT 71.305 151.055 71.475 151.225 ;
        RECT 72.065 151.055 72.235 152.185 ;
        RECT 70.880 150.485 71.135 151.055 ;
        RECT 71.305 150.885 72.235 151.055 ;
        RECT 72.405 151.845 73.415 152.015 ;
        RECT 72.405 151.045 72.575 151.845 ;
        RECT 72.780 151.165 73.055 151.645 ;
        RECT 72.775 150.995 73.055 151.165 ;
        RECT 72.060 150.850 72.235 150.885 ;
        RECT 71.305 150.315 71.635 150.715 ;
        RECT 72.060 150.485 72.590 150.850 ;
        RECT 72.780 150.485 73.055 150.995 ;
        RECT 73.225 150.485 73.415 151.845 ;
        RECT 73.585 151.860 73.755 152.525 ;
        RECT 73.925 152.105 74.095 152.865 ;
        RECT 74.330 152.105 74.845 152.515 ;
        RECT 73.585 151.670 74.335 151.860 ;
        RECT 74.505 151.295 74.845 152.105 ;
        RECT 75.015 151.775 76.225 152.865 ;
        RECT 73.615 151.125 74.845 151.295 ;
        RECT 73.595 150.315 74.105 150.850 ;
        RECT 74.325 150.520 74.570 151.125 ;
        RECT 75.015 151.065 75.535 151.605 ;
        RECT 75.705 151.235 76.225 151.775 ;
        RECT 76.395 151.725 76.780 152.695 ;
        RECT 76.950 152.405 77.275 152.865 ;
        RECT 77.795 152.235 78.075 152.695 ;
        RECT 76.950 152.015 78.075 152.235 ;
        RECT 75.015 150.315 76.225 151.065 ;
        RECT 76.395 151.055 76.675 151.725 ;
        RECT 76.950 151.555 77.400 152.015 ;
        RECT 78.265 151.845 78.665 152.695 ;
        RECT 79.065 152.405 79.335 152.865 ;
        RECT 79.505 152.235 79.790 152.695 ;
        RECT 76.845 151.225 77.400 151.555 ;
        RECT 77.570 151.285 78.665 151.845 ;
        RECT 76.950 151.115 77.400 151.225 ;
        RECT 76.395 150.485 76.780 151.055 ;
        RECT 76.950 150.945 78.075 151.115 ;
        RECT 76.950 150.315 77.275 150.775 ;
        RECT 77.795 150.485 78.075 150.945 ;
        RECT 78.265 150.485 78.665 151.285 ;
        RECT 78.835 152.015 79.790 152.235 ;
        RECT 78.835 151.115 79.045 152.015 ;
        RECT 79.215 151.285 79.905 151.845 ;
        RECT 80.075 151.775 81.745 152.865 ;
        RECT 78.835 150.945 79.790 151.115 ;
        RECT 79.065 150.315 79.335 150.775 ;
        RECT 79.505 150.485 79.790 150.945 ;
        RECT 80.075 151.085 80.825 151.605 ;
        RECT 80.995 151.255 81.745 151.775 ;
        RECT 81.915 151.700 82.205 152.865 ;
        RECT 82.375 152.430 87.720 152.865 ;
        RECT 80.075 150.315 81.745 151.085 ;
        RECT 81.915 150.315 82.205 151.040 ;
        RECT 83.960 150.860 84.300 151.690 ;
        RECT 85.780 151.180 86.130 152.430 ;
        RECT 87.895 151.775 89.105 152.865 ;
        RECT 87.895 151.065 88.415 151.605 ;
        RECT 88.585 151.235 89.105 151.775 ;
        RECT 89.275 152.105 89.790 152.515 ;
        RECT 90.025 152.105 90.195 152.865 ;
        RECT 90.365 152.525 92.395 152.695 ;
        RECT 89.275 151.295 89.615 152.105 ;
        RECT 90.365 151.860 90.535 152.525 ;
        RECT 90.930 152.185 92.055 152.355 ;
        RECT 89.785 151.670 90.535 151.860 ;
        RECT 90.705 151.845 91.715 152.015 ;
        RECT 89.275 151.125 90.505 151.295 ;
        RECT 82.375 150.315 87.720 150.860 ;
        RECT 87.895 150.315 89.105 151.065 ;
        RECT 89.550 150.520 89.795 151.125 ;
        RECT 90.015 150.315 90.525 150.850 ;
        RECT 90.705 150.485 90.895 151.845 ;
        RECT 91.065 150.825 91.340 151.645 ;
        RECT 91.545 151.045 91.715 151.845 ;
        RECT 91.885 151.055 92.055 152.185 ;
        RECT 92.225 151.555 92.395 152.525 ;
        RECT 92.565 151.725 92.735 152.865 ;
        RECT 92.905 151.725 93.240 152.695 ;
        RECT 93.415 151.775 96.005 152.865 ;
        RECT 96.725 152.195 96.895 152.695 ;
        RECT 97.065 152.365 97.395 152.865 ;
        RECT 96.725 152.025 97.390 152.195 ;
        RECT 92.225 151.225 92.420 151.555 ;
        RECT 92.645 151.225 92.900 151.555 ;
        RECT 92.645 151.055 92.815 151.225 ;
        RECT 93.070 151.055 93.240 151.725 ;
        RECT 91.885 150.885 92.815 151.055 ;
        RECT 91.885 150.850 92.060 150.885 ;
        RECT 91.065 150.655 91.345 150.825 ;
        RECT 91.065 150.485 91.340 150.655 ;
        RECT 91.530 150.485 92.060 150.850 ;
        RECT 92.485 150.315 92.815 150.715 ;
        RECT 92.985 150.485 93.240 151.055 ;
        RECT 93.415 151.085 94.625 151.605 ;
        RECT 94.795 151.255 96.005 151.775 ;
        RECT 96.640 151.205 96.990 151.855 ;
        RECT 93.415 150.315 96.005 151.085 ;
        RECT 97.160 151.035 97.390 152.025 ;
        RECT 96.725 150.865 97.390 151.035 ;
        RECT 96.725 150.575 96.895 150.865 ;
        RECT 97.065 150.315 97.395 150.695 ;
        RECT 97.565 150.575 97.750 152.695 ;
        RECT 97.990 152.405 98.255 152.865 ;
        RECT 98.425 152.270 98.675 152.695 ;
        RECT 98.885 152.420 99.990 152.590 ;
        RECT 98.370 152.140 98.675 152.270 ;
        RECT 97.920 150.945 98.200 151.895 ;
        RECT 98.370 151.035 98.540 152.140 ;
        RECT 98.710 151.355 98.950 151.950 ;
        RECT 99.120 151.885 99.650 152.250 ;
        RECT 99.120 151.185 99.290 151.885 ;
        RECT 99.820 151.805 99.990 152.420 ;
        RECT 100.160 152.065 100.330 152.865 ;
        RECT 100.500 152.365 100.750 152.695 ;
        RECT 100.975 152.395 101.860 152.565 ;
        RECT 99.820 151.715 100.330 151.805 ;
        RECT 98.370 150.905 98.595 151.035 ;
        RECT 98.765 150.965 99.290 151.185 ;
        RECT 99.460 151.545 100.330 151.715 ;
        RECT 98.005 150.315 98.255 150.775 ;
        RECT 98.425 150.765 98.595 150.905 ;
        RECT 99.460 150.765 99.630 151.545 ;
        RECT 100.160 151.475 100.330 151.545 ;
        RECT 99.840 151.295 100.040 151.325 ;
        RECT 100.500 151.295 100.670 152.365 ;
        RECT 100.840 151.475 101.030 152.195 ;
        RECT 99.840 150.995 100.670 151.295 ;
        RECT 101.200 151.265 101.520 152.225 ;
        RECT 98.425 150.595 98.760 150.765 ;
        RECT 98.955 150.595 99.630 150.765 ;
        RECT 99.950 150.315 100.320 150.815 ;
        RECT 100.500 150.765 100.670 150.995 ;
        RECT 101.055 150.935 101.520 151.265 ;
        RECT 101.690 151.555 101.860 152.395 ;
        RECT 102.040 152.365 102.355 152.865 ;
        RECT 102.585 152.135 102.925 152.695 ;
        RECT 102.030 151.760 102.925 152.135 ;
        RECT 103.095 151.855 103.265 152.865 ;
        RECT 102.735 151.555 102.925 151.760 ;
        RECT 103.435 151.805 103.765 152.650 ;
        RECT 103.435 151.725 103.825 151.805 ;
        RECT 103.995 151.775 107.505 152.865 ;
        RECT 103.610 151.675 103.825 151.725 ;
        RECT 101.690 151.225 102.565 151.555 ;
        RECT 102.735 151.225 103.485 151.555 ;
        RECT 101.690 150.765 101.860 151.225 ;
        RECT 102.735 151.055 102.935 151.225 ;
        RECT 103.655 151.095 103.825 151.675 ;
        RECT 103.600 151.055 103.825 151.095 ;
        RECT 100.500 150.595 100.905 150.765 ;
        RECT 101.075 150.595 101.860 150.765 ;
        RECT 102.135 150.315 102.345 150.845 ;
        RECT 102.605 150.530 102.935 151.055 ;
        RECT 103.445 150.970 103.825 151.055 ;
        RECT 103.995 151.085 105.645 151.605 ;
        RECT 105.815 151.255 107.505 151.775 ;
        RECT 107.675 151.700 107.965 152.865 ;
        RECT 108.250 152.235 108.535 152.695 ;
        RECT 108.705 152.405 108.975 152.865 ;
        RECT 108.250 152.015 109.205 152.235 ;
        RECT 108.135 151.285 108.825 151.845 ;
        RECT 108.995 151.115 109.205 152.015 ;
        RECT 103.105 150.315 103.275 150.925 ;
        RECT 103.445 150.535 103.775 150.970 ;
        RECT 103.995 150.315 107.505 151.085 ;
        RECT 107.675 150.315 107.965 151.040 ;
        RECT 108.250 150.945 109.205 151.115 ;
        RECT 109.375 151.845 109.775 152.695 ;
        RECT 109.965 152.235 110.245 152.695 ;
        RECT 110.765 152.405 111.090 152.865 ;
        RECT 109.965 152.015 111.090 152.235 ;
        RECT 109.375 151.285 110.470 151.845 ;
        RECT 110.640 151.555 111.090 152.015 ;
        RECT 111.260 151.725 111.645 152.695 ;
        RECT 111.820 151.725 112.140 152.865 ;
        RECT 108.250 150.485 108.535 150.945 ;
        RECT 108.705 150.315 108.975 150.775 ;
        RECT 109.375 150.485 109.775 151.285 ;
        RECT 110.640 151.225 111.195 151.555 ;
        RECT 110.640 151.115 111.090 151.225 ;
        RECT 109.965 150.945 111.090 151.115 ;
        RECT 111.365 151.055 111.645 151.725 ;
        RECT 112.320 151.555 112.515 152.605 ;
        RECT 112.695 152.015 113.025 152.695 ;
        RECT 113.225 152.065 113.480 152.865 ;
        RECT 112.695 151.735 113.045 152.015 ;
        RECT 111.880 151.505 112.140 151.555 ;
        RECT 111.875 151.335 112.140 151.505 ;
        RECT 111.880 151.225 112.140 151.335 ;
        RECT 112.320 151.225 112.705 151.555 ;
        RECT 112.875 151.355 113.045 151.735 ;
        RECT 113.235 151.525 113.480 151.885 ;
        RECT 113.655 151.725 113.935 152.865 ;
        RECT 114.105 151.715 114.435 152.695 ;
        RECT 114.605 151.725 114.865 152.865 ;
        RECT 116.070 152.235 116.355 152.695 ;
        RECT 116.525 152.405 116.795 152.865 ;
        RECT 116.070 152.015 117.025 152.235 ;
        RECT 112.875 151.185 113.395 151.355 ;
        RECT 113.665 151.285 114.000 151.555 ;
        RECT 109.965 150.485 110.245 150.945 ;
        RECT 110.765 150.315 111.090 150.775 ;
        RECT 111.260 150.485 111.645 151.055 ;
        RECT 113.225 151.165 113.395 151.185 ;
        RECT 111.820 150.845 113.035 151.015 ;
        RECT 111.820 150.495 112.110 150.845 ;
        RECT 112.305 150.315 112.635 150.675 ;
        RECT 112.805 150.540 113.035 150.845 ;
        RECT 113.225 150.995 113.425 151.165 ;
        RECT 114.170 151.115 114.340 151.715 ;
        RECT 114.510 151.305 114.845 151.555 ;
        RECT 115.955 151.285 116.645 151.845 ;
        RECT 116.815 151.115 117.025 152.015 ;
        RECT 113.225 150.620 113.395 150.995 ;
        RECT 113.655 150.315 113.965 151.115 ;
        RECT 114.170 150.485 114.865 151.115 ;
        RECT 116.070 150.945 117.025 151.115 ;
        RECT 117.195 151.845 117.595 152.695 ;
        RECT 117.785 152.235 118.065 152.695 ;
        RECT 118.585 152.405 118.910 152.865 ;
        RECT 117.785 152.015 118.910 152.235 ;
        RECT 117.195 151.285 118.290 151.845 ;
        RECT 118.460 151.555 118.910 152.015 ;
        RECT 119.080 151.725 119.465 152.695 ;
        RECT 116.070 150.485 116.355 150.945 ;
        RECT 116.525 150.315 116.795 150.775 ;
        RECT 117.195 150.485 117.595 151.285 ;
        RECT 118.460 151.225 119.015 151.555 ;
        RECT 118.460 151.115 118.910 151.225 ;
        RECT 117.785 150.945 118.910 151.115 ;
        RECT 119.185 151.055 119.465 151.725 ;
        RECT 117.785 150.485 118.065 150.945 ;
        RECT 118.585 150.315 118.910 150.775 ;
        RECT 119.080 150.485 119.465 151.055 ;
        RECT 119.635 152.015 119.895 152.695 ;
        RECT 120.065 152.085 120.315 152.865 ;
        RECT 120.565 152.315 120.815 152.695 ;
        RECT 120.985 152.485 121.340 152.865 ;
        RECT 122.345 152.475 122.680 152.695 ;
        RECT 121.945 152.315 122.175 152.355 ;
        RECT 120.565 152.115 122.175 152.315 ;
        RECT 120.565 152.105 121.400 152.115 ;
        RECT 121.990 152.025 122.175 152.115 ;
        RECT 119.635 150.825 119.805 152.015 ;
        RECT 121.505 151.915 121.835 151.945 ;
        RECT 120.035 151.855 121.835 151.915 ;
        RECT 122.425 151.855 122.680 152.475 ;
        RECT 119.975 151.745 122.680 151.855 ;
        RECT 123.325 151.755 123.620 152.865 ;
        RECT 119.975 151.710 120.175 151.745 ;
        RECT 119.975 151.135 120.145 151.710 ;
        RECT 121.505 151.685 122.680 151.745 ;
        RECT 120.375 151.270 120.785 151.575 ;
        RECT 123.800 151.555 124.050 152.690 ;
        RECT 124.220 151.755 124.480 152.865 ;
        RECT 124.650 151.965 124.910 152.690 ;
        RECT 125.080 152.135 125.340 152.865 ;
        RECT 125.510 151.965 125.770 152.690 ;
        RECT 125.940 152.135 126.200 152.865 ;
        RECT 126.370 151.965 126.630 152.690 ;
        RECT 126.800 152.135 127.060 152.865 ;
        RECT 127.230 151.965 127.490 152.690 ;
        RECT 127.660 152.135 127.955 152.865 ;
        RECT 129.295 152.105 129.810 152.515 ;
        RECT 130.045 152.105 130.215 152.865 ;
        RECT 130.385 152.525 132.415 152.695 ;
        RECT 124.650 151.725 127.960 151.965 ;
        RECT 120.955 151.305 121.285 151.515 ;
        RECT 119.975 151.015 120.245 151.135 ;
        RECT 119.975 150.970 120.820 151.015 ;
        RECT 120.065 150.845 120.820 150.970 ;
        RECT 121.075 150.905 121.285 151.305 ;
        RECT 121.530 151.305 122.005 151.515 ;
        RECT 122.195 151.305 122.685 151.505 ;
        RECT 121.530 150.905 121.750 151.305 ;
        RECT 119.635 150.815 119.865 150.825 ;
        RECT 119.635 150.485 119.895 150.815 ;
        RECT 120.650 150.695 120.820 150.845 ;
        RECT 120.065 150.315 120.395 150.675 ;
        RECT 120.650 150.485 121.950 150.695 ;
        RECT 122.225 150.315 122.680 151.080 ;
        RECT 123.315 150.945 123.630 151.555 ;
        RECT 123.800 151.305 126.820 151.555 ;
        RECT 123.375 150.315 123.620 150.775 ;
        RECT 123.800 150.495 124.050 151.305 ;
        RECT 126.990 151.135 127.960 151.725 ;
        RECT 124.650 150.965 127.960 151.135 ;
        RECT 129.295 151.295 129.635 152.105 ;
        RECT 130.385 151.860 130.555 152.525 ;
        RECT 130.950 152.185 132.075 152.355 ;
        RECT 129.805 151.670 130.555 151.860 ;
        RECT 130.725 151.845 131.735 152.015 ;
        RECT 129.295 151.125 130.525 151.295 ;
        RECT 124.220 150.315 124.480 150.840 ;
        RECT 124.650 150.510 124.910 150.965 ;
        RECT 125.080 150.315 125.340 150.795 ;
        RECT 125.510 150.510 125.770 150.965 ;
        RECT 125.940 150.315 126.200 150.795 ;
        RECT 126.370 150.510 126.630 150.965 ;
        RECT 126.800 150.315 127.060 150.795 ;
        RECT 127.230 150.510 127.490 150.965 ;
        RECT 127.660 150.315 127.960 150.795 ;
        RECT 129.570 150.520 129.815 151.125 ;
        RECT 130.035 150.315 130.545 150.850 ;
        RECT 130.725 150.485 130.915 151.845 ;
        RECT 131.085 150.825 131.360 151.645 ;
        RECT 131.565 151.045 131.735 151.845 ;
        RECT 131.905 151.055 132.075 152.185 ;
        RECT 132.245 151.555 132.415 152.525 ;
        RECT 132.585 151.725 132.755 152.865 ;
        RECT 132.925 151.725 133.260 152.695 ;
        RECT 132.245 151.225 132.440 151.555 ;
        RECT 132.665 151.225 132.920 151.555 ;
        RECT 132.665 151.055 132.835 151.225 ;
        RECT 133.090 151.055 133.260 151.725 ;
        RECT 133.435 151.700 133.725 152.865 ;
        RECT 133.985 152.195 134.155 152.695 ;
        RECT 134.325 152.365 134.655 152.865 ;
        RECT 133.985 152.025 134.650 152.195 ;
        RECT 133.900 151.205 134.250 151.855 ;
        RECT 131.905 150.885 132.835 151.055 ;
        RECT 131.905 150.850 132.080 150.885 ;
        RECT 131.085 150.655 131.365 150.825 ;
        RECT 131.085 150.485 131.360 150.655 ;
        RECT 131.550 150.485 132.080 150.850 ;
        RECT 132.505 150.315 132.835 150.715 ;
        RECT 133.005 150.485 133.260 151.055 ;
        RECT 133.435 150.315 133.725 151.040 ;
        RECT 134.420 151.035 134.650 152.025 ;
        RECT 133.985 150.865 134.650 151.035 ;
        RECT 133.985 150.575 134.155 150.865 ;
        RECT 134.325 150.315 134.655 150.695 ;
        RECT 134.825 150.575 135.010 152.695 ;
        RECT 135.250 152.405 135.515 152.865 ;
        RECT 135.685 152.270 135.935 152.695 ;
        RECT 136.145 152.420 137.250 152.590 ;
        RECT 135.630 152.140 135.935 152.270 ;
        RECT 135.180 150.945 135.460 151.895 ;
        RECT 135.630 151.035 135.800 152.140 ;
        RECT 135.970 151.355 136.210 151.950 ;
        RECT 136.380 151.885 136.910 152.250 ;
        RECT 136.380 151.185 136.550 151.885 ;
        RECT 137.080 151.805 137.250 152.420 ;
        RECT 137.420 152.065 137.590 152.865 ;
        RECT 137.760 152.365 138.010 152.695 ;
        RECT 138.235 152.395 139.120 152.565 ;
        RECT 137.080 151.715 137.590 151.805 ;
        RECT 135.630 150.905 135.855 151.035 ;
        RECT 136.025 150.965 136.550 151.185 ;
        RECT 136.720 151.545 137.590 151.715 ;
        RECT 135.265 150.315 135.515 150.775 ;
        RECT 135.685 150.765 135.855 150.905 ;
        RECT 136.720 150.765 136.890 151.545 ;
        RECT 137.420 151.475 137.590 151.545 ;
        RECT 137.100 151.295 137.300 151.325 ;
        RECT 137.760 151.295 137.930 152.365 ;
        RECT 138.100 151.475 138.290 152.195 ;
        RECT 137.100 150.995 137.930 151.295 ;
        RECT 138.460 151.265 138.780 152.225 ;
        RECT 135.685 150.595 136.020 150.765 ;
        RECT 136.215 150.595 136.890 150.765 ;
        RECT 137.210 150.315 137.580 150.815 ;
        RECT 137.760 150.765 137.930 150.995 ;
        RECT 138.315 150.935 138.780 151.265 ;
        RECT 138.950 151.555 139.120 152.395 ;
        RECT 139.300 152.365 139.615 152.865 ;
        RECT 139.845 152.135 140.185 152.695 ;
        RECT 139.290 151.760 140.185 152.135 ;
        RECT 140.355 151.855 140.525 152.865 ;
        RECT 139.995 151.555 140.185 151.760 ;
        RECT 140.695 151.805 141.025 152.650 ;
        RECT 140.695 151.725 141.085 151.805 ;
        RECT 140.870 151.675 141.085 151.725 ;
        RECT 138.950 151.225 139.825 151.555 ;
        RECT 139.995 151.225 140.745 151.555 ;
        RECT 138.950 150.765 139.120 151.225 ;
        RECT 139.995 151.055 140.195 151.225 ;
        RECT 140.915 151.095 141.085 151.675 ;
        RECT 141.715 151.775 142.925 152.865 ;
        RECT 141.715 151.235 142.235 151.775 ;
        RECT 140.860 151.055 141.085 151.095 ;
        RECT 142.405 151.065 142.925 151.605 ;
        RECT 137.760 150.595 138.165 150.765 ;
        RECT 138.335 150.595 139.120 150.765 ;
        RECT 139.395 150.315 139.605 150.845 ;
        RECT 139.865 150.530 140.195 151.055 ;
        RECT 140.705 150.970 141.085 151.055 ;
        RECT 140.365 150.315 140.535 150.925 ;
        RECT 140.705 150.535 141.035 150.970 ;
        RECT 141.715 150.315 142.925 151.065 ;
        RECT 17.430 150.145 143.010 150.315 ;
        RECT 17.515 149.395 18.725 150.145 ;
        RECT 18.985 149.595 19.155 149.975 ;
        RECT 19.370 149.765 19.700 150.145 ;
        RECT 18.985 149.425 19.700 149.595 ;
        RECT 17.515 148.855 18.035 149.395 ;
        RECT 18.205 148.685 18.725 149.225 ;
        RECT 18.895 148.875 19.250 149.245 ;
        RECT 19.530 149.235 19.700 149.425 ;
        RECT 19.870 149.400 20.125 149.975 ;
        RECT 19.530 148.905 19.785 149.235 ;
        RECT 19.530 148.695 19.700 148.905 ;
        RECT 17.515 147.595 18.725 148.685 ;
        RECT 18.985 148.525 19.700 148.695 ;
        RECT 19.955 148.670 20.125 149.400 ;
        RECT 20.300 149.305 20.560 150.145 ;
        RECT 20.735 149.375 23.325 150.145 ;
        RECT 23.585 149.595 23.755 149.885 ;
        RECT 23.925 149.765 24.255 150.145 ;
        RECT 23.585 149.425 24.250 149.595 ;
        RECT 20.735 148.855 21.945 149.375 ;
        RECT 18.985 147.765 19.155 148.525 ;
        RECT 19.370 147.595 19.700 148.355 ;
        RECT 19.870 147.765 20.125 148.670 ;
        RECT 20.300 147.595 20.560 148.745 ;
        RECT 22.115 148.685 23.325 149.205 ;
        RECT 20.735 147.595 23.325 148.685 ;
        RECT 23.500 148.605 23.850 149.255 ;
        RECT 24.020 148.435 24.250 149.425 ;
        RECT 23.585 148.265 24.250 148.435 ;
        RECT 23.585 147.765 23.755 148.265 ;
        RECT 23.925 147.595 24.255 148.095 ;
        RECT 24.425 147.765 24.610 149.885 ;
        RECT 24.865 149.685 25.115 150.145 ;
        RECT 25.285 149.695 25.620 149.865 ;
        RECT 25.815 149.695 26.490 149.865 ;
        RECT 25.285 149.555 25.455 149.695 ;
        RECT 24.780 148.565 25.060 149.515 ;
        RECT 25.230 149.425 25.455 149.555 ;
        RECT 25.230 148.320 25.400 149.425 ;
        RECT 25.625 149.275 26.150 149.495 ;
        RECT 25.570 148.510 25.810 149.105 ;
        RECT 25.980 148.575 26.150 149.275 ;
        RECT 26.320 148.915 26.490 149.695 ;
        RECT 26.810 149.645 27.180 150.145 ;
        RECT 27.360 149.695 27.765 149.865 ;
        RECT 27.935 149.695 28.720 149.865 ;
        RECT 27.360 149.465 27.530 149.695 ;
        RECT 26.700 149.165 27.530 149.465 ;
        RECT 27.915 149.195 28.380 149.525 ;
        RECT 26.700 149.135 26.900 149.165 ;
        RECT 27.020 148.915 27.190 148.985 ;
        RECT 26.320 148.745 27.190 148.915 ;
        RECT 26.680 148.655 27.190 148.745 ;
        RECT 25.230 148.190 25.535 148.320 ;
        RECT 25.980 148.210 26.510 148.575 ;
        RECT 24.850 147.595 25.115 148.055 ;
        RECT 25.285 147.765 25.535 148.190 ;
        RECT 26.680 148.040 26.850 148.655 ;
        RECT 25.745 147.870 26.850 148.040 ;
        RECT 27.020 147.595 27.190 148.395 ;
        RECT 27.360 148.095 27.530 149.165 ;
        RECT 27.700 148.265 27.890 148.985 ;
        RECT 28.060 148.235 28.380 149.195 ;
        RECT 28.550 149.235 28.720 149.695 ;
        RECT 28.995 149.615 29.205 150.145 ;
        RECT 29.465 149.405 29.795 149.930 ;
        RECT 29.965 149.535 30.135 150.145 ;
        RECT 30.305 149.490 30.635 149.925 ;
        RECT 31.775 149.505 32.115 149.910 ;
        RECT 32.285 149.675 32.455 150.145 ;
        RECT 32.625 149.505 32.875 149.910 ;
        RECT 30.305 149.405 30.685 149.490 ;
        RECT 29.595 149.235 29.795 149.405 ;
        RECT 30.460 149.365 30.685 149.405 ;
        RECT 28.550 148.905 29.425 149.235 ;
        RECT 29.595 148.905 30.345 149.235 ;
        RECT 27.360 147.765 27.610 148.095 ;
        RECT 28.550 148.065 28.720 148.905 ;
        RECT 29.595 148.700 29.785 148.905 ;
        RECT 30.515 148.785 30.685 149.365 ;
        RECT 31.775 149.325 32.875 149.505 ;
        RECT 33.045 149.540 33.295 149.910 ;
        RECT 33.465 149.665 33.910 149.835 ;
        RECT 34.080 149.805 34.300 149.850 ;
        RECT 33.045 149.155 33.215 149.540 ;
        RECT 30.470 148.735 30.685 148.785 ;
        RECT 28.890 148.325 29.785 148.700 ;
        RECT 30.295 148.655 30.685 148.735 ;
        RECT 27.835 147.895 28.720 148.065 ;
        RECT 28.900 147.595 29.215 148.095 ;
        RECT 29.445 147.765 29.785 148.325 ;
        RECT 29.955 147.595 30.125 148.605 ;
        RECT 30.295 147.810 30.625 148.655 ;
        RECT 31.775 148.585 32.120 149.155 ;
        RECT 32.290 148.905 32.850 149.155 ;
        RECT 33.020 148.985 33.215 149.155 ;
        RECT 31.775 147.595 32.120 148.415 ;
        RECT 32.290 147.805 32.465 148.905 ;
        RECT 33.020 148.735 33.190 148.985 ;
        RECT 33.465 148.875 33.635 149.665 ;
        RECT 34.080 149.635 34.305 149.805 ;
        RECT 34.080 149.495 34.300 149.635 ;
        RECT 33.805 149.325 34.300 149.495 ;
        RECT 34.580 149.480 34.750 150.145 ;
        RECT 34.945 149.405 35.285 149.975 ;
        RECT 33.805 149.130 33.980 149.325 ;
        RECT 34.150 148.955 34.600 149.155 ;
        RECT 32.635 148.345 33.190 148.735 ;
        RECT 33.360 148.735 33.635 148.875 ;
        RECT 34.770 148.785 34.940 149.235 ;
        RECT 33.360 148.515 34.375 148.735 ;
        RECT 34.545 148.615 34.940 148.785 ;
        RECT 34.545 148.345 34.715 148.615 ;
        RECT 35.110 148.435 35.285 149.405 ;
        RECT 35.455 149.375 38.965 150.145 ;
        RECT 40.060 149.640 40.395 150.145 ;
        RECT 40.565 149.575 40.805 149.950 ;
        RECT 41.085 149.815 41.255 149.960 ;
        RECT 41.085 149.620 41.460 149.815 ;
        RECT 41.820 149.650 42.215 150.145 ;
        RECT 35.455 148.855 37.105 149.375 ;
        RECT 37.275 148.685 38.965 149.205 ;
        RECT 32.635 148.175 34.715 148.345 ;
        RECT 32.635 147.940 32.965 148.175 ;
        RECT 33.255 147.595 33.655 147.995 ;
        RECT 34.525 147.595 34.855 147.995 ;
        RECT 35.025 147.765 35.285 148.435 ;
        RECT 35.455 147.595 38.965 148.685 ;
        RECT 40.115 148.615 40.415 149.465 ;
        RECT 40.585 149.425 40.805 149.575 ;
        RECT 40.585 149.095 41.120 149.425 ;
        RECT 41.290 149.285 41.460 149.620 ;
        RECT 42.385 149.455 42.625 149.975 ;
        RECT 40.585 148.445 40.820 149.095 ;
        RECT 41.290 148.925 42.275 149.285 ;
        RECT 40.145 148.215 40.820 148.445 ;
        RECT 40.990 148.905 42.275 148.925 ;
        RECT 40.990 148.755 41.850 148.905 ;
        RECT 40.145 147.785 40.315 148.215 ;
        RECT 40.485 147.595 40.815 148.045 ;
        RECT 40.990 147.810 41.275 148.755 ;
        RECT 42.450 148.650 42.625 149.455 ;
        RECT 43.275 149.420 43.565 150.145 ;
        RECT 43.900 149.635 44.140 150.145 ;
        RECT 44.320 149.635 44.600 149.965 ;
        RECT 44.830 149.635 45.045 150.145 ;
        RECT 43.795 148.905 44.150 149.465 ;
        RECT 41.450 148.275 42.145 148.585 ;
        RECT 41.455 147.595 42.140 148.065 ;
        RECT 42.320 147.865 42.625 148.650 ;
        RECT 43.275 147.595 43.565 148.760 ;
        RECT 44.320 148.735 44.490 149.635 ;
        RECT 44.660 148.905 44.925 149.465 ;
        RECT 45.215 149.405 45.830 149.975 ;
        RECT 46.035 149.600 51.380 150.145 ;
        RECT 51.555 149.600 56.900 150.145 ;
        RECT 57.075 149.600 62.420 150.145 ;
        RECT 62.595 149.600 67.940 150.145 ;
        RECT 45.175 148.735 45.345 149.235 ;
        RECT 43.920 148.565 45.345 148.735 ;
        RECT 43.920 148.390 44.310 148.565 ;
        RECT 44.795 147.595 45.125 148.395 ;
        RECT 45.515 148.385 45.830 149.405 ;
        RECT 47.620 148.770 47.960 149.600 ;
        RECT 45.295 147.765 45.830 148.385 ;
        RECT 49.440 148.030 49.790 149.280 ;
        RECT 53.140 148.770 53.480 149.600 ;
        RECT 54.960 148.030 55.310 149.280 ;
        RECT 58.660 148.770 59.000 149.600 ;
        RECT 60.480 148.030 60.830 149.280 ;
        RECT 64.180 148.770 64.520 149.600 ;
        RECT 69.035 149.420 69.325 150.145 ;
        RECT 69.585 149.595 69.755 149.885 ;
        RECT 69.925 149.765 70.255 150.145 ;
        RECT 69.585 149.425 70.250 149.595 ;
        RECT 66.000 148.030 66.350 149.280 ;
        RECT 46.035 147.595 51.380 148.030 ;
        RECT 51.555 147.595 56.900 148.030 ;
        RECT 57.075 147.595 62.420 148.030 ;
        RECT 62.595 147.595 67.940 148.030 ;
        RECT 69.035 147.595 69.325 148.760 ;
        RECT 69.500 148.605 69.850 149.255 ;
        RECT 70.020 148.435 70.250 149.425 ;
        RECT 69.585 148.265 70.250 148.435 ;
        RECT 69.585 147.765 69.755 148.265 ;
        RECT 69.925 147.595 70.255 148.095 ;
        RECT 70.425 147.765 70.610 149.885 ;
        RECT 70.865 149.685 71.115 150.145 ;
        RECT 71.285 149.695 71.620 149.865 ;
        RECT 71.815 149.695 72.490 149.865 ;
        RECT 71.285 149.555 71.455 149.695 ;
        RECT 70.780 148.565 71.060 149.515 ;
        RECT 71.230 149.425 71.455 149.555 ;
        RECT 71.230 148.320 71.400 149.425 ;
        RECT 71.625 149.275 72.150 149.495 ;
        RECT 71.570 148.510 71.810 149.105 ;
        RECT 71.980 148.575 72.150 149.275 ;
        RECT 72.320 148.915 72.490 149.695 ;
        RECT 72.810 149.645 73.180 150.145 ;
        RECT 73.360 149.695 73.765 149.865 ;
        RECT 73.935 149.695 74.720 149.865 ;
        RECT 73.360 149.465 73.530 149.695 ;
        RECT 72.700 149.165 73.530 149.465 ;
        RECT 73.915 149.195 74.380 149.525 ;
        RECT 72.700 149.135 72.900 149.165 ;
        RECT 73.020 148.915 73.190 148.985 ;
        RECT 72.320 148.745 73.190 148.915 ;
        RECT 72.680 148.655 73.190 148.745 ;
        RECT 71.230 148.190 71.535 148.320 ;
        RECT 71.980 148.210 72.510 148.575 ;
        RECT 70.850 147.595 71.115 148.055 ;
        RECT 71.285 147.765 71.535 148.190 ;
        RECT 72.680 148.040 72.850 148.655 ;
        RECT 71.745 147.870 72.850 148.040 ;
        RECT 73.020 147.595 73.190 148.395 ;
        RECT 73.360 148.095 73.530 149.165 ;
        RECT 73.700 148.265 73.890 148.985 ;
        RECT 74.060 148.235 74.380 149.195 ;
        RECT 74.550 149.235 74.720 149.695 ;
        RECT 74.995 149.615 75.205 150.145 ;
        RECT 75.465 149.405 75.795 149.930 ;
        RECT 75.965 149.535 76.135 150.145 ;
        RECT 76.305 149.490 76.635 149.925 ;
        RECT 76.305 149.405 76.685 149.490 ;
        RECT 75.595 149.235 75.795 149.405 ;
        RECT 76.460 149.365 76.685 149.405 ;
        RECT 74.550 148.905 75.425 149.235 ;
        RECT 75.595 148.905 76.345 149.235 ;
        RECT 73.360 147.765 73.610 148.095 ;
        RECT 74.550 148.065 74.720 148.905 ;
        RECT 75.595 148.700 75.785 148.905 ;
        RECT 76.515 148.785 76.685 149.365 ;
        RECT 76.470 148.735 76.685 148.785 ;
        RECT 74.890 148.325 75.785 148.700 ;
        RECT 76.295 148.655 76.685 148.735 ;
        RECT 76.860 149.405 77.115 149.975 ;
        RECT 77.285 149.745 77.615 150.145 ;
        RECT 78.040 149.610 78.570 149.975 ;
        RECT 78.040 149.575 78.215 149.610 ;
        RECT 77.285 149.405 78.215 149.575 ;
        RECT 76.860 148.735 77.030 149.405 ;
        RECT 77.285 149.235 77.455 149.405 ;
        RECT 77.200 148.905 77.455 149.235 ;
        RECT 77.680 148.905 77.875 149.235 ;
        RECT 73.835 147.895 74.720 148.065 ;
        RECT 74.900 147.595 75.215 148.095 ;
        RECT 75.445 147.765 75.785 148.325 ;
        RECT 75.955 147.595 76.125 148.605 ;
        RECT 76.295 147.810 76.625 148.655 ;
        RECT 76.860 147.765 77.195 148.735 ;
        RECT 77.365 147.595 77.535 148.735 ;
        RECT 77.705 147.935 77.875 148.905 ;
        RECT 78.045 148.275 78.215 149.405 ;
        RECT 78.385 148.615 78.555 149.415 ;
        RECT 78.760 149.125 79.035 149.975 ;
        RECT 78.755 148.955 79.035 149.125 ;
        RECT 78.760 148.815 79.035 148.955 ;
        RECT 79.205 148.615 79.395 149.975 ;
        RECT 79.575 149.610 80.085 150.145 ;
        RECT 80.305 149.335 80.550 149.940 ;
        RECT 80.995 149.405 81.380 149.975 ;
        RECT 81.550 149.685 81.875 150.145 ;
        RECT 82.395 149.515 82.675 149.975 ;
        RECT 79.595 149.165 80.825 149.335 ;
        RECT 78.385 148.445 79.395 148.615 ;
        RECT 79.565 148.600 80.315 148.790 ;
        RECT 78.045 148.105 79.170 148.275 ;
        RECT 79.565 147.935 79.735 148.600 ;
        RECT 80.485 148.355 80.825 149.165 ;
        RECT 77.705 147.765 79.735 147.935 ;
        RECT 79.905 147.595 80.075 148.355 ;
        RECT 80.310 147.945 80.825 148.355 ;
        RECT 80.995 148.735 81.275 149.405 ;
        RECT 81.550 149.345 82.675 149.515 ;
        RECT 81.550 149.235 82.000 149.345 ;
        RECT 81.445 148.905 82.000 149.235 ;
        RECT 82.865 149.175 83.265 149.975 ;
        RECT 83.665 149.685 83.935 150.145 ;
        RECT 84.105 149.515 84.390 149.975 ;
        RECT 84.675 149.600 90.020 150.145 ;
        RECT 80.995 147.765 81.380 148.735 ;
        RECT 81.550 148.445 82.000 148.905 ;
        RECT 82.170 148.615 83.265 149.175 ;
        RECT 81.550 148.225 82.675 148.445 ;
        RECT 81.550 147.595 81.875 148.055 ;
        RECT 82.395 147.765 82.675 148.225 ;
        RECT 82.865 147.765 83.265 148.615 ;
        RECT 83.435 149.345 84.390 149.515 ;
        RECT 83.435 148.445 83.645 149.345 ;
        RECT 83.815 148.615 84.505 149.175 ;
        RECT 86.260 148.770 86.600 149.600 ;
        RECT 90.195 149.375 93.705 150.145 ;
        RECT 94.795 149.420 95.085 150.145 ;
        RECT 95.255 149.395 96.465 150.145 ;
        RECT 96.725 149.595 96.895 149.885 ;
        RECT 97.065 149.765 97.395 150.145 ;
        RECT 96.725 149.425 97.390 149.595 ;
        RECT 83.435 148.225 84.390 148.445 ;
        RECT 83.665 147.595 83.935 148.055 ;
        RECT 84.105 147.765 84.390 148.225 ;
        RECT 88.080 148.030 88.430 149.280 ;
        RECT 90.195 148.855 91.845 149.375 ;
        RECT 92.015 148.685 93.705 149.205 ;
        RECT 95.255 148.855 95.775 149.395 ;
        RECT 84.675 147.595 90.020 148.030 ;
        RECT 90.195 147.595 93.705 148.685 ;
        RECT 94.795 147.595 95.085 148.760 ;
        RECT 95.945 148.685 96.465 149.225 ;
        RECT 95.255 147.595 96.465 148.685 ;
        RECT 96.640 148.605 96.990 149.255 ;
        RECT 97.160 148.435 97.390 149.425 ;
        RECT 96.725 148.265 97.390 148.435 ;
        RECT 96.725 147.765 96.895 148.265 ;
        RECT 97.065 147.595 97.395 148.095 ;
        RECT 97.565 147.765 97.750 149.885 ;
        RECT 98.005 149.685 98.255 150.145 ;
        RECT 98.425 149.695 98.760 149.865 ;
        RECT 98.955 149.695 99.630 149.865 ;
        RECT 98.425 149.555 98.595 149.695 ;
        RECT 97.920 148.565 98.200 149.515 ;
        RECT 98.370 149.425 98.595 149.555 ;
        RECT 98.370 148.320 98.540 149.425 ;
        RECT 98.765 149.275 99.290 149.495 ;
        RECT 98.710 148.510 98.950 149.105 ;
        RECT 99.120 148.575 99.290 149.275 ;
        RECT 99.460 148.915 99.630 149.695 ;
        RECT 99.950 149.645 100.320 150.145 ;
        RECT 100.500 149.695 100.905 149.865 ;
        RECT 101.075 149.695 101.860 149.865 ;
        RECT 100.500 149.465 100.670 149.695 ;
        RECT 99.840 149.165 100.670 149.465 ;
        RECT 101.055 149.195 101.520 149.525 ;
        RECT 99.840 149.135 100.040 149.165 ;
        RECT 100.160 148.915 100.330 148.985 ;
        RECT 99.460 148.745 100.330 148.915 ;
        RECT 99.820 148.655 100.330 148.745 ;
        RECT 98.370 148.190 98.675 148.320 ;
        RECT 99.120 148.210 99.650 148.575 ;
        RECT 97.990 147.595 98.255 148.055 ;
        RECT 98.425 147.765 98.675 148.190 ;
        RECT 99.820 148.040 99.990 148.655 ;
        RECT 98.885 147.870 99.990 148.040 ;
        RECT 100.160 147.595 100.330 148.395 ;
        RECT 100.500 148.095 100.670 149.165 ;
        RECT 100.840 148.265 101.030 148.985 ;
        RECT 101.200 148.235 101.520 149.195 ;
        RECT 101.690 149.235 101.860 149.695 ;
        RECT 102.135 149.615 102.345 150.145 ;
        RECT 102.605 149.405 102.935 149.930 ;
        RECT 103.105 149.535 103.275 150.145 ;
        RECT 103.445 149.490 103.775 149.925 ;
        RECT 104.965 149.490 105.295 149.925 ;
        RECT 105.465 149.535 105.635 150.145 ;
        RECT 103.445 149.405 103.825 149.490 ;
        RECT 102.735 149.235 102.935 149.405 ;
        RECT 103.600 149.365 103.825 149.405 ;
        RECT 101.690 148.905 102.565 149.235 ;
        RECT 102.735 148.905 103.485 149.235 ;
        RECT 100.500 147.765 100.750 148.095 ;
        RECT 101.690 148.065 101.860 148.905 ;
        RECT 102.735 148.700 102.925 148.905 ;
        RECT 103.655 148.785 103.825 149.365 ;
        RECT 103.610 148.735 103.825 148.785 ;
        RECT 102.030 148.325 102.925 148.700 ;
        RECT 103.435 148.655 103.825 148.735 ;
        RECT 104.915 149.405 105.295 149.490 ;
        RECT 105.805 149.405 106.135 149.930 ;
        RECT 106.395 149.615 106.605 150.145 ;
        RECT 106.880 149.695 107.665 149.865 ;
        RECT 107.835 149.695 108.240 149.865 ;
        RECT 104.915 149.365 105.140 149.405 ;
        RECT 104.915 148.785 105.085 149.365 ;
        RECT 105.805 149.235 106.005 149.405 ;
        RECT 106.880 149.235 107.050 149.695 ;
        RECT 105.255 148.905 106.005 149.235 ;
        RECT 106.175 148.905 107.050 149.235 ;
        RECT 104.915 148.735 105.130 148.785 ;
        RECT 104.915 148.655 105.305 148.735 ;
        RECT 100.975 147.895 101.860 148.065 ;
        RECT 102.040 147.595 102.355 148.095 ;
        RECT 102.585 147.765 102.925 148.325 ;
        RECT 103.095 147.595 103.265 148.605 ;
        RECT 103.435 147.810 103.765 148.655 ;
        RECT 104.975 147.810 105.305 148.655 ;
        RECT 105.815 148.700 106.005 148.905 ;
        RECT 105.475 147.595 105.645 148.605 ;
        RECT 105.815 148.325 106.710 148.700 ;
        RECT 105.815 147.765 106.155 148.325 ;
        RECT 106.385 147.595 106.700 148.095 ;
        RECT 106.880 148.065 107.050 148.905 ;
        RECT 107.220 149.195 107.685 149.525 ;
        RECT 108.070 149.465 108.240 149.695 ;
        RECT 108.420 149.645 108.790 150.145 ;
        RECT 109.110 149.695 109.785 149.865 ;
        RECT 109.980 149.695 110.315 149.865 ;
        RECT 107.220 148.235 107.540 149.195 ;
        RECT 108.070 149.165 108.900 149.465 ;
        RECT 107.710 148.265 107.900 148.985 ;
        RECT 108.070 148.095 108.240 149.165 ;
        RECT 108.700 149.135 108.900 149.165 ;
        RECT 108.410 148.915 108.580 148.985 ;
        RECT 109.110 148.915 109.280 149.695 ;
        RECT 110.145 149.555 110.315 149.695 ;
        RECT 110.485 149.685 110.735 150.145 ;
        RECT 108.410 148.745 109.280 148.915 ;
        RECT 109.450 149.275 109.975 149.495 ;
        RECT 110.145 149.425 110.370 149.555 ;
        RECT 108.410 148.655 108.920 148.745 ;
        RECT 106.880 147.895 107.765 148.065 ;
        RECT 107.990 147.765 108.240 148.095 ;
        RECT 108.410 147.595 108.580 148.395 ;
        RECT 108.750 148.040 108.920 148.655 ;
        RECT 109.450 148.575 109.620 149.275 ;
        RECT 109.090 148.210 109.620 148.575 ;
        RECT 109.790 148.510 110.030 149.105 ;
        RECT 110.200 148.320 110.370 149.425 ;
        RECT 110.540 148.565 110.820 149.515 ;
        RECT 110.065 148.190 110.370 148.320 ;
        RECT 108.750 147.870 109.855 148.040 ;
        RECT 110.065 147.765 110.315 148.190 ;
        RECT 110.485 147.595 110.750 148.055 ;
        RECT 110.990 147.765 111.175 149.885 ;
        RECT 111.345 149.765 111.675 150.145 ;
        RECT 111.845 149.595 112.015 149.885 ;
        RECT 111.350 149.425 112.015 149.595 ;
        RECT 113.245 149.490 113.575 149.925 ;
        RECT 113.745 149.535 113.915 150.145 ;
        RECT 111.350 148.435 111.580 149.425 ;
        RECT 113.195 149.405 113.575 149.490 ;
        RECT 114.085 149.405 114.415 149.930 ;
        RECT 114.675 149.615 114.885 150.145 ;
        RECT 115.160 149.695 115.945 149.865 ;
        RECT 116.115 149.695 116.520 149.865 ;
        RECT 113.195 149.365 113.420 149.405 ;
        RECT 111.750 148.605 112.100 149.255 ;
        RECT 113.195 148.785 113.365 149.365 ;
        RECT 114.085 149.235 114.285 149.405 ;
        RECT 115.160 149.235 115.330 149.695 ;
        RECT 113.535 148.905 114.285 149.235 ;
        RECT 114.455 148.905 115.330 149.235 ;
        RECT 113.195 148.735 113.410 148.785 ;
        RECT 113.195 148.655 113.585 148.735 ;
        RECT 111.350 148.265 112.015 148.435 ;
        RECT 111.345 147.595 111.675 148.095 ;
        RECT 111.845 147.765 112.015 148.265 ;
        RECT 113.255 147.810 113.585 148.655 ;
        RECT 114.095 148.700 114.285 148.905 ;
        RECT 113.755 147.595 113.925 148.605 ;
        RECT 114.095 148.325 114.990 148.700 ;
        RECT 114.095 147.765 114.435 148.325 ;
        RECT 114.665 147.595 114.980 148.095 ;
        RECT 115.160 148.065 115.330 148.905 ;
        RECT 115.500 149.195 115.965 149.525 ;
        RECT 116.350 149.465 116.520 149.695 ;
        RECT 116.700 149.645 117.070 150.145 ;
        RECT 117.390 149.695 118.065 149.865 ;
        RECT 118.260 149.695 118.595 149.865 ;
        RECT 115.500 148.235 115.820 149.195 ;
        RECT 116.350 149.165 117.180 149.465 ;
        RECT 115.990 148.265 116.180 148.985 ;
        RECT 116.350 148.095 116.520 149.165 ;
        RECT 116.980 149.135 117.180 149.165 ;
        RECT 116.690 148.915 116.860 148.985 ;
        RECT 117.390 148.915 117.560 149.695 ;
        RECT 118.425 149.555 118.595 149.695 ;
        RECT 118.765 149.685 119.015 150.145 ;
        RECT 116.690 148.745 117.560 148.915 ;
        RECT 117.730 149.275 118.255 149.495 ;
        RECT 118.425 149.425 118.650 149.555 ;
        RECT 116.690 148.655 117.200 148.745 ;
        RECT 115.160 147.895 116.045 148.065 ;
        RECT 116.270 147.765 116.520 148.095 ;
        RECT 116.690 147.595 116.860 148.395 ;
        RECT 117.030 148.040 117.200 148.655 ;
        RECT 117.730 148.575 117.900 149.275 ;
        RECT 117.370 148.210 117.900 148.575 ;
        RECT 118.070 148.510 118.310 149.105 ;
        RECT 118.480 148.320 118.650 149.425 ;
        RECT 118.820 148.565 119.100 149.515 ;
        RECT 118.345 148.190 118.650 148.320 ;
        RECT 117.030 147.870 118.135 148.040 ;
        RECT 118.345 147.765 118.595 148.190 ;
        RECT 118.765 147.595 119.030 148.055 ;
        RECT 119.270 147.765 119.455 149.885 ;
        RECT 119.625 149.765 119.955 150.145 ;
        RECT 120.125 149.595 120.295 149.885 ;
        RECT 119.630 149.425 120.295 149.595 ;
        RECT 119.630 148.435 119.860 149.425 ;
        RECT 120.555 149.420 120.845 150.145 ;
        RECT 121.015 149.345 121.325 150.145 ;
        RECT 121.530 149.345 122.225 149.975 ;
        RECT 123.320 149.380 123.775 150.145 ;
        RECT 124.050 149.765 125.350 149.975 ;
        RECT 125.605 149.785 125.935 150.145 ;
        RECT 125.180 149.615 125.350 149.765 ;
        RECT 126.105 149.645 126.365 149.975 ;
        RECT 126.135 149.635 126.365 149.645 ;
        RECT 120.030 148.605 120.380 149.255 ;
        RECT 121.025 148.905 121.360 149.175 ;
        RECT 121.530 148.785 121.700 149.345 ;
        RECT 124.250 149.155 124.470 149.555 ;
        RECT 121.870 148.905 122.205 149.155 ;
        RECT 123.315 148.955 123.805 149.155 ;
        RECT 123.995 148.945 124.470 149.155 ;
        RECT 124.715 149.155 124.925 149.555 ;
        RECT 125.180 149.490 125.935 149.615 ;
        RECT 125.180 149.445 126.025 149.490 ;
        RECT 125.755 149.325 126.025 149.445 ;
        RECT 124.715 148.945 125.045 149.155 ;
        RECT 125.215 148.885 125.625 149.190 ;
        RECT 119.630 148.265 120.295 148.435 ;
        RECT 119.625 147.595 119.955 148.095 ;
        RECT 120.125 147.765 120.295 148.265 ;
        RECT 120.555 147.595 120.845 148.760 ;
        RECT 121.530 148.745 121.705 148.785 ;
        RECT 121.015 147.595 121.295 148.735 ;
        RECT 121.465 147.765 121.795 148.745 ;
        RECT 121.965 147.595 122.225 148.735 ;
        RECT 123.320 148.715 124.495 148.775 ;
        RECT 125.855 148.750 126.025 149.325 ;
        RECT 125.825 148.715 126.025 148.750 ;
        RECT 123.320 148.605 126.025 148.715 ;
        RECT 123.320 147.985 123.575 148.605 ;
        RECT 124.165 148.545 125.965 148.605 ;
        RECT 124.165 148.515 124.495 148.545 ;
        RECT 126.195 148.445 126.365 149.635 ;
        RECT 126.540 149.380 126.995 150.145 ;
        RECT 127.270 149.765 128.570 149.975 ;
        RECT 128.825 149.785 129.155 150.145 ;
        RECT 128.400 149.615 128.570 149.765 ;
        RECT 129.325 149.645 129.585 149.975 ;
        RECT 127.470 149.155 127.690 149.555 ;
        RECT 126.535 148.955 127.025 149.155 ;
        RECT 127.215 148.945 127.690 149.155 ;
        RECT 127.935 149.155 128.145 149.555 ;
        RECT 128.400 149.490 129.155 149.615 ;
        RECT 128.400 149.445 129.245 149.490 ;
        RECT 128.975 149.325 129.245 149.445 ;
        RECT 127.935 148.945 128.265 149.155 ;
        RECT 128.435 148.885 128.845 149.190 ;
        RECT 123.825 148.345 124.010 148.435 ;
        RECT 124.600 148.345 125.435 148.355 ;
        RECT 123.825 148.145 125.435 148.345 ;
        RECT 123.825 148.105 124.055 148.145 ;
        RECT 123.320 147.765 123.655 147.985 ;
        RECT 124.660 147.595 125.015 147.975 ;
        RECT 125.185 147.765 125.435 148.145 ;
        RECT 125.685 147.595 125.935 148.375 ;
        RECT 126.105 147.765 126.365 148.445 ;
        RECT 126.540 148.715 127.715 148.775 ;
        RECT 129.075 148.750 129.245 149.325 ;
        RECT 129.045 148.715 129.245 148.750 ;
        RECT 126.540 148.605 129.245 148.715 ;
        RECT 126.540 147.985 126.795 148.605 ;
        RECT 127.385 148.545 129.185 148.605 ;
        RECT 127.385 148.515 127.715 148.545 ;
        RECT 129.415 148.445 129.585 149.645 ;
        RECT 129.760 149.380 130.215 150.145 ;
        RECT 130.490 149.765 131.790 149.975 ;
        RECT 132.045 149.785 132.375 150.145 ;
        RECT 131.620 149.615 131.790 149.765 ;
        RECT 132.545 149.645 132.805 149.975 ;
        RECT 130.690 149.155 130.910 149.555 ;
        RECT 129.755 148.955 130.245 149.155 ;
        RECT 130.435 148.945 130.910 149.155 ;
        RECT 131.155 149.155 131.365 149.555 ;
        RECT 131.620 149.490 132.375 149.615 ;
        RECT 131.620 149.445 132.465 149.490 ;
        RECT 132.195 149.325 132.465 149.445 ;
        RECT 131.155 148.945 131.485 149.155 ;
        RECT 131.655 148.885 132.065 149.190 ;
        RECT 127.045 148.345 127.230 148.435 ;
        RECT 127.820 148.345 128.655 148.355 ;
        RECT 127.045 148.145 128.655 148.345 ;
        RECT 127.045 148.105 127.275 148.145 ;
        RECT 126.540 147.765 126.875 147.985 ;
        RECT 127.880 147.595 128.235 147.975 ;
        RECT 128.405 147.765 128.655 148.145 ;
        RECT 128.905 147.595 129.155 148.375 ;
        RECT 129.325 147.765 129.585 148.445 ;
        RECT 129.760 148.715 130.935 148.775 ;
        RECT 132.295 148.750 132.465 149.325 ;
        RECT 132.265 148.715 132.465 148.750 ;
        RECT 129.760 148.605 132.465 148.715 ;
        RECT 129.760 147.985 130.015 148.605 ;
        RECT 130.605 148.545 132.405 148.605 ;
        RECT 130.605 148.515 130.935 148.545 ;
        RECT 132.635 148.445 132.805 149.645 ;
        RECT 132.975 149.375 134.645 150.145 ;
        RECT 134.905 149.595 135.075 149.975 ;
        RECT 135.255 149.765 135.585 150.145 ;
        RECT 134.905 149.425 135.570 149.595 ;
        RECT 135.765 149.470 136.025 149.975 ;
        RECT 132.975 148.855 133.725 149.375 ;
        RECT 133.895 148.685 134.645 149.205 ;
        RECT 134.835 148.875 135.165 149.245 ;
        RECT 135.400 149.170 135.570 149.425 ;
        RECT 135.400 148.840 135.685 149.170 ;
        RECT 135.400 148.695 135.570 148.840 ;
        RECT 130.265 148.345 130.450 148.435 ;
        RECT 131.040 148.345 131.875 148.355 ;
        RECT 130.265 148.145 131.875 148.345 ;
        RECT 130.265 148.105 130.495 148.145 ;
        RECT 129.760 147.765 130.095 147.985 ;
        RECT 131.100 147.595 131.455 147.975 ;
        RECT 131.625 147.765 131.875 148.145 ;
        RECT 132.125 147.595 132.375 148.375 ;
        RECT 132.545 147.765 132.805 148.445 ;
        RECT 132.975 147.595 134.645 148.685 ;
        RECT 134.905 148.525 135.570 148.695 ;
        RECT 135.855 148.670 136.025 149.470 ;
        RECT 134.905 147.765 135.075 148.525 ;
        RECT 135.255 147.595 135.585 148.355 ;
        RECT 135.755 147.765 136.025 148.670 ;
        RECT 136.195 149.405 136.580 149.975 ;
        RECT 136.750 149.685 137.075 150.145 ;
        RECT 137.595 149.515 137.875 149.975 ;
        RECT 136.195 148.735 136.475 149.405 ;
        RECT 136.750 149.345 137.875 149.515 ;
        RECT 136.750 149.235 137.200 149.345 ;
        RECT 136.645 148.905 137.200 149.235 ;
        RECT 138.065 149.175 138.465 149.975 ;
        RECT 138.865 149.685 139.135 150.145 ;
        RECT 139.305 149.515 139.590 149.975 ;
        RECT 136.195 147.765 136.580 148.735 ;
        RECT 136.750 148.445 137.200 148.905 ;
        RECT 137.370 148.615 138.465 149.175 ;
        RECT 136.750 148.225 137.875 148.445 ;
        RECT 136.750 147.595 137.075 148.055 ;
        RECT 137.595 147.765 137.875 148.225 ;
        RECT 138.065 147.765 138.465 148.615 ;
        RECT 138.635 149.345 139.590 149.515 ;
        RECT 139.965 149.595 140.135 149.975 ;
        RECT 140.350 149.765 140.680 150.145 ;
        RECT 139.965 149.425 140.680 149.595 ;
        RECT 138.635 148.445 138.845 149.345 ;
        RECT 139.015 148.615 139.705 149.175 ;
        RECT 139.875 148.875 140.230 149.245 ;
        RECT 140.510 149.235 140.680 149.425 ;
        RECT 140.850 149.400 141.105 149.975 ;
        RECT 140.510 148.905 140.765 149.235 ;
        RECT 140.510 148.695 140.680 148.905 ;
        RECT 139.965 148.525 140.680 148.695 ;
        RECT 140.935 148.670 141.105 149.400 ;
        RECT 141.280 149.305 141.540 150.145 ;
        RECT 141.715 149.395 142.925 150.145 ;
        RECT 138.635 148.225 139.590 148.445 ;
        RECT 138.865 147.595 139.135 148.055 ;
        RECT 139.305 147.765 139.590 148.225 ;
        RECT 139.965 147.765 140.135 148.525 ;
        RECT 140.350 147.595 140.680 148.355 ;
        RECT 140.850 147.765 141.105 148.670 ;
        RECT 141.280 147.595 141.540 148.745 ;
        RECT 141.715 148.685 142.235 149.225 ;
        RECT 142.405 148.855 142.925 149.395 ;
        RECT 141.715 147.595 142.925 148.685 ;
        RECT 17.430 147.425 143.010 147.595 ;
        RECT 17.515 146.335 18.725 147.425 ;
        RECT 17.515 145.625 18.035 146.165 ;
        RECT 18.205 145.795 18.725 146.335 ;
        RECT 18.895 146.455 19.165 147.225 ;
        RECT 19.335 146.645 19.665 147.425 ;
        RECT 19.870 146.820 20.055 147.225 ;
        RECT 20.225 147.000 20.560 147.425 ;
        RECT 19.870 146.645 20.535 146.820 ;
        RECT 18.895 146.285 20.025 146.455 ;
        RECT 17.515 144.875 18.725 145.625 ;
        RECT 18.895 145.375 19.065 146.285 ;
        RECT 19.235 145.535 19.595 146.115 ;
        RECT 19.775 145.785 20.025 146.285 ;
        RECT 20.195 145.615 20.535 146.645 ;
        RECT 20.735 146.335 22.405 147.425 ;
        RECT 19.850 145.445 20.535 145.615 ;
        RECT 20.735 145.645 21.485 146.165 ;
        RECT 21.655 145.815 22.405 146.335 ;
        RECT 22.585 146.285 22.915 147.425 ;
        RECT 23.445 146.455 23.775 147.240 ;
        RECT 23.095 146.285 23.775 146.455 ;
        RECT 23.955 146.555 24.230 147.255 ;
        RECT 24.400 146.880 24.655 147.425 ;
        RECT 24.825 146.915 25.305 147.255 ;
        RECT 25.480 146.870 26.085 147.425 ;
        RECT 25.470 146.770 26.085 146.870 ;
        RECT 25.470 146.745 25.655 146.770 ;
        RECT 22.575 145.865 22.925 146.115 ;
        RECT 23.095 145.685 23.265 146.285 ;
        RECT 23.435 145.865 23.785 146.115 ;
        RECT 18.895 145.045 19.155 145.375 ;
        RECT 19.365 144.875 19.640 145.355 ;
        RECT 19.850 145.045 20.055 145.445 ;
        RECT 20.225 144.875 20.560 145.275 ;
        RECT 20.735 144.875 22.405 145.645 ;
        RECT 22.585 144.875 22.855 145.685 ;
        RECT 23.025 145.045 23.355 145.685 ;
        RECT 23.525 144.875 23.765 145.685 ;
        RECT 23.955 145.525 24.125 146.555 ;
        RECT 24.400 146.425 25.155 146.675 ;
        RECT 25.325 146.500 25.655 146.745 ;
        RECT 24.400 146.390 25.170 146.425 ;
        RECT 24.400 146.380 25.185 146.390 ;
        RECT 24.295 146.365 25.190 146.380 ;
        RECT 24.295 146.350 25.210 146.365 ;
        RECT 24.295 146.340 25.230 146.350 ;
        RECT 24.295 146.330 25.255 146.340 ;
        RECT 24.295 146.300 25.325 146.330 ;
        RECT 24.295 146.270 25.345 146.300 ;
        RECT 24.295 146.240 25.365 146.270 ;
        RECT 24.295 146.215 25.395 146.240 ;
        RECT 24.295 146.180 25.430 146.215 ;
        RECT 24.295 146.175 25.460 146.180 ;
        RECT 24.295 145.780 24.525 146.175 ;
        RECT 25.070 146.170 25.460 146.175 ;
        RECT 25.095 146.160 25.460 146.170 ;
        RECT 25.110 146.155 25.460 146.160 ;
        RECT 25.125 146.150 25.460 146.155 ;
        RECT 25.825 146.150 26.085 146.600 ;
        RECT 26.265 146.455 26.595 147.240 ;
        RECT 26.265 146.285 26.945 146.455 ;
        RECT 27.125 146.285 27.455 147.425 ;
        RECT 27.670 146.635 28.205 147.255 ;
        RECT 25.125 146.145 26.085 146.150 ;
        RECT 25.135 146.135 26.085 146.145 ;
        RECT 25.145 146.130 26.085 146.135 ;
        RECT 25.155 146.120 26.085 146.130 ;
        RECT 25.160 146.110 26.085 146.120 ;
        RECT 25.165 146.105 26.085 146.110 ;
        RECT 25.175 146.090 26.085 146.105 ;
        RECT 25.180 146.075 26.085 146.090 ;
        RECT 25.190 146.050 26.085 146.075 ;
        RECT 24.695 145.580 25.025 146.005 ;
        RECT 24.775 145.555 25.025 145.580 ;
        RECT 23.955 145.045 24.215 145.525 ;
        RECT 24.385 144.875 24.635 145.415 ;
        RECT 24.805 145.095 25.025 145.555 ;
        RECT 25.195 145.980 26.085 146.050 ;
        RECT 25.195 145.255 25.365 145.980 ;
        RECT 26.255 145.865 26.605 146.115 ;
        RECT 25.535 145.425 26.085 145.810 ;
        RECT 26.775 145.685 26.945 146.285 ;
        RECT 27.115 145.865 27.465 146.115 ;
        RECT 25.195 145.085 26.085 145.255 ;
        RECT 26.275 144.875 26.515 145.685 ;
        RECT 26.685 145.045 27.015 145.685 ;
        RECT 27.185 144.875 27.455 145.685 ;
        RECT 27.670 145.615 27.985 146.635 ;
        RECT 28.375 146.625 28.705 147.425 ;
        RECT 29.190 146.455 29.580 146.630 ;
        RECT 28.155 146.285 29.580 146.455 ;
        RECT 28.155 145.785 28.325 146.285 ;
        RECT 27.670 145.045 28.285 145.615 ;
        RECT 28.575 145.555 28.840 146.115 ;
        RECT 29.010 145.385 29.180 146.285 ;
        RECT 30.395 146.260 30.685 147.425 ;
        RECT 30.855 146.995 31.195 147.255 ;
        RECT 29.350 145.555 29.705 146.115 ;
        RECT 28.455 144.875 28.670 145.385 ;
        RECT 28.900 145.055 29.180 145.385 ;
        RECT 29.360 144.875 29.600 145.385 ;
        RECT 30.395 144.875 30.685 145.600 ;
        RECT 30.855 145.595 31.115 146.995 ;
        RECT 31.365 146.625 31.695 147.425 ;
        RECT 32.160 146.455 32.410 147.255 ;
        RECT 32.595 146.705 32.925 147.425 ;
        RECT 33.145 146.455 33.395 147.255 ;
        RECT 33.565 147.045 33.900 147.425 ;
        RECT 31.305 146.285 33.495 146.455 ;
        RECT 31.305 146.115 31.620 146.285 ;
        RECT 31.290 145.865 31.620 146.115 ;
        RECT 30.855 145.085 31.195 145.595 ;
        RECT 31.365 144.875 31.635 145.675 ;
        RECT 31.815 145.145 32.095 146.115 ;
        RECT 32.275 145.145 32.575 146.115 ;
        RECT 32.755 145.150 33.105 146.115 ;
        RECT 33.325 145.375 33.495 146.285 ;
        RECT 33.665 145.555 33.905 146.865 ;
        RECT 34.075 146.335 37.585 147.425 ;
        RECT 39.175 146.965 39.390 147.425 ;
        RECT 39.560 146.795 39.890 147.255 ;
        RECT 34.075 145.645 35.725 146.165 ;
        RECT 35.895 145.815 37.585 146.335 ;
        RECT 38.720 146.625 39.890 146.795 ;
        RECT 40.060 146.625 40.310 147.425 ;
        RECT 33.325 145.045 33.820 145.375 ;
        RECT 34.075 144.875 37.585 145.645 ;
        RECT 38.720 145.335 39.090 146.625 ;
        RECT 40.520 146.455 40.800 146.615 ;
        RECT 39.465 146.285 40.800 146.455 ;
        RECT 40.975 146.335 43.565 147.425 ;
        RECT 43.740 147.000 44.075 147.425 ;
        RECT 44.245 146.820 44.430 147.225 ;
        RECT 39.465 146.115 39.635 146.285 ;
        RECT 39.260 145.865 39.635 146.115 ;
        RECT 39.805 145.865 40.280 146.105 ;
        RECT 40.450 145.865 40.800 146.105 ;
        RECT 39.465 145.695 39.635 145.865 ;
        RECT 39.465 145.525 40.800 145.695 ;
        RECT 38.720 145.045 39.470 145.335 ;
        RECT 39.980 144.875 40.310 145.335 ;
        RECT 40.530 145.315 40.800 145.525 ;
        RECT 40.975 145.645 42.185 146.165 ;
        RECT 42.355 145.815 43.565 146.335 ;
        RECT 43.765 146.645 44.430 146.820 ;
        RECT 44.635 146.645 44.965 147.425 ;
        RECT 40.975 144.875 43.565 145.645 ;
        RECT 43.765 145.615 44.105 146.645 ;
        RECT 45.135 146.455 45.405 147.225 ;
        RECT 44.275 146.285 45.405 146.455 ;
        RECT 45.665 146.495 45.835 147.255 ;
        RECT 46.050 146.665 46.380 147.425 ;
        RECT 45.665 146.325 46.380 146.495 ;
        RECT 46.550 146.350 46.805 147.255 ;
        RECT 44.275 145.785 44.525 146.285 ;
        RECT 43.765 145.445 44.450 145.615 ;
        RECT 44.705 145.535 45.065 146.115 ;
        RECT 43.740 144.875 44.075 145.275 ;
        RECT 44.245 145.045 44.450 145.445 ;
        RECT 45.235 145.375 45.405 146.285 ;
        RECT 45.575 145.775 45.930 146.145 ;
        RECT 46.210 146.115 46.380 146.325 ;
        RECT 46.210 145.785 46.465 146.115 ;
        RECT 46.210 145.595 46.380 145.785 ;
        RECT 46.635 145.620 46.805 146.350 ;
        RECT 46.980 146.275 47.240 147.425 ;
        RECT 47.415 146.990 52.760 147.425 ;
        RECT 44.660 144.875 44.935 145.355 ;
        RECT 45.145 145.045 45.405 145.375 ;
        RECT 45.665 145.425 46.380 145.595 ;
        RECT 45.665 145.045 45.835 145.425 ;
        RECT 46.050 144.875 46.380 145.255 ;
        RECT 46.550 145.045 46.805 145.620 ;
        RECT 46.980 144.875 47.240 145.715 ;
        RECT 49.000 145.420 49.340 146.250 ;
        RECT 50.820 145.740 51.170 146.990 ;
        RECT 52.935 146.335 55.525 147.425 ;
        RECT 52.935 145.645 54.145 146.165 ;
        RECT 54.315 145.815 55.525 146.335 ;
        RECT 56.155 146.260 56.445 147.425 ;
        RECT 56.615 146.335 58.285 147.425 ;
        RECT 58.460 147.000 58.795 147.425 ;
        RECT 58.965 146.820 59.150 147.225 ;
        RECT 56.615 145.645 57.365 146.165 ;
        RECT 57.535 145.815 58.285 146.335 ;
        RECT 58.485 146.645 59.150 146.820 ;
        RECT 59.355 146.645 59.685 147.425 ;
        RECT 47.415 144.875 52.760 145.420 ;
        RECT 52.935 144.875 55.525 145.645 ;
        RECT 56.155 144.875 56.445 145.600 ;
        RECT 56.615 144.875 58.285 145.645 ;
        RECT 58.485 145.615 58.825 146.645 ;
        RECT 59.855 146.455 60.125 147.225 ;
        RECT 60.300 147.000 60.635 147.425 ;
        RECT 60.805 146.820 60.990 147.225 ;
        RECT 58.995 146.285 60.125 146.455 ;
        RECT 58.995 145.785 59.245 146.285 ;
        RECT 58.485 145.445 59.170 145.615 ;
        RECT 59.425 145.535 59.785 146.115 ;
        RECT 58.460 144.875 58.795 145.275 ;
        RECT 58.965 145.045 59.170 145.445 ;
        RECT 59.955 145.375 60.125 146.285 ;
        RECT 60.325 146.645 60.990 146.820 ;
        RECT 61.195 146.645 61.525 147.425 ;
        RECT 60.325 145.615 60.665 146.645 ;
        RECT 61.695 146.455 61.965 147.225 ;
        RECT 60.835 146.285 61.965 146.455 ;
        RECT 62.135 146.285 62.415 147.425 ;
        RECT 60.835 145.785 61.085 146.285 ;
        RECT 60.325 145.445 61.010 145.615 ;
        RECT 61.265 145.535 61.625 146.115 ;
        RECT 59.380 144.875 59.655 145.355 ;
        RECT 59.865 145.045 60.125 145.375 ;
        RECT 60.300 144.875 60.635 145.275 ;
        RECT 60.805 145.045 61.010 145.445 ;
        RECT 61.795 145.375 61.965 146.285 ;
        RECT 62.585 146.275 62.915 147.255 ;
        RECT 63.085 146.285 63.345 147.425 ;
        RECT 63.515 146.335 66.105 147.425 ;
        RECT 66.795 146.365 67.125 147.210 ;
        RECT 67.295 146.415 67.465 147.425 ;
        RECT 67.635 146.695 67.975 147.255 ;
        RECT 68.205 146.925 68.520 147.425 ;
        RECT 68.700 146.955 69.585 147.125 ;
        RECT 62.145 145.845 62.480 146.115 ;
        RECT 62.650 145.675 62.820 146.275 ;
        RECT 62.990 145.865 63.325 146.115 ;
        RECT 61.220 144.875 61.495 145.355 ;
        RECT 61.705 145.045 61.965 145.375 ;
        RECT 62.135 144.875 62.445 145.675 ;
        RECT 62.650 145.045 63.345 145.675 ;
        RECT 63.515 145.645 64.725 146.165 ;
        RECT 64.895 145.815 66.105 146.335 ;
        RECT 66.735 146.285 67.125 146.365 ;
        RECT 67.635 146.320 68.530 146.695 ;
        RECT 66.735 146.235 66.950 146.285 ;
        RECT 66.735 145.655 66.905 146.235 ;
        RECT 67.635 146.115 67.825 146.320 ;
        RECT 68.700 146.115 68.870 146.955 ;
        RECT 69.810 146.925 70.060 147.255 ;
        RECT 67.075 145.785 67.825 146.115 ;
        RECT 67.995 145.785 68.870 146.115 ;
        RECT 63.515 144.875 66.105 145.645 ;
        RECT 66.735 145.615 66.960 145.655 ;
        RECT 67.625 145.615 67.825 145.785 ;
        RECT 66.735 145.530 67.115 145.615 ;
        RECT 66.785 145.095 67.115 145.530 ;
        RECT 67.285 144.875 67.455 145.485 ;
        RECT 67.625 145.090 67.955 145.615 ;
        RECT 68.215 144.875 68.425 145.405 ;
        RECT 68.700 145.325 68.870 145.785 ;
        RECT 69.040 145.825 69.360 146.785 ;
        RECT 69.530 146.035 69.720 146.755 ;
        RECT 69.890 145.855 70.060 146.925 ;
        RECT 70.230 146.625 70.400 147.425 ;
        RECT 70.570 146.980 71.675 147.150 ;
        RECT 70.570 146.365 70.740 146.980 ;
        RECT 71.885 146.830 72.135 147.255 ;
        RECT 72.305 146.965 72.570 147.425 ;
        RECT 70.910 146.445 71.440 146.810 ;
        RECT 71.885 146.700 72.190 146.830 ;
        RECT 70.230 146.275 70.740 146.365 ;
        RECT 70.230 146.105 71.100 146.275 ;
        RECT 70.230 146.035 70.400 146.105 ;
        RECT 70.520 145.855 70.720 145.885 ;
        RECT 69.040 145.495 69.505 145.825 ;
        RECT 69.890 145.555 70.720 145.855 ;
        RECT 69.890 145.325 70.060 145.555 ;
        RECT 68.700 145.155 69.485 145.325 ;
        RECT 69.655 145.155 70.060 145.325 ;
        RECT 70.240 144.875 70.610 145.375 ;
        RECT 70.930 145.325 71.100 146.105 ;
        RECT 71.270 145.745 71.440 146.445 ;
        RECT 71.610 145.915 71.850 146.510 ;
        RECT 71.270 145.525 71.795 145.745 ;
        RECT 72.020 145.595 72.190 146.700 ;
        RECT 71.965 145.465 72.190 145.595 ;
        RECT 72.360 145.505 72.640 146.455 ;
        RECT 71.965 145.325 72.135 145.465 ;
        RECT 70.930 145.155 71.605 145.325 ;
        RECT 71.800 145.155 72.135 145.325 ;
        RECT 72.305 144.875 72.555 145.335 ;
        RECT 72.810 145.135 72.995 147.255 ;
        RECT 73.165 146.925 73.495 147.425 ;
        RECT 73.665 146.755 73.835 147.255 ;
        RECT 73.170 146.585 73.835 146.755 ;
        RECT 73.170 145.595 73.400 146.585 ;
        RECT 73.570 145.765 73.920 146.415 ;
        RECT 74.100 146.285 74.435 147.255 ;
        RECT 74.605 146.285 74.775 147.425 ;
        RECT 74.945 147.085 76.975 147.255 ;
        RECT 74.100 145.615 74.270 146.285 ;
        RECT 74.945 146.115 75.115 147.085 ;
        RECT 74.440 145.785 74.695 146.115 ;
        RECT 74.920 145.785 75.115 146.115 ;
        RECT 75.285 146.745 76.410 146.915 ;
        RECT 74.525 145.615 74.695 145.785 ;
        RECT 75.285 145.615 75.455 146.745 ;
        RECT 73.170 145.425 73.835 145.595 ;
        RECT 73.165 144.875 73.495 145.255 ;
        RECT 73.665 145.135 73.835 145.425 ;
        RECT 74.100 145.045 74.355 145.615 ;
        RECT 74.525 145.445 75.455 145.615 ;
        RECT 75.625 146.405 76.635 146.575 ;
        RECT 75.625 145.605 75.795 146.405 ;
        RECT 76.000 145.725 76.275 146.205 ;
        RECT 75.995 145.555 76.275 145.725 ;
        RECT 75.280 145.410 75.455 145.445 ;
        RECT 74.525 144.875 74.855 145.275 ;
        RECT 75.280 145.045 75.810 145.410 ;
        RECT 76.000 145.045 76.275 145.555 ;
        RECT 76.445 145.045 76.635 146.405 ;
        RECT 76.805 146.420 76.975 147.085 ;
        RECT 77.145 146.665 77.315 147.425 ;
        RECT 77.550 146.665 78.065 147.075 ;
        RECT 76.805 146.230 77.555 146.420 ;
        RECT 77.725 145.855 78.065 146.665 ;
        RECT 78.290 146.555 78.575 147.425 ;
        RECT 78.745 146.795 79.005 147.255 ;
        RECT 79.180 146.965 79.435 147.425 ;
        RECT 79.605 146.795 79.865 147.255 ;
        RECT 78.745 146.625 79.865 146.795 ;
        RECT 80.035 146.625 80.345 147.425 ;
        RECT 78.745 146.375 79.005 146.625 ;
        RECT 80.515 146.455 80.825 147.255 ;
        RECT 76.835 145.685 78.065 145.855 ;
        RECT 78.250 146.205 79.005 146.375 ;
        RECT 79.795 146.285 80.825 146.455 ;
        RECT 78.250 145.695 78.655 146.205 ;
        RECT 79.795 146.035 79.965 146.285 ;
        RECT 78.825 145.865 79.965 146.035 ;
        RECT 76.815 144.875 77.325 145.410 ;
        RECT 77.545 145.080 77.790 145.685 ;
        RECT 78.250 145.525 79.900 145.695 ;
        RECT 80.135 145.545 80.485 146.115 ;
        RECT 78.295 144.875 78.575 145.355 ;
        RECT 78.745 145.135 79.005 145.525 ;
        RECT 79.180 144.875 79.435 145.355 ;
        RECT 79.605 145.135 79.900 145.525 ;
        RECT 80.655 145.375 80.825 146.285 ;
        RECT 81.915 146.260 82.205 147.425 ;
        RECT 82.375 146.335 84.045 147.425 ;
        RECT 82.375 145.645 83.125 146.165 ;
        RECT 83.295 145.815 84.045 146.335 ;
        RECT 84.220 146.285 84.555 147.255 ;
        RECT 84.725 146.285 84.895 147.425 ;
        RECT 85.065 147.085 87.095 147.255 ;
        RECT 80.080 144.875 80.355 145.355 ;
        RECT 80.525 145.045 80.825 145.375 ;
        RECT 81.915 144.875 82.205 145.600 ;
        RECT 82.375 144.875 84.045 145.645 ;
        RECT 84.220 145.615 84.390 146.285 ;
        RECT 85.065 146.115 85.235 147.085 ;
        RECT 84.560 145.785 84.815 146.115 ;
        RECT 85.040 145.785 85.235 146.115 ;
        RECT 85.405 146.745 86.530 146.915 ;
        RECT 84.645 145.615 84.815 145.785 ;
        RECT 85.405 145.615 85.575 146.745 ;
        RECT 84.220 145.045 84.475 145.615 ;
        RECT 84.645 145.445 85.575 145.615 ;
        RECT 85.745 146.405 86.755 146.575 ;
        RECT 85.745 145.605 85.915 146.405 ;
        RECT 85.400 145.410 85.575 145.445 ;
        RECT 84.645 144.875 84.975 145.275 ;
        RECT 85.400 145.045 85.930 145.410 ;
        RECT 86.120 145.385 86.395 146.205 ;
        RECT 86.115 145.215 86.395 145.385 ;
        RECT 86.120 145.045 86.395 145.215 ;
        RECT 86.565 145.045 86.755 146.405 ;
        RECT 86.925 146.420 87.095 147.085 ;
        RECT 87.265 146.665 87.435 147.425 ;
        RECT 87.670 146.665 88.185 147.075 ;
        RECT 86.925 146.230 87.675 146.420 ;
        RECT 87.845 145.855 88.185 146.665 ;
        RECT 88.470 146.795 88.755 147.255 ;
        RECT 88.925 146.965 89.195 147.425 ;
        RECT 88.470 146.575 89.425 146.795 ;
        RECT 86.955 145.685 88.185 145.855 ;
        RECT 88.355 145.845 89.045 146.405 ;
        RECT 86.935 144.875 87.445 145.410 ;
        RECT 87.665 145.080 87.910 145.685 ;
        RECT 89.215 145.675 89.425 146.575 ;
        RECT 88.470 145.505 89.425 145.675 ;
        RECT 89.595 146.405 89.995 147.255 ;
        RECT 90.185 146.795 90.465 147.255 ;
        RECT 90.985 146.965 91.310 147.425 ;
        RECT 90.185 146.575 91.310 146.795 ;
        RECT 89.595 145.845 90.690 146.405 ;
        RECT 90.860 146.115 91.310 146.575 ;
        RECT 91.480 146.285 91.865 147.255 ;
        RECT 92.035 146.990 97.380 147.425 ;
        RECT 88.470 145.045 88.755 145.505 ;
        RECT 88.925 144.875 89.195 145.335 ;
        RECT 89.595 145.045 89.995 145.845 ;
        RECT 90.860 145.785 91.415 146.115 ;
        RECT 90.860 145.675 91.310 145.785 ;
        RECT 90.185 145.505 91.310 145.675 ;
        RECT 91.585 145.615 91.865 146.285 ;
        RECT 90.185 145.045 90.465 145.505 ;
        RECT 90.985 144.875 91.310 145.335 ;
        RECT 91.480 145.045 91.865 145.615 ;
        RECT 93.620 145.420 93.960 146.250 ;
        RECT 95.440 145.740 95.790 146.990 ;
        RECT 97.555 146.335 98.765 147.425 ;
        RECT 97.555 145.625 98.075 146.165 ;
        RECT 98.245 145.795 98.765 146.335 ;
        RECT 98.940 146.285 99.275 147.255 ;
        RECT 99.445 146.285 99.615 147.425 ;
        RECT 99.785 147.085 101.815 147.255 ;
        RECT 92.035 144.875 97.380 145.420 ;
        RECT 97.555 144.875 98.765 145.625 ;
        RECT 98.940 145.615 99.110 146.285 ;
        RECT 99.785 146.115 99.955 147.085 ;
        RECT 99.280 145.785 99.535 146.115 ;
        RECT 99.760 145.785 99.955 146.115 ;
        RECT 100.125 146.745 101.250 146.915 ;
        RECT 99.365 145.615 99.535 145.785 ;
        RECT 100.125 145.615 100.295 146.745 ;
        RECT 98.940 145.045 99.195 145.615 ;
        RECT 99.365 145.445 100.295 145.615 ;
        RECT 100.465 146.405 101.475 146.575 ;
        RECT 100.465 145.605 100.635 146.405 ;
        RECT 100.840 145.725 101.115 146.205 ;
        RECT 100.835 145.555 101.115 145.725 ;
        RECT 100.120 145.410 100.295 145.445 ;
        RECT 99.365 144.875 99.695 145.275 ;
        RECT 100.120 145.045 100.650 145.410 ;
        RECT 100.840 145.045 101.115 145.555 ;
        RECT 101.285 145.045 101.475 146.405 ;
        RECT 101.645 146.420 101.815 147.085 ;
        RECT 101.985 146.665 102.155 147.425 ;
        RECT 102.390 146.665 102.905 147.075 ;
        RECT 101.645 146.230 102.395 146.420 ;
        RECT 102.565 145.855 102.905 146.665 ;
        RECT 101.675 145.685 102.905 145.855 ;
        RECT 103.080 146.285 103.415 147.255 ;
        RECT 103.585 146.285 103.755 147.425 ;
        RECT 103.925 147.085 105.955 147.255 ;
        RECT 101.655 144.875 102.165 145.410 ;
        RECT 102.385 145.080 102.630 145.685 ;
        RECT 103.080 145.615 103.250 146.285 ;
        RECT 103.925 146.115 104.095 147.085 ;
        RECT 103.420 145.785 103.675 146.115 ;
        RECT 103.900 145.785 104.095 146.115 ;
        RECT 104.265 146.745 105.390 146.915 ;
        RECT 103.505 145.615 103.675 145.785 ;
        RECT 104.265 145.615 104.435 146.745 ;
        RECT 103.080 145.045 103.335 145.615 ;
        RECT 103.505 145.445 104.435 145.615 ;
        RECT 104.605 146.405 105.615 146.575 ;
        RECT 104.605 145.605 104.775 146.405 ;
        RECT 104.260 145.410 104.435 145.445 ;
        RECT 103.505 144.875 103.835 145.275 ;
        RECT 104.260 145.045 104.790 145.410 ;
        RECT 104.980 145.385 105.255 146.205 ;
        RECT 104.975 145.215 105.255 145.385 ;
        RECT 104.980 145.045 105.255 145.215 ;
        RECT 105.425 145.045 105.615 146.405 ;
        RECT 105.785 146.420 105.955 147.085 ;
        RECT 106.125 146.665 106.295 147.425 ;
        RECT 106.530 146.665 107.045 147.075 ;
        RECT 105.785 146.230 106.535 146.420 ;
        RECT 106.705 145.855 107.045 146.665 ;
        RECT 107.675 146.260 107.965 147.425 ;
        RECT 108.710 146.795 108.995 147.255 ;
        RECT 109.165 146.965 109.435 147.425 ;
        RECT 108.710 146.575 109.665 146.795 ;
        RECT 105.815 145.685 107.045 145.855 ;
        RECT 108.595 145.845 109.285 146.405 ;
        RECT 105.795 144.875 106.305 145.410 ;
        RECT 106.525 145.080 106.770 145.685 ;
        RECT 109.455 145.675 109.665 146.575 ;
        RECT 107.675 144.875 107.965 145.600 ;
        RECT 108.710 145.505 109.665 145.675 ;
        RECT 109.835 146.405 110.235 147.255 ;
        RECT 110.425 146.795 110.705 147.255 ;
        RECT 111.225 146.965 111.550 147.425 ;
        RECT 110.425 146.575 111.550 146.795 ;
        RECT 109.835 145.845 110.930 146.405 ;
        RECT 111.100 146.115 111.550 146.575 ;
        RECT 111.720 146.285 112.105 147.255 ;
        RECT 112.315 146.285 112.545 147.425 ;
        RECT 108.710 145.045 108.995 145.505 ;
        RECT 109.165 144.875 109.435 145.335 ;
        RECT 109.835 145.045 110.235 145.845 ;
        RECT 111.100 145.785 111.655 146.115 ;
        RECT 111.100 145.675 111.550 145.785 ;
        RECT 110.425 145.505 111.550 145.675 ;
        RECT 111.825 145.615 112.105 146.285 ;
        RECT 112.715 146.275 113.045 147.255 ;
        RECT 113.215 146.285 113.425 147.425 ;
        RECT 114.575 146.285 114.835 147.425 ;
        RECT 115.005 146.275 115.335 147.255 ;
        RECT 115.505 146.285 115.785 147.425 ;
        RECT 115.955 146.335 119.465 147.425 ;
        RECT 112.295 145.865 112.625 146.115 ;
        RECT 110.425 145.045 110.705 145.505 ;
        RECT 111.225 144.875 111.550 145.335 ;
        RECT 111.720 145.045 112.105 145.615 ;
        RECT 112.315 144.875 112.545 145.695 ;
        RECT 112.795 145.675 113.045 146.275 ;
        RECT 114.595 145.865 114.930 146.115 ;
        RECT 112.715 145.045 113.045 145.675 ;
        RECT 113.215 144.875 113.425 145.695 ;
        RECT 115.100 145.675 115.270 146.275 ;
        RECT 115.440 145.845 115.775 146.115 ;
        RECT 114.575 145.045 115.270 145.675 ;
        RECT 115.475 144.875 115.785 145.675 ;
        RECT 115.955 145.645 117.605 146.165 ;
        RECT 117.775 145.815 119.465 146.335 ;
        RECT 119.635 146.665 120.150 147.075 ;
        RECT 120.385 146.665 120.555 147.425 ;
        RECT 120.725 147.085 122.755 147.255 ;
        RECT 119.635 145.855 119.975 146.665 ;
        RECT 120.725 146.420 120.895 147.085 ;
        RECT 121.290 146.745 122.415 146.915 ;
        RECT 120.145 146.230 120.895 146.420 ;
        RECT 121.065 146.405 122.075 146.575 ;
        RECT 119.635 145.685 120.865 145.855 ;
        RECT 115.955 144.875 119.465 145.645 ;
        RECT 119.910 145.080 120.155 145.685 ;
        RECT 120.375 144.875 120.885 145.410 ;
        RECT 121.065 145.045 121.255 146.405 ;
        RECT 121.425 146.065 121.700 146.205 ;
        RECT 121.425 145.895 121.705 146.065 ;
        RECT 121.425 145.045 121.700 145.895 ;
        RECT 121.905 145.605 122.075 146.405 ;
        RECT 122.245 145.615 122.415 146.745 ;
        RECT 122.585 146.115 122.755 147.085 ;
        RECT 122.925 146.285 123.095 147.425 ;
        RECT 123.265 146.285 123.600 147.255 ;
        RECT 122.585 145.785 122.780 146.115 ;
        RECT 123.005 145.785 123.260 146.115 ;
        RECT 123.005 145.615 123.175 145.785 ;
        RECT 123.430 145.615 123.600 146.285 ;
        RECT 123.780 146.275 124.040 147.425 ;
        RECT 124.215 146.350 124.470 147.255 ;
        RECT 124.640 146.665 124.970 147.425 ;
        RECT 125.185 146.495 125.355 147.255 ;
        RECT 126.165 146.755 126.335 147.255 ;
        RECT 126.505 146.925 126.835 147.425 ;
        RECT 126.165 146.585 126.830 146.755 ;
        RECT 122.245 145.445 123.175 145.615 ;
        RECT 122.245 145.410 122.420 145.445 ;
        RECT 121.890 145.045 122.420 145.410 ;
        RECT 122.845 144.875 123.175 145.275 ;
        RECT 123.345 145.045 123.600 145.615 ;
        RECT 123.780 144.875 124.040 145.715 ;
        RECT 124.215 145.620 124.385 146.350 ;
        RECT 124.640 146.325 125.355 146.495 ;
        RECT 124.640 146.115 124.810 146.325 ;
        RECT 124.555 145.785 124.810 146.115 ;
        RECT 124.215 145.045 124.470 145.620 ;
        RECT 124.640 145.595 124.810 145.785 ;
        RECT 125.090 145.775 125.445 146.145 ;
        RECT 126.080 145.765 126.430 146.415 ;
        RECT 126.600 145.595 126.830 146.585 ;
        RECT 124.640 145.425 125.355 145.595 ;
        RECT 124.640 144.875 124.970 145.255 ;
        RECT 125.185 145.045 125.355 145.425 ;
        RECT 126.165 145.425 126.830 145.595 ;
        RECT 126.165 145.135 126.335 145.425 ;
        RECT 126.505 144.875 126.835 145.255 ;
        RECT 127.005 145.135 127.190 147.255 ;
        RECT 127.430 146.965 127.695 147.425 ;
        RECT 127.865 146.830 128.115 147.255 ;
        RECT 128.325 146.980 129.430 147.150 ;
        RECT 127.810 146.700 128.115 146.830 ;
        RECT 127.360 145.505 127.640 146.455 ;
        RECT 127.810 145.595 127.980 146.700 ;
        RECT 128.150 145.915 128.390 146.510 ;
        RECT 128.560 146.445 129.090 146.810 ;
        RECT 128.560 145.745 128.730 146.445 ;
        RECT 129.260 146.365 129.430 146.980 ;
        RECT 129.600 146.625 129.770 147.425 ;
        RECT 129.940 146.925 130.190 147.255 ;
        RECT 130.415 146.955 131.300 147.125 ;
        RECT 129.260 146.275 129.770 146.365 ;
        RECT 127.810 145.465 128.035 145.595 ;
        RECT 128.205 145.525 128.730 145.745 ;
        RECT 128.900 146.105 129.770 146.275 ;
        RECT 127.445 144.875 127.695 145.335 ;
        RECT 127.865 145.325 128.035 145.465 ;
        RECT 128.900 145.325 129.070 146.105 ;
        RECT 129.600 146.035 129.770 146.105 ;
        RECT 129.280 145.855 129.480 145.885 ;
        RECT 129.940 145.855 130.110 146.925 ;
        RECT 130.280 146.035 130.470 146.755 ;
        RECT 129.280 145.555 130.110 145.855 ;
        RECT 130.640 145.825 130.960 146.785 ;
        RECT 127.865 145.155 128.200 145.325 ;
        RECT 128.395 145.155 129.070 145.325 ;
        RECT 129.390 144.875 129.760 145.375 ;
        RECT 129.940 145.325 130.110 145.555 ;
        RECT 130.495 145.495 130.960 145.825 ;
        RECT 131.130 146.115 131.300 146.955 ;
        RECT 131.480 146.925 131.795 147.425 ;
        RECT 132.025 146.695 132.365 147.255 ;
        RECT 131.470 146.320 132.365 146.695 ;
        RECT 132.535 146.415 132.705 147.425 ;
        RECT 132.175 146.115 132.365 146.320 ;
        RECT 132.875 146.365 133.205 147.210 ;
        RECT 132.875 146.285 133.265 146.365 ;
        RECT 133.050 146.235 133.265 146.285 ;
        RECT 133.435 146.260 133.725 147.425 ;
        RECT 133.895 146.285 134.280 147.255 ;
        RECT 134.450 146.965 134.775 147.425 ;
        RECT 135.295 146.795 135.575 147.255 ;
        RECT 134.450 146.575 135.575 146.795 ;
        RECT 131.130 145.785 132.005 146.115 ;
        RECT 132.175 145.785 132.925 146.115 ;
        RECT 131.130 145.325 131.300 145.785 ;
        RECT 132.175 145.615 132.375 145.785 ;
        RECT 133.095 145.655 133.265 146.235 ;
        RECT 133.040 145.615 133.265 145.655 ;
        RECT 129.940 145.155 130.345 145.325 ;
        RECT 130.515 145.155 131.300 145.325 ;
        RECT 131.575 144.875 131.785 145.405 ;
        RECT 132.045 145.090 132.375 145.615 ;
        RECT 132.885 145.530 133.265 145.615 ;
        RECT 133.895 145.615 134.175 146.285 ;
        RECT 134.450 146.115 134.900 146.575 ;
        RECT 135.765 146.405 136.165 147.255 ;
        RECT 136.565 146.965 136.835 147.425 ;
        RECT 137.005 146.795 137.290 147.255 ;
        RECT 134.345 145.785 134.900 146.115 ;
        RECT 135.070 145.845 136.165 146.405 ;
        RECT 134.450 145.675 134.900 145.785 ;
        RECT 132.545 144.875 132.715 145.485 ;
        RECT 132.885 145.095 133.215 145.530 ;
        RECT 133.435 144.875 133.725 145.600 ;
        RECT 133.895 145.045 134.280 145.615 ;
        RECT 134.450 145.505 135.575 145.675 ;
        RECT 134.450 144.875 134.775 145.335 ;
        RECT 135.295 145.045 135.575 145.505 ;
        RECT 135.765 145.045 136.165 145.845 ;
        RECT 136.335 146.575 137.290 146.795 ;
        RECT 136.335 145.675 136.545 146.575 ;
        RECT 138.125 146.495 138.295 147.255 ;
        RECT 138.510 146.665 138.840 147.425 ;
        RECT 136.715 145.845 137.405 146.405 ;
        RECT 138.125 146.325 138.840 146.495 ;
        RECT 139.010 146.350 139.265 147.255 ;
        RECT 138.035 145.775 138.390 146.145 ;
        RECT 138.670 146.115 138.840 146.325 ;
        RECT 138.670 145.785 138.925 146.115 ;
        RECT 136.335 145.505 137.290 145.675 ;
        RECT 138.670 145.595 138.840 145.785 ;
        RECT 139.095 145.620 139.265 146.350 ;
        RECT 139.440 146.275 139.700 147.425 ;
        RECT 139.965 146.495 140.135 147.255 ;
        RECT 140.350 146.665 140.680 147.425 ;
        RECT 139.965 146.325 140.680 146.495 ;
        RECT 140.850 146.350 141.105 147.255 ;
        RECT 139.875 145.775 140.230 146.145 ;
        RECT 140.510 146.115 140.680 146.325 ;
        RECT 140.510 145.785 140.765 146.115 ;
        RECT 136.565 144.875 136.835 145.335 ;
        RECT 137.005 145.045 137.290 145.505 ;
        RECT 138.125 145.425 138.840 145.595 ;
        RECT 138.125 145.045 138.295 145.425 ;
        RECT 138.510 144.875 138.840 145.255 ;
        RECT 139.010 145.045 139.265 145.620 ;
        RECT 139.440 144.875 139.700 145.715 ;
        RECT 140.510 145.595 140.680 145.785 ;
        RECT 140.935 145.620 141.105 146.350 ;
        RECT 141.280 146.275 141.540 147.425 ;
        RECT 141.715 146.335 142.925 147.425 ;
        RECT 141.715 145.795 142.235 146.335 ;
        RECT 139.965 145.425 140.680 145.595 ;
        RECT 139.965 145.045 140.135 145.425 ;
        RECT 140.350 144.875 140.680 145.255 ;
        RECT 140.850 145.045 141.105 145.620 ;
        RECT 141.280 144.875 141.540 145.715 ;
        RECT 142.405 145.625 142.925 146.165 ;
        RECT 141.715 144.875 142.925 145.625 ;
        RECT 17.430 144.705 143.010 144.875 ;
        RECT 17.515 143.955 18.725 144.705 ;
        RECT 17.515 143.415 18.035 143.955 ;
        RECT 18.895 143.935 20.565 144.705 ;
        RECT 20.735 144.055 20.995 144.535 ;
        RECT 21.165 144.245 21.495 144.705 ;
        RECT 21.685 144.065 21.885 144.485 ;
        RECT 18.205 143.245 18.725 143.785 ;
        RECT 18.895 143.415 19.645 143.935 ;
        RECT 19.815 143.245 20.565 143.765 ;
        RECT 17.515 142.155 18.725 143.245 ;
        RECT 18.895 142.155 20.565 143.245 ;
        RECT 20.735 143.025 20.905 144.055 ;
        RECT 21.075 143.365 21.305 143.795 ;
        RECT 21.475 143.545 21.885 144.065 ;
        RECT 22.055 144.220 22.845 144.485 ;
        RECT 22.055 143.365 22.310 144.220 ;
        RECT 23.025 143.885 23.355 144.305 ;
        RECT 23.525 143.885 23.785 144.705 ;
        RECT 24.040 144.205 24.535 144.535 ;
        RECT 23.025 143.795 23.275 143.885 ;
        RECT 22.480 143.545 23.275 143.795 ;
        RECT 21.075 143.195 22.865 143.365 ;
        RECT 20.735 142.325 21.010 143.025 ;
        RECT 21.180 142.900 21.895 143.195 ;
        RECT 22.115 142.835 22.445 143.025 ;
        RECT 21.220 142.155 21.435 142.700 ;
        RECT 21.605 142.325 22.080 142.665 ;
        RECT 22.250 142.660 22.445 142.835 ;
        RECT 22.615 142.830 22.865 143.195 ;
        RECT 22.250 142.155 22.865 142.660 ;
        RECT 23.105 142.325 23.275 143.545 ;
        RECT 23.445 142.835 23.785 143.715 ;
        RECT 23.955 142.715 24.195 144.025 ;
        RECT 24.365 143.295 24.535 144.205 ;
        RECT 24.755 143.465 25.105 144.430 ;
        RECT 25.285 143.465 25.585 144.435 ;
        RECT 25.765 143.465 26.045 144.435 ;
        RECT 26.225 143.905 26.495 144.705 ;
        RECT 26.665 143.985 27.005 144.495 ;
        RECT 27.265 144.155 27.435 144.445 ;
        RECT 27.605 144.325 27.935 144.705 ;
        RECT 27.265 143.985 27.930 144.155 ;
        RECT 26.240 143.465 26.570 143.715 ;
        RECT 26.240 143.295 26.555 143.465 ;
        RECT 24.365 143.125 26.555 143.295 ;
        RECT 23.525 142.155 23.785 142.665 ;
        RECT 23.960 142.155 24.295 142.535 ;
        RECT 24.465 142.325 24.715 143.125 ;
        RECT 24.935 142.155 25.265 142.875 ;
        RECT 25.450 142.325 25.700 143.125 ;
        RECT 26.165 142.155 26.495 142.955 ;
        RECT 26.745 142.585 27.005 143.985 ;
        RECT 27.180 143.165 27.530 143.815 ;
        RECT 27.700 142.995 27.930 143.985 ;
        RECT 26.665 142.325 27.005 142.585 ;
        RECT 27.265 142.825 27.930 142.995 ;
        RECT 27.265 142.325 27.435 142.825 ;
        RECT 27.605 142.155 27.935 142.655 ;
        RECT 28.105 142.325 28.290 144.445 ;
        RECT 28.545 144.245 28.795 144.705 ;
        RECT 28.965 144.255 29.300 144.425 ;
        RECT 29.495 144.255 30.170 144.425 ;
        RECT 28.965 144.115 29.135 144.255 ;
        RECT 28.460 143.125 28.740 144.075 ;
        RECT 28.910 143.985 29.135 144.115 ;
        RECT 28.910 142.880 29.080 143.985 ;
        RECT 29.305 143.835 29.830 144.055 ;
        RECT 29.250 143.070 29.490 143.665 ;
        RECT 29.660 143.135 29.830 143.835 ;
        RECT 30.000 143.475 30.170 144.255 ;
        RECT 30.490 144.205 30.860 144.705 ;
        RECT 31.040 144.255 31.445 144.425 ;
        RECT 31.615 144.255 32.400 144.425 ;
        RECT 31.040 144.025 31.210 144.255 ;
        RECT 30.380 143.725 31.210 144.025 ;
        RECT 31.595 143.755 32.060 144.085 ;
        RECT 30.380 143.695 30.580 143.725 ;
        RECT 30.700 143.475 30.870 143.545 ;
        RECT 30.000 143.305 30.870 143.475 ;
        RECT 30.360 143.215 30.870 143.305 ;
        RECT 28.910 142.750 29.215 142.880 ;
        RECT 29.660 142.770 30.190 143.135 ;
        RECT 28.530 142.155 28.795 142.615 ;
        RECT 28.965 142.325 29.215 142.750 ;
        RECT 30.360 142.600 30.530 143.215 ;
        RECT 29.425 142.430 30.530 142.600 ;
        RECT 30.700 142.155 30.870 142.955 ;
        RECT 31.040 142.655 31.210 143.725 ;
        RECT 31.380 142.825 31.570 143.545 ;
        RECT 31.740 142.795 32.060 143.755 ;
        RECT 32.230 143.795 32.400 144.255 ;
        RECT 32.675 144.175 32.885 144.705 ;
        RECT 33.145 143.965 33.475 144.490 ;
        RECT 33.645 144.095 33.815 144.705 ;
        RECT 33.985 144.050 34.315 144.485 ;
        RECT 33.985 143.965 34.365 144.050 ;
        RECT 33.275 143.795 33.475 143.965 ;
        RECT 34.140 143.925 34.365 143.965 ;
        RECT 32.230 143.465 33.105 143.795 ;
        RECT 33.275 143.465 34.025 143.795 ;
        RECT 31.040 142.325 31.290 142.655 ;
        RECT 32.230 142.625 32.400 143.465 ;
        RECT 33.275 143.260 33.465 143.465 ;
        RECT 34.195 143.345 34.365 143.925 ;
        RECT 34.575 143.885 34.805 144.705 ;
        RECT 34.975 143.905 35.305 144.535 ;
        RECT 34.555 143.465 34.885 143.715 ;
        RECT 34.150 143.295 34.365 143.345 ;
        RECT 35.055 143.305 35.305 143.905 ;
        RECT 35.475 143.885 35.685 144.705 ;
        RECT 36.845 143.895 37.115 144.705 ;
        RECT 37.285 143.895 37.615 144.535 ;
        RECT 37.785 143.895 38.025 144.705 ;
        RECT 38.220 143.940 38.675 144.705 ;
        RECT 38.950 144.325 40.250 144.535 ;
        RECT 40.505 144.345 40.835 144.705 ;
        RECT 40.080 144.175 40.250 144.325 ;
        RECT 41.005 144.205 41.265 144.535 ;
        RECT 36.835 143.465 37.185 143.715 ;
        RECT 32.570 142.885 33.465 143.260 ;
        RECT 33.975 143.215 34.365 143.295 ;
        RECT 31.515 142.455 32.400 142.625 ;
        RECT 32.580 142.155 32.895 142.655 ;
        RECT 33.125 142.325 33.465 142.885 ;
        RECT 33.635 142.155 33.805 143.165 ;
        RECT 33.975 142.370 34.305 143.215 ;
        RECT 34.575 142.155 34.805 143.295 ;
        RECT 34.975 142.325 35.305 143.305 ;
        RECT 37.355 143.295 37.525 143.895 ;
        RECT 39.150 143.715 39.370 144.115 ;
        RECT 37.695 143.465 38.045 143.715 ;
        RECT 38.215 143.515 38.705 143.715 ;
        RECT 38.895 143.505 39.370 143.715 ;
        RECT 39.615 143.715 39.825 144.115 ;
        RECT 40.080 144.050 40.835 144.175 ;
        RECT 40.080 144.005 40.925 144.050 ;
        RECT 40.655 143.885 40.925 144.005 ;
        RECT 39.615 143.505 39.945 143.715 ;
        RECT 40.115 143.445 40.525 143.750 ;
        RECT 35.475 142.155 35.685 143.295 ;
        RECT 36.845 142.155 37.175 143.295 ;
        RECT 37.355 143.125 38.035 143.295 ;
        RECT 37.705 142.340 38.035 143.125 ;
        RECT 38.220 143.275 39.395 143.335 ;
        RECT 40.755 143.310 40.925 143.885 ;
        RECT 40.725 143.275 40.925 143.310 ;
        RECT 38.220 143.165 40.925 143.275 ;
        RECT 38.220 142.545 38.475 143.165 ;
        RECT 39.065 143.105 40.865 143.165 ;
        RECT 39.065 143.075 39.395 143.105 ;
        RECT 41.095 143.005 41.265 144.205 ;
        RECT 41.435 143.935 43.105 144.705 ;
        RECT 43.275 143.980 43.565 144.705 ;
        RECT 43.735 144.315 44.995 144.495 ;
        RECT 41.435 143.415 42.185 143.935 ;
        RECT 42.355 143.245 43.105 143.765 ;
        RECT 38.725 142.905 38.910 142.995 ;
        RECT 39.500 142.905 40.335 142.915 ;
        RECT 38.725 142.705 40.335 142.905 ;
        RECT 38.725 142.665 38.955 142.705 ;
        RECT 38.220 142.325 38.555 142.545 ;
        RECT 39.560 142.155 39.915 142.535 ;
        RECT 40.085 142.325 40.335 142.705 ;
        RECT 40.585 142.155 40.835 142.935 ;
        RECT 41.005 142.325 41.265 143.005 ;
        RECT 41.435 142.155 43.105 143.245 ;
        RECT 43.275 142.155 43.565 143.320 ;
        RECT 43.735 142.800 43.975 144.125 ;
        RECT 44.145 143.965 44.495 144.145 ;
        RECT 44.665 144.095 44.995 144.315 ;
        RECT 45.185 144.265 45.355 144.705 ;
        RECT 45.525 144.095 45.865 144.510 ;
        RECT 46.035 144.160 51.380 144.705 ;
        RECT 44.665 143.965 45.865 144.095 ;
        RECT 44.145 142.955 44.315 143.965 ;
        RECT 44.835 143.925 45.865 143.965 ;
        RECT 44.485 143.375 44.655 143.795 ;
        RECT 44.870 143.545 45.235 143.715 ;
        RECT 44.485 143.125 44.885 143.375 ;
        RECT 45.055 143.345 45.235 143.545 ;
        RECT 45.405 143.515 45.865 143.715 ;
        RECT 45.055 143.175 45.375 143.345 ;
        RECT 44.145 142.745 44.985 142.955 ;
        RECT 43.785 142.155 43.995 142.615 ;
        RECT 44.485 142.325 44.985 142.745 ;
        RECT 45.175 142.385 45.375 143.175 ;
        RECT 45.545 142.155 45.865 143.335 ;
        RECT 47.620 143.330 47.960 144.160 ;
        RECT 51.555 143.935 54.145 144.705 ;
        RECT 54.365 144.050 54.695 144.485 ;
        RECT 54.865 144.095 55.035 144.705 ;
        RECT 54.315 143.965 54.695 144.050 ;
        RECT 55.205 143.965 55.535 144.490 ;
        RECT 55.795 144.175 56.005 144.705 ;
        RECT 56.280 144.255 57.065 144.425 ;
        RECT 57.235 144.255 57.640 144.425 ;
        RECT 49.440 142.590 49.790 143.840 ;
        RECT 51.555 143.415 52.765 143.935 ;
        RECT 54.315 143.925 54.540 143.965 ;
        RECT 52.935 143.245 54.145 143.765 ;
        RECT 46.035 142.155 51.380 142.590 ;
        RECT 51.555 142.155 54.145 143.245 ;
        RECT 54.315 143.345 54.485 143.925 ;
        RECT 55.205 143.795 55.405 143.965 ;
        RECT 56.280 143.795 56.450 144.255 ;
        RECT 54.655 143.465 55.405 143.795 ;
        RECT 55.575 143.465 56.450 143.795 ;
        RECT 54.315 143.295 54.530 143.345 ;
        RECT 54.315 143.215 54.705 143.295 ;
        RECT 54.375 142.370 54.705 143.215 ;
        RECT 55.215 143.260 55.405 143.465 ;
        RECT 54.875 142.155 55.045 143.165 ;
        RECT 55.215 142.885 56.110 143.260 ;
        RECT 55.215 142.325 55.555 142.885 ;
        RECT 55.785 142.155 56.100 142.655 ;
        RECT 56.280 142.625 56.450 143.465 ;
        RECT 56.620 143.755 57.085 144.085 ;
        RECT 57.470 144.025 57.640 144.255 ;
        RECT 57.820 144.205 58.190 144.705 ;
        RECT 58.510 144.255 59.185 144.425 ;
        RECT 59.380 144.255 59.715 144.425 ;
        RECT 56.620 142.795 56.940 143.755 ;
        RECT 57.470 143.725 58.300 144.025 ;
        RECT 57.110 142.825 57.300 143.545 ;
        RECT 57.470 142.655 57.640 143.725 ;
        RECT 58.100 143.695 58.300 143.725 ;
        RECT 57.810 143.475 57.980 143.545 ;
        RECT 58.510 143.475 58.680 144.255 ;
        RECT 59.545 144.115 59.715 144.255 ;
        RECT 59.885 144.245 60.135 144.705 ;
        RECT 57.810 143.305 58.680 143.475 ;
        RECT 58.850 143.835 59.375 144.055 ;
        RECT 59.545 143.985 59.770 144.115 ;
        RECT 57.810 143.215 58.320 143.305 ;
        RECT 56.280 142.455 57.165 142.625 ;
        RECT 57.390 142.325 57.640 142.655 ;
        RECT 57.810 142.155 57.980 142.955 ;
        RECT 58.150 142.600 58.320 143.215 ;
        RECT 58.850 143.135 59.020 143.835 ;
        RECT 58.490 142.770 59.020 143.135 ;
        RECT 59.190 143.070 59.430 143.665 ;
        RECT 59.600 142.880 59.770 143.985 ;
        RECT 59.940 143.125 60.220 144.075 ;
        RECT 59.465 142.750 59.770 142.880 ;
        RECT 58.150 142.430 59.255 142.600 ;
        RECT 59.465 142.325 59.715 142.750 ;
        RECT 59.885 142.155 60.150 142.615 ;
        RECT 60.390 142.325 60.575 144.445 ;
        RECT 60.745 144.325 61.075 144.705 ;
        RECT 61.245 144.155 61.415 144.445 ;
        RECT 60.750 143.985 61.415 144.155 ;
        RECT 61.765 144.155 61.935 144.445 ;
        RECT 62.105 144.325 62.435 144.705 ;
        RECT 61.765 143.985 62.430 144.155 ;
        RECT 60.750 142.995 60.980 143.985 ;
        RECT 61.150 143.165 61.500 143.815 ;
        RECT 61.680 143.165 62.030 143.815 ;
        RECT 62.200 142.995 62.430 143.985 ;
        RECT 60.750 142.825 61.415 142.995 ;
        RECT 60.745 142.155 61.075 142.655 ;
        RECT 61.245 142.325 61.415 142.825 ;
        RECT 61.765 142.825 62.430 142.995 ;
        RECT 61.765 142.325 61.935 142.825 ;
        RECT 62.105 142.155 62.435 142.655 ;
        RECT 62.605 142.325 62.790 144.445 ;
        RECT 63.045 144.245 63.295 144.705 ;
        RECT 63.465 144.255 63.800 144.425 ;
        RECT 63.995 144.255 64.670 144.425 ;
        RECT 63.465 144.115 63.635 144.255 ;
        RECT 62.960 143.125 63.240 144.075 ;
        RECT 63.410 143.985 63.635 144.115 ;
        RECT 63.410 142.880 63.580 143.985 ;
        RECT 63.805 143.835 64.330 144.055 ;
        RECT 63.750 143.070 63.990 143.665 ;
        RECT 64.160 143.135 64.330 143.835 ;
        RECT 64.500 143.475 64.670 144.255 ;
        RECT 64.990 144.205 65.360 144.705 ;
        RECT 65.540 144.255 65.945 144.425 ;
        RECT 66.115 144.255 66.900 144.425 ;
        RECT 65.540 144.025 65.710 144.255 ;
        RECT 64.880 143.725 65.710 144.025 ;
        RECT 66.095 143.755 66.560 144.085 ;
        RECT 64.880 143.695 65.080 143.725 ;
        RECT 65.200 143.475 65.370 143.545 ;
        RECT 64.500 143.305 65.370 143.475 ;
        RECT 64.860 143.215 65.370 143.305 ;
        RECT 63.410 142.750 63.715 142.880 ;
        RECT 64.160 142.770 64.690 143.135 ;
        RECT 63.030 142.155 63.295 142.615 ;
        RECT 63.465 142.325 63.715 142.750 ;
        RECT 64.860 142.600 65.030 143.215 ;
        RECT 63.925 142.430 65.030 142.600 ;
        RECT 65.200 142.155 65.370 142.955 ;
        RECT 65.540 142.655 65.710 143.725 ;
        RECT 65.880 142.825 66.070 143.545 ;
        RECT 66.240 142.795 66.560 143.755 ;
        RECT 66.730 143.795 66.900 144.255 ;
        RECT 67.175 144.175 67.385 144.705 ;
        RECT 67.645 143.965 67.975 144.490 ;
        RECT 68.145 144.095 68.315 144.705 ;
        RECT 68.485 144.050 68.815 144.485 ;
        RECT 68.485 143.965 68.865 144.050 ;
        RECT 69.035 143.980 69.325 144.705 ;
        RECT 69.975 144.195 70.215 144.705 ;
        RECT 67.775 143.795 67.975 143.965 ;
        RECT 68.640 143.925 68.865 143.965 ;
        RECT 66.730 143.465 67.605 143.795 ;
        RECT 67.775 143.465 68.525 143.795 ;
        RECT 65.540 142.325 65.790 142.655 ;
        RECT 66.730 142.625 66.900 143.465 ;
        RECT 67.775 143.260 67.965 143.465 ;
        RECT 68.695 143.345 68.865 143.925 ;
        RECT 69.960 143.465 70.215 144.025 ;
        RECT 70.385 143.965 70.715 144.500 ;
        RECT 70.930 143.965 71.100 144.705 ;
        RECT 71.310 144.055 71.640 144.525 ;
        RECT 71.810 144.225 71.980 144.705 ;
        RECT 72.150 144.055 72.480 144.525 ;
        RECT 72.650 144.225 72.820 144.705 ;
        RECT 68.650 143.295 68.865 143.345 ;
        RECT 67.070 142.885 67.965 143.260 ;
        RECT 68.475 143.215 68.865 143.295 ;
        RECT 66.015 142.455 66.900 142.625 ;
        RECT 67.080 142.155 67.395 142.655 ;
        RECT 67.625 142.325 67.965 142.885 ;
        RECT 68.135 142.155 68.305 143.165 ;
        RECT 68.475 142.370 68.805 143.215 ;
        RECT 69.035 142.155 69.325 143.320 ;
        RECT 70.385 143.295 70.565 143.965 ;
        RECT 71.310 143.885 73.005 144.055 ;
        RECT 73.225 144.050 73.555 144.485 ;
        RECT 73.725 144.095 73.895 144.705 ;
        RECT 70.735 143.465 71.110 143.795 ;
        RECT 71.280 143.545 72.490 143.715 ;
        RECT 71.280 143.295 71.485 143.545 ;
        RECT 72.660 143.295 73.005 143.885 ;
        RECT 70.025 143.125 71.485 143.295 ;
        RECT 72.150 143.125 73.005 143.295 ;
        RECT 73.175 143.965 73.555 144.050 ;
        RECT 74.065 143.965 74.395 144.490 ;
        RECT 74.655 144.175 74.865 144.705 ;
        RECT 75.140 144.255 75.925 144.425 ;
        RECT 76.095 144.255 76.500 144.425 ;
        RECT 73.175 143.925 73.400 143.965 ;
        RECT 73.175 143.345 73.345 143.925 ;
        RECT 74.065 143.795 74.265 143.965 ;
        RECT 75.140 143.795 75.310 144.255 ;
        RECT 73.515 143.465 74.265 143.795 ;
        RECT 74.435 143.465 75.310 143.795 ;
        RECT 73.175 143.295 73.390 143.345 ;
        RECT 73.175 143.215 73.565 143.295 ;
        RECT 70.025 142.325 70.385 143.125 ;
        RECT 72.150 142.955 72.480 143.125 ;
        RECT 70.930 142.155 71.100 142.955 ;
        RECT 71.310 142.785 72.480 142.955 ;
        RECT 71.310 142.325 71.640 142.785 ;
        RECT 71.810 142.155 71.980 142.615 ;
        RECT 72.150 142.325 72.480 142.785 ;
        RECT 72.650 142.155 72.820 142.955 ;
        RECT 73.235 142.370 73.565 143.215 ;
        RECT 74.075 143.260 74.265 143.465 ;
        RECT 73.735 142.155 73.905 143.165 ;
        RECT 74.075 142.885 74.970 143.260 ;
        RECT 74.075 142.325 74.415 142.885 ;
        RECT 74.645 142.155 74.960 142.655 ;
        RECT 75.140 142.625 75.310 143.465 ;
        RECT 75.480 143.755 75.945 144.085 ;
        RECT 76.330 144.025 76.500 144.255 ;
        RECT 76.680 144.205 77.050 144.705 ;
        RECT 77.370 144.255 78.045 144.425 ;
        RECT 78.240 144.255 78.575 144.425 ;
        RECT 75.480 142.795 75.800 143.755 ;
        RECT 76.330 143.725 77.160 144.025 ;
        RECT 75.970 142.825 76.160 143.545 ;
        RECT 76.330 142.655 76.500 143.725 ;
        RECT 76.960 143.695 77.160 143.725 ;
        RECT 76.670 143.475 76.840 143.545 ;
        RECT 77.370 143.475 77.540 144.255 ;
        RECT 78.405 144.115 78.575 144.255 ;
        RECT 78.745 144.245 78.995 144.705 ;
        RECT 76.670 143.305 77.540 143.475 ;
        RECT 77.710 143.835 78.235 144.055 ;
        RECT 78.405 143.985 78.630 144.115 ;
        RECT 76.670 143.215 77.180 143.305 ;
        RECT 75.140 142.455 76.025 142.625 ;
        RECT 76.250 142.325 76.500 142.655 ;
        RECT 76.670 142.155 76.840 142.955 ;
        RECT 77.010 142.600 77.180 143.215 ;
        RECT 77.710 143.135 77.880 143.835 ;
        RECT 77.350 142.770 77.880 143.135 ;
        RECT 78.050 143.070 78.290 143.665 ;
        RECT 78.460 142.880 78.630 143.985 ;
        RECT 78.800 143.125 79.080 144.075 ;
        RECT 78.325 142.750 78.630 142.880 ;
        RECT 77.010 142.430 78.115 142.600 ;
        RECT 78.325 142.325 78.575 142.750 ;
        RECT 78.745 142.155 79.010 142.615 ;
        RECT 79.250 142.325 79.435 144.445 ;
        RECT 79.605 144.325 79.935 144.705 ;
        RECT 80.105 144.155 80.275 144.445 ;
        RECT 79.610 143.985 80.275 144.155 ;
        RECT 80.625 144.155 80.795 144.445 ;
        RECT 80.965 144.325 81.295 144.705 ;
        RECT 80.625 143.985 81.290 144.155 ;
        RECT 79.610 142.995 79.840 143.985 ;
        RECT 80.010 143.165 80.360 143.815 ;
        RECT 80.540 143.165 80.890 143.815 ;
        RECT 81.060 142.995 81.290 143.985 ;
        RECT 79.610 142.825 80.275 142.995 ;
        RECT 79.605 142.155 79.935 142.655 ;
        RECT 80.105 142.325 80.275 142.825 ;
        RECT 80.625 142.825 81.290 142.995 ;
        RECT 80.625 142.325 80.795 142.825 ;
        RECT 80.965 142.155 81.295 142.655 ;
        RECT 81.465 142.325 81.650 144.445 ;
        RECT 81.905 144.245 82.155 144.705 ;
        RECT 82.325 144.255 82.660 144.425 ;
        RECT 82.855 144.255 83.530 144.425 ;
        RECT 82.325 144.115 82.495 144.255 ;
        RECT 81.820 143.125 82.100 144.075 ;
        RECT 82.270 143.985 82.495 144.115 ;
        RECT 82.270 142.880 82.440 143.985 ;
        RECT 82.665 143.835 83.190 144.055 ;
        RECT 82.610 143.070 82.850 143.665 ;
        RECT 83.020 143.135 83.190 143.835 ;
        RECT 83.360 143.475 83.530 144.255 ;
        RECT 83.850 144.205 84.220 144.705 ;
        RECT 84.400 144.255 84.805 144.425 ;
        RECT 84.975 144.255 85.760 144.425 ;
        RECT 84.400 144.025 84.570 144.255 ;
        RECT 83.740 143.725 84.570 144.025 ;
        RECT 84.955 143.755 85.420 144.085 ;
        RECT 83.740 143.695 83.940 143.725 ;
        RECT 84.060 143.475 84.230 143.545 ;
        RECT 83.360 143.305 84.230 143.475 ;
        RECT 83.720 143.215 84.230 143.305 ;
        RECT 82.270 142.750 82.575 142.880 ;
        RECT 83.020 142.770 83.550 143.135 ;
        RECT 81.890 142.155 82.155 142.615 ;
        RECT 82.325 142.325 82.575 142.750 ;
        RECT 83.720 142.600 83.890 143.215 ;
        RECT 82.785 142.430 83.890 142.600 ;
        RECT 84.060 142.155 84.230 142.955 ;
        RECT 84.400 142.655 84.570 143.725 ;
        RECT 84.740 142.825 84.930 143.545 ;
        RECT 85.100 142.795 85.420 143.755 ;
        RECT 85.590 143.795 85.760 144.255 ;
        RECT 86.035 144.175 86.245 144.705 ;
        RECT 86.505 143.965 86.835 144.490 ;
        RECT 87.005 144.095 87.175 144.705 ;
        RECT 87.345 144.050 87.675 144.485 ;
        RECT 87.345 143.965 87.725 144.050 ;
        RECT 86.635 143.795 86.835 143.965 ;
        RECT 87.500 143.925 87.725 143.965 ;
        RECT 85.590 143.465 86.465 143.795 ;
        RECT 86.635 143.465 87.385 143.795 ;
        RECT 84.400 142.325 84.650 142.655 ;
        RECT 85.590 142.625 85.760 143.465 ;
        RECT 86.635 143.260 86.825 143.465 ;
        RECT 87.555 143.345 87.725 143.925 ;
        RECT 87.510 143.295 87.725 143.345 ;
        RECT 85.930 142.885 86.825 143.260 ;
        RECT 87.335 143.215 87.725 143.295 ;
        RECT 87.900 143.965 88.155 144.535 ;
        RECT 88.325 144.305 88.655 144.705 ;
        RECT 89.080 144.170 89.610 144.535 ;
        RECT 89.800 144.365 90.075 144.535 ;
        RECT 89.795 144.195 90.075 144.365 ;
        RECT 89.080 144.135 89.255 144.170 ;
        RECT 88.325 143.965 89.255 144.135 ;
        RECT 87.900 143.295 88.070 143.965 ;
        RECT 88.325 143.795 88.495 143.965 ;
        RECT 88.240 143.465 88.495 143.795 ;
        RECT 88.720 143.465 88.915 143.795 ;
        RECT 84.875 142.455 85.760 142.625 ;
        RECT 85.940 142.155 86.255 142.655 ;
        RECT 86.485 142.325 86.825 142.885 ;
        RECT 86.995 142.155 87.165 143.165 ;
        RECT 87.335 142.370 87.665 143.215 ;
        RECT 87.900 142.325 88.235 143.295 ;
        RECT 88.405 142.155 88.575 143.295 ;
        RECT 88.745 142.495 88.915 143.465 ;
        RECT 89.085 142.835 89.255 143.965 ;
        RECT 89.425 143.175 89.595 143.975 ;
        RECT 89.800 143.375 90.075 144.195 ;
        RECT 90.245 143.175 90.435 144.535 ;
        RECT 90.615 144.170 91.125 144.705 ;
        RECT 91.345 143.895 91.590 144.500 ;
        RECT 92.035 143.935 94.625 144.705 ;
        RECT 94.795 143.980 95.085 144.705 ;
        RECT 95.260 143.965 95.515 144.535 ;
        RECT 95.685 144.305 96.015 144.705 ;
        RECT 96.440 144.170 96.970 144.535 ;
        RECT 96.440 144.135 96.615 144.170 ;
        RECT 95.685 143.965 96.615 144.135 ;
        RECT 90.635 143.725 91.865 143.895 ;
        RECT 89.425 143.005 90.435 143.175 ;
        RECT 90.605 143.160 91.355 143.350 ;
        RECT 89.085 142.665 90.210 142.835 ;
        RECT 90.605 142.495 90.775 143.160 ;
        RECT 91.525 142.915 91.865 143.725 ;
        RECT 92.035 143.415 93.245 143.935 ;
        RECT 93.415 143.245 94.625 143.765 ;
        RECT 88.745 142.325 90.775 142.495 ;
        RECT 90.945 142.155 91.115 142.915 ;
        RECT 91.350 142.505 91.865 142.915 ;
        RECT 92.035 142.155 94.625 143.245 ;
        RECT 94.795 142.155 95.085 143.320 ;
        RECT 95.260 143.295 95.430 143.965 ;
        RECT 95.685 143.795 95.855 143.965 ;
        RECT 95.600 143.465 95.855 143.795 ;
        RECT 96.080 143.465 96.275 143.795 ;
        RECT 95.260 142.325 95.595 143.295 ;
        RECT 95.765 142.155 95.935 143.295 ;
        RECT 96.105 142.495 96.275 143.465 ;
        RECT 96.445 142.835 96.615 143.965 ;
        RECT 96.785 143.175 96.955 143.975 ;
        RECT 97.160 143.685 97.435 144.535 ;
        RECT 97.155 143.515 97.435 143.685 ;
        RECT 97.160 143.375 97.435 143.515 ;
        RECT 97.605 143.175 97.795 144.535 ;
        RECT 97.975 144.170 98.485 144.705 ;
        RECT 98.705 143.895 98.950 144.500 ;
        RECT 99.395 143.965 99.780 144.535 ;
        RECT 99.950 144.245 100.275 144.705 ;
        RECT 100.795 144.075 101.075 144.535 ;
        RECT 97.995 143.725 99.225 143.895 ;
        RECT 96.785 143.005 97.795 143.175 ;
        RECT 97.965 143.160 98.715 143.350 ;
        RECT 96.445 142.665 97.570 142.835 ;
        RECT 97.965 142.495 98.135 143.160 ;
        RECT 98.885 142.915 99.225 143.725 ;
        RECT 96.105 142.325 98.135 142.495 ;
        RECT 98.305 142.155 98.475 142.915 ;
        RECT 98.710 142.505 99.225 142.915 ;
        RECT 99.395 143.295 99.675 143.965 ;
        RECT 99.950 143.905 101.075 144.075 ;
        RECT 99.950 143.795 100.400 143.905 ;
        RECT 99.845 143.465 100.400 143.795 ;
        RECT 101.265 143.735 101.665 144.535 ;
        RECT 102.065 144.245 102.335 144.705 ;
        RECT 102.505 144.075 102.790 144.535 ;
        RECT 103.075 144.160 108.420 144.705 ;
        RECT 108.595 144.160 113.940 144.705 ;
        RECT 114.115 144.160 119.460 144.705 ;
        RECT 99.395 142.325 99.780 143.295 ;
        RECT 99.950 143.005 100.400 143.465 ;
        RECT 100.570 143.175 101.665 143.735 ;
        RECT 99.950 142.785 101.075 143.005 ;
        RECT 99.950 142.155 100.275 142.615 ;
        RECT 100.795 142.325 101.075 142.785 ;
        RECT 101.265 142.325 101.665 143.175 ;
        RECT 101.835 143.905 102.790 144.075 ;
        RECT 101.835 143.005 102.045 143.905 ;
        RECT 102.215 143.175 102.905 143.735 ;
        RECT 104.660 143.330 105.000 144.160 ;
        RECT 101.835 142.785 102.790 143.005 ;
        RECT 102.065 142.155 102.335 142.615 ;
        RECT 102.505 142.325 102.790 142.785 ;
        RECT 106.480 142.590 106.830 143.840 ;
        RECT 110.180 143.330 110.520 144.160 ;
        RECT 112.000 142.590 112.350 143.840 ;
        RECT 115.700 143.330 116.040 144.160 ;
        RECT 120.555 143.980 120.845 144.705 ;
        RECT 121.935 143.905 122.245 144.705 ;
        RECT 122.450 143.905 123.145 144.535 ;
        RECT 123.315 143.935 126.825 144.705 ;
        RECT 126.995 143.955 128.205 144.705 ;
        RECT 128.380 143.965 128.635 144.535 ;
        RECT 128.805 144.305 129.135 144.705 ;
        RECT 129.560 144.170 130.090 144.535 ;
        RECT 130.280 144.365 130.555 144.535 ;
        RECT 130.275 144.195 130.555 144.365 ;
        RECT 129.560 144.135 129.735 144.170 ;
        RECT 128.805 143.965 129.735 144.135 ;
        RECT 122.450 143.855 122.625 143.905 ;
        RECT 117.520 142.590 117.870 143.840 ;
        RECT 121.945 143.465 122.280 143.735 ;
        RECT 103.075 142.155 108.420 142.590 ;
        RECT 108.595 142.155 113.940 142.590 ;
        RECT 114.115 142.155 119.460 142.590 ;
        RECT 120.555 142.155 120.845 143.320 ;
        RECT 122.450 143.305 122.620 143.855 ;
        RECT 122.790 143.465 123.125 143.715 ;
        RECT 123.315 143.415 124.965 143.935 ;
        RECT 121.935 142.155 122.215 143.295 ;
        RECT 122.385 142.325 122.715 143.305 ;
        RECT 122.885 142.155 123.145 143.295 ;
        RECT 125.135 143.245 126.825 143.765 ;
        RECT 126.995 143.415 127.515 143.955 ;
        RECT 127.685 143.245 128.205 143.785 ;
        RECT 123.315 142.155 126.825 143.245 ;
        RECT 126.995 142.155 128.205 143.245 ;
        RECT 128.380 143.295 128.550 143.965 ;
        RECT 128.805 143.795 128.975 143.965 ;
        RECT 128.720 143.465 128.975 143.795 ;
        RECT 129.200 143.465 129.395 143.795 ;
        RECT 128.380 142.325 128.715 143.295 ;
        RECT 128.885 142.155 129.055 143.295 ;
        RECT 129.225 142.495 129.395 143.465 ;
        RECT 129.565 142.835 129.735 143.965 ;
        RECT 129.905 143.175 130.075 143.975 ;
        RECT 130.280 143.375 130.555 144.195 ;
        RECT 130.725 143.175 130.915 144.535 ;
        RECT 131.095 144.170 131.605 144.705 ;
        RECT 131.825 143.895 132.070 144.500 ;
        RECT 132.515 143.935 136.025 144.705 ;
        RECT 136.745 144.155 136.915 144.535 ;
        RECT 137.095 144.325 137.425 144.705 ;
        RECT 136.745 143.985 137.410 144.155 ;
        RECT 137.605 144.030 137.865 144.535 ;
        RECT 131.115 143.725 132.345 143.895 ;
        RECT 129.905 143.005 130.915 143.175 ;
        RECT 131.085 143.160 131.835 143.350 ;
        RECT 129.565 142.665 130.690 142.835 ;
        RECT 131.085 142.495 131.255 143.160 ;
        RECT 132.005 142.915 132.345 143.725 ;
        RECT 132.515 143.415 134.165 143.935 ;
        RECT 134.335 143.245 136.025 143.765 ;
        RECT 136.675 143.435 137.005 143.805 ;
        RECT 137.240 143.730 137.410 143.985 ;
        RECT 137.240 143.400 137.525 143.730 ;
        RECT 137.240 143.255 137.410 143.400 ;
        RECT 129.225 142.325 131.255 142.495 ;
        RECT 131.425 142.155 131.595 142.915 ;
        RECT 131.830 142.505 132.345 142.915 ;
        RECT 132.515 142.155 136.025 143.245 ;
        RECT 136.745 143.085 137.410 143.255 ;
        RECT 137.695 143.230 137.865 144.030 ;
        RECT 138.035 143.935 141.545 144.705 ;
        RECT 141.715 143.955 142.925 144.705 ;
        RECT 138.035 143.415 139.685 143.935 ;
        RECT 139.855 143.245 141.545 143.765 ;
        RECT 136.745 142.325 136.915 143.085 ;
        RECT 137.095 142.155 137.425 142.915 ;
        RECT 137.595 142.325 137.865 143.230 ;
        RECT 138.035 142.155 141.545 143.245 ;
        RECT 141.715 143.245 142.235 143.785 ;
        RECT 142.405 143.415 142.925 143.955 ;
        RECT 141.715 142.155 142.925 143.245 ;
        RECT 17.430 141.985 143.010 142.155 ;
        RECT 17.515 140.895 18.725 141.985 ;
        RECT 18.895 140.895 20.565 141.985 ;
        RECT 20.825 141.315 20.995 141.815 ;
        RECT 21.165 141.485 21.495 141.985 ;
        RECT 20.825 141.145 21.490 141.315 ;
        RECT 17.515 140.185 18.035 140.725 ;
        RECT 18.205 140.355 18.725 140.895 ;
        RECT 18.895 140.205 19.645 140.725 ;
        RECT 19.815 140.375 20.565 140.895 ;
        RECT 20.740 140.325 21.090 140.975 ;
        RECT 17.515 139.435 18.725 140.185 ;
        RECT 18.895 139.435 20.565 140.205 ;
        RECT 21.260 140.155 21.490 141.145 ;
        RECT 20.825 139.985 21.490 140.155 ;
        RECT 20.825 139.695 20.995 139.985 ;
        RECT 21.165 139.435 21.495 139.815 ;
        RECT 21.665 139.695 21.850 141.815 ;
        RECT 22.090 141.525 22.355 141.985 ;
        RECT 22.525 141.390 22.775 141.815 ;
        RECT 22.985 141.540 24.090 141.710 ;
        RECT 22.470 141.260 22.775 141.390 ;
        RECT 22.020 140.065 22.300 141.015 ;
        RECT 22.470 140.155 22.640 141.260 ;
        RECT 22.810 140.475 23.050 141.070 ;
        RECT 23.220 141.005 23.750 141.370 ;
        RECT 23.220 140.305 23.390 141.005 ;
        RECT 23.920 140.925 24.090 141.540 ;
        RECT 24.260 141.185 24.430 141.985 ;
        RECT 24.600 141.485 24.850 141.815 ;
        RECT 25.075 141.515 25.960 141.685 ;
        RECT 23.920 140.835 24.430 140.925 ;
        RECT 22.470 140.025 22.695 140.155 ;
        RECT 22.865 140.085 23.390 140.305 ;
        RECT 23.560 140.665 24.430 140.835 ;
        RECT 22.105 139.435 22.355 139.895 ;
        RECT 22.525 139.885 22.695 140.025 ;
        RECT 23.560 139.885 23.730 140.665 ;
        RECT 24.260 140.595 24.430 140.665 ;
        RECT 23.940 140.415 24.140 140.445 ;
        RECT 24.600 140.415 24.770 141.485 ;
        RECT 24.940 140.595 25.130 141.315 ;
        RECT 23.940 140.115 24.770 140.415 ;
        RECT 25.300 140.385 25.620 141.345 ;
        RECT 22.525 139.715 22.860 139.885 ;
        RECT 23.055 139.715 23.730 139.885 ;
        RECT 24.050 139.435 24.420 139.935 ;
        RECT 24.600 139.885 24.770 140.115 ;
        RECT 25.155 140.055 25.620 140.385 ;
        RECT 25.790 140.675 25.960 141.515 ;
        RECT 26.140 141.485 26.455 141.985 ;
        RECT 26.685 141.255 27.025 141.815 ;
        RECT 26.130 140.880 27.025 141.255 ;
        RECT 27.195 140.975 27.365 141.985 ;
        RECT 26.835 140.675 27.025 140.880 ;
        RECT 27.535 140.925 27.865 141.770 ;
        RECT 28.095 141.265 28.555 141.815 ;
        RECT 28.745 141.265 29.075 141.985 ;
        RECT 27.535 140.845 27.925 140.925 ;
        RECT 27.710 140.795 27.925 140.845 ;
        RECT 25.790 140.345 26.665 140.675 ;
        RECT 26.835 140.345 27.585 140.675 ;
        RECT 25.790 139.885 25.960 140.345 ;
        RECT 26.835 140.175 27.035 140.345 ;
        RECT 27.755 140.215 27.925 140.795 ;
        RECT 27.700 140.175 27.925 140.215 ;
        RECT 24.600 139.715 25.005 139.885 ;
        RECT 25.175 139.715 25.960 139.885 ;
        RECT 26.235 139.435 26.445 139.965 ;
        RECT 26.705 139.650 27.035 140.175 ;
        RECT 27.545 140.090 27.925 140.175 ;
        RECT 27.205 139.435 27.375 140.045 ;
        RECT 27.545 139.655 27.875 140.090 ;
        RECT 28.095 139.895 28.345 141.265 ;
        RECT 29.275 141.095 29.575 141.645 ;
        RECT 29.745 141.315 30.025 141.985 ;
        RECT 28.635 140.925 29.575 141.095 ;
        RECT 28.635 140.675 28.805 140.925 ;
        RECT 29.945 140.675 30.210 141.035 ;
        RECT 30.395 140.820 30.685 141.985 ;
        RECT 30.855 140.845 31.115 141.985 ;
        RECT 31.285 140.835 31.615 141.815 ;
        RECT 31.785 140.845 32.065 141.985 ;
        RECT 32.235 140.845 32.495 141.985 ;
        RECT 32.735 141.475 34.350 141.805 ;
        RECT 31.375 140.795 31.550 140.835 ;
        RECT 28.515 140.345 28.805 140.675 ;
        RECT 28.975 140.425 29.315 140.675 ;
        RECT 29.535 140.425 30.210 140.675 ;
        RECT 30.875 140.425 31.210 140.675 ;
        RECT 28.635 140.255 28.805 140.345 ;
        RECT 28.635 140.065 30.025 140.255 ;
        RECT 31.380 140.235 31.550 140.795 ;
        RECT 32.745 140.675 32.915 141.235 ;
        RECT 33.175 141.135 34.350 141.305 ;
        RECT 34.520 141.185 34.800 141.985 ;
        RECT 33.175 140.845 33.505 141.135 ;
        RECT 34.180 141.015 34.350 141.135 ;
        RECT 33.675 140.675 33.920 140.965 ;
        RECT 34.180 140.845 34.840 141.015 ;
        RECT 35.010 140.845 35.285 141.815 ;
        RECT 35.660 141.015 35.990 141.815 ;
        RECT 36.160 141.185 36.490 141.985 ;
        RECT 36.790 141.015 37.120 141.815 ;
        RECT 37.765 141.185 38.015 141.985 ;
        RECT 35.660 140.845 38.095 141.015 ;
        RECT 38.285 140.845 38.455 141.985 ;
        RECT 38.625 140.845 38.965 141.815 ;
        RECT 34.670 140.675 34.840 140.845 ;
        RECT 31.720 140.405 32.055 140.675 ;
        RECT 32.240 140.425 32.575 140.675 ;
        RECT 32.745 140.345 33.460 140.675 ;
        RECT 33.675 140.345 34.500 140.675 ;
        RECT 34.670 140.345 34.945 140.675 ;
        RECT 32.745 140.255 32.995 140.345 ;
        RECT 28.095 139.605 28.655 139.895 ;
        RECT 28.825 139.435 29.075 139.895 ;
        RECT 29.695 139.705 30.025 140.065 ;
        RECT 30.395 139.435 30.685 140.160 ;
        RECT 30.855 139.605 31.550 140.235 ;
        RECT 31.755 139.435 32.065 140.235 ;
        RECT 32.235 139.435 32.495 140.255 ;
        RECT 32.665 139.835 32.995 140.255 ;
        RECT 34.670 140.175 34.840 140.345 ;
        RECT 33.175 140.005 34.840 140.175 ;
        RECT 35.115 140.110 35.285 140.845 ;
        RECT 35.455 140.425 35.805 140.675 ;
        RECT 35.990 140.215 36.160 140.845 ;
        RECT 36.330 140.425 36.660 140.625 ;
        RECT 36.830 140.425 37.160 140.625 ;
        RECT 37.330 140.425 37.750 140.625 ;
        RECT 37.925 140.595 38.095 140.845 ;
        RECT 37.925 140.425 38.620 140.595 ;
        RECT 38.790 140.285 38.965 140.845 ;
        RECT 33.175 139.605 33.435 140.005 ;
        RECT 33.605 139.435 33.935 139.835 ;
        RECT 34.105 139.655 34.275 140.005 ;
        RECT 34.445 139.435 34.820 139.835 ;
        RECT 35.010 139.765 35.285 140.110 ;
        RECT 35.660 139.605 36.160 140.215 ;
        RECT 36.790 140.085 38.015 140.255 ;
        RECT 38.735 140.235 38.965 140.285 ;
        RECT 36.790 139.605 37.120 140.085 ;
        RECT 37.290 139.435 37.515 139.895 ;
        RECT 37.685 139.605 38.015 140.085 ;
        RECT 38.205 139.435 38.455 140.235 ;
        RECT 38.625 139.605 38.965 140.235 ;
        RECT 39.135 141.115 39.410 141.815 ;
        RECT 39.620 141.440 39.835 141.985 ;
        RECT 40.005 141.475 40.480 141.815 ;
        RECT 40.650 141.480 41.265 141.985 ;
        RECT 40.650 141.305 40.845 141.480 ;
        RECT 39.135 140.085 39.305 141.115 ;
        RECT 39.580 140.945 40.295 141.240 ;
        RECT 40.515 141.115 40.845 141.305 ;
        RECT 41.015 140.945 41.265 141.310 ;
        RECT 39.475 140.775 41.265 140.945 ;
        RECT 39.475 140.345 39.705 140.775 ;
        RECT 39.135 139.605 39.395 140.085 ;
        RECT 39.875 140.075 40.285 140.595 ;
        RECT 39.565 139.435 39.895 139.895 ;
        RECT 40.085 139.655 40.285 140.075 ;
        RECT 40.455 139.920 40.710 140.775 ;
        RECT 41.505 140.595 41.675 141.815 ;
        RECT 41.925 141.475 42.185 141.985 ;
        RECT 40.880 140.345 41.675 140.595 ;
        RECT 41.845 140.425 42.185 141.305 ;
        RECT 42.360 141.185 42.675 141.985 ;
        RECT 42.940 141.630 44.020 141.800 ;
        RECT 42.940 141.015 43.110 141.630 ;
        RECT 41.425 140.255 41.675 140.345 ;
        RECT 40.455 139.655 41.245 139.920 ;
        RECT 41.425 139.835 41.755 140.255 ;
        RECT 41.925 139.435 42.185 140.255 ;
        RECT 42.355 140.005 42.625 141.015 ;
        RECT 42.795 140.845 43.110 141.015 ;
        RECT 42.795 140.175 42.965 140.845 ;
        RECT 43.280 140.675 43.515 141.355 ;
        RECT 43.685 140.845 44.020 141.630 ;
        RECT 44.195 140.895 46.785 141.985 ;
        RECT 43.135 140.345 43.515 140.675 ;
        RECT 43.685 140.345 44.020 140.675 ;
        RECT 44.195 140.205 45.405 140.725 ;
        RECT 45.575 140.375 46.785 140.895 ;
        RECT 47.435 141.095 47.695 141.805 ;
        RECT 47.865 141.275 48.195 141.985 ;
        RECT 48.365 141.095 48.595 141.805 ;
        RECT 47.435 140.855 48.595 141.095 ;
        RECT 48.775 141.075 49.045 141.805 ;
        RECT 49.225 141.255 49.565 141.985 ;
        RECT 48.775 140.855 49.545 141.075 ;
        RECT 47.425 140.345 47.725 140.675 ;
        RECT 47.905 140.365 48.430 140.675 ;
        RECT 48.610 140.365 49.075 140.675 ;
        RECT 42.795 140.005 44.020 140.175 ;
        RECT 42.425 139.435 42.755 139.835 ;
        RECT 42.925 139.735 43.095 140.005 ;
        RECT 43.265 139.435 43.595 139.835 ;
        RECT 43.765 139.735 44.020 140.005 ;
        RECT 44.195 139.435 46.785 140.205 ;
        RECT 47.435 139.435 47.725 140.165 ;
        RECT 47.905 139.725 48.135 140.365 ;
        RECT 49.255 140.185 49.545 140.855 ;
        RECT 48.315 139.985 49.545 140.185 ;
        RECT 48.315 139.615 48.625 139.985 ;
        RECT 48.805 139.435 49.475 139.805 ;
        RECT 49.735 139.615 49.995 141.805 ;
        RECT 50.175 140.895 53.685 141.985 ;
        RECT 53.855 141.430 54.460 141.985 ;
        RECT 54.635 141.475 55.115 141.815 ;
        RECT 55.285 141.440 55.540 141.985 ;
        RECT 53.855 141.330 54.470 141.430 ;
        RECT 54.285 141.305 54.470 141.330 ;
        RECT 50.175 140.205 51.825 140.725 ;
        RECT 51.995 140.375 53.685 140.895 ;
        RECT 53.855 140.710 54.115 141.160 ;
        RECT 54.285 141.060 54.615 141.305 ;
        RECT 54.785 140.985 55.540 141.235 ;
        RECT 55.710 141.115 55.985 141.815 ;
        RECT 54.770 140.950 55.540 140.985 ;
        RECT 54.755 140.940 55.540 140.950 ;
        RECT 54.750 140.925 55.645 140.940 ;
        RECT 54.730 140.910 55.645 140.925 ;
        RECT 54.710 140.900 55.645 140.910 ;
        RECT 54.685 140.890 55.645 140.900 ;
        RECT 54.615 140.860 55.645 140.890 ;
        RECT 54.595 140.830 55.645 140.860 ;
        RECT 54.575 140.800 55.645 140.830 ;
        RECT 54.545 140.775 55.645 140.800 ;
        RECT 54.510 140.740 55.645 140.775 ;
        RECT 54.480 140.735 55.645 140.740 ;
        RECT 54.480 140.730 54.870 140.735 ;
        RECT 54.480 140.720 54.845 140.730 ;
        RECT 54.480 140.715 54.830 140.720 ;
        RECT 54.480 140.710 54.815 140.715 ;
        RECT 53.855 140.705 54.815 140.710 ;
        RECT 53.855 140.695 54.805 140.705 ;
        RECT 53.855 140.690 54.795 140.695 ;
        RECT 53.855 140.680 54.785 140.690 ;
        RECT 53.855 140.670 54.780 140.680 ;
        RECT 53.855 140.665 54.775 140.670 ;
        RECT 53.855 140.650 54.765 140.665 ;
        RECT 53.855 140.635 54.760 140.650 ;
        RECT 53.855 140.610 54.750 140.635 ;
        RECT 53.855 140.540 54.745 140.610 ;
        RECT 50.175 139.435 53.685 140.205 ;
        RECT 53.855 139.985 54.405 140.370 ;
        RECT 54.575 139.815 54.745 140.540 ;
        RECT 53.855 139.645 54.745 139.815 ;
        RECT 54.915 140.140 55.245 140.565 ;
        RECT 55.415 140.340 55.645 140.735 ;
        RECT 54.915 139.655 55.135 140.140 ;
        RECT 55.815 140.085 55.985 141.115 ;
        RECT 56.155 140.820 56.445 141.985 ;
        RECT 56.705 141.315 56.875 141.815 ;
        RECT 57.045 141.485 57.375 141.985 ;
        RECT 56.705 141.145 57.370 141.315 ;
        RECT 56.620 140.325 56.970 140.975 ;
        RECT 55.305 139.435 55.555 139.975 ;
        RECT 55.725 139.605 55.985 140.085 ;
        RECT 56.155 139.435 56.445 140.160 ;
        RECT 57.140 140.155 57.370 141.145 ;
        RECT 56.705 139.985 57.370 140.155 ;
        RECT 56.705 139.695 56.875 139.985 ;
        RECT 57.045 139.435 57.375 139.815 ;
        RECT 57.545 139.695 57.730 141.815 ;
        RECT 57.970 141.525 58.235 141.985 ;
        RECT 58.405 141.390 58.655 141.815 ;
        RECT 58.865 141.540 59.970 141.710 ;
        RECT 58.350 141.260 58.655 141.390 ;
        RECT 57.900 140.065 58.180 141.015 ;
        RECT 58.350 140.155 58.520 141.260 ;
        RECT 58.690 140.475 58.930 141.070 ;
        RECT 59.100 141.005 59.630 141.370 ;
        RECT 59.100 140.305 59.270 141.005 ;
        RECT 59.800 140.925 59.970 141.540 ;
        RECT 60.140 141.185 60.310 141.985 ;
        RECT 60.480 141.485 60.730 141.815 ;
        RECT 60.955 141.515 61.840 141.685 ;
        RECT 59.800 140.835 60.310 140.925 ;
        RECT 58.350 140.025 58.575 140.155 ;
        RECT 58.745 140.085 59.270 140.305 ;
        RECT 59.440 140.665 60.310 140.835 ;
        RECT 57.985 139.435 58.235 139.895 ;
        RECT 58.405 139.885 58.575 140.025 ;
        RECT 59.440 139.885 59.610 140.665 ;
        RECT 60.140 140.595 60.310 140.665 ;
        RECT 59.820 140.415 60.020 140.445 ;
        RECT 60.480 140.415 60.650 141.485 ;
        RECT 60.820 140.595 61.010 141.315 ;
        RECT 59.820 140.115 60.650 140.415 ;
        RECT 61.180 140.385 61.500 141.345 ;
        RECT 58.405 139.715 58.740 139.885 ;
        RECT 58.935 139.715 59.610 139.885 ;
        RECT 59.930 139.435 60.300 139.935 ;
        RECT 60.480 139.885 60.650 140.115 ;
        RECT 61.035 140.055 61.500 140.385 ;
        RECT 61.670 140.675 61.840 141.515 ;
        RECT 62.020 141.485 62.335 141.985 ;
        RECT 62.565 141.255 62.905 141.815 ;
        RECT 62.010 140.880 62.905 141.255 ;
        RECT 63.075 140.975 63.245 141.985 ;
        RECT 62.715 140.675 62.905 140.880 ;
        RECT 63.415 140.925 63.745 141.770 ;
        RECT 63.415 140.845 63.805 140.925 ;
        RECT 63.975 140.895 67.485 141.985 ;
        RECT 68.575 141.430 69.180 141.985 ;
        RECT 69.355 141.475 69.835 141.815 ;
        RECT 70.005 141.440 70.260 141.985 ;
        RECT 68.575 141.330 69.190 141.430 ;
        RECT 69.005 141.305 69.190 141.330 ;
        RECT 63.590 140.795 63.805 140.845 ;
        RECT 61.670 140.345 62.545 140.675 ;
        RECT 62.715 140.345 63.465 140.675 ;
        RECT 61.670 139.885 61.840 140.345 ;
        RECT 62.715 140.175 62.915 140.345 ;
        RECT 63.635 140.215 63.805 140.795 ;
        RECT 63.580 140.175 63.805 140.215 ;
        RECT 60.480 139.715 60.885 139.885 ;
        RECT 61.055 139.715 61.840 139.885 ;
        RECT 62.115 139.435 62.325 139.965 ;
        RECT 62.585 139.650 62.915 140.175 ;
        RECT 63.425 140.090 63.805 140.175 ;
        RECT 63.975 140.205 65.625 140.725 ;
        RECT 65.795 140.375 67.485 140.895 ;
        RECT 68.575 140.710 68.835 141.160 ;
        RECT 69.005 141.060 69.335 141.305 ;
        RECT 69.505 140.985 70.260 141.235 ;
        RECT 70.430 141.115 70.705 141.815 ;
        RECT 69.490 140.950 70.260 140.985 ;
        RECT 69.475 140.940 70.260 140.950 ;
        RECT 69.470 140.925 70.365 140.940 ;
        RECT 69.450 140.910 70.365 140.925 ;
        RECT 69.430 140.900 70.365 140.910 ;
        RECT 69.405 140.890 70.365 140.900 ;
        RECT 69.335 140.860 70.365 140.890 ;
        RECT 69.315 140.830 70.365 140.860 ;
        RECT 69.295 140.800 70.365 140.830 ;
        RECT 69.265 140.775 70.365 140.800 ;
        RECT 69.230 140.740 70.365 140.775 ;
        RECT 69.200 140.735 70.365 140.740 ;
        RECT 69.200 140.730 69.590 140.735 ;
        RECT 69.200 140.720 69.565 140.730 ;
        RECT 69.200 140.715 69.550 140.720 ;
        RECT 69.200 140.710 69.535 140.715 ;
        RECT 68.575 140.705 69.535 140.710 ;
        RECT 68.575 140.695 69.525 140.705 ;
        RECT 68.575 140.690 69.515 140.695 ;
        RECT 68.575 140.680 69.505 140.690 ;
        RECT 68.575 140.670 69.500 140.680 ;
        RECT 68.575 140.665 69.495 140.670 ;
        RECT 68.575 140.650 69.485 140.665 ;
        RECT 68.575 140.635 69.480 140.650 ;
        RECT 68.575 140.610 69.470 140.635 ;
        RECT 68.575 140.540 69.465 140.610 ;
        RECT 63.085 139.435 63.255 140.045 ;
        RECT 63.425 139.655 63.755 140.090 ;
        RECT 63.975 139.435 67.485 140.205 ;
        RECT 68.575 139.985 69.125 140.370 ;
        RECT 69.295 139.815 69.465 140.540 ;
        RECT 68.575 139.645 69.465 139.815 ;
        RECT 69.635 140.140 69.965 140.565 ;
        RECT 70.135 140.340 70.365 140.735 ;
        RECT 69.635 139.655 69.855 140.140 ;
        RECT 70.535 140.085 70.705 141.115 ;
        RECT 70.025 139.435 70.275 139.975 ;
        RECT 70.445 139.605 70.705 140.085 ;
        RECT 70.875 140.795 71.215 141.815 ;
        RECT 71.385 140.795 72.075 141.985 ;
        RECT 72.245 141.015 72.575 141.815 ;
        RECT 72.745 141.185 72.915 141.985 ;
        RECT 73.085 141.355 73.415 141.815 ;
        RECT 73.585 141.525 73.755 141.985 ;
        RECT 73.925 141.355 74.255 141.815 ;
        RECT 73.085 141.015 74.255 141.355 ;
        RECT 74.425 141.185 74.595 141.985 ;
        RECT 74.765 141.015 75.095 141.815 ;
        RECT 75.265 141.185 75.955 141.985 ;
        RECT 76.125 141.015 76.455 141.815 ;
        RECT 76.625 141.185 76.795 141.985 ;
        RECT 76.965 141.015 77.295 141.815 ;
        RECT 72.245 140.795 77.295 141.015 ;
        RECT 77.465 140.795 77.795 141.985 ;
        RECT 78.235 140.845 78.620 141.815 ;
        RECT 78.790 141.525 79.115 141.985 ;
        RECT 79.635 141.355 79.915 141.815 ;
        RECT 78.790 141.135 79.915 141.355 ;
        RECT 70.875 140.255 71.050 140.795 ;
        RECT 71.220 140.425 71.570 140.625 ;
        RECT 71.795 140.425 73.415 140.625 ;
        RECT 73.585 140.425 73.890 140.795 ;
        RECT 74.060 140.425 75.270 140.625 ;
        RECT 75.535 140.455 77.290 140.625 ;
        RECT 75.580 140.425 77.290 140.455 ;
        RECT 71.795 140.255 72.075 140.425 ;
        RECT 73.585 140.255 73.755 140.425 ;
        RECT 70.875 140.065 72.075 140.255 ;
        RECT 70.875 139.605 71.215 140.065 ;
        RECT 72.245 139.985 73.755 140.255 ;
        RECT 73.925 140.065 77.295 140.255 ;
        RECT 73.925 139.985 75.515 140.065 ;
        RECT 71.385 139.435 71.635 139.895 ;
        RECT 71.825 139.605 75.515 139.815 ;
        RECT 75.705 139.435 75.955 139.895 ;
        RECT 76.125 139.605 76.455 140.065 ;
        RECT 76.625 139.435 76.795 139.895 ;
        RECT 76.965 139.605 77.295 140.065 ;
        RECT 77.465 139.435 77.795 140.255 ;
        RECT 78.235 140.175 78.515 140.845 ;
        RECT 78.790 140.675 79.240 141.135 ;
        RECT 80.105 140.965 80.505 141.815 ;
        RECT 80.905 141.525 81.175 141.985 ;
        RECT 81.345 141.355 81.630 141.815 ;
        RECT 78.685 140.345 79.240 140.675 ;
        RECT 79.410 140.405 80.505 140.965 ;
        RECT 78.790 140.235 79.240 140.345 ;
        RECT 78.235 139.605 78.620 140.175 ;
        RECT 78.790 140.065 79.915 140.235 ;
        RECT 78.790 139.435 79.115 139.895 ;
        RECT 79.635 139.605 79.915 140.065 ;
        RECT 80.105 139.605 80.505 140.405 ;
        RECT 80.675 141.135 81.630 141.355 ;
        RECT 80.675 140.235 80.885 141.135 ;
        RECT 81.055 140.405 81.745 140.965 ;
        RECT 81.915 140.820 82.205 141.985 ;
        RECT 83.355 140.925 83.685 141.770 ;
        RECT 83.855 140.975 84.025 141.985 ;
        RECT 84.195 141.255 84.535 141.815 ;
        RECT 84.765 141.485 85.080 141.985 ;
        RECT 85.260 141.515 86.145 141.685 ;
        RECT 83.295 140.845 83.685 140.925 ;
        RECT 84.195 140.880 85.090 141.255 ;
        RECT 83.295 140.795 83.510 140.845 ;
        RECT 80.675 140.065 81.630 140.235 ;
        RECT 83.295 140.215 83.465 140.795 ;
        RECT 84.195 140.675 84.385 140.880 ;
        RECT 85.260 140.675 85.430 141.515 ;
        RECT 86.370 141.485 86.620 141.815 ;
        RECT 83.635 140.345 84.385 140.675 ;
        RECT 84.555 140.345 85.430 140.675 ;
        RECT 83.295 140.175 83.520 140.215 ;
        RECT 84.185 140.175 84.385 140.345 ;
        RECT 80.905 139.435 81.175 139.895 ;
        RECT 81.345 139.605 81.630 140.065 ;
        RECT 81.915 139.435 82.205 140.160 ;
        RECT 83.295 140.090 83.675 140.175 ;
        RECT 83.345 139.655 83.675 140.090 ;
        RECT 83.845 139.435 84.015 140.045 ;
        RECT 84.185 139.650 84.515 140.175 ;
        RECT 84.775 139.435 84.985 139.965 ;
        RECT 85.260 139.885 85.430 140.345 ;
        RECT 85.600 140.385 85.920 141.345 ;
        RECT 86.090 140.595 86.280 141.315 ;
        RECT 86.450 140.415 86.620 141.485 ;
        RECT 86.790 141.185 86.960 141.985 ;
        RECT 87.130 141.540 88.235 141.710 ;
        RECT 87.130 140.925 87.300 141.540 ;
        RECT 88.445 141.390 88.695 141.815 ;
        RECT 88.865 141.525 89.130 141.985 ;
        RECT 87.470 141.005 88.000 141.370 ;
        RECT 88.445 141.260 88.750 141.390 ;
        RECT 86.790 140.835 87.300 140.925 ;
        RECT 86.790 140.665 87.660 140.835 ;
        RECT 86.790 140.595 86.960 140.665 ;
        RECT 87.080 140.415 87.280 140.445 ;
        RECT 85.600 140.055 86.065 140.385 ;
        RECT 86.450 140.115 87.280 140.415 ;
        RECT 86.450 139.885 86.620 140.115 ;
        RECT 85.260 139.715 86.045 139.885 ;
        RECT 86.215 139.715 86.620 139.885 ;
        RECT 86.800 139.435 87.170 139.935 ;
        RECT 87.490 139.885 87.660 140.665 ;
        RECT 87.830 140.305 88.000 141.005 ;
        RECT 88.170 140.475 88.410 141.070 ;
        RECT 87.830 140.085 88.355 140.305 ;
        RECT 88.580 140.155 88.750 141.260 ;
        RECT 88.525 140.025 88.750 140.155 ;
        RECT 88.920 140.065 89.200 141.015 ;
        RECT 88.525 139.885 88.695 140.025 ;
        RECT 87.490 139.715 88.165 139.885 ;
        RECT 88.360 139.715 88.695 139.885 ;
        RECT 88.865 139.435 89.115 139.895 ;
        RECT 89.370 139.695 89.555 141.815 ;
        RECT 89.725 141.485 90.055 141.985 ;
        RECT 90.225 141.315 90.395 141.815 ;
        RECT 89.730 141.145 90.395 141.315 ;
        RECT 90.745 141.315 90.915 141.815 ;
        RECT 91.085 141.485 91.415 141.985 ;
        RECT 90.745 141.145 91.410 141.315 ;
        RECT 89.730 140.155 89.960 141.145 ;
        RECT 90.130 140.325 90.480 140.975 ;
        RECT 90.660 140.325 91.010 140.975 ;
        RECT 91.180 140.155 91.410 141.145 ;
        RECT 89.730 139.985 90.395 140.155 ;
        RECT 89.725 139.435 90.055 139.815 ;
        RECT 90.225 139.695 90.395 139.985 ;
        RECT 90.745 139.985 91.410 140.155 ;
        RECT 90.745 139.695 90.915 139.985 ;
        RECT 91.085 139.435 91.415 139.815 ;
        RECT 91.585 139.695 91.770 141.815 ;
        RECT 92.010 141.525 92.275 141.985 ;
        RECT 92.445 141.390 92.695 141.815 ;
        RECT 92.905 141.540 94.010 141.710 ;
        RECT 92.390 141.260 92.695 141.390 ;
        RECT 91.940 140.065 92.220 141.015 ;
        RECT 92.390 140.155 92.560 141.260 ;
        RECT 92.730 140.475 92.970 141.070 ;
        RECT 93.140 141.005 93.670 141.370 ;
        RECT 93.140 140.305 93.310 141.005 ;
        RECT 93.840 140.925 94.010 141.540 ;
        RECT 94.180 141.185 94.350 141.985 ;
        RECT 94.520 141.485 94.770 141.815 ;
        RECT 94.995 141.515 95.880 141.685 ;
        RECT 93.840 140.835 94.350 140.925 ;
        RECT 92.390 140.025 92.615 140.155 ;
        RECT 92.785 140.085 93.310 140.305 ;
        RECT 93.480 140.665 94.350 140.835 ;
        RECT 92.025 139.435 92.275 139.895 ;
        RECT 92.445 139.885 92.615 140.025 ;
        RECT 93.480 139.885 93.650 140.665 ;
        RECT 94.180 140.595 94.350 140.665 ;
        RECT 93.860 140.415 94.060 140.445 ;
        RECT 94.520 140.415 94.690 141.485 ;
        RECT 94.860 140.595 95.050 141.315 ;
        RECT 93.860 140.115 94.690 140.415 ;
        RECT 95.220 140.385 95.540 141.345 ;
        RECT 92.445 139.715 92.780 139.885 ;
        RECT 92.975 139.715 93.650 139.885 ;
        RECT 93.970 139.435 94.340 139.935 ;
        RECT 94.520 139.885 94.690 140.115 ;
        RECT 95.075 140.055 95.540 140.385 ;
        RECT 95.710 140.675 95.880 141.515 ;
        RECT 96.060 141.485 96.375 141.985 ;
        RECT 96.605 141.255 96.945 141.815 ;
        RECT 96.050 140.880 96.945 141.255 ;
        RECT 97.115 140.975 97.285 141.985 ;
        RECT 96.755 140.675 96.945 140.880 ;
        RECT 97.455 140.925 97.785 141.770 ;
        RECT 99.025 141.315 99.195 141.815 ;
        RECT 99.365 141.485 99.695 141.985 ;
        RECT 99.025 141.145 99.690 141.315 ;
        RECT 97.455 140.845 97.845 140.925 ;
        RECT 97.630 140.795 97.845 140.845 ;
        RECT 95.710 140.345 96.585 140.675 ;
        RECT 96.755 140.345 97.505 140.675 ;
        RECT 95.710 139.885 95.880 140.345 ;
        RECT 96.755 140.175 96.955 140.345 ;
        RECT 97.675 140.215 97.845 140.795 ;
        RECT 98.940 140.325 99.290 140.975 ;
        RECT 97.620 140.175 97.845 140.215 ;
        RECT 94.520 139.715 94.925 139.885 ;
        RECT 95.095 139.715 95.880 139.885 ;
        RECT 96.155 139.435 96.365 139.965 ;
        RECT 96.625 139.650 96.955 140.175 ;
        RECT 97.465 140.090 97.845 140.175 ;
        RECT 99.460 140.155 99.690 141.145 ;
        RECT 97.125 139.435 97.295 140.045 ;
        RECT 97.465 139.655 97.795 140.090 ;
        RECT 99.025 139.985 99.690 140.155 ;
        RECT 99.025 139.695 99.195 139.985 ;
        RECT 99.365 139.435 99.695 139.815 ;
        RECT 99.865 139.695 100.050 141.815 ;
        RECT 100.290 141.525 100.555 141.985 ;
        RECT 100.725 141.390 100.975 141.815 ;
        RECT 101.185 141.540 102.290 141.710 ;
        RECT 100.670 141.260 100.975 141.390 ;
        RECT 100.220 140.065 100.500 141.015 ;
        RECT 100.670 140.155 100.840 141.260 ;
        RECT 101.010 140.475 101.250 141.070 ;
        RECT 101.420 141.005 101.950 141.370 ;
        RECT 101.420 140.305 101.590 141.005 ;
        RECT 102.120 140.925 102.290 141.540 ;
        RECT 102.460 141.185 102.630 141.985 ;
        RECT 102.800 141.485 103.050 141.815 ;
        RECT 103.275 141.515 104.160 141.685 ;
        RECT 102.120 140.835 102.630 140.925 ;
        RECT 100.670 140.025 100.895 140.155 ;
        RECT 101.065 140.085 101.590 140.305 ;
        RECT 101.760 140.665 102.630 140.835 ;
        RECT 100.305 139.435 100.555 139.895 ;
        RECT 100.725 139.885 100.895 140.025 ;
        RECT 101.760 139.885 101.930 140.665 ;
        RECT 102.460 140.595 102.630 140.665 ;
        RECT 102.140 140.415 102.340 140.445 ;
        RECT 102.800 140.415 102.970 141.485 ;
        RECT 103.140 140.595 103.330 141.315 ;
        RECT 102.140 140.115 102.970 140.415 ;
        RECT 103.500 140.385 103.820 141.345 ;
        RECT 100.725 139.715 101.060 139.885 ;
        RECT 101.255 139.715 101.930 139.885 ;
        RECT 102.250 139.435 102.620 139.935 ;
        RECT 102.800 139.885 102.970 140.115 ;
        RECT 103.355 140.055 103.820 140.385 ;
        RECT 103.990 140.675 104.160 141.515 ;
        RECT 104.340 141.485 104.655 141.985 ;
        RECT 104.885 141.255 105.225 141.815 ;
        RECT 104.330 140.880 105.225 141.255 ;
        RECT 105.395 140.975 105.565 141.985 ;
        RECT 105.035 140.675 105.225 140.880 ;
        RECT 105.735 140.925 106.065 141.770 ;
        RECT 105.735 140.845 106.125 140.925 ;
        RECT 106.295 140.895 107.505 141.985 ;
        RECT 105.910 140.795 106.125 140.845 ;
        RECT 103.990 140.345 104.865 140.675 ;
        RECT 105.035 140.345 105.785 140.675 ;
        RECT 103.990 139.885 104.160 140.345 ;
        RECT 105.035 140.175 105.235 140.345 ;
        RECT 105.955 140.215 106.125 140.795 ;
        RECT 105.900 140.175 106.125 140.215 ;
        RECT 102.800 139.715 103.205 139.885 ;
        RECT 103.375 139.715 104.160 139.885 ;
        RECT 104.435 139.435 104.645 139.965 ;
        RECT 104.905 139.650 105.235 140.175 ;
        RECT 105.745 140.090 106.125 140.175 ;
        RECT 106.295 140.185 106.815 140.725 ;
        RECT 106.985 140.355 107.505 140.895 ;
        RECT 107.675 140.820 107.965 141.985 ;
        RECT 108.135 140.845 108.520 141.815 ;
        RECT 108.690 141.525 109.015 141.985 ;
        RECT 109.535 141.355 109.815 141.815 ;
        RECT 108.690 141.135 109.815 141.355 ;
        RECT 105.405 139.435 105.575 140.045 ;
        RECT 105.745 139.655 106.075 140.090 ;
        RECT 106.295 139.435 107.505 140.185 ;
        RECT 108.135 140.175 108.415 140.845 ;
        RECT 108.690 140.675 109.140 141.135 ;
        RECT 110.005 140.965 110.405 141.815 ;
        RECT 110.805 141.525 111.075 141.985 ;
        RECT 111.245 141.355 111.530 141.815 ;
        RECT 108.585 140.345 109.140 140.675 ;
        RECT 109.310 140.405 110.405 140.965 ;
        RECT 108.690 140.235 109.140 140.345 ;
        RECT 107.675 139.435 107.965 140.160 ;
        RECT 108.135 139.605 108.520 140.175 ;
        RECT 108.690 140.065 109.815 140.235 ;
        RECT 108.690 139.435 109.015 139.895 ;
        RECT 109.535 139.605 109.815 140.065 ;
        RECT 110.005 139.605 110.405 140.405 ;
        RECT 110.575 141.135 111.530 141.355 ;
        RECT 110.575 140.235 110.785 141.135 ;
        RECT 110.955 140.405 111.645 140.965 ;
        RECT 111.815 140.845 112.200 141.815 ;
        RECT 112.370 141.525 112.695 141.985 ;
        RECT 113.215 141.355 113.495 141.815 ;
        RECT 112.370 141.135 113.495 141.355 ;
        RECT 110.575 140.065 111.530 140.235 ;
        RECT 110.805 139.435 111.075 139.895 ;
        RECT 111.245 139.605 111.530 140.065 ;
        RECT 111.815 140.175 112.095 140.845 ;
        RECT 112.370 140.675 112.820 141.135 ;
        RECT 113.685 140.965 114.085 141.815 ;
        RECT 114.485 141.525 114.755 141.985 ;
        RECT 114.925 141.355 115.210 141.815 ;
        RECT 112.265 140.345 112.820 140.675 ;
        RECT 112.990 140.405 114.085 140.965 ;
        RECT 112.370 140.235 112.820 140.345 ;
        RECT 111.815 139.605 112.200 140.175 ;
        RECT 112.370 140.065 113.495 140.235 ;
        RECT 112.370 139.435 112.695 139.895 ;
        RECT 113.215 139.605 113.495 140.065 ;
        RECT 113.685 139.605 114.085 140.405 ;
        RECT 114.255 141.135 115.210 141.355 ;
        RECT 114.255 140.235 114.465 141.135 ;
        RECT 115.700 141.015 116.030 141.815 ;
        RECT 116.200 141.185 116.530 141.985 ;
        RECT 116.830 141.015 117.160 141.815 ;
        RECT 117.805 141.185 118.055 141.985 ;
        RECT 114.635 140.405 115.325 140.965 ;
        RECT 115.700 140.845 118.135 141.015 ;
        RECT 118.325 140.845 118.495 141.985 ;
        RECT 118.665 140.845 119.005 141.815 ;
        RECT 115.495 140.425 115.845 140.675 ;
        RECT 114.255 140.065 115.210 140.235 ;
        RECT 116.030 140.215 116.200 140.845 ;
        RECT 116.370 140.425 116.700 140.625 ;
        RECT 116.870 140.425 117.200 140.625 ;
        RECT 117.370 140.425 117.790 140.625 ;
        RECT 117.965 140.595 118.135 140.845 ;
        RECT 117.965 140.425 118.660 140.595 ;
        RECT 114.485 139.435 114.755 139.895 ;
        RECT 114.925 139.605 115.210 140.065 ;
        RECT 115.700 139.605 116.200 140.215 ;
        RECT 116.830 140.085 118.055 140.255 ;
        RECT 118.830 140.235 119.005 140.845 ;
        RECT 116.830 139.605 117.160 140.085 ;
        RECT 117.330 139.435 117.555 139.895 ;
        RECT 117.725 139.605 118.055 140.085 ;
        RECT 118.245 139.435 118.495 140.235 ;
        RECT 118.665 139.605 119.005 140.235 ;
        RECT 119.210 141.195 119.745 141.815 ;
        RECT 119.210 140.175 119.525 141.195 ;
        RECT 119.915 141.185 120.245 141.985 ;
        RECT 121.475 141.550 126.820 141.985 ;
        RECT 126.995 141.550 132.340 141.985 ;
        RECT 120.730 141.015 121.120 141.190 ;
        RECT 119.695 140.845 121.120 141.015 ;
        RECT 119.695 140.345 119.865 140.845 ;
        RECT 119.210 139.605 119.825 140.175 ;
        RECT 120.115 140.115 120.380 140.675 ;
        RECT 120.550 139.945 120.720 140.845 ;
        RECT 120.890 140.115 121.245 140.675 ;
        RECT 123.060 139.980 123.400 140.810 ;
        RECT 124.880 140.300 125.230 141.550 ;
        RECT 128.580 139.980 128.920 140.810 ;
        RECT 130.400 140.300 130.750 141.550 ;
        RECT 133.435 140.820 133.725 141.985 ;
        RECT 133.985 141.315 134.155 141.815 ;
        RECT 134.325 141.485 134.655 141.985 ;
        RECT 133.985 141.145 134.650 141.315 ;
        RECT 133.900 140.325 134.250 140.975 ;
        RECT 119.995 139.435 120.210 139.945 ;
        RECT 120.440 139.615 120.720 139.945 ;
        RECT 120.900 139.435 121.140 139.945 ;
        RECT 121.475 139.435 126.820 139.980 ;
        RECT 126.995 139.435 132.340 139.980 ;
        RECT 133.435 139.435 133.725 140.160 ;
        RECT 134.420 140.155 134.650 141.145 ;
        RECT 133.985 139.985 134.650 140.155 ;
        RECT 133.985 139.695 134.155 139.985 ;
        RECT 134.325 139.435 134.655 139.815 ;
        RECT 134.825 139.695 135.010 141.815 ;
        RECT 135.250 141.525 135.515 141.985 ;
        RECT 135.685 141.390 135.935 141.815 ;
        RECT 136.145 141.540 137.250 141.710 ;
        RECT 135.630 141.260 135.935 141.390 ;
        RECT 135.180 140.065 135.460 141.015 ;
        RECT 135.630 140.155 135.800 141.260 ;
        RECT 135.970 140.475 136.210 141.070 ;
        RECT 136.380 141.005 136.910 141.370 ;
        RECT 136.380 140.305 136.550 141.005 ;
        RECT 137.080 140.925 137.250 141.540 ;
        RECT 137.420 141.185 137.590 141.985 ;
        RECT 137.760 141.485 138.010 141.815 ;
        RECT 138.235 141.515 139.120 141.685 ;
        RECT 137.080 140.835 137.590 140.925 ;
        RECT 135.630 140.025 135.855 140.155 ;
        RECT 136.025 140.085 136.550 140.305 ;
        RECT 136.720 140.665 137.590 140.835 ;
        RECT 135.265 139.435 135.515 139.895 ;
        RECT 135.685 139.885 135.855 140.025 ;
        RECT 136.720 139.885 136.890 140.665 ;
        RECT 137.420 140.595 137.590 140.665 ;
        RECT 137.100 140.415 137.300 140.445 ;
        RECT 137.760 140.415 137.930 141.485 ;
        RECT 138.100 140.595 138.290 141.315 ;
        RECT 137.100 140.115 137.930 140.415 ;
        RECT 138.460 140.385 138.780 141.345 ;
        RECT 135.685 139.715 136.020 139.885 ;
        RECT 136.215 139.715 136.890 139.885 ;
        RECT 137.210 139.435 137.580 139.935 ;
        RECT 137.760 139.885 137.930 140.115 ;
        RECT 138.315 140.055 138.780 140.385 ;
        RECT 138.950 140.675 139.120 141.515 ;
        RECT 139.300 141.485 139.615 141.985 ;
        RECT 139.845 141.255 140.185 141.815 ;
        RECT 139.290 140.880 140.185 141.255 ;
        RECT 140.355 140.975 140.525 141.985 ;
        RECT 139.995 140.675 140.185 140.880 ;
        RECT 140.695 140.925 141.025 141.770 ;
        RECT 140.695 140.845 141.085 140.925 ;
        RECT 140.870 140.795 141.085 140.845 ;
        RECT 138.950 140.345 139.825 140.675 ;
        RECT 139.995 140.345 140.745 140.675 ;
        RECT 138.950 139.885 139.120 140.345 ;
        RECT 139.995 140.175 140.195 140.345 ;
        RECT 140.915 140.215 141.085 140.795 ;
        RECT 141.715 140.895 142.925 141.985 ;
        RECT 141.715 140.355 142.235 140.895 ;
        RECT 140.860 140.175 141.085 140.215 ;
        RECT 142.405 140.185 142.925 140.725 ;
        RECT 137.760 139.715 138.165 139.885 ;
        RECT 138.335 139.715 139.120 139.885 ;
        RECT 139.395 139.435 139.605 139.965 ;
        RECT 139.865 139.650 140.195 140.175 ;
        RECT 140.705 140.090 141.085 140.175 ;
        RECT 140.365 139.435 140.535 140.045 ;
        RECT 140.705 139.655 141.035 140.090 ;
        RECT 141.715 139.435 142.925 140.185 ;
        RECT 17.430 139.265 143.010 139.435 ;
        RECT 17.515 138.515 18.725 139.265 ;
        RECT 19.905 138.715 20.075 139.005 ;
        RECT 20.245 138.885 20.575 139.265 ;
        RECT 19.905 138.545 20.570 138.715 ;
        RECT 17.515 137.975 18.035 138.515 ;
        RECT 18.205 137.805 18.725 138.345 ;
        RECT 17.515 136.715 18.725 137.805 ;
        RECT 19.820 137.725 20.170 138.375 ;
        RECT 20.340 137.555 20.570 138.545 ;
        RECT 19.905 137.385 20.570 137.555 ;
        RECT 19.905 136.885 20.075 137.385 ;
        RECT 20.245 136.715 20.575 137.215 ;
        RECT 20.745 136.885 20.930 139.005 ;
        RECT 21.185 138.805 21.435 139.265 ;
        RECT 21.605 138.815 21.940 138.985 ;
        RECT 22.135 138.815 22.810 138.985 ;
        RECT 21.605 138.675 21.775 138.815 ;
        RECT 21.100 137.685 21.380 138.635 ;
        RECT 21.550 138.545 21.775 138.675 ;
        RECT 21.550 137.440 21.720 138.545 ;
        RECT 21.945 138.395 22.470 138.615 ;
        RECT 21.890 137.630 22.130 138.225 ;
        RECT 22.300 137.695 22.470 138.395 ;
        RECT 22.640 138.035 22.810 138.815 ;
        RECT 23.130 138.765 23.500 139.265 ;
        RECT 23.680 138.815 24.085 138.985 ;
        RECT 24.255 138.815 25.040 138.985 ;
        RECT 23.680 138.585 23.850 138.815 ;
        RECT 23.020 138.285 23.850 138.585 ;
        RECT 24.235 138.315 24.700 138.645 ;
        RECT 23.020 138.255 23.220 138.285 ;
        RECT 23.340 138.035 23.510 138.105 ;
        RECT 22.640 137.865 23.510 138.035 ;
        RECT 23.000 137.775 23.510 137.865 ;
        RECT 21.550 137.310 21.855 137.440 ;
        RECT 22.300 137.330 22.830 137.695 ;
        RECT 21.170 136.715 21.435 137.175 ;
        RECT 21.605 136.885 21.855 137.310 ;
        RECT 23.000 137.160 23.170 137.775 ;
        RECT 22.065 136.990 23.170 137.160 ;
        RECT 23.340 136.715 23.510 137.515 ;
        RECT 23.680 137.215 23.850 138.285 ;
        RECT 24.020 137.385 24.210 138.105 ;
        RECT 24.380 137.355 24.700 138.315 ;
        RECT 24.870 138.355 25.040 138.815 ;
        RECT 25.315 138.735 25.525 139.265 ;
        RECT 25.785 138.525 26.115 139.050 ;
        RECT 26.285 138.655 26.455 139.265 ;
        RECT 26.625 138.610 26.955 139.045 ;
        RECT 26.625 138.525 27.005 138.610 ;
        RECT 25.915 138.355 26.115 138.525 ;
        RECT 26.780 138.485 27.005 138.525 ;
        RECT 24.870 138.025 25.745 138.355 ;
        RECT 25.915 138.025 26.665 138.355 ;
        RECT 23.680 136.885 23.930 137.215 ;
        RECT 24.870 137.185 25.040 138.025 ;
        RECT 25.915 137.820 26.105 138.025 ;
        RECT 26.835 137.905 27.005 138.485 ;
        RECT 27.195 138.455 27.435 139.265 ;
        RECT 27.605 138.455 27.935 139.095 ;
        RECT 28.105 138.455 28.375 139.265 ;
        RECT 28.575 138.455 28.815 139.265 ;
        RECT 28.985 138.455 29.315 139.095 ;
        RECT 29.485 138.455 29.755 139.265 ;
        RECT 29.935 138.720 35.280 139.265 ;
        RECT 27.175 138.025 27.525 138.275 ;
        RECT 26.790 137.855 27.005 137.905 ;
        RECT 27.695 137.855 27.865 138.455 ;
        RECT 28.035 138.025 28.385 138.275 ;
        RECT 28.555 138.025 28.905 138.275 ;
        RECT 29.075 137.855 29.245 138.455 ;
        RECT 29.415 138.025 29.765 138.275 ;
        RECT 31.520 137.890 31.860 138.720 ;
        RECT 36.415 138.445 36.645 139.265 ;
        RECT 36.815 138.465 37.145 139.095 ;
        RECT 25.210 137.445 26.105 137.820 ;
        RECT 26.615 137.775 27.005 137.855 ;
        RECT 24.155 137.015 25.040 137.185 ;
        RECT 25.220 136.715 25.535 137.215 ;
        RECT 25.765 136.885 26.105 137.445 ;
        RECT 26.275 136.715 26.445 137.725 ;
        RECT 26.615 136.930 26.945 137.775 ;
        RECT 27.185 137.685 27.865 137.855 ;
        RECT 27.185 136.900 27.515 137.685 ;
        RECT 28.045 136.715 28.375 137.855 ;
        RECT 28.565 137.685 29.245 137.855 ;
        RECT 28.565 136.900 28.895 137.685 ;
        RECT 29.425 136.715 29.755 137.855 ;
        RECT 33.340 137.150 33.690 138.400 ;
        RECT 36.395 138.025 36.725 138.275 ;
        RECT 36.895 137.865 37.145 138.465 ;
        RECT 37.315 138.445 37.525 139.265 ;
        RECT 37.755 138.465 38.450 139.095 ;
        RECT 38.655 138.465 38.965 139.265 ;
        RECT 39.225 138.695 39.395 139.095 ;
        RECT 39.635 138.865 39.965 139.265 ;
        RECT 40.235 138.925 41.640 139.095 ;
        RECT 40.235 138.695 40.405 138.925 ;
        RECT 39.225 138.525 40.405 138.695 ;
        RECT 41.470 138.695 41.640 138.925 ;
        RECT 41.810 138.885 42.140 139.265 ;
        RECT 37.775 138.025 38.110 138.275 ;
        RECT 38.280 137.905 38.450 138.465 ;
        RECT 40.575 138.355 40.765 138.585 ;
        RECT 38.620 138.025 38.955 138.295 ;
        RECT 39.195 138.025 39.380 138.355 ;
        RECT 39.635 138.025 40.110 138.355 ;
        RECT 40.420 138.025 40.765 138.355 ;
        RECT 41.025 138.025 41.220 138.600 ;
        RECT 41.470 138.525 42.165 138.695 ;
        RECT 42.335 138.680 42.645 139.095 ;
        RECT 41.995 138.355 42.165 138.525 ;
        RECT 41.490 138.025 41.825 138.355 ;
        RECT 41.995 138.025 42.305 138.355 ;
        RECT 38.275 137.865 38.450 137.905 ;
        RECT 29.935 136.715 35.280 137.150 ;
        RECT 36.415 136.715 36.645 137.855 ;
        RECT 36.815 136.885 37.145 137.865 ;
        RECT 37.315 136.715 37.525 137.855 ;
        RECT 37.755 136.715 38.015 137.855 ;
        RECT 38.185 136.885 38.515 137.865 ;
        RECT 41.995 137.855 42.165 138.025 ;
        RECT 38.685 136.715 38.965 137.855 ;
        RECT 39.225 137.685 42.165 137.855 ;
        RECT 39.225 136.885 39.395 137.685 ;
        RECT 42.475 137.565 42.645 138.680 ;
        RECT 43.275 138.540 43.565 139.265 ;
        RECT 43.735 138.885 44.625 139.055 ;
        RECT 43.735 138.330 44.285 138.715 ;
        RECT 44.455 138.160 44.625 138.885 ;
        RECT 43.735 138.090 44.625 138.160 ;
        RECT 44.795 138.560 45.015 139.045 ;
        RECT 45.185 138.725 45.435 139.265 ;
        RECT 45.605 138.615 45.865 139.095 ;
        RECT 44.795 138.135 45.125 138.560 ;
        RECT 43.735 138.065 44.630 138.090 ;
        RECT 43.735 138.050 44.640 138.065 ;
        RECT 43.735 138.035 44.645 138.050 ;
        RECT 43.735 138.030 44.655 138.035 ;
        RECT 43.735 138.020 44.660 138.030 ;
        RECT 43.735 138.010 44.665 138.020 ;
        RECT 43.735 138.005 44.675 138.010 ;
        RECT 43.735 137.995 44.685 138.005 ;
        RECT 43.735 137.990 44.695 137.995 ;
        RECT 40.155 137.345 41.715 137.515 ;
        RECT 40.155 136.885 40.405 137.345 ;
        RECT 40.605 136.715 41.275 137.095 ;
        RECT 41.465 136.885 41.715 137.345 ;
        RECT 41.890 136.715 42.135 137.175 ;
        RECT 42.305 136.925 42.645 137.565 ;
        RECT 43.275 136.715 43.565 137.880 ;
        RECT 43.735 137.540 43.995 137.990 ;
        RECT 44.360 137.985 44.695 137.990 ;
        RECT 44.360 137.980 44.710 137.985 ;
        RECT 44.360 137.970 44.725 137.980 ;
        RECT 44.360 137.965 44.750 137.970 ;
        RECT 45.295 137.965 45.525 138.360 ;
        RECT 44.360 137.960 45.525 137.965 ;
        RECT 44.390 137.925 45.525 137.960 ;
        RECT 44.425 137.900 45.525 137.925 ;
        RECT 44.455 137.870 45.525 137.900 ;
        RECT 44.475 137.840 45.525 137.870 ;
        RECT 44.495 137.810 45.525 137.840 ;
        RECT 44.565 137.800 45.525 137.810 ;
        RECT 44.590 137.790 45.525 137.800 ;
        RECT 44.610 137.775 45.525 137.790 ;
        RECT 44.630 137.760 45.525 137.775 ;
        RECT 44.635 137.750 45.420 137.760 ;
        RECT 44.650 137.715 45.420 137.750 ;
        RECT 44.165 137.395 44.495 137.640 ;
        RECT 44.665 137.465 45.420 137.715 ;
        RECT 45.695 137.585 45.865 138.615 ;
        RECT 46.035 138.515 47.245 139.265 ;
        RECT 47.425 138.670 47.675 139.095 ;
        RECT 47.845 138.840 48.175 139.265 ;
        RECT 48.345 138.845 49.435 139.095 ;
        RECT 49.625 138.845 50.715 139.095 ;
        RECT 48.345 138.670 48.515 138.845 ;
        RECT 46.035 137.975 46.555 138.515 ;
        RECT 47.425 138.500 48.515 138.670 ;
        RECT 48.685 138.505 50.375 138.675 ;
        RECT 50.545 138.670 50.715 138.845 ;
        RECT 50.885 138.840 51.215 139.265 ;
        RECT 51.385 138.670 51.705 139.095 ;
        RECT 46.725 137.805 47.245 138.345 ;
        RECT 47.480 138.245 48.110 138.275 ;
        RECT 47.475 138.075 48.110 138.245 ;
        RECT 48.400 138.075 49.030 138.275 ;
        RECT 49.200 137.865 49.490 138.505 ;
        RECT 50.545 138.500 51.705 138.670 ;
        RECT 52.105 138.585 52.275 138.960 ;
        RECT 52.075 138.415 52.275 138.585 ;
        RECT 52.465 138.735 52.695 139.040 ;
        RECT 52.865 138.905 53.195 139.265 ;
        RECT 53.390 138.735 53.680 139.085 ;
        RECT 52.465 138.565 53.680 138.735 ;
        RECT 53.855 138.465 54.550 139.095 ;
        RECT 54.755 138.465 55.065 139.265 ;
        RECT 55.440 138.485 55.940 139.095 ;
        RECT 52.105 138.395 52.275 138.415 ;
        RECT 49.775 138.075 50.430 138.275 ;
        RECT 50.720 138.245 51.830 138.275 ;
        RECT 50.695 138.075 51.830 138.245 ;
        RECT 52.105 138.225 52.625 138.395 ;
        RECT 44.165 137.370 44.350 137.395 ;
        RECT 43.735 137.270 44.350 137.370 ;
        RECT 43.735 136.715 44.340 137.270 ;
        RECT 44.515 136.885 44.995 137.225 ;
        RECT 45.165 136.715 45.420 137.260 ;
        RECT 45.590 136.885 45.865 137.585 ;
        RECT 46.035 136.715 47.245 137.805 ;
        RECT 47.425 137.695 49.490 137.865 ;
        RECT 47.425 136.885 47.675 137.695 ;
        RECT 47.845 137.055 48.095 137.525 ;
        RECT 48.265 137.225 48.595 137.695 ;
        RECT 48.765 137.055 48.935 137.525 ;
        RECT 49.105 137.225 49.490 137.695 ;
        RECT 49.705 137.695 51.635 137.865 ;
        RECT 52.020 137.695 52.265 138.055 ;
        RECT 52.455 137.845 52.625 138.225 ;
        RECT 52.795 138.025 53.180 138.355 ;
        RECT 53.360 138.025 53.620 138.355 ;
        RECT 53.875 138.025 54.210 138.275 ;
        RECT 49.705 137.055 49.955 137.695 ;
        RECT 47.845 136.885 49.955 137.055 ;
        RECT 50.125 136.715 50.295 137.525 ;
        RECT 50.465 136.885 50.795 137.695 ;
        RECT 50.965 136.715 51.135 137.525 ;
        RECT 51.305 136.885 51.635 137.695 ;
        RECT 52.455 137.565 52.805 137.845 ;
        RECT 52.020 136.715 52.275 137.515 ;
        RECT 52.475 136.885 52.805 137.565 ;
        RECT 52.985 136.975 53.180 138.025 ;
        RECT 54.380 137.865 54.550 138.465 ;
        RECT 54.720 138.025 55.055 138.295 ;
        RECT 55.235 138.025 55.585 138.275 ;
        RECT 53.360 136.715 53.680 137.855 ;
        RECT 53.855 136.715 54.115 137.855 ;
        RECT 54.285 136.885 54.615 137.865 ;
        RECT 55.770 137.855 55.940 138.485 ;
        RECT 56.570 138.615 56.900 139.095 ;
        RECT 57.070 138.805 57.295 139.265 ;
        RECT 57.465 138.615 57.795 139.095 ;
        RECT 56.570 138.445 57.795 138.615 ;
        RECT 57.985 138.465 58.235 139.265 ;
        RECT 58.405 138.465 58.745 139.095 ;
        RECT 58.915 138.885 59.805 139.055 ;
        RECT 56.110 138.075 56.440 138.275 ;
        RECT 56.610 138.075 56.940 138.275 ;
        RECT 57.110 138.075 57.530 138.275 ;
        RECT 57.705 138.105 58.400 138.275 ;
        RECT 57.705 137.855 57.875 138.105 ;
        RECT 58.570 137.855 58.745 138.465 ;
        RECT 58.915 138.330 59.465 138.715 ;
        RECT 59.635 138.160 59.805 138.885 ;
        RECT 54.785 136.715 55.065 137.855 ;
        RECT 55.440 137.685 57.875 137.855 ;
        RECT 55.440 136.885 55.770 137.685 ;
        RECT 55.940 136.715 56.270 137.515 ;
        RECT 56.570 136.885 56.900 137.685 ;
        RECT 57.545 136.715 57.795 137.515 ;
        RECT 58.065 136.715 58.235 137.855 ;
        RECT 58.405 136.885 58.745 137.855 ;
        RECT 58.915 138.090 59.805 138.160 ;
        RECT 59.975 138.560 60.195 139.045 ;
        RECT 60.365 138.725 60.615 139.265 ;
        RECT 60.785 138.615 61.045 139.095 ;
        RECT 59.975 138.135 60.305 138.560 ;
        RECT 58.915 138.065 59.810 138.090 ;
        RECT 58.915 138.050 59.820 138.065 ;
        RECT 58.915 138.035 59.825 138.050 ;
        RECT 58.915 138.030 59.835 138.035 ;
        RECT 58.915 138.020 59.840 138.030 ;
        RECT 58.915 138.010 59.845 138.020 ;
        RECT 58.915 138.005 59.855 138.010 ;
        RECT 58.915 137.995 59.865 138.005 ;
        RECT 58.915 137.990 59.875 137.995 ;
        RECT 58.915 137.540 59.175 137.990 ;
        RECT 59.540 137.985 59.875 137.990 ;
        RECT 59.540 137.980 59.890 137.985 ;
        RECT 59.540 137.970 59.905 137.980 ;
        RECT 59.540 137.965 59.930 137.970 ;
        RECT 60.475 137.965 60.705 138.360 ;
        RECT 59.540 137.960 60.705 137.965 ;
        RECT 59.570 137.925 60.705 137.960 ;
        RECT 59.605 137.900 60.705 137.925 ;
        RECT 59.635 137.870 60.705 137.900 ;
        RECT 59.655 137.840 60.705 137.870 ;
        RECT 59.675 137.810 60.705 137.840 ;
        RECT 59.745 137.800 60.705 137.810 ;
        RECT 59.770 137.790 60.705 137.800 ;
        RECT 59.790 137.775 60.705 137.790 ;
        RECT 59.810 137.760 60.705 137.775 ;
        RECT 59.815 137.750 60.600 137.760 ;
        RECT 59.830 137.715 60.600 137.750 ;
        RECT 59.345 137.395 59.675 137.640 ;
        RECT 59.845 137.465 60.600 137.715 ;
        RECT 60.875 137.585 61.045 138.615 ;
        RECT 61.235 138.455 61.475 139.265 ;
        RECT 61.645 138.455 61.975 139.095 ;
        RECT 62.145 138.455 62.415 139.265 ;
        RECT 62.595 138.720 67.940 139.265 ;
        RECT 61.215 138.025 61.565 138.275 ;
        RECT 61.735 137.855 61.905 138.455 ;
        RECT 62.075 138.025 62.425 138.275 ;
        RECT 64.180 137.890 64.520 138.720 ;
        RECT 69.035 138.540 69.325 139.265 ;
        RECT 69.495 138.515 70.705 139.265 ;
        RECT 59.345 137.370 59.530 137.395 ;
        RECT 58.915 137.270 59.530 137.370 ;
        RECT 58.915 136.715 59.520 137.270 ;
        RECT 59.695 136.885 60.175 137.225 ;
        RECT 60.345 136.715 60.600 137.260 ;
        RECT 60.770 136.885 61.045 137.585 ;
        RECT 61.225 137.685 61.905 137.855 ;
        RECT 61.225 136.900 61.555 137.685 ;
        RECT 62.085 136.715 62.415 137.855 ;
        RECT 66.000 137.150 66.350 138.400 ;
        RECT 69.495 137.975 70.015 138.515 ;
        RECT 70.875 138.445 71.135 139.265 ;
        RECT 71.305 138.445 71.635 138.865 ;
        RECT 71.815 138.780 72.605 139.045 ;
        RECT 71.385 138.355 71.635 138.445 ;
        RECT 62.595 136.715 67.940 137.150 ;
        RECT 69.035 136.715 69.325 137.880 ;
        RECT 70.185 137.805 70.705 138.345 ;
        RECT 69.495 136.715 70.705 137.805 ;
        RECT 70.875 137.395 71.215 138.275 ;
        RECT 71.385 138.105 72.180 138.355 ;
        RECT 70.875 136.715 71.135 137.225 ;
        RECT 71.385 136.885 71.555 138.105 ;
        RECT 72.350 137.925 72.605 138.780 ;
        RECT 72.775 138.625 72.975 139.045 ;
        RECT 73.165 138.805 73.495 139.265 ;
        RECT 72.775 138.105 73.185 138.625 ;
        RECT 73.665 138.615 73.925 139.095 ;
        RECT 74.095 138.885 74.985 139.055 ;
        RECT 73.355 137.925 73.585 138.355 ;
        RECT 71.795 137.755 73.585 137.925 ;
        RECT 71.795 137.390 72.045 137.755 ;
        RECT 72.215 137.395 72.545 137.585 ;
        RECT 72.765 137.460 73.480 137.755 ;
        RECT 73.755 137.585 73.925 138.615 ;
        RECT 74.095 138.330 74.645 138.715 ;
        RECT 74.815 138.160 74.985 138.885 ;
        RECT 72.215 137.220 72.410 137.395 ;
        RECT 71.795 136.715 72.410 137.220 ;
        RECT 72.580 136.885 73.055 137.225 ;
        RECT 73.225 136.715 73.440 137.260 ;
        RECT 73.650 136.885 73.925 137.585 ;
        RECT 74.095 138.090 74.985 138.160 ;
        RECT 75.155 138.585 75.375 139.045 ;
        RECT 75.545 138.725 75.795 139.265 ;
        RECT 75.965 138.615 76.225 139.095 ;
        RECT 75.155 138.560 75.405 138.585 ;
        RECT 75.155 138.135 75.485 138.560 ;
        RECT 74.095 138.065 74.990 138.090 ;
        RECT 74.095 138.050 75.000 138.065 ;
        RECT 74.095 138.035 75.005 138.050 ;
        RECT 74.095 138.030 75.015 138.035 ;
        RECT 74.095 138.020 75.020 138.030 ;
        RECT 74.095 138.010 75.025 138.020 ;
        RECT 74.095 138.005 75.035 138.010 ;
        RECT 74.095 137.995 75.045 138.005 ;
        RECT 74.095 137.990 75.055 137.995 ;
        RECT 74.095 137.540 74.355 137.990 ;
        RECT 74.720 137.985 75.055 137.990 ;
        RECT 74.720 137.980 75.070 137.985 ;
        RECT 74.720 137.970 75.085 137.980 ;
        RECT 74.720 137.965 75.110 137.970 ;
        RECT 75.655 137.965 75.885 138.360 ;
        RECT 74.720 137.960 75.885 137.965 ;
        RECT 74.750 137.925 75.885 137.960 ;
        RECT 74.785 137.900 75.885 137.925 ;
        RECT 74.815 137.870 75.885 137.900 ;
        RECT 74.835 137.840 75.885 137.870 ;
        RECT 74.855 137.810 75.885 137.840 ;
        RECT 74.925 137.800 75.885 137.810 ;
        RECT 74.950 137.790 75.885 137.800 ;
        RECT 74.970 137.775 75.885 137.790 ;
        RECT 74.990 137.760 75.885 137.775 ;
        RECT 74.995 137.750 75.780 137.760 ;
        RECT 75.010 137.715 75.780 137.750 ;
        RECT 74.525 137.395 74.855 137.640 ;
        RECT 75.025 137.465 75.780 137.715 ;
        RECT 76.055 137.585 76.225 138.615 ;
        RECT 76.455 138.445 76.665 139.265 ;
        RECT 76.835 138.465 77.165 139.095 ;
        RECT 76.835 137.865 77.085 138.465 ;
        RECT 77.335 138.445 77.565 139.265 ;
        RECT 78.235 138.755 78.540 139.265 ;
        RECT 77.255 138.025 77.585 138.275 ;
        RECT 78.235 138.025 78.550 138.585 ;
        RECT 78.720 138.275 78.970 139.085 ;
        RECT 79.140 138.740 79.400 139.265 ;
        RECT 79.580 138.275 79.830 139.085 ;
        RECT 80.000 138.705 80.260 139.265 ;
        RECT 80.430 138.615 80.690 139.070 ;
        RECT 80.860 138.785 81.120 139.265 ;
        RECT 81.290 138.615 81.550 139.070 ;
        RECT 81.720 138.785 81.980 139.265 ;
        RECT 82.150 138.615 82.410 139.070 ;
        RECT 82.580 138.785 82.825 139.265 ;
        RECT 82.995 138.615 83.270 139.070 ;
        RECT 83.440 138.785 83.685 139.265 ;
        RECT 83.855 138.615 84.115 139.070 ;
        RECT 84.295 138.785 84.545 139.265 ;
        RECT 84.715 138.615 84.975 139.070 ;
        RECT 85.155 138.785 85.405 139.265 ;
        RECT 85.575 138.615 85.835 139.070 ;
        RECT 86.015 138.785 86.275 139.265 ;
        RECT 86.445 138.615 86.705 139.070 ;
        RECT 86.875 138.785 87.175 139.265 ;
        RECT 87.525 138.715 87.695 139.005 ;
        RECT 87.865 138.885 88.195 139.265 ;
        RECT 80.430 138.445 87.175 138.615 ;
        RECT 87.525 138.545 88.190 138.715 ;
        RECT 78.720 138.025 85.840 138.275 ;
        RECT 74.525 137.370 74.710 137.395 ;
        RECT 74.095 137.270 74.710 137.370 ;
        RECT 74.095 136.715 74.700 137.270 ;
        RECT 74.875 136.885 75.355 137.225 ;
        RECT 75.525 136.715 75.780 137.260 ;
        RECT 75.950 136.885 76.225 137.585 ;
        RECT 76.455 136.715 76.665 137.855 ;
        RECT 76.835 136.885 77.165 137.865 ;
        RECT 77.335 136.715 77.565 137.855 ;
        RECT 78.245 136.715 78.540 137.525 ;
        RECT 78.720 136.885 78.965 138.025 ;
        RECT 79.140 136.715 79.400 137.525 ;
        RECT 79.580 136.890 79.830 138.025 ;
        RECT 86.010 137.855 87.175 138.445 ;
        RECT 80.430 137.630 87.175 137.855 ;
        RECT 87.440 137.725 87.790 138.375 ;
        RECT 80.430 137.615 85.835 137.630 ;
        RECT 80.000 136.720 80.260 137.515 ;
        RECT 80.430 136.890 80.690 137.615 ;
        RECT 80.860 136.720 81.120 137.445 ;
        RECT 81.290 136.890 81.550 137.615 ;
        RECT 81.720 136.720 81.980 137.445 ;
        RECT 82.150 136.890 82.410 137.615 ;
        RECT 82.580 136.720 82.840 137.445 ;
        RECT 83.010 136.890 83.270 137.615 ;
        RECT 83.440 136.720 83.685 137.445 ;
        RECT 83.855 136.890 84.115 137.615 ;
        RECT 84.300 136.720 84.545 137.445 ;
        RECT 84.715 136.890 84.975 137.615 ;
        RECT 85.160 136.720 85.405 137.445 ;
        RECT 85.575 136.890 85.835 137.615 ;
        RECT 86.020 136.720 86.275 137.445 ;
        RECT 86.445 136.890 86.735 137.630 ;
        RECT 87.960 137.555 88.190 138.545 ;
        RECT 80.000 136.715 86.275 136.720 ;
        RECT 86.905 136.715 87.175 137.460 ;
        RECT 87.525 137.385 88.190 137.555 ;
        RECT 87.525 136.885 87.695 137.385 ;
        RECT 87.865 136.715 88.195 137.215 ;
        RECT 88.365 136.885 88.550 139.005 ;
        RECT 88.805 138.805 89.055 139.265 ;
        RECT 89.225 138.815 89.560 138.985 ;
        RECT 89.755 138.815 90.430 138.985 ;
        RECT 89.225 138.675 89.395 138.815 ;
        RECT 88.720 137.685 89.000 138.635 ;
        RECT 89.170 138.545 89.395 138.675 ;
        RECT 89.170 137.440 89.340 138.545 ;
        RECT 89.565 138.395 90.090 138.615 ;
        RECT 89.510 137.630 89.750 138.225 ;
        RECT 89.920 137.695 90.090 138.395 ;
        RECT 90.260 138.035 90.430 138.815 ;
        RECT 90.750 138.765 91.120 139.265 ;
        RECT 91.300 138.815 91.705 138.985 ;
        RECT 91.875 138.815 92.660 138.985 ;
        RECT 91.300 138.585 91.470 138.815 ;
        RECT 90.640 138.285 91.470 138.585 ;
        RECT 91.855 138.315 92.320 138.645 ;
        RECT 90.640 138.255 90.840 138.285 ;
        RECT 90.960 138.035 91.130 138.105 ;
        RECT 90.260 137.865 91.130 138.035 ;
        RECT 90.620 137.775 91.130 137.865 ;
        RECT 89.170 137.310 89.475 137.440 ;
        RECT 89.920 137.330 90.450 137.695 ;
        RECT 88.790 136.715 89.055 137.175 ;
        RECT 89.225 136.885 89.475 137.310 ;
        RECT 90.620 137.160 90.790 137.775 ;
        RECT 89.685 136.990 90.790 137.160 ;
        RECT 90.960 136.715 91.130 137.515 ;
        RECT 91.300 137.215 91.470 138.285 ;
        RECT 91.640 137.385 91.830 138.105 ;
        RECT 92.000 137.355 92.320 138.315 ;
        RECT 92.490 138.355 92.660 138.815 ;
        RECT 92.935 138.735 93.145 139.265 ;
        RECT 93.405 138.525 93.735 139.050 ;
        RECT 93.905 138.655 94.075 139.265 ;
        RECT 94.245 138.610 94.575 139.045 ;
        RECT 94.245 138.525 94.625 138.610 ;
        RECT 94.795 138.540 95.085 139.265 ;
        RECT 93.535 138.355 93.735 138.525 ;
        RECT 94.400 138.485 94.625 138.525 ;
        RECT 92.490 138.025 93.365 138.355 ;
        RECT 93.535 138.025 94.285 138.355 ;
        RECT 91.300 136.885 91.550 137.215 ;
        RECT 92.490 137.185 92.660 138.025 ;
        RECT 93.535 137.820 93.725 138.025 ;
        RECT 94.455 137.905 94.625 138.485 ;
        RECT 95.255 138.495 96.925 139.265 ;
        RECT 97.645 138.715 97.815 139.005 ;
        RECT 97.985 138.885 98.315 139.265 ;
        RECT 97.645 138.545 98.310 138.715 ;
        RECT 95.255 137.975 96.005 138.495 ;
        RECT 94.410 137.855 94.625 137.905 ;
        RECT 92.830 137.445 93.725 137.820 ;
        RECT 94.235 137.775 94.625 137.855 ;
        RECT 91.775 137.015 92.660 137.185 ;
        RECT 92.840 136.715 93.155 137.215 ;
        RECT 93.385 136.885 93.725 137.445 ;
        RECT 93.895 136.715 94.065 137.725 ;
        RECT 94.235 136.930 94.565 137.775 ;
        RECT 94.795 136.715 95.085 137.880 ;
        RECT 96.175 137.805 96.925 138.325 ;
        RECT 95.255 136.715 96.925 137.805 ;
        RECT 97.560 137.725 97.910 138.375 ;
        RECT 98.080 137.555 98.310 138.545 ;
        RECT 97.645 137.385 98.310 137.555 ;
        RECT 97.645 136.885 97.815 137.385 ;
        RECT 97.985 136.715 98.315 137.215 ;
        RECT 98.485 136.885 98.670 139.005 ;
        RECT 98.925 138.805 99.175 139.265 ;
        RECT 99.345 138.815 99.680 138.985 ;
        RECT 99.875 138.815 100.550 138.985 ;
        RECT 99.345 138.675 99.515 138.815 ;
        RECT 98.840 137.685 99.120 138.635 ;
        RECT 99.290 138.545 99.515 138.675 ;
        RECT 99.290 137.440 99.460 138.545 ;
        RECT 99.685 138.395 100.210 138.615 ;
        RECT 99.630 137.630 99.870 138.225 ;
        RECT 100.040 137.695 100.210 138.395 ;
        RECT 100.380 138.035 100.550 138.815 ;
        RECT 100.870 138.765 101.240 139.265 ;
        RECT 101.420 138.815 101.825 138.985 ;
        RECT 101.995 138.815 102.780 138.985 ;
        RECT 101.420 138.585 101.590 138.815 ;
        RECT 100.760 138.285 101.590 138.585 ;
        RECT 101.975 138.315 102.440 138.645 ;
        RECT 100.760 138.255 100.960 138.285 ;
        RECT 101.080 138.035 101.250 138.105 ;
        RECT 100.380 137.865 101.250 138.035 ;
        RECT 100.740 137.775 101.250 137.865 ;
        RECT 99.290 137.310 99.595 137.440 ;
        RECT 100.040 137.330 100.570 137.695 ;
        RECT 98.910 136.715 99.175 137.175 ;
        RECT 99.345 136.885 99.595 137.310 ;
        RECT 100.740 137.160 100.910 137.775 ;
        RECT 99.805 136.990 100.910 137.160 ;
        RECT 101.080 136.715 101.250 137.515 ;
        RECT 101.420 137.215 101.590 138.285 ;
        RECT 101.760 137.385 101.950 138.105 ;
        RECT 102.120 137.355 102.440 138.315 ;
        RECT 102.610 138.355 102.780 138.815 ;
        RECT 103.055 138.735 103.265 139.265 ;
        RECT 103.525 138.525 103.855 139.050 ;
        RECT 104.025 138.655 104.195 139.265 ;
        RECT 104.365 138.610 104.695 139.045 ;
        RECT 104.365 138.525 104.745 138.610 ;
        RECT 103.655 138.355 103.855 138.525 ;
        RECT 104.520 138.485 104.745 138.525 ;
        RECT 102.610 138.025 103.485 138.355 ;
        RECT 103.655 138.025 104.405 138.355 ;
        RECT 101.420 136.885 101.670 137.215 ;
        RECT 102.610 137.185 102.780 138.025 ;
        RECT 103.655 137.820 103.845 138.025 ;
        RECT 104.575 137.905 104.745 138.485 ;
        RECT 104.530 137.855 104.745 137.905 ;
        RECT 102.950 137.445 103.845 137.820 ;
        RECT 104.355 137.775 104.745 137.855 ;
        RECT 104.920 138.525 105.175 139.095 ;
        RECT 105.345 138.865 105.675 139.265 ;
        RECT 106.100 138.730 106.630 139.095 ;
        RECT 106.820 138.925 107.095 139.095 ;
        RECT 106.815 138.755 107.095 138.925 ;
        RECT 106.100 138.695 106.275 138.730 ;
        RECT 105.345 138.525 106.275 138.695 ;
        RECT 104.920 137.855 105.090 138.525 ;
        RECT 105.345 138.355 105.515 138.525 ;
        RECT 105.260 138.025 105.515 138.355 ;
        RECT 105.740 138.025 105.935 138.355 ;
        RECT 101.895 137.015 102.780 137.185 ;
        RECT 102.960 136.715 103.275 137.215 ;
        RECT 103.505 136.885 103.845 137.445 ;
        RECT 104.015 136.715 104.185 137.725 ;
        RECT 104.355 136.930 104.685 137.775 ;
        RECT 104.920 136.885 105.255 137.855 ;
        RECT 105.425 136.715 105.595 137.855 ;
        RECT 105.765 137.055 105.935 138.025 ;
        RECT 106.105 137.395 106.275 138.525 ;
        RECT 106.445 137.735 106.615 138.535 ;
        RECT 106.820 137.935 107.095 138.755 ;
        RECT 107.265 137.735 107.455 139.095 ;
        RECT 107.635 138.730 108.145 139.265 ;
        RECT 108.365 138.455 108.610 139.060 ;
        RECT 109.060 138.525 109.315 139.095 ;
        RECT 109.485 138.865 109.815 139.265 ;
        RECT 110.240 138.730 110.770 139.095 ;
        RECT 110.960 138.925 111.235 139.095 ;
        RECT 110.955 138.755 111.235 138.925 ;
        RECT 110.240 138.695 110.415 138.730 ;
        RECT 109.485 138.525 110.415 138.695 ;
        RECT 107.655 138.285 108.885 138.455 ;
        RECT 106.445 137.565 107.455 137.735 ;
        RECT 107.625 137.720 108.375 137.910 ;
        RECT 106.105 137.225 107.230 137.395 ;
        RECT 107.625 137.055 107.795 137.720 ;
        RECT 108.545 137.475 108.885 138.285 ;
        RECT 105.765 136.885 107.795 137.055 ;
        RECT 107.965 136.715 108.135 137.475 ;
        RECT 108.370 137.065 108.885 137.475 ;
        RECT 109.060 137.855 109.230 138.525 ;
        RECT 109.485 138.355 109.655 138.525 ;
        RECT 109.400 138.025 109.655 138.355 ;
        RECT 109.880 138.025 110.075 138.355 ;
        RECT 109.060 136.885 109.395 137.855 ;
        RECT 109.565 136.715 109.735 137.855 ;
        RECT 109.905 137.055 110.075 138.025 ;
        RECT 110.245 137.395 110.415 138.525 ;
        RECT 110.585 137.735 110.755 138.535 ;
        RECT 110.960 137.935 111.235 138.755 ;
        RECT 111.405 137.735 111.595 139.095 ;
        RECT 111.775 138.730 112.285 139.265 ;
        RECT 112.505 138.455 112.750 139.060 ;
        RECT 113.285 138.715 113.455 139.005 ;
        RECT 113.625 138.885 113.955 139.265 ;
        RECT 113.285 138.545 113.950 138.715 ;
        RECT 111.795 138.285 113.025 138.455 ;
        RECT 110.585 137.565 111.595 137.735 ;
        RECT 111.765 137.720 112.515 137.910 ;
        RECT 110.245 137.225 111.370 137.395 ;
        RECT 111.765 137.055 111.935 137.720 ;
        RECT 112.685 137.475 113.025 138.285 ;
        RECT 113.200 137.725 113.550 138.375 ;
        RECT 113.720 137.555 113.950 138.545 ;
        RECT 109.905 136.885 111.935 137.055 ;
        RECT 112.105 136.715 112.275 137.475 ;
        RECT 112.510 137.065 113.025 137.475 ;
        RECT 113.285 137.385 113.950 137.555 ;
        RECT 113.285 136.885 113.455 137.385 ;
        RECT 113.625 136.715 113.955 137.215 ;
        RECT 114.125 136.885 114.310 139.005 ;
        RECT 114.565 138.805 114.815 139.265 ;
        RECT 114.985 138.815 115.320 138.985 ;
        RECT 115.515 138.815 116.190 138.985 ;
        RECT 114.985 138.675 115.155 138.815 ;
        RECT 114.480 137.685 114.760 138.635 ;
        RECT 114.930 138.545 115.155 138.675 ;
        RECT 114.930 137.440 115.100 138.545 ;
        RECT 115.325 138.395 115.850 138.615 ;
        RECT 115.270 137.630 115.510 138.225 ;
        RECT 115.680 137.695 115.850 138.395 ;
        RECT 116.020 138.035 116.190 138.815 ;
        RECT 116.510 138.765 116.880 139.265 ;
        RECT 117.060 138.815 117.465 138.985 ;
        RECT 117.635 138.815 118.420 138.985 ;
        RECT 117.060 138.585 117.230 138.815 ;
        RECT 116.400 138.285 117.230 138.585 ;
        RECT 117.615 138.315 118.080 138.645 ;
        RECT 116.400 138.255 116.600 138.285 ;
        RECT 116.720 138.035 116.890 138.105 ;
        RECT 116.020 137.865 116.890 138.035 ;
        RECT 116.380 137.775 116.890 137.865 ;
        RECT 114.930 137.310 115.235 137.440 ;
        RECT 115.680 137.330 116.210 137.695 ;
        RECT 114.550 136.715 114.815 137.175 ;
        RECT 114.985 136.885 115.235 137.310 ;
        RECT 116.380 137.160 116.550 137.775 ;
        RECT 115.445 136.990 116.550 137.160 ;
        RECT 116.720 136.715 116.890 137.515 ;
        RECT 117.060 137.215 117.230 138.285 ;
        RECT 117.400 137.385 117.590 138.105 ;
        RECT 117.760 137.355 118.080 138.315 ;
        RECT 118.250 138.355 118.420 138.815 ;
        RECT 118.695 138.735 118.905 139.265 ;
        RECT 119.165 138.525 119.495 139.050 ;
        RECT 119.665 138.655 119.835 139.265 ;
        RECT 120.005 138.610 120.335 139.045 ;
        RECT 120.005 138.525 120.385 138.610 ;
        RECT 120.555 138.540 120.845 139.265 ;
        RECT 121.105 138.715 121.275 139.005 ;
        RECT 121.445 138.885 121.775 139.265 ;
        RECT 121.105 138.545 121.770 138.715 ;
        RECT 119.295 138.355 119.495 138.525 ;
        RECT 120.160 138.485 120.385 138.525 ;
        RECT 118.250 138.025 119.125 138.355 ;
        RECT 119.295 138.025 120.045 138.355 ;
        RECT 117.060 136.885 117.310 137.215 ;
        RECT 118.250 137.185 118.420 138.025 ;
        RECT 119.295 137.820 119.485 138.025 ;
        RECT 120.215 137.905 120.385 138.485 ;
        RECT 120.170 137.855 120.385 137.905 ;
        RECT 118.590 137.445 119.485 137.820 ;
        RECT 119.995 137.775 120.385 137.855 ;
        RECT 117.535 137.015 118.420 137.185 ;
        RECT 118.600 136.715 118.915 137.215 ;
        RECT 119.145 136.885 119.485 137.445 ;
        RECT 119.655 136.715 119.825 137.725 ;
        RECT 119.995 136.930 120.325 137.775 ;
        RECT 120.555 136.715 120.845 137.880 ;
        RECT 121.020 137.725 121.370 138.375 ;
        RECT 121.540 137.555 121.770 138.545 ;
        RECT 121.105 137.385 121.770 137.555 ;
        RECT 121.105 136.885 121.275 137.385 ;
        RECT 121.445 136.715 121.775 137.215 ;
        RECT 121.945 136.885 122.130 139.005 ;
        RECT 122.385 138.805 122.635 139.265 ;
        RECT 122.805 138.815 123.140 138.985 ;
        RECT 123.335 138.815 124.010 138.985 ;
        RECT 122.805 138.675 122.975 138.815 ;
        RECT 122.300 137.685 122.580 138.635 ;
        RECT 122.750 138.545 122.975 138.675 ;
        RECT 122.750 137.440 122.920 138.545 ;
        RECT 123.145 138.395 123.670 138.615 ;
        RECT 123.090 137.630 123.330 138.225 ;
        RECT 123.500 137.695 123.670 138.395 ;
        RECT 123.840 138.035 124.010 138.815 ;
        RECT 124.330 138.765 124.700 139.265 ;
        RECT 124.880 138.815 125.285 138.985 ;
        RECT 125.455 138.815 126.240 138.985 ;
        RECT 124.880 138.585 125.050 138.815 ;
        RECT 124.220 138.285 125.050 138.585 ;
        RECT 125.435 138.315 125.900 138.645 ;
        RECT 124.220 138.255 124.420 138.285 ;
        RECT 124.540 138.035 124.710 138.105 ;
        RECT 123.840 137.865 124.710 138.035 ;
        RECT 124.200 137.775 124.710 137.865 ;
        RECT 122.750 137.310 123.055 137.440 ;
        RECT 123.500 137.330 124.030 137.695 ;
        RECT 122.370 136.715 122.635 137.175 ;
        RECT 122.805 136.885 123.055 137.310 ;
        RECT 124.200 137.160 124.370 137.775 ;
        RECT 123.265 136.990 124.370 137.160 ;
        RECT 124.540 136.715 124.710 137.515 ;
        RECT 124.880 137.215 125.050 138.285 ;
        RECT 125.220 137.385 125.410 138.105 ;
        RECT 125.580 137.355 125.900 138.315 ;
        RECT 126.070 138.355 126.240 138.815 ;
        RECT 126.515 138.735 126.725 139.265 ;
        RECT 126.985 138.525 127.315 139.050 ;
        RECT 127.485 138.655 127.655 139.265 ;
        RECT 127.825 138.610 128.155 139.045 ;
        RECT 127.825 138.525 128.205 138.610 ;
        RECT 127.115 138.355 127.315 138.525 ;
        RECT 127.980 138.485 128.205 138.525 ;
        RECT 126.070 138.025 126.945 138.355 ;
        RECT 127.115 138.025 127.865 138.355 ;
        RECT 124.880 136.885 125.130 137.215 ;
        RECT 126.070 137.185 126.240 138.025 ;
        RECT 127.115 137.820 127.305 138.025 ;
        RECT 128.035 137.905 128.205 138.485 ;
        RECT 128.375 138.495 130.045 139.265 ;
        RECT 128.375 137.975 129.125 138.495 ;
        RECT 130.420 138.485 130.920 139.095 ;
        RECT 127.990 137.855 128.205 137.905 ;
        RECT 126.410 137.445 127.305 137.820 ;
        RECT 127.815 137.775 128.205 137.855 ;
        RECT 129.295 137.805 130.045 138.325 ;
        RECT 130.215 138.025 130.565 138.275 ;
        RECT 130.750 137.855 130.920 138.485 ;
        RECT 131.550 138.615 131.880 139.095 ;
        RECT 132.050 138.805 132.275 139.265 ;
        RECT 132.445 138.615 132.775 139.095 ;
        RECT 131.550 138.445 132.775 138.615 ;
        RECT 132.965 138.465 133.215 139.265 ;
        RECT 133.385 138.465 133.725 139.095 ;
        RECT 134.060 138.755 134.300 139.265 ;
        RECT 134.480 138.755 134.760 139.085 ;
        RECT 134.990 138.755 135.205 139.265 ;
        RECT 131.090 138.075 131.420 138.275 ;
        RECT 131.590 138.075 131.920 138.275 ;
        RECT 132.090 138.075 132.510 138.275 ;
        RECT 132.685 138.105 133.380 138.275 ;
        RECT 132.685 137.855 132.855 138.105 ;
        RECT 133.550 137.855 133.725 138.465 ;
        RECT 133.955 138.025 134.310 138.585 ;
        RECT 134.480 137.855 134.650 138.755 ;
        RECT 134.820 138.025 135.085 138.585 ;
        RECT 135.375 138.525 135.990 139.095 ;
        RECT 135.335 137.855 135.505 138.355 ;
        RECT 125.355 137.015 126.240 137.185 ;
        RECT 126.420 136.715 126.735 137.215 ;
        RECT 126.965 136.885 127.305 137.445 ;
        RECT 127.475 136.715 127.645 137.725 ;
        RECT 127.815 136.930 128.145 137.775 ;
        RECT 128.375 136.715 130.045 137.805 ;
        RECT 130.420 137.685 132.855 137.855 ;
        RECT 130.420 136.885 130.750 137.685 ;
        RECT 130.920 136.715 131.250 137.515 ;
        RECT 131.550 136.885 131.880 137.685 ;
        RECT 132.525 136.715 132.775 137.515 ;
        RECT 133.045 136.715 133.215 137.855 ;
        RECT 133.385 136.885 133.725 137.855 ;
        RECT 134.080 137.685 135.505 137.855 ;
        RECT 134.080 137.510 134.470 137.685 ;
        RECT 134.955 136.715 135.285 137.515 ;
        RECT 135.675 137.505 135.990 138.525 ;
        RECT 136.195 138.495 137.865 139.265 ;
        RECT 138.125 138.715 138.295 139.095 ;
        RECT 138.510 138.885 138.840 139.265 ;
        RECT 138.125 138.545 138.840 138.715 ;
        RECT 136.195 137.975 136.945 138.495 ;
        RECT 137.115 137.805 137.865 138.325 ;
        RECT 138.035 137.995 138.390 138.365 ;
        RECT 138.670 138.355 138.840 138.545 ;
        RECT 139.010 138.520 139.265 139.095 ;
        RECT 138.670 138.025 138.925 138.355 ;
        RECT 138.670 137.815 138.840 138.025 ;
        RECT 135.455 136.885 135.990 137.505 ;
        RECT 136.195 136.715 137.865 137.805 ;
        RECT 138.125 137.645 138.840 137.815 ;
        RECT 139.095 137.790 139.265 138.520 ;
        RECT 139.440 138.425 139.700 139.265 ;
        RECT 139.965 138.715 140.135 139.095 ;
        RECT 140.350 138.885 140.680 139.265 ;
        RECT 139.965 138.545 140.680 138.715 ;
        RECT 139.875 137.995 140.230 138.365 ;
        RECT 140.510 138.355 140.680 138.545 ;
        RECT 140.850 138.520 141.105 139.095 ;
        RECT 140.510 138.025 140.765 138.355 ;
        RECT 138.125 136.885 138.295 137.645 ;
        RECT 138.510 136.715 138.840 137.475 ;
        RECT 139.010 136.885 139.265 137.790 ;
        RECT 139.440 136.715 139.700 137.865 ;
        RECT 140.510 137.815 140.680 138.025 ;
        RECT 139.965 137.645 140.680 137.815 ;
        RECT 140.935 137.790 141.105 138.520 ;
        RECT 141.280 138.425 141.540 139.265 ;
        RECT 141.715 138.515 142.925 139.265 ;
        RECT 139.965 136.885 140.135 137.645 ;
        RECT 140.350 136.715 140.680 137.475 ;
        RECT 140.850 136.885 141.105 137.790 ;
        RECT 141.280 136.715 141.540 137.865 ;
        RECT 141.715 137.805 142.235 138.345 ;
        RECT 142.405 137.975 142.925 138.515 ;
        RECT 141.715 136.715 142.925 137.805 ;
        RECT 17.430 136.545 143.010 136.715 ;
        RECT 17.515 135.455 18.725 136.545 ;
        RECT 18.895 135.455 22.405 136.545 ;
        RECT 17.515 134.745 18.035 135.285 ;
        RECT 18.205 134.915 18.725 135.455 ;
        RECT 18.895 134.765 20.545 135.285 ;
        RECT 20.715 134.935 22.405 135.455 ;
        RECT 22.575 135.675 22.850 136.375 ;
        RECT 23.020 136.000 23.275 136.545 ;
        RECT 23.445 136.035 23.925 136.375 ;
        RECT 24.100 135.990 24.705 136.545 ;
        RECT 24.875 136.110 30.220 136.545 ;
        RECT 24.090 135.890 24.705 135.990 ;
        RECT 24.090 135.865 24.275 135.890 ;
        RECT 17.515 133.995 18.725 134.745 ;
        RECT 18.895 133.995 22.405 134.765 ;
        RECT 22.575 134.645 22.745 135.675 ;
        RECT 23.020 135.545 23.775 135.795 ;
        RECT 23.945 135.620 24.275 135.865 ;
        RECT 23.020 135.510 23.790 135.545 ;
        RECT 23.020 135.500 23.805 135.510 ;
        RECT 22.915 135.485 23.810 135.500 ;
        RECT 22.915 135.470 23.830 135.485 ;
        RECT 22.915 135.460 23.850 135.470 ;
        RECT 22.915 135.450 23.875 135.460 ;
        RECT 22.915 135.420 23.945 135.450 ;
        RECT 22.915 135.390 23.965 135.420 ;
        RECT 22.915 135.360 23.985 135.390 ;
        RECT 22.915 135.335 24.015 135.360 ;
        RECT 22.915 135.300 24.050 135.335 ;
        RECT 22.915 135.295 24.080 135.300 ;
        RECT 22.915 134.900 23.145 135.295 ;
        RECT 23.690 135.290 24.080 135.295 ;
        RECT 23.715 135.280 24.080 135.290 ;
        RECT 23.730 135.275 24.080 135.280 ;
        RECT 23.745 135.270 24.080 135.275 ;
        RECT 24.445 135.270 24.705 135.720 ;
        RECT 23.745 135.265 24.705 135.270 ;
        RECT 23.755 135.255 24.705 135.265 ;
        RECT 23.765 135.250 24.705 135.255 ;
        RECT 23.775 135.240 24.705 135.250 ;
        RECT 23.780 135.230 24.705 135.240 ;
        RECT 23.785 135.225 24.705 135.230 ;
        RECT 23.795 135.210 24.705 135.225 ;
        RECT 23.800 135.195 24.705 135.210 ;
        RECT 23.810 135.170 24.705 135.195 ;
        RECT 23.315 134.700 23.645 135.125 ;
        RECT 22.575 134.165 22.835 134.645 ;
        RECT 23.005 133.995 23.255 134.535 ;
        RECT 23.425 134.215 23.645 134.700 ;
        RECT 23.815 135.100 24.705 135.170 ;
        RECT 23.815 134.375 23.985 135.100 ;
        RECT 24.155 134.545 24.705 134.930 ;
        RECT 26.460 134.540 26.800 135.370 ;
        RECT 28.280 134.860 28.630 136.110 ;
        RECT 30.395 135.380 30.685 136.545 ;
        RECT 30.855 136.110 36.200 136.545 ;
        RECT 23.815 134.205 24.705 134.375 ;
        RECT 24.875 133.995 30.220 134.540 ;
        RECT 30.395 133.995 30.685 134.720 ;
        RECT 32.440 134.540 32.780 135.370 ;
        RECT 34.260 134.860 34.610 136.110 ;
        RECT 36.375 135.455 37.585 136.545 ;
        RECT 36.375 134.745 36.895 135.285 ;
        RECT 37.065 134.915 37.585 135.455 ;
        RECT 37.755 134.980 38.105 136.375 ;
        RECT 38.275 135.745 38.680 136.545 ;
        RECT 38.850 136.205 40.385 136.375 ;
        RECT 38.850 135.575 39.020 136.205 ;
        RECT 38.275 135.405 39.020 135.575 ;
        RECT 30.855 133.995 36.200 134.540 ;
        RECT 36.375 133.995 37.585 134.745 ;
        RECT 37.755 134.165 38.025 134.980 ;
        RECT 38.275 134.905 38.445 135.405 ;
        RECT 39.190 135.235 39.460 135.980 ;
        RECT 38.615 134.905 38.950 135.235 ;
        RECT 39.120 134.905 39.460 135.235 ;
        RECT 39.650 135.235 39.885 135.980 ;
        RECT 40.055 135.575 40.385 136.205 ;
        RECT 40.570 135.745 40.805 136.545 ;
        RECT 40.975 135.575 41.265 136.375 ;
        RECT 41.635 135.875 41.915 136.545 ;
        RECT 42.085 135.655 42.385 136.205 ;
        RECT 42.585 135.825 42.915 136.545 ;
        RECT 43.105 135.825 43.565 136.375 ;
        RECT 40.055 135.405 41.265 135.575 ;
        RECT 39.650 134.905 39.940 135.235 ;
        RECT 40.110 134.905 40.510 135.235 ;
        RECT 40.680 134.735 40.850 135.405 ;
        RECT 41.450 135.235 41.715 135.595 ;
        RECT 42.085 135.485 43.025 135.655 ;
        RECT 42.855 135.235 43.025 135.485 ;
        RECT 41.020 134.905 41.265 135.235 ;
        RECT 41.450 134.985 42.125 135.235 ;
        RECT 42.345 134.985 42.685 135.235 ;
        RECT 42.855 134.905 43.145 135.235 ;
        RECT 42.855 134.815 43.025 134.905 ;
        RECT 38.195 133.995 38.865 134.735 ;
        RECT 39.035 134.565 40.430 134.735 ;
        RECT 39.035 134.220 39.330 134.565 ;
        RECT 39.510 133.995 39.885 134.395 ;
        RECT 40.100 134.220 40.430 134.565 ;
        RECT 40.680 134.165 41.265 134.735 ;
        RECT 41.635 134.625 43.025 134.815 ;
        RECT 41.635 134.265 41.965 134.625 ;
        RECT 43.315 134.455 43.565 135.825 ;
        RECT 43.735 135.455 46.325 136.545 ;
        RECT 42.585 133.995 42.835 134.455 ;
        RECT 43.005 134.165 43.565 134.455 ;
        RECT 43.735 134.765 44.945 135.285 ;
        RECT 45.115 134.935 46.325 135.455 ;
        RECT 46.495 135.405 46.765 136.375 ;
        RECT 46.975 135.745 47.255 136.545 ;
        RECT 47.425 136.035 49.080 136.325 ;
        RECT 47.490 135.695 49.080 135.865 ;
        RECT 47.490 135.575 47.660 135.695 ;
        RECT 46.935 135.405 47.660 135.575 ;
        RECT 43.735 133.995 46.325 134.765 ;
        RECT 46.495 134.670 46.665 135.405 ;
        RECT 46.935 135.235 47.105 135.405 ;
        RECT 46.835 134.905 47.105 135.235 ;
        RECT 47.275 134.905 47.680 135.235 ;
        RECT 47.850 134.905 48.560 135.525 ;
        RECT 48.760 135.405 49.080 135.695 ;
        RECT 49.255 135.405 49.515 136.375 ;
        RECT 49.710 136.135 50.040 136.545 ;
        RECT 50.240 135.955 50.410 136.375 ;
        RECT 50.625 136.135 51.295 136.545 ;
        RECT 51.530 135.955 51.700 136.375 ;
        RECT 52.005 136.105 52.335 136.545 ;
        RECT 49.685 135.785 51.700 135.955 ;
        RECT 52.505 135.925 52.680 136.375 ;
        RECT 46.935 134.735 47.105 134.905 ;
        RECT 46.495 134.325 46.765 134.670 ;
        RECT 46.935 134.565 48.545 134.735 ;
        RECT 48.730 134.665 49.080 135.235 ;
        RECT 49.255 134.715 49.425 135.405 ;
        RECT 49.685 135.235 49.855 135.785 ;
        RECT 49.595 134.905 49.855 135.235 ;
        RECT 46.955 133.995 47.335 134.395 ;
        RECT 47.505 134.215 47.675 134.565 ;
        RECT 47.845 133.995 48.175 134.395 ;
        RECT 48.375 134.215 48.545 134.565 ;
        RECT 48.745 133.995 49.075 134.495 ;
        RECT 49.255 134.250 49.595 134.715 ;
        RECT 50.025 134.575 50.365 135.605 ;
        RECT 50.555 135.185 50.825 135.605 ;
        RECT 50.555 135.015 50.865 135.185 ;
        RECT 49.260 134.205 49.595 134.250 ;
        RECT 49.765 133.995 50.095 134.375 ;
        RECT 50.555 134.330 50.825 135.015 ;
        RECT 51.050 134.330 51.330 135.605 ;
        RECT 51.530 134.495 51.700 135.785 ;
        RECT 52.050 135.755 52.680 135.925 ;
        RECT 52.050 135.235 52.220 135.755 ;
        RECT 51.870 134.905 52.220 135.235 ;
        RECT 52.400 134.905 52.765 135.585 ;
        RECT 52.050 134.735 52.220 134.905 ;
        RECT 52.050 134.565 52.680 134.735 ;
        RECT 51.530 134.165 51.760 134.495 ;
        RECT 52.005 133.995 52.335 134.375 ;
        RECT 52.505 134.165 52.680 134.565 ;
        RECT 52.935 134.275 53.215 136.375 ;
        RECT 53.405 135.785 54.190 136.545 ;
        RECT 54.585 135.715 54.970 136.375 ;
        RECT 54.585 135.615 54.995 135.715 ;
        RECT 53.385 135.405 54.995 135.615 ;
        RECT 55.295 135.525 55.495 136.315 ;
        RECT 53.385 134.805 53.660 135.405 ;
        RECT 55.165 135.355 55.495 135.525 ;
        RECT 55.665 135.365 55.985 136.545 ;
        RECT 56.155 135.380 56.445 136.545 ;
        RECT 56.625 135.935 56.955 136.365 ;
        RECT 57.135 136.105 57.330 136.545 ;
        RECT 57.500 135.935 57.830 136.365 ;
        RECT 56.625 135.765 57.830 135.935 ;
        RECT 56.625 135.435 57.520 135.765 ;
        RECT 58.000 135.595 58.275 136.365 ;
        RECT 58.455 136.110 63.800 136.545 ;
        RECT 63.975 136.110 69.320 136.545 ;
        RECT 57.690 135.405 58.275 135.595 ;
        RECT 55.165 135.235 55.345 135.355 ;
        RECT 53.830 134.985 54.185 135.235 ;
        RECT 54.380 135.185 54.845 135.235 ;
        RECT 54.375 135.015 54.845 135.185 ;
        RECT 54.380 134.985 54.845 135.015 ;
        RECT 55.015 134.985 55.345 135.235 ;
        RECT 55.520 134.985 55.985 135.185 ;
        RECT 56.630 134.905 56.925 135.235 ;
        RECT 57.105 134.905 57.520 135.235 ;
        RECT 53.385 134.625 54.635 134.805 ;
        RECT 54.270 134.555 54.635 134.625 ;
        RECT 54.805 134.605 55.985 134.775 ;
        RECT 53.445 133.995 53.615 134.455 ;
        RECT 54.805 134.385 55.135 134.605 ;
        RECT 53.885 134.205 55.135 134.385 ;
        RECT 55.305 133.995 55.475 134.435 ;
        RECT 55.645 134.190 55.985 134.605 ;
        RECT 56.155 133.995 56.445 134.720 ;
        RECT 56.625 133.995 56.925 134.725 ;
        RECT 57.105 134.285 57.335 134.905 ;
        RECT 57.690 134.735 57.865 135.405 ;
        RECT 57.535 134.555 57.865 134.735 ;
        RECT 58.035 134.585 58.275 135.235 ;
        RECT 57.535 134.175 57.760 134.555 ;
        RECT 60.040 134.540 60.380 135.370 ;
        RECT 61.860 134.860 62.210 136.110 ;
        RECT 65.560 134.540 65.900 135.370 ;
        RECT 67.380 134.860 67.730 136.110 ;
        RECT 69.495 135.455 72.085 136.545 ;
        RECT 69.495 134.765 70.705 135.285 ;
        RECT 70.875 134.935 72.085 135.455 ;
        RECT 72.255 135.825 72.715 136.375 ;
        RECT 72.905 135.825 73.235 136.545 ;
        RECT 57.930 133.995 58.260 134.385 ;
        RECT 58.455 133.995 63.800 134.540 ;
        RECT 63.975 133.995 69.320 134.540 ;
        RECT 69.495 133.995 72.085 134.765 ;
        RECT 72.255 134.455 72.505 135.825 ;
        RECT 73.435 135.655 73.735 136.205 ;
        RECT 73.905 135.875 74.185 136.545 ;
        RECT 72.795 135.485 73.735 135.655 ;
        RECT 72.795 135.235 72.965 135.485 ;
        RECT 74.105 135.235 74.370 135.595 ;
        RECT 74.555 135.455 77.145 136.545 ;
        RECT 72.675 134.905 72.965 135.235 ;
        RECT 73.135 134.985 73.475 135.235 ;
        RECT 73.695 134.985 74.370 135.235 ;
        RECT 72.795 134.815 72.965 134.905 ;
        RECT 72.795 134.625 74.185 134.815 ;
        RECT 72.255 134.165 72.815 134.455 ;
        RECT 72.985 133.995 73.235 134.455 ;
        RECT 73.855 134.265 74.185 134.625 ;
        RECT 74.555 134.765 75.765 135.285 ;
        RECT 75.935 134.935 77.145 135.455 ;
        RECT 77.775 135.785 78.290 136.195 ;
        RECT 78.525 135.785 78.695 136.545 ;
        RECT 78.865 136.205 80.895 136.375 ;
        RECT 77.775 134.975 78.115 135.785 ;
        RECT 78.865 135.540 79.035 136.205 ;
        RECT 79.430 135.865 80.555 136.035 ;
        RECT 78.285 135.350 79.035 135.540 ;
        RECT 79.205 135.525 80.215 135.695 ;
        RECT 77.775 134.805 79.005 134.975 ;
        RECT 74.555 133.995 77.145 134.765 ;
        RECT 78.050 134.200 78.295 134.805 ;
        RECT 78.515 133.995 79.025 134.530 ;
        RECT 79.205 134.165 79.395 135.525 ;
        RECT 79.565 135.185 79.840 135.325 ;
        RECT 79.565 135.015 79.845 135.185 ;
        RECT 79.565 134.165 79.840 135.015 ;
        RECT 80.045 134.725 80.215 135.525 ;
        RECT 80.385 134.735 80.555 135.865 ;
        RECT 80.725 135.235 80.895 136.205 ;
        RECT 81.065 135.405 81.235 136.545 ;
        RECT 81.405 135.405 81.740 136.375 ;
        RECT 80.725 134.905 80.920 135.235 ;
        RECT 81.145 134.905 81.400 135.235 ;
        RECT 81.145 134.735 81.315 134.905 ;
        RECT 81.570 134.735 81.740 135.405 ;
        RECT 81.915 135.380 82.205 136.545 ;
        RECT 82.375 135.455 85.885 136.545 ;
        RECT 80.385 134.565 81.315 134.735 ;
        RECT 80.385 134.530 80.560 134.565 ;
        RECT 80.030 134.165 80.560 134.530 ;
        RECT 80.985 133.995 81.315 134.395 ;
        RECT 81.485 134.165 81.740 134.735 ;
        RECT 82.375 134.765 84.025 135.285 ;
        RECT 84.195 134.935 85.885 135.455 ;
        RECT 86.055 135.785 86.570 136.195 ;
        RECT 86.805 135.785 86.975 136.545 ;
        RECT 87.145 136.205 89.175 136.375 ;
        RECT 86.055 134.975 86.395 135.785 ;
        RECT 87.145 135.540 87.315 136.205 ;
        RECT 87.710 135.865 88.835 136.035 ;
        RECT 86.565 135.350 87.315 135.540 ;
        RECT 87.485 135.525 88.495 135.695 ;
        RECT 86.055 134.805 87.285 134.975 ;
        RECT 81.915 133.995 82.205 134.720 ;
        RECT 82.375 133.995 85.885 134.765 ;
        RECT 86.330 134.200 86.575 134.805 ;
        RECT 86.795 133.995 87.305 134.530 ;
        RECT 87.485 134.165 87.675 135.525 ;
        RECT 87.845 134.505 88.120 135.325 ;
        RECT 88.325 134.725 88.495 135.525 ;
        RECT 88.665 134.735 88.835 135.865 ;
        RECT 89.005 135.235 89.175 136.205 ;
        RECT 89.345 135.405 89.515 136.545 ;
        RECT 89.685 135.405 90.020 136.375 ;
        RECT 89.005 134.905 89.200 135.235 ;
        RECT 89.425 134.905 89.680 135.235 ;
        RECT 89.425 134.735 89.595 134.905 ;
        RECT 89.850 134.735 90.020 135.405 ;
        RECT 88.665 134.565 89.595 134.735 ;
        RECT 88.665 134.530 88.840 134.565 ;
        RECT 87.845 134.335 88.125 134.505 ;
        RECT 87.845 134.165 88.120 134.335 ;
        RECT 88.310 134.165 88.840 134.530 ;
        RECT 89.265 133.995 89.595 134.395 ;
        RECT 89.765 134.165 90.020 134.735 ;
        RECT 90.195 135.405 90.580 136.375 ;
        RECT 90.750 136.085 91.075 136.545 ;
        RECT 91.595 135.915 91.875 136.375 ;
        RECT 90.750 135.695 91.875 135.915 ;
        RECT 90.195 134.735 90.475 135.405 ;
        RECT 90.750 135.235 91.200 135.695 ;
        RECT 92.065 135.525 92.465 136.375 ;
        RECT 92.865 136.085 93.135 136.545 ;
        RECT 93.305 135.915 93.590 136.375 ;
        RECT 90.645 134.905 91.200 135.235 ;
        RECT 91.370 134.965 92.465 135.525 ;
        RECT 90.750 134.795 91.200 134.905 ;
        RECT 90.195 134.165 90.580 134.735 ;
        RECT 90.750 134.625 91.875 134.795 ;
        RECT 90.750 133.995 91.075 134.455 ;
        RECT 91.595 134.165 91.875 134.625 ;
        RECT 92.065 134.165 92.465 134.965 ;
        RECT 92.635 135.695 93.590 135.915 ;
        RECT 92.635 134.795 92.845 135.695 ;
        RECT 93.015 134.965 93.705 135.525 ;
        RECT 93.875 135.455 97.385 136.545 ;
        RECT 97.645 135.875 97.815 136.375 ;
        RECT 97.985 136.045 98.315 136.545 ;
        RECT 97.645 135.705 98.310 135.875 ;
        RECT 92.635 134.625 93.590 134.795 ;
        RECT 92.865 133.995 93.135 134.455 ;
        RECT 93.305 134.165 93.590 134.625 ;
        RECT 93.875 134.765 95.525 135.285 ;
        RECT 95.695 134.935 97.385 135.455 ;
        RECT 97.560 134.885 97.910 135.535 ;
        RECT 93.875 133.995 97.385 134.765 ;
        RECT 98.080 134.715 98.310 135.705 ;
        RECT 97.645 134.545 98.310 134.715 ;
        RECT 97.645 134.255 97.815 134.545 ;
        RECT 97.985 133.995 98.315 134.375 ;
        RECT 98.485 134.255 98.670 136.375 ;
        RECT 98.910 136.085 99.175 136.545 ;
        RECT 99.345 135.950 99.595 136.375 ;
        RECT 99.805 136.100 100.910 136.270 ;
        RECT 99.290 135.820 99.595 135.950 ;
        RECT 98.840 134.625 99.120 135.575 ;
        RECT 99.290 134.715 99.460 135.820 ;
        RECT 99.630 135.035 99.870 135.630 ;
        RECT 100.040 135.565 100.570 135.930 ;
        RECT 100.040 134.865 100.210 135.565 ;
        RECT 100.740 135.485 100.910 136.100 ;
        RECT 101.080 135.745 101.250 136.545 ;
        RECT 101.420 136.045 101.670 136.375 ;
        RECT 101.895 136.075 102.780 136.245 ;
        RECT 100.740 135.395 101.250 135.485 ;
        RECT 99.290 134.585 99.515 134.715 ;
        RECT 99.685 134.645 100.210 134.865 ;
        RECT 100.380 135.225 101.250 135.395 ;
        RECT 98.925 133.995 99.175 134.455 ;
        RECT 99.345 134.445 99.515 134.585 ;
        RECT 100.380 134.445 100.550 135.225 ;
        RECT 101.080 135.155 101.250 135.225 ;
        RECT 100.760 134.975 100.960 135.005 ;
        RECT 101.420 134.975 101.590 136.045 ;
        RECT 101.760 135.155 101.950 135.875 ;
        RECT 100.760 134.675 101.590 134.975 ;
        RECT 102.120 134.945 102.440 135.905 ;
        RECT 99.345 134.275 99.680 134.445 ;
        RECT 99.875 134.275 100.550 134.445 ;
        RECT 100.870 133.995 101.240 134.495 ;
        RECT 101.420 134.445 101.590 134.675 ;
        RECT 101.975 134.615 102.440 134.945 ;
        RECT 102.610 135.235 102.780 136.075 ;
        RECT 102.960 136.045 103.275 136.545 ;
        RECT 103.505 135.815 103.845 136.375 ;
        RECT 102.950 135.440 103.845 135.815 ;
        RECT 104.015 135.535 104.185 136.545 ;
        RECT 103.655 135.235 103.845 135.440 ;
        RECT 104.355 135.485 104.685 136.330 ;
        RECT 104.355 135.405 104.745 135.485 ;
        RECT 104.915 135.455 107.505 136.545 ;
        RECT 104.530 135.355 104.745 135.405 ;
        RECT 102.610 134.905 103.485 135.235 ;
        RECT 103.655 134.905 104.405 135.235 ;
        RECT 102.610 134.445 102.780 134.905 ;
        RECT 103.655 134.735 103.855 134.905 ;
        RECT 104.575 134.775 104.745 135.355 ;
        RECT 104.520 134.735 104.745 134.775 ;
        RECT 101.420 134.275 101.825 134.445 ;
        RECT 101.995 134.275 102.780 134.445 ;
        RECT 103.055 133.995 103.265 134.525 ;
        RECT 103.525 134.210 103.855 134.735 ;
        RECT 104.365 134.650 104.745 134.735 ;
        RECT 104.915 134.765 106.125 135.285 ;
        RECT 106.295 134.935 107.505 135.455 ;
        RECT 107.675 135.380 107.965 136.545 ;
        RECT 108.135 135.405 108.520 136.375 ;
        RECT 108.690 136.085 109.015 136.545 ;
        RECT 109.535 135.915 109.815 136.375 ;
        RECT 108.690 135.695 109.815 135.915 ;
        RECT 104.025 133.995 104.195 134.605 ;
        RECT 104.365 134.215 104.695 134.650 ;
        RECT 104.915 133.995 107.505 134.765 ;
        RECT 108.135 134.735 108.415 135.405 ;
        RECT 108.690 135.235 109.140 135.695 ;
        RECT 110.005 135.525 110.405 136.375 ;
        RECT 110.805 136.085 111.075 136.545 ;
        RECT 111.245 135.915 111.530 136.375 ;
        RECT 108.585 134.905 109.140 135.235 ;
        RECT 109.310 134.965 110.405 135.525 ;
        RECT 108.690 134.795 109.140 134.905 ;
        RECT 107.675 133.995 107.965 134.720 ;
        RECT 108.135 134.165 108.520 134.735 ;
        RECT 108.690 134.625 109.815 134.795 ;
        RECT 108.690 133.995 109.015 134.455 ;
        RECT 109.535 134.165 109.815 134.625 ;
        RECT 110.005 134.165 110.405 134.965 ;
        RECT 110.575 135.695 111.530 135.915 ;
        RECT 110.575 134.795 110.785 135.695 ;
        RECT 110.955 134.965 111.645 135.525 ;
        RECT 112.735 135.405 113.075 136.375 ;
        RECT 113.245 135.405 113.415 136.545 ;
        RECT 113.685 135.745 113.935 136.545 ;
        RECT 114.580 135.575 114.910 136.375 ;
        RECT 115.210 135.745 115.540 136.545 ;
        RECT 115.710 135.575 116.040 136.375 ;
        RECT 116.505 135.875 116.675 136.375 ;
        RECT 116.845 136.045 117.175 136.545 ;
        RECT 116.505 135.705 117.170 135.875 ;
        RECT 113.605 135.405 116.040 135.575 ;
        RECT 112.735 134.795 112.910 135.405 ;
        RECT 113.605 135.155 113.775 135.405 ;
        RECT 113.080 134.985 113.775 135.155 ;
        RECT 113.950 134.985 114.370 135.185 ;
        RECT 114.540 134.985 114.870 135.185 ;
        RECT 115.040 134.985 115.370 135.185 ;
        RECT 110.575 134.625 111.530 134.795 ;
        RECT 110.805 133.995 111.075 134.455 ;
        RECT 111.245 134.165 111.530 134.625 ;
        RECT 112.735 134.165 113.075 134.795 ;
        RECT 113.245 133.995 113.495 134.795 ;
        RECT 113.685 134.645 114.910 134.815 ;
        RECT 113.685 134.165 114.015 134.645 ;
        RECT 114.185 133.995 114.410 134.455 ;
        RECT 114.580 134.165 114.910 134.645 ;
        RECT 115.540 134.775 115.710 135.405 ;
        RECT 115.895 134.985 116.245 135.235 ;
        RECT 116.420 134.885 116.770 135.535 ;
        RECT 115.540 134.165 116.040 134.775 ;
        RECT 116.940 134.715 117.170 135.705 ;
        RECT 116.505 134.545 117.170 134.715 ;
        RECT 116.505 134.255 116.675 134.545 ;
        RECT 116.845 133.995 117.175 134.375 ;
        RECT 117.345 134.255 117.530 136.375 ;
        RECT 117.770 136.085 118.035 136.545 ;
        RECT 118.205 135.950 118.455 136.375 ;
        RECT 118.665 136.100 119.770 136.270 ;
        RECT 118.150 135.820 118.455 135.950 ;
        RECT 117.700 134.625 117.980 135.575 ;
        RECT 118.150 134.715 118.320 135.820 ;
        RECT 118.490 135.035 118.730 135.630 ;
        RECT 118.900 135.565 119.430 135.930 ;
        RECT 118.900 134.865 119.070 135.565 ;
        RECT 119.600 135.485 119.770 136.100 ;
        RECT 119.940 135.745 120.110 136.545 ;
        RECT 120.280 136.045 120.530 136.375 ;
        RECT 120.755 136.075 121.640 136.245 ;
        RECT 119.600 135.395 120.110 135.485 ;
        RECT 118.150 134.585 118.375 134.715 ;
        RECT 118.545 134.645 119.070 134.865 ;
        RECT 119.240 135.225 120.110 135.395 ;
        RECT 117.785 133.995 118.035 134.455 ;
        RECT 118.205 134.445 118.375 134.585 ;
        RECT 119.240 134.445 119.410 135.225 ;
        RECT 119.940 135.155 120.110 135.225 ;
        RECT 119.620 134.975 119.820 135.005 ;
        RECT 120.280 134.975 120.450 136.045 ;
        RECT 120.620 135.155 120.810 135.875 ;
        RECT 119.620 134.675 120.450 134.975 ;
        RECT 120.980 134.945 121.300 135.905 ;
        RECT 118.205 134.275 118.540 134.445 ;
        RECT 118.735 134.275 119.410 134.445 ;
        RECT 119.730 133.995 120.100 134.495 ;
        RECT 120.280 134.445 120.450 134.675 ;
        RECT 120.835 134.615 121.300 134.945 ;
        RECT 121.470 135.235 121.640 136.075 ;
        RECT 121.820 136.045 122.135 136.545 ;
        RECT 122.365 135.815 122.705 136.375 ;
        RECT 121.810 135.440 122.705 135.815 ;
        RECT 122.875 135.535 123.045 136.545 ;
        RECT 122.515 135.235 122.705 135.440 ;
        RECT 123.215 135.485 123.545 136.330 ;
        RECT 123.960 135.575 124.350 135.750 ;
        RECT 124.835 135.745 125.165 136.545 ;
        RECT 125.335 135.755 125.870 136.375 ;
        RECT 123.215 135.405 123.605 135.485 ;
        RECT 123.960 135.405 125.385 135.575 ;
        RECT 123.390 135.355 123.605 135.405 ;
        RECT 121.470 134.905 122.345 135.235 ;
        RECT 122.515 134.905 123.265 135.235 ;
        RECT 121.470 134.445 121.640 134.905 ;
        RECT 122.515 134.735 122.715 134.905 ;
        RECT 123.435 134.775 123.605 135.355 ;
        RECT 123.380 134.735 123.605 134.775 ;
        RECT 120.280 134.275 120.685 134.445 ;
        RECT 120.855 134.275 121.640 134.445 ;
        RECT 121.915 133.995 122.125 134.525 ;
        RECT 122.385 134.210 122.715 134.735 ;
        RECT 123.225 134.650 123.605 134.735 ;
        RECT 123.835 134.675 124.190 135.235 ;
        RECT 122.885 133.995 123.055 134.605 ;
        RECT 123.225 134.215 123.555 134.650 ;
        RECT 124.360 134.505 124.530 135.405 ;
        RECT 124.700 134.675 124.965 135.235 ;
        RECT 125.215 134.905 125.385 135.405 ;
        RECT 125.555 134.735 125.870 135.755 ;
        RECT 126.075 135.455 127.285 136.545 ;
        RECT 123.940 133.995 124.180 134.505 ;
        RECT 124.360 134.175 124.640 134.505 ;
        RECT 124.870 133.995 125.085 134.505 ;
        RECT 125.255 134.165 125.870 134.735 ;
        RECT 126.075 134.745 126.595 135.285 ;
        RECT 126.765 134.915 127.285 135.455 ;
        RECT 127.640 135.575 128.030 135.750 ;
        RECT 128.515 135.745 128.845 136.545 ;
        RECT 129.015 135.755 129.550 136.375 ;
        RECT 127.640 135.405 129.065 135.575 ;
        RECT 126.075 133.995 127.285 134.745 ;
        RECT 127.515 134.675 127.870 135.235 ;
        RECT 128.040 134.505 128.210 135.405 ;
        RECT 128.380 134.675 128.645 135.235 ;
        RECT 128.895 134.905 129.065 135.405 ;
        RECT 129.235 134.735 129.550 135.755 ;
        RECT 129.960 135.575 130.290 136.375 ;
        RECT 130.460 135.745 130.790 136.545 ;
        RECT 131.090 135.575 131.420 136.375 ;
        RECT 132.065 135.745 132.315 136.545 ;
        RECT 129.960 135.405 132.395 135.575 ;
        RECT 132.585 135.405 132.755 136.545 ;
        RECT 132.925 135.405 133.265 136.375 ;
        RECT 129.755 134.985 130.105 135.235 ;
        RECT 130.290 134.775 130.460 135.405 ;
        RECT 130.630 134.985 130.960 135.185 ;
        RECT 131.130 134.985 131.460 135.185 ;
        RECT 131.630 134.985 132.050 135.185 ;
        RECT 132.225 135.155 132.395 135.405 ;
        RECT 132.225 134.985 132.920 135.155 ;
        RECT 133.090 134.845 133.265 135.405 ;
        RECT 133.435 135.380 133.725 136.545 ;
        RECT 133.985 135.875 134.155 136.375 ;
        RECT 134.325 136.045 134.655 136.545 ;
        RECT 133.985 135.705 134.650 135.875 ;
        RECT 133.900 134.885 134.250 135.535 ;
        RECT 127.620 133.995 127.860 134.505 ;
        RECT 128.040 134.175 128.320 134.505 ;
        RECT 128.550 133.995 128.765 134.505 ;
        RECT 128.935 134.165 129.550 134.735 ;
        RECT 129.960 134.165 130.460 134.775 ;
        RECT 131.090 134.645 132.315 134.815 ;
        RECT 133.035 134.795 133.265 134.845 ;
        RECT 131.090 134.165 131.420 134.645 ;
        RECT 131.590 133.995 131.815 134.455 ;
        RECT 131.985 134.165 132.315 134.645 ;
        RECT 132.505 133.995 132.755 134.795 ;
        RECT 132.925 134.165 133.265 134.795 ;
        RECT 133.435 133.995 133.725 134.720 ;
        RECT 134.420 134.715 134.650 135.705 ;
        RECT 133.985 134.545 134.650 134.715 ;
        RECT 133.985 134.255 134.155 134.545 ;
        RECT 134.325 133.995 134.655 134.375 ;
        RECT 134.825 134.255 135.010 136.375 ;
        RECT 135.250 136.085 135.515 136.545 ;
        RECT 135.685 135.950 135.935 136.375 ;
        RECT 136.145 136.100 137.250 136.270 ;
        RECT 135.630 135.820 135.935 135.950 ;
        RECT 135.180 134.625 135.460 135.575 ;
        RECT 135.630 134.715 135.800 135.820 ;
        RECT 135.970 135.035 136.210 135.630 ;
        RECT 136.380 135.565 136.910 135.930 ;
        RECT 136.380 134.865 136.550 135.565 ;
        RECT 137.080 135.485 137.250 136.100 ;
        RECT 137.420 135.745 137.590 136.545 ;
        RECT 137.760 136.045 138.010 136.375 ;
        RECT 138.235 136.075 139.120 136.245 ;
        RECT 137.080 135.395 137.590 135.485 ;
        RECT 135.630 134.585 135.855 134.715 ;
        RECT 136.025 134.645 136.550 134.865 ;
        RECT 136.720 135.225 137.590 135.395 ;
        RECT 135.265 133.995 135.515 134.455 ;
        RECT 135.685 134.445 135.855 134.585 ;
        RECT 136.720 134.445 136.890 135.225 ;
        RECT 137.420 135.155 137.590 135.225 ;
        RECT 137.100 134.975 137.300 135.005 ;
        RECT 137.760 134.975 137.930 136.045 ;
        RECT 138.100 135.155 138.290 135.875 ;
        RECT 137.100 134.675 137.930 134.975 ;
        RECT 138.460 134.945 138.780 135.905 ;
        RECT 135.685 134.275 136.020 134.445 ;
        RECT 136.215 134.275 136.890 134.445 ;
        RECT 137.210 133.995 137.580 134.495 ;
        RECT 137.760 134.445 137.930 134.675 ;
        RECT 138.315 134.615 138.780 134.945 ;
        RECT 138.950 135.235 139.120 136.075 ;
        RECT 139.300 136.045 139.615 136.545 ;
        RECT 139.845 135.815 140.185 136.375 ;
        RECT 139.290 135.440 140.185 135.815 ;
        RECT 140.355 135.535 140.525 136.545 ;
        RECT 139.995 135.235 140.185 135.440 ;
        RECT 140.695 135.485 141.025 136.330 ;
        RECT 140.695 135.405 141.085 135.485 ;
        RECT 140.870 135.355 141.085 135.405 ;
        RECT 138.950 134.905 139.825 135.235 ;
        RECT 139.995 134.905 140.745 135.235 ;
        RECT 138.950 134.445 139.120 134.905 ;
        RECT 139.995 134.735 140.195 134.905 ;
        RECT 140.915 134.775 141.085 135.355 ;
        RECT 141.715 135.455 142.925 136.545 ;
        RECT 141.715 134.915 142.235 135.455 ;
        RECT 140.860 134.735 141.085 134.775 ;
        RECT 142.405 134.745 142.925 135.285 ;
        RECT 137.760 134.275 138.165 134.445 ;
        RECT 138.335 134.275 139.120 134.445 ;
        RECT 139.395 133.995 139.605 134.525 ;
        RECT 139.865 134.210 140.195 134.735 ;
        RECT 140.705 134.650 141.085 134.735 ;
        RECT 140.365 133.995 140.535 134.605 ;
        RECT 140.705 134.215 141.035 134.650 ;
        RECT 141.715 133.995 142.925 134.745 ;
        RECT 17.430 133.825 143.010 133.995 ;
        RECT 17.515 133.075 18.725 133.825 ;
        RECT 18.895 133.280 24.240 133.825 ;
        RECT 17.515 132.535 18.035 133.075 ;
        RECT 18.205 132.365 18.725 132.905 ;
        RECT 20.480 132.450 20.820 133.280 ;
        RECT 24.415 133.055 26.085 133.825 ;
        RECT 17.515 131.275 18.725 132.365 ;
        RECT 22.300 131.710 22.650 132.960 ;
        RECT 24.415 132.535 25.165 133.055 ;
        RECT 26.265 133.015 26.535 133.825 ;
        RECT 26.705 133.015 27.035 133.655 ;
        RECT 27.205 133.015 27.445 133.825 ;
        RECT 27.635 133.280 32.980 133.825 ;
        RECT 25.335 132.365 26.085 132.885 ;
        RECT 26.255 132.585 26.605 132.835 ;
        RECT 26.775 132.415 26.945 133.015 ;
        RECT 27.115 132.585 27.465 132.835 ;
        RECT 29.220 132.450 29.560 133.280 ;
        RECT 33.155 133.055 36.665 133.825 ;
        RECT 37.385 133.485 37.555 133.520 ;
        RECT 37.355 133.315 37.555 133.485 ;
        RECT 18.895 131.275 24.240 131.710 ;
        RECT 24.415 131.275 26.085 132.365 ;
        RECT 26.265 131.275 26.595 132.415 ;
        RECT 26.775 132.245 27.455 132.415 ;
        RECT 27.125 131.460 27.455 132.245 ;
        RECT 31.040 131.710 31.390 132.960 ;
        RECT 33.155 132.535 34.805 133.055 ;
        RECT 37.385 132.955 37.555 133.315 ;
        RECT 37.745 133.295 37.975 133.600 ;
        RECT 38.145 133.465 38.475 133.825 ;
        RECT 38.670 133.295 38.960 133.645 ;
        RECT 37.745 133.125 38.960 133.295 ;
        RECT 39.145 133.095 39.445 133.825 ;
        RECT 34.975 132.365 36.665 132.885 ;
        RECT 37.385 132.785 37.905 132.955 ;
        RECT 39.625 132.915 39.855 133.535 ;
        RECT 40.055 133.265 40.280 133.645 ;
        RECT 40.450 133.435 40.780 133.825 ;
        RECT 40.055 133.085 40.385 133.265 ;
        RECT 27.635 131.275 32.980 131.710 ;
        RECT 33.155 131.275 36.665 132.365 ;
        RECT 37.300 132.255 37.545 132.615 ;
        RECT 37.735 132.405 37.905 132.785 ;
        RECT 38.075 132.585 38.460 132.915 ;
        RECT 38.640 132.805 38.900 132.915 ;
        RECT 38.640 132.635 38.905 132.805 ;
        RECT 38.640 132.585 38.900 132.635 ;
        RECT 39.150 132.585 39.445 132.915 ;
        RECT 39.625 132.585 40.040 132.915 ;
        RECT 37.735 132.125 38.085 132.405 ;
        RECT 37.300 131.275 37.555 132.075 ;
        RECT 37.755 131.445 38.085 132.125 ;
        RECT 38.265 131.535 38.460 132.585 ;
        RECT 40.210 132.415 40.385 133.085 ;
        RECT 40.555 132.585 40.795 133.235 ;
        RECT 40.975 133.055 42.645 133.825 ;
        RECT 43.275 133.100 43.565 133.825 ;
        RECT 43.735 133.280 49.080 133.825 ;
        RECT 50.340 133.315 50.580 133.825 ;
        RECT 50.760 133.315 51.040 133.645 ;
        RECT 51.270 133.315 51.485 133.825 ;
        RECT 40.975 132.535 41.725 133.055 ;
        RECT 38.640 131.275 38.960 132.415 ;
        RECT 39.145 132.055 40.040 132.385 ;
        RECT 40.210 132.225 40.795 132.415 ;
        RECT 41.895 132.365 42.645 132.885 ;
        RECT 45.320 132.450 45.660 133.280 ;
        RECT 39.145 131.885 40.350 132.055 ;
        RECT 39.145 131.455 39.475 131.885 ;
        RECT 39.655 131.275 39.850 131.715 ;
        RECT 40.020 131.455 40.350 131.885 ;
        RECT 40.520 131.455 40.795 132.225 ;
        RECT 40.975 131.275 42.645 132.365 ;
        RECT 43.275 131.275 43.565 132.440 ;
        RECT 47.140 131.710 47.490 132.960 ;
        RECT 50.235 132.585 50.590 133.145 ;
        RECT 50.760 132.415 50.930 133.315 ;
        RECT 51.100 132.585 51.365 133.145 ;
        RECT 51.655 133.085 52.270 133.655 ;
        RECT 51.615 132.415 51.785 132.915 ;
        RECT 50.360 132.245 51.785 132.415 ;
        RECT 50.360 132.070 50.750 132.245 ;
        RECT 43.735 131.275 49.080 131.710 ;
        RECT 51.235 131.275 51.565 132.075 ;
        RECT 51.955 132.065 52.270 133.085 ;
        RECT 51.735 131.445 52.270 132.065 ;
        RECT 52.510 133.085 53.125 133.655 ;
        RECT 53.295 133.315 53.510 133.825 ;
        RECT 53.740 133.315 54.020 133.645 ;
        RECT 54.200 133.315 54.440 133.825 ;
        RECT 55.695 133.445 56.585 133.615 ;
        RECT 52.510 132.065 52.825 133.085 ;
        RECT 52.995 132.415 53.165 132.915 ;
        RECT 53.415 132.585 53.680 133.145 ;
        RECT 53.850 132.415 54.020 133.315 ;
        RECT 54.190 132.585 54.545 133.145 ;
        RECT 55.695 132.890 56.245 133.275 ;
        RECT 56.415 132.720 56.585 133.445 ;
        RECT 55.695 132.650 56.585 132.720 ;
        RECT 56.755 133.120 56.975 133.605 ;
        RECT 57.145 133.285 57.395 133.825 ;
        RECT 57.565 133.175 57.825 133.655 ;
        RECT 56.755 132.695 57.085 133.120 ;
        RECT 55.695 132.625 56.590 132.650 ;
        RECT 55.695 132.610 56.600 132.625 ;
        RECT 55.695 132.595 56.605 132.610 ;
        RECT 55.695 132.590 56.615 132.595 ;
        RECT 55.695 132.580 56.620 132.590 ;
        RECT 55.695 132.570 56.625 132.580 ;
        RECT 55.695 132.565 56.635 132.570 ;
        RECT 55.695 132.555 56.645 132.565 ;
        RECT 55.695 132.550 56.655 132.555 ;
        RECT 52.995 132.245 54.420 132.415 ;
        RECT 52.510 131.445 53.045 132.065 ;
        RECT 53.215 131.275 53.545 132.075 ;
        RECT 54.030 132.070 54.420 132.245 ;
        RECT 55.695 132.100 55.955 132.550 ;
        RECT 56.320 132.545 56.655 132.550 ;
        RECT 56.320 132.540 56.670 132.545 ;
        RECT 56.320 132.530 56.685 132.540 ;
        RECT 56.320 132.525 56.710 132.530 ;
        RECT 57.255 132.525 57.485 132.920 ;
        RECT 56.320 132.520 57.485 132.525 ;
        RECT 56.350 132.485 57.485 132.520 ;
        RECT 56.385 132.460 57.485 132.485 ;
        RECT 56.415 132.430 57.485 132.460 ;
        RECT 56.435 132.400 57.485 132.430 ;
        RECT 56.455 132.370 57.485 132.400 ;
        RECT 56.525 132.360 57.485 132.370 ;
        RECT 56.550 132.350 57.485 132.360 ;
        RECT 56.570 132.335 57.485 132.350 ;
        RECT 56.590 132.320 57.485 132.335 ;
        RECT 56.595 132.310 57.380 132.320 ;
        RECT 56.610 132.275 57.380 132.310 ;
        RECT 56.125 131.955 56.455 132.200 ;
        RECT 56.625 132.025 57.380 132.275 ;
        RECT 57.655 132.145 57.825 133.175 ;
        RECT 58.045 133.170 58.375 133.605 ;
        RECT 58.545 133.215 58.715 133.825 ;
        RECT 57.995 133.085 58.375 133.170 ;
        RECT 58.885 133.085 59.215 133.610 ;
        RECT 59.475 133.295 59.685 133.825 ;
        RECT 59.960 133.375 60.745 133.545 ;
        RECT 60.915 133.375 61.320 133.545 ;
        RECT 57.995 133.045 58.220 133.085 ;
        RECT 57.995 132.465 58.165 133.045 ;
        RECT 58.885 132.915 59.085 133.085 ;
        RECT 59.960 132.915 60.130 133.375 ;
        RECT 58.335 132.585 59.085 132.915 ;
        RECT 59.255 132.585 60.130 132.915 ;
        RECT 57.995 132.415 58.210 132.465 ;
        RECT 57.995 132.335 58.385 132.415 ;
        RECT 56.125 131.930 56.310 131.955 ;
        RECT 55.695 131.830 56.310 131.930 ;
        RECT 55.695 131.275 56.300 131.830 ;
        RECT 56.475 131.445 56.955 131.785 ;
        RECT 57.125 131.275 57.380 131.820 ;
        RECT 57.550 131.445 57.825 132.145 ;
        RECT 58.055 131.490 58.385 132.335 ;
        RECT 58.895 132.380 59.085 132.585 ;
        RECT 58.555 131.275 58.725 132.285 ;
        RECT 58.895 132.005 59.790 132.380 ;
        RECT 58.895 131.445 59.235 132.005 ;
        RECT 59.465 131.275 59.780 131.775 ;
        RECT 59.960 131.745 60.130 132.585 ;
        RECT 60.300 132.875 60.765 133.205 ;
        RECT 61.150 133.145 61.320 133.375 ;
        RECT 61.500 133.325 61.870 133.825 ;
        RECT 62.190 133.375 62.865 133.545 ;
        RECT 63.060 133.375 63.395 133.545 ;
        RECT 60.300 131.915 60.620 132.875 ;
        RECT 61.150 132.845 61.980 133.145 ;
        RECT 60.790 131.945 60.980 132.665 ;
        RECT 61.150 131.775 61.320 132.845 ;
        RECT 61.780 132.815 61.980 132.845 ;
        RECT 61.490 132.595 61.660 132.665 ;
        RECT 62.190 132.595 62.360 133.375 ;
        RECT 63.225 133.235 63.395 133.375 ;
        RECT 63.565 133.365 63.815 133.825 ;
        RECT 61.490 132.425 62.360 132.595 ;
        RECT 62.530 132.955 63.055 133.175 ;
        RECT 63.225 133.105 63.450 133.235 ;
        RECT 61.490 132.335 62.000 132.425 ;
        RECT 59.960 131.575 60.845 131.745 ;
        RECT 61.070 131.445 61.320 131.775 ;
        RECT 61.490 131.275 61.660 132.075 ;
        RECT 61.830 131.720 62.000 132.335 ;
        RECT 62.530 132.255 62.700 132.955 ;
        RECT 62.170 131.890 62.700 132.255 ;
        RECT 62.870 132.190 63.110 132.785 ;
        RECT 63.280 132.000 63.450 133.105 ;
        RECT 63.620 132.245 63.900 133.195 ;
        RECT 63.145 131.870 63.450 132.000 ;
        RECT 61.830 131.550 62.935 131.720 ;
        RECT 63.145 131.445 63.395 131.870 ;
        RECT 63.565 131.275 63.830 131.735 ;
        RECT 64.070 131.445 64.255 133.565 ;
        RECT 64.425 133.445 64.755 133.825 ;
        RECT 64.925 133.275 65.095 133.565 ;
        RECT 64.430 133.105 65.095 133.275 ;
        RECT 64.430 132.115 64.660 133.105 ;
        RECT 65.355 133.055 68.865 133.825 ;
        RECT 69.035 133.100 69.325 133.825 ;
        RECT 70.505 133.275 70.675 133.565 ;
        RECT 70.845 133.445 71.175 133.825 ;
        RECT 70.505 133.105 71.170 133.275 ;
        RECT 64.830 132.285 65.180 132.935 ;
        RECT 65.355 132.535 67.005 133.055 ;
        RECT 67.175 132.365 68.865 132.885 ;
        RECT 64.430 131.945 65.095 132.115 ;
        RECT 64.425 131.275 64.755 131.775 ;
        RECT 64.925 131.445 65.095 131.945 ;
        RECT 65.355 131.275 68.865 132.365 ;
        RECT 69.035 131.275 69.325 132.440 ;
        RECT 70.420 132.285 70.770 132.935 ;
        RECT 70.940 132.115 71.170 133.105 ;
        RECT 70.505 131.945 71.170 132.115 ;
        RECT 70.505 131.445 70.675 131.945 ;
        RECT 70.845 131.275 71.175 131.775 ;
        RECT 71.345 131.445 71.530 133.565 ;
        RECT 71.785 133.365 72.035 133.825 ;
        RECT 72.205 133.375 72.540 133.545 ;
        RECT 72.735 133.375 73.410 133.545 ;
        RECT 72.205 133.235 72.375 133.375 ;
        RECT 71.700 132.245 71.980 133.195 ;
        RECT 72.150 133.105 72.375 133.235 ;
        RECT 72.150 132.000 72.320 133.105 ;
        RECT 72.545 132.955 73.070 133.175 ;
        RECT 72.490 132.190 72.730 132.785 ;
        RECT 72.900 132.255 73.070 132.955 ;
        RECT 73.240 132.595 73.410 133.375 ;
        RECT 73.730 133.325 74.100 133.825 ;
        RECT 74.280 133.375 74.685 133.545 ;
        RECT 74.855 133.375 75.640 133.545 ;
        RECT 74.280 133.145 74.450 133.375 ;
        RECT 73.620 132.845 74.450 133.145 ;
        RECT 74.835 132.875 75.300 133.205 ;
        RECT 73.620 132.815 73.820 132.845 ;
        RECT 73.940 132.595 74.110 132.665 ;
        RECT 73.240 132.425 74.110 132.595 ;
        RECT 73.600 132.335 74.110 132.425 ;
        RECT 72.150 131.870 72.455 132.000 ;
        RECT 72.900 131.890 73.430 132.255 ;
        RECT 71.770 131.275 72.035 131.735 ;
        RECT 72.205 131.445 72.455 131.870 ;
        RECT 73.600 131.720 73.770 132.335 ;
        RECT 72.665 131.550 73.770 131.720 ;
        RECT 73.940 131.275 74.110 132.075 ;
        RECT 74.280 131.775 74.450 132.845 ;
        RECT 74.620 131.945 74.810 132.665 ;
        RECT 74.980 131.915 75.300 132.875 ;
        RECT 75.470 132.915 75.640 133.375 ;
        RECT 75.915 133.295 76.125 133.825 ;
        RECT 76.385 133.085 76.715 133.610 ;
        RECT 76.885 133.215 77.055 133.825 ;
        RECT 77.225 133.170 77.555 133.605 ;
        RECT 77.775 133.280 83.120 133.825 ;
        RECT 83.295 133.280 88.640 133.825 ;
        RECT 88.815 133.280 94.160 133.825 ;
        RECT 77.225 133.085 77.605 133.170 ;
        RECT 76.515 132.915 76.715 133.085 ;
        RECT 77.380 133.045 77.605 133.085 ;
        RECT 75.470 132.585 76.345 132.915 ;
        RECT 76.515 132.585 77.265 132.915 ;
        RECT 74.280 131.445 74.530 131.775 ;
        RECT 75.470 131.745 75.640 132.585 ;
        RECT 76.515 132.380 76.705 132.585 ;
        RECT 77.435 132.465 77.605 133.045 ;
        RECT 77.390 132.415 77.605 132.465 ;
        RECT 79.360 132.450 79.700 133.280 ;
        RECT 75.810 132.005 76.705 132.380 ;
        RECT 77.215 132.335 77.605 132.415 ;
        RECT 74.755 131.575 75.640 131.745 ;
        RECT 75.820 131.275 76.135 131.775 ;
        RECT 76.365 131.445 76.705 132.005 ;
        RECT 76.875 131.275 77.045 132.285 ;
        RECT 77.215 131.490 77.545 132.335 ;
        RECT 81.180 131.710 81.530 132.960 ;
        RECT 84.880 132.450 85.220 133.280 ;
        RECT 86.700 131.710 87.050 132.960 ;
        RECT 90.400 132.450 90.740 133.280 ;
        RECT 94.795 133.100 95.085 133.825 ;
        RECT 95.255 133.280 100.600 133.825 ;
        RECT 92.220 131.710 92.570 132.960 ;
        RECT 96.840 132.450 97.180 133.280 ;
        RECT 101.240 133.085 101.495 133.655 ;
        RECT 101.665 133.425 101.995 133.825 ;
        RECT 102.420 133.290 102.950 133.655 ;
        RECT 103.140 133.485 103.415 133.655 ;
        RECT 103.135 133.315 103.415 133.485 ;
        RECT 102.420 133.255 102.595 133.290 ;
        RECT 101.665 133.085 102.595 133.255 ;
        RECT 77.775 131.275 83.120 131.710 ;
        RECT 83.295 131.275 88.640 131.710 ;
        RECT 88.815 131.275 94.160 131.710 ;
        RECT 94.795 131.275 95.085 132.440 ;
        RECT 98.660 131.710 99.010 132.960 ;
        RECT 101.240 132.415 101.410 133.085 ;
        RECT 101.665 132.915 101.835 133.085 ;
        RECT 101.580 132.585 101.835 132.915 ;
        RECT 102.060 132.585 102.255 132.915 ;
        RECT 95.255 131.275 100.600 131.710 ;
        RECT 101.240 131.445 101.575 132.415 ;
        RECT 101.745 131.275 101.915 132.415 ;
        RECT 102.085 131.615 102.255 132.585 ;
        RECT 102.425 131.955 102.595 133.085 ;
        RECT 102.765 132.295 102.935 133.095 ;
        RECT 103.140 132.495 103.415 133.315 ;
        RECT 103.585 132.295 103.775 133.655 ;
        RECT 103.955 133.290 104.465 133.825 ;
        RECT 104.685 133.015 104.930 133.620 ;
        RECT 105.375 133.055 108.885 133.825 ;
        RECT 103.975 132.845 105.205 133.015 ;
        RECT 102.765 132.125 103.775 132.295 ;
        RECT 103.945 132.280 104.695 132.470 ;
        RECT 102.425 131.785 103.550 131.955 ;
        RECT 103.945 131.615 104.115 132.280 ;
        RECT 104.865 132.035 105.205 132.845 ;
        RECT 105.375 132.535 107.025 133.055 ;
        RECT 107.195 132.365 108.885 132.885 ;
        RECT 102.085 131.445 104.115 131.615 ;
        RECT 104.285 131.275 104.455 132.035 ;
        RECT 104.690 131.625 105.205 132.035 ;
        RECT 105.375 131.275 108.885 132.365 ;
        RECT 109.520 132.225 109.855 133.645 ;
        RECT 110.035 133.455 110.780 133.825 ;
        RECT 111.345 133.285 111.600 133.645 ;
        RECT 111.780 133.455 112.110 133.825 ;
        RECT 112.290 133.285 112.515 133.645 ;
        RECT 110.030 133.095 112.515 133.285 ;
        RECT 110.030 132.405 110.255 133.095 ;
        RECT 112.735 133.055 114.405 133.825 ;
        RECT 110.455 132.585 110.735 132.915 ;
        RECT 110.915 132.585 111.490 132.915 ;
        RECT 111.670 132.585 112.105 132.915 ;
        RECT 112.285 132.585 112.555 132.915 ;
        RECT 112.735 132.535 113.485 133.055 ;
        RECT 114.780 133.045 115.280 133.655 ;
        RECT 110.030 132.225 112.525 132.405 ;
        RECT 113.655 132.365 114.405 132.885 ;
        RECT 114.575 132.585 114.925 132.835 ;
        RECT 115.110 132.415 115.280 133.045 ;
        RECT 115.910 133.175 116.240 133.655 ;
        RECT 116.410 133.365 116.635 133.825 ;
        RECT 116.805 133.175 117.135 133.655 ;
        RECT 115.910 133.005 117.135 133.175 ;
        RECT 117.325 133.025 117.575 133.825 ;
        RECT 117.745 133.025 118.085 133.655 ;
        RECT 115.450 132.635 115.780 132.835 ;
        RECT 115.950 132.635 116.280 132.835 ;
        RECT 116.450 132.635 116.870 132.835 ;
        RECT 117.045 132.665 117.740 132.835 ;
        RECT 117.045 132.415 117.215 132.665 ;
        RECT 117.910 132.415 118.085 133.025 ;
        RECT 109.520 131.455 109.785 132.225 ;
        RECT 109.955 131.275 110.285 131.995 ;
        RECT 110.475 131.815 111.665 132.045 ;
        RECT 110.475 131.455 110.735 131.815 ;
        RECT 110.905 131.275 111.235 131.645 ;
        RECT 111.405 131.455 111.665 131.815 ;
        RECT 112.235 131.455 112.525 132.225 ;
        RECT 112.735 131.275 114.405 132.365 ;
        RECT 114.780 132.245 117.215 132.415 ;
        RECT 114.780 131.445 115.110 132.245 ;
        RECT 115.280 131.275 115.610 132.075 ;
        RECT 115.910 131.445 116.240 132.245 ;
        RECT 116.885 131.275 117.135 132.075 ;
        RECT 117.405 131.275 117.575 132.415 ;
        RECT 117.745 131.445 118.085 132.415 ;
        RECT 118.290 133.085 118.905 133.655 ;
        RECT 119.075 133.315 119.290 133.825 ;
        RECT 119.520 133.315 119.800 133.645 ;
        RECT 119.980 133.315 120.220 133.825 ;
        RECT 118.290 132.065 118.605 133.085 ;
        RECT 118.775 132.415 118.945 132.915 ;
        RECT 119.195 132.585 119.460 133.145 ;
        RECT 119.630 132.415 119.800 133.315 ;
        RECT 119.970 132.585 120.325 133.145 ;
        RECT 120.555 133.100 120.845 133.825 ;
        RECT 121.015 133.280 126.360 133.825 ;
        RECT 122.600 132.450 122.940 133.280 ;
        RECT 126.535 133.055 128.205 133.825 ;
        RECT 128.835 133.325 129.095 133.655 ;
        RECT 129.265 133.465 129.595 133.825 ;
        RECT 129.850 133.445 131.150 133.655 ;
        RECT 118.775 132.245 120.200 132.415 ;
        RECT 118.290 131.445 118.825 132.065 ;
        RECT 118.995 131.275 119.325 132.075 ;
        RECT 119.810 132.070 120.200 132.245 ;
        RECT 120.555 131.275 120.845 132.440 ;
        RECT 124.420 131.710 124.770 132.960 ;
        RECT 126.535 132.535 127.285 133.055 ;
        RECT 127.455 132.365 128.205 132.885 ;
        RECT 121.015 131.275 126.360 131.710 ;
        RECT 126.535 131.275 128.205 132.365 ;
        RECT 128.835 132.125 129.005 133.325 ;
        RECT 129.850 133.295 130.020 133.445 ;
        RECT 129.265 133.170 130.020 133.295 ;
        RECT 129.175 133.125 130.020 133.170 ;
        RECT 129.175 133.005 129.445 133.125 ;
        RECT 129.175 132.430 129.345 133.005 ;
        RECT 129.575 132.565 129.985 132.870 ;
        RECT 130.275 132.835 130.485 133.235 ;
        RECT 130.155 132.625 130.485 132.835 ;
        RECT 130.730 132.835 130.950 133.235 ;
        RECT 131.425 133.060 131.880 133.825 ;
        RECT 132.145 133.275 132.315 133.565 ;
        RECT 132.485 133.445 132.815 133.825 ;
        RECT 132.145 133.105 132.810 133.275 ;
        RECT 130.730 132.625 131.205 132.835 ;
        RECT 131.395 132.635 131.885 132.835 ;
        RECT 129.175 132.395 129.375 132.430 ;
        RECT 130.705 132.395 131.880 132.455 ;
        RECT 129.175 132.285 131.880 132.395 ;
        RECT 132.060 132.285 132.410 132.935 ;
        RECT 129.235 132.225 131.035 132.285 ;
        RECT 130.705 132.195 131.035 132.225 ;
        RECT 128.835 131.445 129.095 132.125 ;
        RECT 129.265 131.275 129.515 132.055 ;
        RECT 129.765 132.025 130.600 132.035 ;
        RECT 131.190 132.025 131.375 132.115 ;
        RECT 129.765 131.825 131.375 132.025 ;
        RECT 129.765 131.445 130.015 131.825 ;
        RECT 131.145 131.785 131.375 131.825 ;
        RECT 131.625 131.665 131.880 132.285 ;
        RECT 132.580 132.115 132.810 133.105 ;
        RECT 130.185 131.275 130.540 131.655 ;
        RECT 131.545 131.445 131.880 131.665 ;
        RECT 132.145 131.945 132.810 132.115 ;
        RECT 132.145 131.445 132.315 131.945 ;
        RECT 132.485 131.275 132.815 131.775 ;
        RECT 132.985 131.445 133.170 133.565 ;
        RECT 133.425 133.365 133.675 133.825 ;
        RECT 133.845 133.375 134.180 133.545 ;
        RECT 134.375 133.375 135.050 133.545 ;
        RECT 133.845 133.235 134.015 133.375 ;
        RECT 133.340 132.245 133.620 133.195 ;
        RECT 133.790 133.105 134.015 133.235 ;
        RECT 133.790 132.000 133.960 133.105 ;
        RECT 134.185 132.955 134.710 133.175 ;
        RECT 134.130 132.190 134.370 132.785 ;
        RECT 134.540 132.255 134.710 132.955 ;
        RECT 134.880 132.595 135.050 133.375 ;
        RECT 135.370 133.325 135.740 133.825 ;
        RECT 135.920 133.375 136.325 133.545 ;
        RECT 136.495 133.375 137.280 133.545 ;
        RECT 135.920 133.145 136.090 133.375 ;
        RECT 135.260 132.845 136.090 133.145 ;
        RECT 136.475 132.875 136.940 133.205 ;
        RECT 135.260 132.815 135.460 132.845 ;
        RECT 135.580 132.595 135.750 132.665 ;
        RECT 134.880 132.425 135.750 132.595 ;
        RECT 135.240 132.335 135.750 132.425 ;
        RECT 133.790 131.870 134.095 132.000 ;
        RECT 134.540 131.890 135.070 132.255 ;
        RECT 133.410 131.275 133.675 131.735 ;
        RECT 133.845 131.445 134.095 131.870 ;
        RECT 135.240 131.720 135.410 132.335 ;
        RECT 134.305 131.550 135.410 131.720 ;
        RECT 135.580 131.275 135.750 132.075 ;
        RECT 135.920 131.775 136.090 132.845 ;
        RECT 136.260 131.945 136.450 132.665 ;
        RECT 136.620 131.915 136.940 132.875 ;
        RECT 137.110 132.915 137.280 133.375 ;
        RECT 137.555 133.295 137.765 133.825 ;
        RECT 138.025 133.085 138.355 133.610 ;
        RECT 138.525 133.215 138.695 133.825 ;
        RECT 138.865 133.170 139.195 133.605 ;
        RECT 139.965 133.275 140.135 133.655 ;
        RECT 140.350 133.445 140.680 133.825 ;
        RECT 138.865 133.085 139.245 133.170 ;
        RECT 139.965 133.105 140.680 133.275 ;
        RECT 138.155 132.915 138.355 133.085 ;
        RECT 139.020 133.045 139.245 133.085 ;
        RECT 137.110 132.585 137.985 132.915 ;
        RECT 138.155 132.585 138.905 132.915 ;
        RECT 135.920 131.445 136.170 131.775 ;
        RECT 137.110 131.745 137.280 132.585 ;
        RECT 138.155 132.380 138.345 132.585 ;
        RECT 139.075 132.465 139.245 133.045 ;
        RECT 139.875 132.555 140.230 132.925 ;
        RECT 140.510 132.915 140.680 133.105 ;
        RECT 140.850 133.080 141.105 133.655 ;
        RECT 140.510 132.585 140.765 132.915 ;
        RECT 139.030 132.415 139.245 132.465 ;
        RECT 137.450 132.005 138.345 132.380 ;
        RECT 138.855 132.335 139.245 132.415 ;
        RECT 140.510 132.375 140.680 132.585 ;
        RECT 136.395 131.575 137.280 131.745 ;
        RECT 137.460 131.275 137.775 131.775 ;
        RECT 138.005 131.445 138.345 132.005 ;
        RECT 138.515 131.275 138.685 132.285 ;
        RECT 138.855 131.490 139.185 132.335 ;
        RECT 139.965 132.205 140.680 132.375 ;
        RECT 140.935 132.350 141.105 133.080 ;
        RECT 141.280 132.985 141.540 133.825 ;
        RECT 141.715 133.075 142.925 133.825 ;
        RECT 139.965 131.445 140.135 132.205 ;
        RECT 140.350 131.275 140.680 132.035 ;
        RECT 140.850 131.445 141.105 132.350 ;
        RECT 141.280 131.275 141.540 132.425 ;
        RECT 141.715 132.365 142.235 132.905 ;
        RECT 142.405 132.535 142.925 133.075 ;
        RECT 141.715 131.275 142.925 132.365 ;
        RECT 17.430 131.105 143.010 131.275 ;
        RECT 17.515 130.015 18.725 131.105 ;
        RECT 18.895 130.015 22.405 131.105 ;
        RECT 17.515 129.305 18.035 129.845 ;
        RECT 18.205 129.475 18.725 130.015 ;
        RECT 18.895 129.325 20.545 129.845 ;
        RECT 20.715 129.495 22.405 130.015 ;
        RECT 22.575 130.675 22.915 130.935 ;
        RECT 17.515 128.555 18.725 129.305 ;
        RECT 18.895 128.555 22.405 129.325 ;
        RECT 22.575 129.275 22.835 130.675 ;
        RECT 23.085 130.305 23.415 131.105 ;
        RECT 23.880 130.135 24.130 130.935 ;
        RECT 24.315 130.385 24.645 131.105 ;
        RECT 24.865 130.135 25.115 130.935 ;
        RECT 25.285 130.725 25.620 131.105 ;
        RECT 23.025 129.965 25.215 130.135 ;
        RECT 23.025 129.795 23.340 129.965 ;
        RECT 23.010 129.545 23.340 129.795 ;
        RECT 22.575 128.765 22.915 129.275 ;
        RECT 23.085 128.555 23.355 129.355 ;
        RECT 23.535 128.825 23.815 129.795 ;
        RECT 23.995 128.825 24.295 129.795 ;
        RECT 24.475 128.830 24.825 129.795 ;
        RECT 25.045 129.055 25.215 129.965 ;
        RECT 25.385 129.235 25.625 130.545 ;
        RECT 25.830 130.315 26.365 130.935 ;
        RECT 25.830 129.295 26.145 130.315 ;
        RECT 26.535 130.305 26.865 131.105 ;
        RECT 27.350 130.135 27.740 130.310 ;
        RECT 26.315 129.965 27.740 130.135 ;
        RECT 28.095 130.235 28.370 130.935 ;
        RECT 28.540 130.560 28.795 131.105 ;
        RECT 28.965 130.595 29.445 130.935 ;
        RECT 29.620 130.550 30.225 131.105 ;
        RECT 29.610 130.450 30.225 130.550 ;
        RECT 29.610 130.425 29.795 130.450 ;
        RECT 26.315 129.465 26.485 129.965 ;
        RECT 25.045 128.725 25.540 129.055 ;
        RECT 25.830 128.725 26.445 129.295 ;
        RECT 26.735 129.235 27.000 129.795 ;
        RECT 27.170 129.065 27.340 129.965 ;
        RECT 27.510 129.235 27.865 129.795 ;
        RECT 28.095 129.205 28.265 130.235 ;
        RECT 28.540 130.105 29.295 130.355 ;
        RECT 29.465 130.180 29.795 130.425 ;
        RECT 28.540 130.070 29.310 130.105 ;
        RECT 28.540 130.060 29.325 130.070 ;
        RECT 28.435 130.045 29.330 130.060 ;
        RECT 28.435 130.030 29.350 130.045 ;
        RECT 28.435 130.020 29.370 130.030 ;
        RECT 28.435 130.010 29.395 130.020 ;
        RECT 28.435 129.980 29.465 130.010 ;
        RECT 28.435 129.950 29.485 129.980 ;
        RECT 28.435 129.920 29.505 129.950 ;
        RECT 28.435 129.895 29.535 129.920 ;
        RECT 28.435 129.860 29.570 129.895 ;
        RECT 28.435 129.855 29.600 129.860 ;
        RECT 28.435 129.460 28.665 129.855 ;
        RECT 29.210 129.850 29.600 129.855 ;
        RECT 29.235 129.840 29.600 129.850 ;
        RECT 29.250 129.835 29.600 129.840 ;
        RECT 29.265 129.830 29.600 129.835 ;
        RECT 29.965 129.830 30.225 130.280 ;
        RECT 30.395 129.940 30.685 131.105 ;
        RECT 30.865 130.135 31.195 130.920 ;
        RECT 30.865 129.965 31.545 130.135 ;
        RECT 31.725 129.965 32.055 131.105 ;
        RECT 32.235 130.670 37.580 131.105 ;
        RECT 29.265 129.825 30.225 129.830 ;
        RECT 29.275 129.815 30.225 129.825 ;
        RECT 29.285 129.810 30.225 129.815 ;
        RECT 29.295 129.800 30.225 129.810 ;
        RECT 29.300 129.790 30.225 129.800 ;
        RECT 29.305 129.785 30.225 129.790 ;
        RECT 29.315 129.770 30.225 129.785 ;
        RECT 29.320 129.755 30.225 129.770 ;
        RECT 29.330 129.730 30.225 129.755 ;
        RECT 28.835 129.260 29.165 129.685 ;
        RECT 26.615 128.555 26.830 129.065 ;
        RECT 27.060 128.735 27.340 129.065 ;
        RECT 27.520 128.555 27.760 129.065 ;
        RECT 28.095 128.725 28.355 129.205 ;
        RECT 28.525 128.555 28.775 129.095 ;
        RECT 28.945 128.775 29.165 129.260 ;
        RECT 29.335 129.660 30.225 129.730 ;
        RECT 29.335 128.935 29.505 129.660 ;
        RECT 30.855 129.545 31.205 129.795 ;
        RECT 29.675 129.105 30.225 129.490 ;
        RECT 31.375 129.365 31.545 129.965 ;
        RECT 31.715 129.545 32.065 129.795 ;
        RECT 29.335 128.765 30.225 128.935 ;
        RECT 30.395 128.555 30.685 129.280 ;
        RECT 30.875 128.555 31.115 129.365 ;
        RECT 31.285 128.725 31.615 129.365 ;
        RECT 31.785 128.555 32.055 129.365 ;
        RECT 33.820 129.100 34.160 129.930 ;
        RECT 35.640 129.420 35.990 130.670 ;
        RECT 37.765 130.155 38.040 130.925 ;
        RECT 38.210 130.495 38.540 130.925 ;
        RECT 38.710 130.665 38.905 131.105 ;
        RECT 39.085 130.495 39.415 130.925 ;
        RECT 39.595 130.670 44.940 131.105 ;
        RECT 45.115 130.670 50.460 131.105 ;
        RECT 38.210 130.325 39.415 130.495 ;
        RECT 37.765 129.965 38.350 130.155 ;
        RECT 38.520 129.995 39.415 130.325 ;
        RECT 37.765 129.145 38.005 129.795 ;
        RECT 38.175 129.295 38.350 129.965 ;
        RECT 38.520 129.465 38.935 129.795 ;
        RECT 39.115 129.465 39.410 129.795 ;
        RECT 38.175 129.115 38.505 129.295 ;
        RECT 32.235 128.555 37.580 129.100 ;
        RECT 37.780 128.555 38.110 128.945 ;
        RECT 38.280 128.735 38.505 129.115 ;
        RECT 38.705 128.845 38.935 129.465 ;
        RECT 39.115 128.555 39.415 129.285 ;
        RECT 41.180 129.100 41.520 129.930 ;
        RECT 43.000 129.420 43.350 130.670 ;
        RECT 46.700 129.100 47.040 129.930 ;
        RECT 48.520 129.420 48.870 130.670 ;
        RECT 50.635 130.015 53.225 131.105 ;
        RECT 50.635 129.325 51.845 129.845 ;
        RECT 52.015 129.495 53.225 130.015 ;
        RECT 53.405 130.135 53.735 130.920 ;
        RECT 53.405 129.965 54.085 130.135 ;
        RECT 54.265 129.965 54.595 131.105 ;
        RECT 54.785 130.135 55.115 130.920 ;
        RECT 54.785 129.965 55.465 130.135 ;
        RECT 55.645 129.965 55.975 131.105 ;
        RECT 53.395 129.545 53.745 129.795 ;
        RECT 53.915 129.365 54.085 129.965 ;
        RECT 54.255 129.545 54.605 129.795 ;
        RECT 54.775 129.545 55.125 129.795 ;
        RECT 55.295 129.365 55.465 129.965 ;
        RECT 56.155 129.940 56.445 131.105 ;
        RECT 56.615 130.005 56.935 130.935 ;
        RECT 57.115 130.425 57.515 130.935 ;
        RECT 57.685 130.595 57.855 131.105 ;
        RECT 58.025 130.425 58.355 130.935 ;
        RECT 57.115 130.255 58.355 130.425 ;
        RECT 58.525 130.255 58.695 131.105 ;
        RECT 59.285 130.255 59.665 130.935 ;
        RECT 59.835 130.670 65.180 131.105 ;
        RECT 56.615 129.835 57.245 130.005 ;
        RECT 55.635 129.545 55.985 129.795 ;
        RECT 39.595 128.555 44.940 129.100 ;
        RECT 45.115 128.555 50.460 129.100 ;
        RECT 50.635 128.555 53.225 129.325 ;
        RECT 53.415 128.555 53.655 129.365 ;
        RECT 53.825 128.725 54.155 129.365 ;
        RECT 54.325 128.555 54.595 129.365 ;
        RECT 54.795 128.555 55.035 129.365 ;
        RECT 55.205 128.725 55.535 129.365 ;
        RECT 55.705 128.555 55.975 129.365 ;
        RECT 56.155 128.555 56.445 129.280 ;
        RECT 56.615 128.555 56.905 129.390 ;
        RECT 57.075 128.955 57.245 129.835 ;
        RECT 58.020 129.915 59.325 130.085 ;
        RECT 57.415 129.295 57.645 129.795 ;
        RECT 58.020 129.715 58.190 129.915 ;
        RECT 57.815 129.545 58.190 129.715 ;
        RECT 58.360 129.545 58.910 129.745 ;
        RECT 59.080 129.465 59.325 129.915 ;
        RECT 59.495 129.295 59.665 130.255 ;
        RECT 57.415 129.125 59.665 129.295 ;
        RECT 57.075 128.785 58.030 128.955 ;
        RECT 58.445 128.555 58.775 128.945 ;
        RECT 58.945 128.805 59.115 129.125 ;
        RECT 61.420 129.100 61.760 129.930 ;
        RECT 63.240 129.420 63.590 130.670 ;
        RECT 65.355 130.015 67.945 131.105 ;
        RECT 68.665 130.435 68.835 130.935 ;
        RECT 69.005 130.605 69.335 131.105 ;
        RECT 68.665 130.265 69.330 130.435 ;
        RECT 65.355 129.325 66.565 129.845 ;
        RECT 66.735 129.495 67.945 130.015 ;
        RECT 68.580 129.445 68.930 130.095 ;
        RECT 59.285 128.555 59.615 128.945 ;
        RECT 59.835 128.555 65.180 129.100 ;
        RECT 65.355 128.555 67.945 129.325 ;
        RECT 69.100 129.275 69.330 130.265 ;
        RECT 68.665 129.105 69.330 129.275 ;
        RECT 68.665 128.815 68.835 129.105 ;
        RECT 69.005 128.555 69.335 128.935 ;
        RECT 69.505 128.815 69.690 130.935 ;
        RECT 69.930 130.645 70.195 131.105 ;
        RECT 70.365 130.510 70.615 130.935 ;
        RECT 70.825 130.660 71.930 130.830 ;
        RECT 70.310 130.380 70.615 130.510 ;
        RECT 69.860 129.185 70.140 130.135 ;
        RECT 70.310 129.275 70.480 130.380 ;
        RECT 70.650 129.595 70.890 130.190 ;
        RECT 71.060 130.125 71.590 130.490 ;
        RECT 71.060 129.425 71.230 130.125 ;
        RECT 71.760 130.045 71.930 130.660 ;
        RECT 72.100 130.305 72.270 131.105 ;
        RECT 72.440 130.605 72.690 130.935 ;
        RECT 72.915 130.635 73.800 130.805 ;
        RECT 71.760 129.955 72.270 130.045 ;
        RECT 70.310 129.145 70.535 129.275 ;
        RECT 70.705 129.205 71.230 129.425 ;
        RECT 71.400 129.785 72.270 129.955 ;
        RECT 69.945 128.555 70.195 129.015 ;
        RECT 70.365 129.005 70.535 129.145 ;
        RECT 71.400 129.005 71.570 129.785 ;
        RECT 72.100 129.715 72.270 129.785 ;
        RECT 71.780 129.535 71.980 129.565 ;
        RECT 72.440 129.535 72.610 130.605 ;
        RECT 72.780 129.715 72.970 130.435 ;
        RECT 71.780 129.235 72.610 129.535 ;
        RECT 73.140 129.505 73.460 130.465 ;
        RECT 70.365 128.835 70.700 129.005 ;
        RECT 70.895 128.835 71.570 129.005 ;
        RECT 71.890 128.555 72.260 129.055 ;
        RECT 72.440 129.005 72.610 129.235 ;
        RECT 72.995 129.175 73.460 129.505 ;
        RECT 73.630 129.795 73.800 130.635 ;
        RECT 73.980 130.605 74.295 131.105 ;
        RECT 74.525 130.375 74.865 130.935 ;
        RECT 73.970 130.000 74.865 130.375 ;
        RECT 75.035 130.095 75.205 131.105 ;
        RECT 74.675 129.795 74.865 130.000 ;
        RECT 75.375 130.045 75.705 130.890 ;
        RECT 75.875 130.190 76.045 131.105 ;
        RECT 75.375 129.965 75.765 130.045 ;
        RECT 75.550 129.915 75.765 129.965 ;
        RECT 73.630 129.465 74.505 129.795 ;
        RECT 74.675 129.465 75.425 129.795 ;
        RECT 73.630 129.005 73.800 129.465 ;
        RECT 74.675 129.295 74.875 129.465 ;
        RECT 75.595 129.335 75.765 129.915 ;
        RECT 75.540 129.295 75.765 129.335 ;
        RECT 72.440 128.835 72.845 129.005 ;
        RECT 73.015 128.835 73.800 129.005 ;
        RECT 74.075 128.555 74.285 129.085 ;
        RECT 74.545 128.770 74.875 129.295 ;
        RECT 75.385 129.210 75.765 129.295 ;
        RECT 76.400 129.965 76.735 130.935 ;
        RECT 76.905 129.965 77.075 131.105 ;
        RECT 77.245 130.765 79.275 130.935 ;
        RECT 76.400 129.295 76.570 129.965 ;
        RECT 77.245 129.795 77.415 130.765 ;
        RECT 76.740 129.465 76.995 129.795 ;
        RECT 77.220 129.465 77.415 129.795 ;
        RECT 77.585 130.425 78.710 130.595 ;
        RECT 76.825 129.295 76.995 129.465 ;
        RECT 77.585 129.295 77.755 130.425 ;
        RECT 75.045 128.555 75.215 129.165 ;
        RECT 75.385 128.775 75.715 129.210 ;
        RECT 75.885 128.555 76.055 129.070 ;
        RECT 76.400 128.725 76.655 129.295 ;
        RECT 76.825 129.125 77.755 129.295 ;
        RECT 77.925 130.085 78.935 130.255 ;
        RECT 77.925 129.285 78.095 130.085 ;
        RECT 78.300 129.745 78.575 129.885 ;
        RECT 78.295 129.575 78.575 129.745 ;
        RECT 77.580 129.090 77.755 129.125 ;
        RECT 76.825 128.555 77.155 128.955 ;
        RECT 77.580 128.725 78.110 129.090 ;
        RECT 78.300 128.725 78.575 129.575 ;
        RECT 78.745 128.725 78.935 130.085 ;
        RECT 79.105 130.100 79.275 130.765 ;
        RECT 79.445 130.345 79.615 131.105 ;
        RECT 79.850 130.345 80.365 130.755 ;
        RECT 79.105 129.910 79.855 130.100 ;
        RECT 80.025 129.535 80.365 130.345 ;
        RECT 80.535 130.015 81.745 131.105 ;
        RECT 79.135 129.365 80.365 129.535 ;
        RECT 79.115 128.555 79.625 129.090 ;
        RECT 79.845 128.760 80.090 129.365 ;
        RECT 80.535 129.305 81.055 129.845 ;
        RECT 81.225 129.475 81.745 130.015 ;
        RECT 81.915 129.940 82.205 131.105 ;
        RECT 82.465 130.435 82.635 130.935 ;
        RECT 82.805 130.605 83.135 131.105 ;
        RECT 82.465 130.265 83.130 130.435 ;
        RECT 82.380 129.445 82.730 130.095 ;
        RECT 80.535 128.555 81.745 129.305 ;
        RECT 81.915 128.555 82.205 129.280 ;
        RECT 82.900 129.275 83.130 130.265 ;
        RECT 82.465 129.105 83.130 129.275 ;
        RECT 82.465 128.815 82.635 129.105 ;
        RECT 82.805 128.555 83.135 128.935 ;
        RECT 83.305 128.815 83.490 130.935 ;
        RECT 83.730 130.645 83.995 131.105 ;
        RECT 84.165 130.510 84.415 130.935 ;
        RECT 84.625 130.660 85.730 130.830 ;
        RECT 84.110 130.380 84.415 130.510 ;
        RECT 83.660 129.185 83.940 130.135 ;
        RECT 84.110 129.275 84.280 130.380 ;
        RECT 84.450 129.595 84.690 130.190 ;
        RECT 84.860 130.125 85.390 130.490 ;
        RECT 84.860 129.425 85.030 130.125 ;
        RECT 85.560 130.045 85.730 130.660 ;
        RECT 85.900 130.305 86.070 131.105 ;
        RECT 86.240 130.605 86.490 130.935 ;
        RECT 86.715 130.635 87.600 130.805 ;
        RECT 85.560 129.955 86.070 130.045 ;
        RECT 84.110 129.145 84.335 129.275 ;
        RECT 84.505 129.205 85.030 129.425 ;
        RECT 85.200 129.785 86.070 129.955 ;
        RECT 83.745 128.555 83.995 129.015 ;
        RECT 84.165 129.005 84.335 129.145 ;
        RECT 85.200 129.005 85.370 129.785 ;
        RECT 85.900 129.715 86.070 129.785 ;
        RECT 85.580 129.535 85.780 129.565 ;
        RECT 86.240 129.535 86.410 130.605 ;
        RECT 86.580 129.715 86.770 130.435 ;
        RECT 85.580 129.235 86.410 129.535 ;
        RECT 86.940 129.505 87.260 130.465 ;
        RECT 84.165 128.835 84.500 129.005 ;
        RECT 84.695 128.835 85.370 129.005 ;
        RECT 85.690 128.555 86.060 129.055 ;
        RECT 86.240 129.005 86.410 129.235 ;
        RECT 86.795 129.175 87.260 129.505 ;
        RECT 87.430 129.795 87.600 130.635 ;
        RECT 87.780 130.605 88.095 131.105 ;
        RECT 88.325 130.375 88.665 130.935 ;
        RECT 87.770 130.000 88.665 130.375 ;
        RECT 88.835 130.095 89.005 131.105 ;
        RECT 88.475 129.795 88.665 130.000 ;
        RECT 89.175 130.045 89.505 130.890 ;
        RECT 89.675 130.190 89.845 131.105 ;
        RECT 89.175 129.965 89.565 130.045 ;
        RECT 89.350 129.915 89.565 129.965 ;
        RECT 87.430 129.465 88.305 129.795 ;
        RECT 88.475 129.465 89.225 129.795 ;
        RECT 87.430 129.005 87.600 129.465 ;
        RECT 88.475 129.295 88.675 129.465 ;
        RECT 89.395 129.335 89.565 129.915 ;
        RECT 89.340 129.295 89.565 129.335 ;
        RECT 86.240 128.835 86.645 129.005 ;
        RECT 86.815 128.835 87.600 129.005 ;
        RECT 87.875 128.555 88.085 129.085 ;
        RECT 88.345 128.770 88.675 129.295 ;
        RECT 89.185 129.210 89.565 129.295 ;
        RECT 90.200 129.965 90.535 130.935 ;
        RECT 90.705 129.965 90.875 131.105 ;
        RECT 91.045 130.765 93.075 130.935 ;
        RECT 90.200 129.295 90.370 129.965 ;
        RECT 91.045 129.795 91.215 130.765 ;
        RECT 90.540 129.465 90.795 129.795 ;
        RECT 91.020 129.465 91.215 129.795 ;
        RECT 91.385 130.425 92.510 130.595 ;
        RECT 90.625 129.295 90.795 129.465 ;
        RECT 91.385 129.295 91.555 130.425 ;
        RECT 88.845 128.555 89.015 129.165 ;
        RECT 89.185 128.775 89.515 129.210 ;
        RECT 89.685 128.555 89.855 129.070 ;
        RECT 90.200 128.725 90.455 129.295 ;
        RECT 90.625 129.125 91.555 129.295 ;
        RECT 91.725 130.085 92.735 130.255 ;
        RECT 91.725 129.285 91.895 130.085 ;
        RECT 91.380 129.090 91.555 129.125 ;
        RECT 90.625 128.555 90.955 128.955 ;
        RECT 91.380 128.725 91.910 129.090 ;
        RECT 92.100 129.065 92.375 129.885 ;
        RECT 92.095 128.895 92.375 129.065 ;
        RECT 92.100 128.725 92.375 128.895 ;
        RECT 92.545 128.725 92.735 130.085 ;
        RECT 92.905 130.100 93.075 130.765 ;
        RECT 93.245 130.345 93.415 131.105 ;
        RECT 93.650 130.345 94.165 130.755 ;
        RECT 92.905 129.910 93.655 130.100 ;
        RECT 93.825 129.535 94.165 130.345 ;
        RECT 94.335 130.015 97.845 131.105 ;
        RECT 92.935 129.365 94.165 129.535 ;
        RECT 92.915 128.555 93.425 129.090 ;
        RECT 93.645 128.760 93.890 129.365 ;
        RECT 94.335 129.325 95.985 129.845 ;
        RECT 96.155 129.495 97.845 130.015 ;
        RECT 98.480 129.965 98.815 130.935 ;
        RECT 98.985 129.965 99.155 131.105 ;
        RECT 99.325 130.765 101.355 130.935 ;
        RECT 94.335 128.555 97.845 129.325 ;
        RECT 98.480 129.295 98.650 129.965 ;
        RECT 99.325 129.795 99.495 130.765 ;
        RECT 98.820 129.465 99.075 129.795 ;
        RECT 99.300 129.465 99.495 129.795 ;
        RECT 99.665 130.425 100.790 130.595 ;
        RECT 98.905 129.295 99.075 129.465 ;
        RECT 99.665 129.295 99.835 130.425 ;
        RECT 98.480 128.725 98.735 129.295 ;
        RECT 98.905 129.125 99.835 129.295 ;
        RECT 100.005 130.085 101.015 130.255 ;
        RECT 100.005 129.285 100.175 130.085 ;
        RECT 100.380 129.405 100.655 129.885 ;
        RECT 100.375 129.235 100.655 129.405 ;
        RECT 99.660 129.090 99.835 129.125 ;
        RECT 98.905 128.555 99.235 128.955 ;
        RECT 99.660 128.725 100.190 129.090 ;
        RECT 100.380 128.725 100.655 129.235 ;
        RECT 100.825 128.725 101.015 130.085 ;
        RECT 101.185 130.100 101.355 130.765 ;
        RECT 101.525 130.345 101.695 131.105 ;
        RECT 101.930 130.345 102.445 130.755 ;
        RECT 101.185 129.910 101.935 130.100 ;
        RECT 102.105 129.535 102.445 130.345 ;
        RECT 101.215 129.365 102.445 129.535 ;
        RECT 102.615 129.965 103.000 130.935 ;
        RECT 103.170 130.645 103.495 131.105 ;
        RECT 104.015 130.475 104.295 130.935 ;
        RECT 103.170 130.255 104.295 130.475 ;
        RECT 101.195 128.555 101.705 129.090 ;
        RECT 101.925 128.760 102.170 129.365 ;
        RECT 102.615 129.295 102.895 129.965 ;
        RECT 103.170 129.795 103.620 130.255 ;
        RECT 104.485 130.085 104.885 130.935 ;
        RECT 105.285 130.645 105.555 131.105 ;
        RECT 105.725 130.475 106.010 130.935 ;
        RECT 103.065 129.465 103.620 129.795 ;
        RECT 103.790 129.525 104.885 130.085 ;
        RECT 103.170 129.355 103.620 129.465 ;
        RECT 102.615 128.725 103.000 129.295 ;
        RECT 103.170 129.185 104.295 129.355 ;
        RECT 103.170 128.555 103.495 129.015 ;
        RECT 104.015 128.725 104.295 129.185 ;
        RECT 104.485 128.725 104.885 129.525 ;
        RECT 105.055 130.255 106.010 130.475 ;
        RECT 105.055 129.355 105.265 130.255 ;
        RECT 105.435 129.525 106.125 130.085 ;
        RECT 106.295 130.015 107.505 131.105 ;
        RECT 105.055 129.185 106.010 129.355 ;
        RECT 105.285 128.555 105.555 129.015 ;
        RECT 105.725 128.725 106.010 129.185 ;
        RECT 106.295 129.305 106.815 129.845 ;
        RECT 106.985 129.475 107.505 130.015 ;
        RECT 107.675 129.940 107.965 131.105 ;
        RECT 108.135 130.015 110.725 131.105 ;
        RECT 108.135 129.325 109.345 129.845 ;
        RECT 109.515 129.495 110.725 130.015 ;
        RECT 111.360 130.155 111.625 130.925 ;
        RECT 111.795 130.385 112.125 131.105 ;
        RECT 112.315 130.565 112.575 130.925 ;
        RECT 112.745 130.735 113.075 131.105 ;
        RECT 113.245 130.565 113.505 130.925 ;
        RECT 112.315 130.335 113.505 130.565 ;
        RECT 114.075 130.155 114.365 130.925 ;
        RECT 106.295 128.555 107.505 129.305 ;
        RECT 107.675 128.555 107.965 129.280 ;
        RECT 108.135 128.555 110.725 129.325 ;
        RECT 111.360 128.735 111.695 130.155 ;
        RECT 111.870 129.975 114.365 130.155 ;
        RECT 114.580 130.155 114.845 130.925 ;
        RECT 115.015 130.385 115.345 131.105 ;
        RECT 115.535 130.565 115.795 130.925 ;
        RECT 115.965 130.735 116.295 131.105 ;
        RECT 116.465 130.565 116.725 130.925 ;
        RECT 115.535 130.335 116.725 130.565 ;
        RECT 117.295 130.155 117.585 130.925 ;
        RECT 111.870 129.285 112.095 129.975 ;
        RECT 112.295 129.465 112.575 129.795 ;
        RECT 112.755 129.465 113.330 129.795 ;
        RECT 113.510 129.465 113.945 129.795 ;
        RECT 114.125 129.465 114.395 129.795 ;
        RECT 111.870 129.095 114.355 129.285 ;
        RECT 111.875 128.555 112.620 128.925 ;
        RECT 113.185 128.735 113.440 129.095 ;
        RECT 113.620 128.555 113.950 128.925 ;
        RECT 114.130 128.735 114.355 129.095 ;
        RECT 114.580 128.735 114.915 130.155 ;
        RECT 115.090 129.975 117.585 130.155 ;
        RECT 117.830 130.315 118.365 130.935 ;
        RECT 115.090 129.285 115.315 129.975 ;
        RECT 115.515 129.465 115.795 129.795 ;
        RECT 115.975 129.465 116.550 129.795 ;
        RECT 116.730 129.465 117.165 129.795 ;
        RECT 117.345 129.465 117.615 129.795 ;
        RECT 117.830 129.295 118.145 130.315 ;
        RECT 118.535 130.305 118.865 131.105 ;
        RECT 119.350 130.135 119.740 130.310 ;
        RECT 118.315 129.965 119.740 130.135 ;
        RECT 120.095 130.015 121.765 131.105 ;
        RECT 118.315 129.465 118.485 129.965 ;
        RECT 115.090 129.095 117.575 129.285 ;
        RECT 115.095 128.555 115.840 128.925 ;
        RECT 116.405 128.735 116.660 129.095 ;
        RECT 116.840 128.555 117.170 128.925 ;
        RECT 117.350 128.735 117.575 129.095 ;
        RECT 117.830 128.725 118.445 129.295 ;
        RECT 118.735 129.235 119.000 129.795 ;
        RECT 119.170 129.065 119.340 129.965 ;
        RECT 119.510 129.235 119.865 129.795 ;
        RECT 120.095 129.325 120.845 129.845 ;
        RECT 121.015 129.495 121.765 130.015 ;
        RECT 121.935 130.255 122.195 130.935 ;
        RECT 122.365 130.325 122.615 131.105 ;
        RECT 122.865 130.555 123.115 130.935 ;
        RECT 123.285 130.725 123.640 131.105 ;
        RECT 124.645 130.715 124.980 130.935 ;
        RECT 124.245 130.555 124.475 130.595 ;
        RECT 122.865 130.355 124.475 130.555 ;
        RECT 122.865 130.345 123.700 130.355 ;
        RECT 124.290 130.265 124.475 130.355 ;
        RECT 118.615 128.555 118.830 129.065 ;
        RECT 119.060 128.735 119.340 129.065 ;
        RECT 119.520 128.555 119.760 129.065 ;
        RECT 120.095 128.555 121.765 129.325 ;
        RECT 121.935 129.055 122.105 130.255 ;
        RECT 123.805 130.155 124.135 130.185 ;
        RECT 122.335 130.095 124.135 130.155 ;
        RECT 124.725 130.095 124.980 130.715 ;
        RECT 125.155 130.670 130.500 131.105 ;
        RECT 122.275 129.985 124.980 130.095 ;
        RECT 122.275 129.950 122.475 129.985 ;
        RECT 122.275 129.375 122.445 129.950 ;
        RECT 123.805 129.925 124.980 129.985 ;
        RECT 122.675 129.510 123.085 129.815 ;
        RECT 123.255 129.545 123.585 129.755 ;
        RECT 122.275 129.255 122.545 129.375 ;
        RECT 122.275 129.210 123.120 129.255 ;
        RECT 122.365 129.085 123.120 129.210 ;
        RECT 123.375 129.145 123.585 129.545 ;
        RECT 123.830 129.545 124.305 129.755 ;
        RECT 124.495 129.545 124.985 129.745 ;
        RECT 123.830 129.145 124.050 129.545 ;
        RECT 121.935 128.725 122.195 129.055 ;
        RECT 122.950 128.935 123.120 129.085 ;
        RECT 122.365 128.555 122.695 128.915 ;
        RECT 122.950 128.725 124.250 128.935 ;
        RECT 124.525 128.555 124.980 129.320 ;
        RECT 126.740 129.100 127.080 129.930 ;
        RECT 128.560 129.420 128.910 130.670 ;
        RECT 131.320 130.135 131.710 130.310 ;
        RECT 132.195 130.305 132.525 131.105 ;
        RECT 132.695 130.315 133.230 130.935 ;
        RECT 131.320 129.965 132.745 130.135 ;
        RECT 131.195 129.235 131.550 129.795 ;
        RECT 125.155 128.555 130.500 129.100 ;
        RECT 131.720 129.065 131.890 129.965 ;
        RECT 132.060 129.235 132.325 129.795 ;
        RECT 132.575 129.465 132.745 129.965 ;
        RECT 132.915 129.295 133.230 130.315 ;
        RECT 133.435 129.940 133.725 131.105 ;
        RECT 134.100 130.135 134.430 130.935 ;
        RECT 134.600 130.305 134.930 131.105 ;
        RECT 135.230 130.135 135.560 130.935 ;
        RECT 136.205 130.305 136.455 131.105 ;
        RECT 134.100 129.965 136.535 130.135 ;
        RECT 136.725 129.965 136.895 131.105 ;
        RECT 137.065 129.965 137.405 130.935 ;
        RECT 133.895 129.545 134.245 129.795 ;
        RECT 134.430 129.335 134.600 129.965 ;
        RECT 134.770 129.545 135.100 129.745 ;
        RECT 135.270 129.545 135.600 129.745 ;
        RECT 135.770 129.545 136.190 129.745 ;
        RECT 136.365 129.715 136.535 129.965 ;
        RECT 136.365 129.545 137.060 129.715 ;
        RECT 131.300 128.555 131.540 129.065 ;
        RECT 131.720 128.735 132.000 129.065 ;
        RECT 132.230 128.555 132.445 129.065 ;
        RECT 132.615 128.725 133.230 129.295 ;
        RECT 133.435 128.555 133.725 129.280 ;
        RECT 134.100 128.725 134.600 129.335 ;
        RECT 135.230 129.205 136.455 129.375 ;
        RECT 137.230 129.355 137.405 129.965 ;
        RECT 135.230 128.725 135.560 129.205 ;
        RECT 135.730 128.555 135.955 129.015 ;
        RECT 136.125 128.725 136.455 129.205 ;
        RECT 136.645 128.555 136.895 129.355 ;
        RECT 137.065 128.725 137.405 129.355 ;
        RECT 137.575 130.255 137.835 130.935 ;
        RECT 138.005 130.325 138.255 131.105 ;
        RECT 138.505 130.555 138.755 130.935 ;
        RECT 138.925 130.725 139.280 131.105 ;
        RECT 140.285 130.715 140.620 130.935 ;
        RECT 139.885 130.555 140.115 130.595 ;
        RECT 138.505 130.355 140.115 130.555 ;
        RECT 138.505 130.345 139.340 130.355 ;
        RECT 139.930 130.265 140.115 130.355 ;
        RECT 137.575 129.055 137.745 130.255 ;
        RECT 139.445 130.155 139.775 130.185 ;
        RECT 137.975 130.095 139.775 130.155 ;
        RECT 140.365 130.095 140.620 130.715 ;
        RECT 137.915 129.985 140.620 130.095 ;
        RECT 137.915 129.950 138.115 129.985 ;
        RECT 137.915 129.375 138.085 129.950 ;
        RECT 139.445 129.925 140.620 129.985 ;
        RECT 141.715 130.015 142.925 131.105 ;
        RECT 138.315 129.510 138.725 129.815 ;
        RECT 138.895 129.545 139.225 129.755 ;
        RECT 137.915 129.255 138.185 129.375 ;
        RECT 137.915 129.210 138.760 129.255 ;
        RECT 138.005 129.085 138.760 129.210 ;
        RECT 139.015 129.145 139.225 129.545 ;
        RECT 139.470 129.545 139.945 129.755 ;
        RECT 140.135 129.545 140.625 129.745 ;
        RECT 139.470 129.145 139.690 129.545 ;
        RECT 141.715 129.475 142.235 130.015 ;
        RECT 137.575 128.725 137.835 129.055 ;
        RECT 138.590 128.935 138.760 129.085 ;
        RECT 138.005 128.555 138.335 128.915 ;
        RECT 138.590 128.725 139.890 128.935 ;
        RECT 140.165 128.555 140.620 129.320 ;
        RECT 142.405 129.305 142.925 129.845 ;
        RECT 141.715 128.555 142.925 129.305 ;
        RECT 17.430 128.385 143.010 128.555 ;
        RECT 17.515 127.635 18.725 128.385 ;
        RECT 17.515 127.095 18.035 127.635 ;
        RECT 18.895 127.585 19.205 128.385 ;
        RECT 19.410 127.585 20.105 128.215 ;
        RECT 20.365 127.835 20.535 128.125 ;
        RECT 20.705 128.005 21.035 128.385 ;
        RECT 20.365 127.665 21.030 127.835 ;
        RECT 18.205 126.925 18.725 127.465 ;
        RECT 18.905 127.145 19.240 127.415 ;
        RECT 19.410 126.985 19.580 127.585 ;
        RECT 19.750 127.145 20.085 127.395 ;
        RECT 17.515 125.835 18.725 126.925 ;
        RECT 18.895 125.835 19.175 126.975 ;
        RECT 19.345 126.005 19.675 126.985 ;
        RECT 19.845 125.835 20.105 126.975 ;
        RECT 20.280 126.845 20.630 127.495 ;
        RECT 20.800 126.675 21.030 127.665 ;
        RECT 20.365 126.505 21.030 126.675 ;
        RECT 20.365 126.005 20.535 126.505 ;
        RECT 20.705 125.835 21.035 126.335 ;
        RECT 21.205 126.005 21.390 128.125 ;
        RECT 21.645 127.925 21.895 128.385 ;
        RECT 22.065 127.935 22.400 128.105 ;
        RECT 22.595 127.935 23.270 128.105 ;
        RECT 22.065 127.795 22.235 127.935 ;
        RECT 21.560 126.805 21.840 127.755 ;
        RECT 22.010 127.665 22.235 127.795 ;
        RECT 22.010 126.560 22.180 127.665 ;
        RECT 22.405 127.515 22.930 127.735 ;
        RECT 22.350 126.750 22.590 127.345 ;
        RECT 22.760 126.815 22.930 127.515 ;
        RECT 23.100 127.155 23.270 127.935 ;
        RECT 23.590 127.885 23.960 128.385 ;
        RECT 24.140 127.935 24.545 128.105 ;
        RECT 24.715 127.935 25.500 128.105 ;
        RECT 24.140 127.705 24.310 127.935 ;
        RECT 23.480 127.405 24.310 127.705 ;
        RECT 24.695 127.435 25.160 127.765 ;
        RECT 23.480 127.375 23.680 127.405 ;
        RECT 23.800 127.155 23.970 127.225 ;
        RECT 23.100 126.985 23.970 127.155 ;
        RECT 23.460 126.895 23.970 126.985 ;
        RECT 22.010 126.430 22.315 126.560 ;
        RECT 22.760 126.450 23.290 126.815 ;
        RECT 21.630 125.835 21.895 126.295 ;
        RECT 22.065 126.005 22.315 126.430 ;
        RECT 23.460 126.280 23.630 126.895 ;
        RECT 22.525 126.110 23.630 126.280 ;
        RECT 23.800 125.835 23.970 126.635 ;
        RECT 24.140 126.335 24.310 127.405 ;
        RECT 24.480 126.505 24.670 127.225 ;
        RECT 24.840 126.475 25.160 127.435 ;
        RECT 25.330 127.475 25.500 127.935 ;
        RECT 25.775 127.855 25.985 128.385 ;
        RECT 26.245 127.645 26.575 128.170 ;
        RECT 26.745 127.775 26.915 128.385 ;
        RECT 27.085 127.730 27.415 128.165 ;
        RECT 27.635 127.735 27.895 128.215 ;
        RECT 28.065 127.845 28.315 128.385 ;
        RECT 27.085 127.645 27.465 127.730 ;
        RECT 26.375 127.475 26.575 127.645 ;
        RECT 27.240 127.605 27.465 127.645 ;
        RECT 25.330 127.145 26.205 127.475 ;
        RECT 26.375 127.145 27.125 127.475 ;
        RECT 24.140 126.005 24.390 126.335 ;
        RECT 25.330 126.305 25.500 127.145 ;
        RECT 26.375 126.940 26.565 127.145 ;
        RECT 27.295 127.025 27.465 127.605 ;
        RECT 27.250 126.975 27.465 127.025 ;
        RECT 25.670 126.565 26.565 126.940 ;
        RECT 27.075 126.895 27.465 126.975 ;
        RECT 24.615 126.135 25.500 126.305 ;
        RECT 25.680 125.835 25.995 126.335 ;
        RECT 26.225 126.005 26.565 126.565 ;
        RECT 26.735 125.835 26.905 126.845 ;
        RECT 27.075 126.050 27.405 126.895 ;
        RECT 27.635 126.705 27.805 127.735 ;
        RECT 28.485 127.680 28.705 128.165 ;
        RECT 27.975 127.085 28.205 127.480 ;
        RECT 28.375 127.255 28.705 127.680 ;
        RECT 28.875 128.005 29.765 128.175 ;
        RECT 28.875 127.280 29.045 128.005 ;
        RECT 30.020 127.885 30.515 128.215 ;
        RECT 29.215 127.450 29.765 127.835 ;
        RECT 28.875 127.210 29.765 127.280 ;
        RECT 28.870 127.185 29.765 127.210 ;
        RECT 28.860 127.170 29.765 127.185 ;
        RECT 28.855 127.155 29.765 127.170 ;
        RECT 28.845 127.150 29.765 127.155 ;
        RECT 28.840 127.140 29.765 127.150 ;
        RECT 28.835 127.130 29.765 127.140 ;
        RECT 28.825 127.125 29.765 127.130 ;
        RECT 28.815 127.115 29.765 127.125 ;
        RECT 28.805 127.110 29.765 127.115 ;
        RECT 28.805 127.105 29.140 127.110 ;
        RECT 28.790 127.100 29.140 127.105 ;
        RECT 28.775 127.090 29.140 127.100 ;
        RECT 28.750 127.085 29.140 127.090 ;
        RECT 27.975 127.080 29.140 127.085 ;
        RECT 27.975 127.045 29.110 127.080 ;
        RECT 27.975 127.020 29.075 127.045 ;
        RECT 27.975 126.990 29.045 127.020 ;
        RECT 27.975 126.960 29.025 126.990 ;
        RECT 27.975 126.930 29.005 126.960 ;
        RECT 27.975 126.920 28.935 126.930 ;
        RECT 27.975 126.910 28.910 126.920 ;
        RECT 27.975 126.895 28.890 126.910 ;
        RECT 27.975 126.880 28.870 126.895 ;
        RECT 28.080 126.870 28.865 126.880 ;
        RECT 28.080 126.835 28.850 126.870 ;
        RECT 27.635 126.005 27.910 126.705 ;
        RECT 28.080 126.585 28.835 126.835 ;
        RECT 29.005 126.515 29.335 126.760 ;
        RECT 29.505 126.660 29.765 127.110 ;
        RECT 29.150 126.490 29.335 126.515 ;
        RECT 29.150 126.390 29.765 126.490 ;
        RECT 29.935 126.395 30.175 127.705 ;
        RECT 30.345 126.975 30.515 127.885 ;
        RECT 30.735 127.145 31.085 128.110 ;
        RECT 31.265 127.145 31.565 128.115 ;
        RECT 31.745 127.145 32.025 128.115 ;
        RECT 32.205 127.585 32.475 128.385 ;
        RECT 32.645 127.665 32.985 128.175 ;
        RECT 32.220 127.145 32.550 127.395 ;
        RECT 32.220 126.975 32.535 127.145 ;
        RECT 30.345 126.805 32.535 126.975 ;
        RECT 28.080 125.835 28.335 126.380 ;
        RECT 28.505 126.005 28.985 126.345 ;
        RECT 29.160 125.835 29.765 126.390 ;
        RECT 29.940 125.835 30.275 126.215 ;
        RECT 30.445 126.005 30.695 126.805 ;
        RECT 30.915 125.835 31.245 126.555 ;
        RECT 31.430 126.005 31.680 126.805 ;
        RECT 32.145 125.835 32.475 126.635 ;
        RECT 32.725 126.265 32.985 127.665 ;
        RECT 33.165 127.655 33.465 128.385 ;
        RECT 33.645 127.475 33.875 128.095 ;
        RECT 34.075 127.825 34.300 128.205 ;
        RECT 34.470 127.995 34.800 128.385 ;
        RECT 34.075 127.645 34.405 127.825 ;
        RECT 33.170 127.145 33.465 127.475 ;
        RECT 33.645 127.145 34.060 127.475 ;
        RECT 34.230 126.975 34.405 127.645 ;
        RECT 34.575 127.145 34.815 127.795 ;
        RECT 34.995 127.755 35.335 128.215 ;
        RECT 35.505 127.925 35.675 128.385 ;
        RECT 36.305 127.950 36.665 128.215 ;
        RECT 36.310 127.945 36.665 127.950 ;
        RECT 36.315 127.935 36.665 127.945 ;
        RECT 36.320 127.930 36.665 127.935 ;
        RECT 36.325 127.920 36.665 127.930 ;
        RECT 36.905 127.925 37.075 128.385 ;
        RECT 36.330 127.915 36.665 127.920 ;
        RECT 36.340 127.905 36.665 127.915 ;
        RECT 36.350 127.895 36.665 127.905 ;
        RECT 35.845 127.755 36.175 127.835 ;
        RECT 34.995 127.565 36.175 127.755 ;
        RECT 36.365 127.755 36.665 127.895 ;
        RECT 36.365 127.565 37.075 127.755 ;
        RECT 34.995 127.195 35.325 127.395 ;
        RECT 35.635 127.375 35.965 127.395 ;
        RECT 35.515 127.195 35.965 127.375 ;
        RECT 32.645 126.005 32.985 126.265 ;
        RECT 33.165 126.615 34.060 126.945 ;
        RECT 34.230 126.785 34.815 126.975 ;
        RECT 34.995 126.855 35.225 127.195 ;
        RECT 33.165 126.445 34.370 126.615 ;
        RECT 33.165 126.015 33.495 126.445 ;
        RECT 33.675 125.835 33.870 126.275 ;
        RECT 34.040 126.015 34.370 126.445 ;
        RECT 34.540 126.015 34.815 126.785 ;
        RECT 35.005 125.835 35.335 126.555 ;
        RECT 35.515 126.080 35.730 127.195 ;
        RECT 36.135 127.165 36.605 127.395 ;
        RECT 36.790 126.995 37.075 127.565 ;
        RECT 37.245 127.440 37.585 128.215 ;
        RECT 37.755 127.775 38.095 128.190 ;
        RECT 38.265 127.945 38.435 128.385 ;
        RECT 38.605 127.995 39.855 128.175 ;
        RECT 38.605 127.775 38.935 127.995 ;
        RECT 40.125 127.925 40.295 128.385 ;
        RECT 37.755 127.605 38.935 127.775 ;
        RECT 39.105 127.755 39.470 127.825 ;
        RECT 39.105 127.575 40.355 127.755 ;
        RECT 35.925 126.780 37.075 126.995 ;
        RECT 35.925 126.005 36.255 126.780 ;
        RECT 36.425 125.835 37.135 126.610 ;
        RECT 37.305 126.005 37.585 127.440 ;
        RECT 37.755 127.195 38.220 127.395 ;
        RECT 38.395 127.145 38.725 127.395 ;
        RECT 38.895 127.365 39.360 127.395 ;
        RECT 38.895 127.195 39.365 127.365 ;
        RECT 38.895 127.145 39.360 127.195 ;
        RECT 39.555 127.145 39.910 127.395 ;
        RECT 38.395 127.025 38.575 127.145 ;
        RECT 37.755 125.835 38.075 127.015 ;
        RECT 38.245 126.855 38.575 127.025 ;
        RECT 40.080 126.975 40.355 127.575 ;
        RECT 38.245 126.065 38.445 126.855 ;
        RECT 38.745 126.765 40.355 126.975 ;
        RECT 38.745 126.665 39.155 126.765 ;
        RECT 38.770 126.005 39.155 126.665 ;
        RECT 39.550 125.835 40.335 126.595 ;
        RECT 40.525 126.005 40.805 128.105 ;
        RECT 40.975 127.615 42.645 128.385 ;
        RECT 43.275 127.660 43.565 128.385 ;
        RECT 43.735 127.840 49.080 128.385 ;
        RECT 50.260 127.885 50.755 128.215 ;
        RECT 40.975 127.095 41.725 127.615 ;
        RECT 41.895 126.925 42.645 127.445 ;
        RECT 45.320 127.010 45.660 127.840 ;
        RECT 40.975 125.835 42.645 126.925 ;
        RECT 43.275 125.835 43.565 127.000 ;
        RECT 47.140 126.270 47.490 127.520 ;
        RECT 50.175 126.395 50.415 127.705 ;
        RECT 50.585 126.975 50.755 127.885 ;
        RECT 50.975 127.145 51.325 128.110 ;
        RECT 51.505 127.145 51.805 128.115 ;
        RECT 51.985 127.145 52.265 128.115 ;
        RECT 52.445 127.585 52.715 128.385 ;
        RECT 52.885 127.665 53.225 128.175 ;
        RECT 53.445 127.730 53.775 128.165 ;
        RECT 53.945 127.775 54.115 128.385 ;
        RECT 52.460 127.145 52.790 127.395 ;
        RECT 52.460 126.975 52.775 127.145 ;
        RECT 50.585 126.805 52.775 126.975 ;
        RECT 43.735 125.835 49.080 126.270 ;
        RECT 50.180 125.835 50.515 126.215 ;
        RECT 50.685 126.005 50.935 126.805 ;
        RECT 51.155 125.835 51.485 126.555 ;
        RECT 51.670 126.005 51.920 126.805 ;
        RECT 52.385 125.835 52.715 126.635 ;
        RECT 52.965 126.265 53.225 127.665 ;
        RECT 53.395 127.645 53.775 127.730 ;
        RECT 54.285 127.645 54.615 128.170 ;
        RECT 54.875 127.855 55.085 128.385 ;
        RECT 55.360 127.935 56.145 128.105 ;
        RECT 56.315 127.935 56.720 128.105 ;
        RECT 53.395 127.605 53.620 127.645 ;
        RECT 53.395 127.025 53.565 127.605 ;
        RECT 54.285 127.475 54.485 127.645 ;
        RECT 55.360 127.475 55.530 127.935 ;
        RECT 53.735 127.145 54.485 127.475 ;
        RECT 54.655 127.145 55.530 127.475 ;
        RECT 53.395 126.975 53.610 127.025 ;
        RECT 53.395 126.895 53.785 126.975 ;
        RECT 52.885 126.005 53.225 126.265 ;
        RECT 53.455 126.050 53.785 126.895 ;
        RECT 54.295 126.940 54.485 127.145 ;
        RECT 53.955 125.835 54.125 126.845 ;
        RECT 54.295 126.565 55.190 126.940 ;
        RECT 54.295 126.005 54.635 126.565 ;
        RECT 54.865 125.835 55.180 126.335 ;
        RECT 55.360 126.305 55.530 127.145 ;
        RECT 55.700 127.435 56.165 127.765 ;
        RECT 56.550 127.705 56.720 127.935 ;
        RECT 56.900 127.885 57.270 128.385 ;
        RECT 57.590 127.935 58.265 128.105 ;
        RECT 58.460 127.935 58.795 128.105 ;
        RECT 55.700 126.475 56.020 127.435 ;
        RECT 56.550 127.405 57.380 127.705 ;
        RECT 56.190 126.505 56.380 127.225 ;
        RECT 56.550 126.335 56.720 127.405 ;
        RECT 57.180 127.375 57.380 127.405 ;
        RECT 56.890 127.155 57.060 127.225 ;
        RECT 57.590 127.155 57.760 127.935 ;
        RECT 58.625 127.795 58.795 127.935 ;
        RECT 58.965 127.925 59.215 128.385 ;
        RECT 56.890 126.985 57.760 127.155 ;
        RECT 57.930 127.515 58.455 127.735 ;
        RECT 58.625 127.665 58.850 127.795 ;
        RECT 56.890 126.895 57.400 126.985 ;
        RECT 55.360 126.135 56.245 126.305 ;
        RECT 56.470 126.005 56.720 126.335 ;
        RECT 56.890 125.835 57.060 126.635 ;
        RECT 57.230 126.280 57.400 126.895 ;
        RECT 57.930 126.815 58.100 127.515 ;
        RECT 57.570 126.450 58.100 126.815 ;
        RECT 58.270 126.750 58.510 127.345 ;
        RECT 58.680 126.560 58.850 127.665 ;
        RECT 59.020 126.805 59.300 127.755 ;
        RECT 58.545 126.430 58.850 126.560 ;
        RECT 57.230 126.110 58.335 126.280 ;
        RECT 58.545 126.005 58.795 126.430 ;
        RECT 58.965 125.835 59.230 126.295 ;
        RECT 59.470 126.005 59.655 128.125 ;
        RECT 59.825 128.005 60.155 128.385 ;
        RECT 60.325 127.835 60.495 128.125 ;
        RECT 60.755 127.840 66.100 128.385 ;
        RECT 59.830 127.665 60.495 127.835 ;
        RECT 59.830 126.675 60.060 127.665 ;
        RECT 60.230 126.845 60.580 127.495 ;
        RECT 62.340 127.010 62.680 127.840 ;
        RECT 66.275 127.615 68.865 128.385 ;
        RECT 69.035 127.660 69.325 128.385 ;
        RECT 69.585 127.835 69.755 128.125 ;
        RECT 69.925 128.005 70.255 128.385 ;
        RECT 69.585 127.665 70.250 127.835 ;
        RECT 59.830 126.505 60.495 126.675 ;
        RECT 59.825 125.835 60.155 126.335 ;
        RECT 60.325 126.005 60.495 126.505 ;
        RECT 64.160 126.270 64.510 127.520 ;
        RECT 66.275 127.095 67.485 127.615 ;
        RECT 67.655 126.925 68.865 127.445 ;
        RECT 60.755 125.835 66.100 126.270 ;
        RECT 66.275 125.835 68.865 126.925 ;
        RECT 69.035 125.835 69.325 127.000 ;
        RECT 69.500 126.845 69.850 127.495 ;
        RECT 70.020 126.675 70.250 127.665 ;
        RECT 69.585 126.505 70.250 126.675 ;
        RECT 69.585 126.005 69.755 126.505 ;
        RECT 69.925 125.835 70.255 126.335 ;
        RECT 70.425 126.005 70.610 128.125 ;
        RECT 70.865 127.925 71.115 128.385 ;
        RECT 71.285 127.935 71.620 128.105 ;
        RECT 71.815 127.935 72.490 128.105 ;
        RECT 71.285 127.795 71.455 127.935 ;
        RECT 70.780 126.805 71.060 127.755 ;
        RECT 71.230 127.665 71.455 127.795 ;
        RECT 71.230 126.560 71.400 127.665 ;
        RECT 71.625 127.515 72.150 127.735 ;
        RECT 71.570 126.750 71.810 127.345 ;
        RECT 71.980 126.815 72.150 127.515 ;
        RECT 72.320 127.155 72.490 127.935 ;
        RECT 72.810 127.885 73.180 128.385 ;
        RECT 73.360 127.935 73.765 128.105 ;
        RECT 73.935 127.935 74.720 128.105 ;
        RECT 73.360 127.705 73.530 127.935 ;
        RECT 72.700 127.405 73.530 127.705 ;
        RECT 73.915 127.435 74.380 127.765 ;
        RECT 72.700 127.375 72.900 127.405 ;
        RECT 73.020 127.155 73.190 127.225 ;
        RECT 72.320 126.985 73.190 127.155 ;
        RECT 72.680 126.895 73.190 126.985 ;
        RECT 71.230 126.430 71.535 126.560 ;
        RECT 71.980 126.450 72.510 126.815 ;
        RECT 70.850 125.835 71.115 126.295 ;
        RECT 71.285 126.005 71.535 126.430 ;
        RECT 72.680 126.280 72.850 126.895 ;
        RECT 71.745 126.110 72.850 126.280 ;
        RECT 73.020 125.835 73.190 126.635 ;
        RECT 73.360 126.335 73.530 127.405 ;
        RECT 73.700 126.505 73.890 127.225 ;
        RECT 74.060 126.475 74.380 127.435 ;
        RECT 74.550 127.475 74.720 127.935 ;
        RECT 74.995 127.855 75.205 128.385 ;
        RECT 75.465 127.645 75.795 128.170 ;
        RECT 75.965 127.775 76.135 128.385 ;
        RECT 76.305 127.730 76.635 128.165 ;
        RECT 76.305 127.645 76.685 127.730 ;
        RECT 75.595 127.475 75.795 127.645 ;
        RECT 76.460 127.605 76.685 127.645 ;
        RECT 74.550 127.145 75.425 127.475 ;
        RECT 75.595 127.145 76.345 127.475 ;
        RECT 73.360 126.005 73.610 126.335 ;
        RECT 74.550 126.305 74.720 127.145 ;
        RECT 75.595 126.940 75.785 127.145 ;
        RECT 76.515 127.025 76.685 127.605 ;
        RECT 76.875 127.575 77.115 128.385 ;
        RECT 77.285 127.575 77.615 128.215 ;
        RECT 77.785 127.575 78.055 128.385 ;
        RECT 76.855 127.145 77.205 127.395 ;
        RECT 76.470 126.975 76.685 127.025 ;
        RECT 77.375 126.975 77.545 127.575 ;
        RECT 78.235 127.565 78.495 128.385 ;
        RECT 78.665 127.565 78.995 127.985 ;
        RECT 79.175 127.900 79.965 128.165 ;
        RECT 78.745 127.475 78.995 127.565 ;
        RECT 77.715 127.145 78.065 127.395 ;
        RECT 74.890 126.565 75.785 126.940 ;
        RECT 76.295 126.895 76.685 126.975 ;
        RECT 73.835 126.135 74.720 126.305 ;
        RECT 74.900 125.835 75.215 126.335 ;
        RECT 75.445 126.005 75.785 126.565 ;
        RECT 75.955 125.835 76.125 126.845 ;
        RECT 76.295 126.050 76.625 126.895 ;
        RECT 76.865 126.805 77.545 126.975 ;
        RECT 76.865 126.020 77.195 126.805 ;
        RECT 77.725 125.835 78.055 126.975 ;
        RECT 78.235 126.515 78.575 127.395 ;
        RECT 78.745 127.225 79.540 127.475 ;
        RECT 78.235 125.835 78.495 126.345 ;
        RECT 78.745 126.005 78.915 127.225 ;
        RECT 79.710 127.045 79.965 127.900 ;
        RECT 80.135 127.745 80.335 128.165 ;
        RECT 80.525 127.925 80.855 128.385 ;
        RECT 80.135 127.225 80.545 127.745 ;
        RECT 81.025 127.735 81.285 128.215 ;
        RECT 80.715 127.045 80.945 127.475 ;
        RECT 79.155 126.875 80.945 127.045 ;
        RECT 79.155 126.510 79.405 126.875 ;
        RECT 79.575 126.515 79.905 126.705 ;
        RECT 80.125 126.580 80.840 126.875 ;
        RECT 81.115 126.705 81.285 127.735 ;
        RECT 81.730 127.575 81.975 128.180 ;
        RECT 82.195 127.850 82.705 128.385 ;
        RECT 79.575 126.340 79.770 126.515 ;
        RECT 79.155 125.835 79.770 126.340 ;
        RECT 79.940 126.005 80.415 126.345 ;
        RECT 80.585 125.835 80.800 126.380 ;
        RECT 81.010 126.005 81.285 126.705 ;
        RECT 81.455 127.405 82.685 127.575 ;
        RECT 81.455 126.595 81.795 127.405 ;
        RECT 81.965 126.840 82.715 127.030 ;
        RECT 81.455 126.185 81.970 126.595 ;
        RECT 82.205 125.835 82.375 126.595 ;
        RECT 82.545 126.175 82.715 126.840 ;
        RECT 82.885 126.855 83.075 128.215 ;
        RECT 83.245 127.365 83.520 128.215 ;
        RECT 83.710 127.850 84.240 128.215 ;
        RECT 84.665 127.985 84.995 128.385 ;
        RECT 84.065 127.815 84.240 127.850 ;
        RECT 83.245 127.195 83.525 127.365 ;
        RECT 83.245 127.055 83.520 127.195 ;
        RECT 83.725 126.855 83.895 127.655 ;
        RECT 82.885 126.685 83.895 126.855 ;
        RECT 84.065 127.645 84.995 127.815 ;
        RECT 85.165 127.645 85.420 128.215 ;
        RECT 85.685 127.835 85.855 128.125 ;
        RECT 86.025 128.005 86.355 128.385 ;
        RECT 85.685 127.665 86.350 127.835 ;
        RECT 84.065 126.515 84.235 127.645 ;
        RECT 84.825 127.475 84.995 127.645 ;
        RECT 83.110 126.345 84.235 126.515 ;
        RECT 84.405 127.145 84.600 127.475 ;
        RECT 84.825 127.145 85.080 127.475 ;
        RECT 84.405 126.175 84.575 127.145 ;
        RECT 85.250 126.975 85.420 127.645 ;
        RECT 82.545 126.005 84.575 126.175 ;
        RECT 84.745 125.835 84.915 126.975 ;
        RECT 85.085 126.005 85.420 126.975 ;
        RECT 85.600 126.845 85.950 127.495 ;
        RECT 86.120 126.675 86.350 127.665 ;
        RECT 85.685 126.505 86.350 126.675 ;
        RECT 85.685 126.005 85.855 126.505 ;
        RECT 86.025 125.835 86.355 126.335 ;
        RECT 86.525 126.005 86.710 128.125 ;
        RECT 86.965 127.925 87.215 128.385 ;
        RECT 87.385 127.935 87.720 128.105 ;
        RECT 87.915 127.935 88.590 128.105 ;
        RECT 87.385 127.795 87.555 127.935 ;
        RECT 86.880 126.805 87.160 127.755 ;
        RECT 87.330 127.665 87.555 127.795 ;
        RECT 87.330 126.560 87.500 127.665 ;
        RECT 87.725 127.515 88.250 127.735 ;
        RECT 87.670 126.750 87.910 127.345 ;
        RECT 88.080 126.815 88.250 127.515 ;
        RECT 88.420 127.155 88.590 127.935 ;
        RECT 88.910 127.885 89.280 128.385 ;
        RECT 89.460 127.935 89.865 128.105 ;
        RECT 90.035 127.935 90.820 128.105 ;
        RECT 89.460 127.705 89.630 127.935 ;
        RECT 88.800 127.405 89.630 127.705 ;
        RECT 90.015 127.435 90.480 127.765 ;
        RECT 88.800 127.375 89.000 127.405 ;
        RECT 89.120 127.155 89.290 127.225 ;
        RECT 88.420 126.985 89.290 127.155 ;
        RECT 88.780 126.895 89.290 126.985 ;
        RECT 87.330 126.430 87.635 126.560 ;
        RECT 88.080 126.450 88.610 126.815 ;
        RECT 86.950 125.835 87.215 126.295 ;
        RECT 87.385 126.005 87.635 126.430 ;
        RECT 88.780 126.280 88.950 126.895 ;
        RECT 87.845 126.110 88.950 126.280 ;
        RECT 89.120 125.835 89.290 126.635 ;
        RECT 89.460 126.335 89.630 127.405 ;
        RECT 89.800 126.505 89.990 127.225 ;
        RECT 90.160 126.475 90.480 127.435 ;
        RECT 90.650 127.475 90.820 127.935 ;
        RECT 91.095 127.855 91.305 128.385 ;
        RECT 91.565 127.645 91.895 128.170 ;
        RECT 92.065 127.775 92.235 128.385 ;
        RECT 92.405 127.730 92.735 128.165 ;
        RECT 92.905 127.870 93.075 128.385 ;
        RECT 92.405 127.645 92.785 127.730 ;
        RECT 91.695 127.475 91.895 127.645 ;
        RECT 92.560 127.605 92.785 127.645 ;
        RECT 90.650 127.145 91.525 127.475 ;
        RECT 91.695 127.145 92.445 127.475 ;
        RECT 89.460 126.005 89.710 126.335 ;
        RECT 90.650 126.305 90.820 127.145 ;
        RECT 91.695 126.940 91.885 127.145 ;
        RECT 92.615 127.025 92.785 127.605 ;
        RECT 93.415 127.635 94.625 128.385 ;
        RECT 94.795 127.660 95.085 128.385 ;
        RECT 93.415 127.095 93.935 127.635 ;
        RECT 95.255 127.615 96.925 128.385 ;
        RECT 97.185 127.835 97.355 128.125 ;
        RECT 97.525 128.005 97.855 128.385 ;
        RECT 97.185 127.665 97.850 127.835 ;
        RECT 92.570 126.975 92.785 127.025 ;
        RECT 90.990 126.565 91.885 126.940 ;
        RECT 92.395 126.895 92.785 126.975 ;
        RECT 94.105 126.925 94.625 127.465 ;
        RECT 95.255 127.095 96.005 127.615 ;
        RECT 89.935 126.135 90.820 126.305 ;
        RECT 91.000 125.835 91.315 126.335 ;
        RECT 91.545 126.005 91.885 126.565 ;
        RECT 92.055 125.835 92.225 126.845 ;
        RECT 92.395 126.050 92.725 126.895 ;
        RECT 92.895 125.835 93.065 126.750 ;
        RECT 93.415 125.835 94.625 126.925 ;
        RECT 94.795 125.835 95.085 127.000 ;
        RECT 96.175 126.925 96.925 127.445 ;
        RECT 95.255 125.835 96.925 126.925 ;
        RECT 97.100 126.845 97.450 127.495 ;
        RECT 97.620 126.675 97.850 127.665 ;
        RECT 97.185 126.505 97.850 126.675 ;
        RECT 97.185 126.005 97.355 126.505 ;
        RECT 97.525 125.835 97.855 126.335 ;
        RECT 98.025 126.005 98.210 128.125 ;
        RECT 98.465 127.925 98.715 128.385 ;
        RECT 98.885 127.935 99.220 128.105 ;
        RECT 99.415 127.935 100.090 128.105 ;
        RECT 98.885 127.795 99.055 127.935 ;
        RECT 98.380 126.805 98.660 127.755 ;
        RECT 98.830 127.665 99.055 127.795 ;
        RECT 98.830 126.560 99.000 127.665 ;
        RECT 99.225 127.515 99.750 127.735 ;
        RECT 99.170 126.750 99.410 127.345 ;
        RECT 99.580 126.815 99.750 127.515 ;
        RECT 99.920 127.155 100.090 127.935 ;
        RECT 100.410 127.885 100.780 128.385 ;
        RECT 100.960 127.935 101.365 128.105 ;
        RECT 101.535 127.935 102.320 128.105 ;
        RECT 100.960 127.705 101.130 127.935 ;
        RECT 100.300 127.405 101.130 127.705 ;
        RECT 101.515 127.435 101.980 127.765 ;
        RECT 100.300 127.375 100.500 127.405 ;
        RECT 100.620 127.155 100.790 127.225 ;
        RECT 99.920 126.985 100.790 127.155 ;
        RECT 100.280 126.895 100.790 126.985 ;
        RECT 98.830 126.430 99.135 126.560 ;
        RECT 99.580 126.450 100.110 126.815 ;
        RECT 98.450 125.835 98.715 126.295 ;
        RECT 98.885 126.005 99.135 126.430 ;
        RECT 100.280 126.280 100.450 126.895 ;
        RECT 99.345 126.110 100.450 126.280 ;
        RECT 100.620 125.835 100.790 126.635 ;
        RECT 100.960 126.335 101.130 127.405 ;
        RECT 101.300 126.505 101.490 127.225 ;
        RECT 101.660 126.475 101.980 127.435 ;
        RECT 102.150 127.475 102.320 127.935 ;
        RECT 102.595 127.855 102.805 128.385 ;
        RECT 103.065 127.645 103.395 128.170 ;
        RECT 103.565 127.775 103.735 128.385 ;
        RECT 103.905 127.730 104.235 128.165 ;
        RECT 103.905 127.645 104.285 127.730 ;
        RECT 103.195 127.475 103.395 127.645 ;
        RECT 104.060 127.605 104.285 127.645 ;
        RECT 102.150 127.145 103.025 127.475 ;
        RECT 103.195 127.145 103.945 127.475 ;
        RECT 100.960 126.005 101.210 126.335 ;
        RECT 102.150 126.305 102.320 127.145 ;
        RECT 103.195 126.940 103.385 127.145 ;
        RECT 104.115 127.025 104.285 127.605 ;
        RECT 104.070 126.975 104.285 127.025 ;
        RECT 102.490 126.565 103.385 126.940 ;
        RECT 103.895 126.895 104.285 126.975 ;
        RECT 104.460 127.645 104.715 128.215 ;
        RECT 104.885 127.985 105.215 128.385 ;
        RECT 105.640 127.850 106.170 128.215 ;
        RECT 105.640 127.815 105.815 127.850 ;
        RECT 104.885 127.645 105.815 127.815 ;
        RECT 104.460 126.975 104.630 127.645 ;
        RECT 104.885 127.475 105.055 127.645 ;
        RECT 104.800 127.145 105.055 127.475 ;
        RECT 105.280 127.145 105.475 127.475 ;
        RECT 101.435 126.135 102.320 126.305 ;
        RECT 102.500 125.835 102.815 126.335 ;
        RECT 103.045 126.005 103.385 126.565 ;
        RECT 103.555 125.835 103.725 126.845 ;
        RECT 103.895 126.050 104.225 126.895 ;
        RECT 104.460 126.005 104.795 126.975 ;
        RECT 104.965 125.835 105.135 126.975 ;
        RECT 105.305 126.175 105.475 127.145 ;
        RECT 105.645 126.515 105.815 127.645 ;
        RECT 105.985 126.855 106.155 127.655 ;
        RECT 106.360 127.365 106.635 128.215 ;
        RECT 106.355 127.195 106.635 127.365 ;
        RECT 106.360 127.055 106.635 127.195 ;
        RECT 106.805 126.855 106.995 128.215 ;
        RECT 107.175 127.850 107.685 128.385 ;
        RECT 107.905 127.575 108.150 128.180 ;
        RECT 108.595 127.635 109.805 128.385 ;
        RECT 110.065 127.835 110.235 128.125 ;
        RECT 110.405 128.005 110.735 128.385 ;
        RECT 110.065 127.665 110.730 127.835 ;
        RECT 107.195 127.405 108.425 127.575 ;
        RECT 105.985 126.685 106.995 126.855 ;
        RECT 107.165 126.840 107.915 127.030 ;
        RECT 105.645 126.345 106.770 126.515 ;
        RECT 107.165 126.175 107.335 126.840 ;
        RECT 108.085 126.595 108.425 127.405 ;
        RECT 108.595 127.095 109.115 127.635 ;
        RECT 109.285 126.925 109.805 127.465 ;
        RECT 105.305 126.005 107.335 126.175 ;
        RECT 107.505 125.835 107.675 126.595 ;
        RECT 107.910 126.185 108.425 126.595 ;
        RECT 108.595 125.835 109.805 126.925 ;
        RECT 109.980 126.845 110.330 127.495 ;
        RECT 110.500 126.675 110.730 127.665 ;
        RECT 110.065 126.505 110.730 126.675 ;
        RECT 110.065 126.005 110.235 126.505 ;
        RECT 110.405 125.835 110.735 126.335 ;
        RECT 110.905 126.005 111.090 128.125 ;
        RECT 111.345 127.925 111.595 128.385 ;
        RECT 111.765 127.935 112.100 128.105 ;
        RECT 112.295 127.935 112.970 128.105 ;
        RECT 111.765 127.795 111.935 127.935 ;
        RECT 111.260 126.805 111.540 127.755 ;
        RECT 111.710 127.665 111.935 127.795 ;
        RECT 111.710 126.560 111.880 127.665 ;
        RECT 112.105 127.515 112.630 127.735 ;
        RECT 112.050 126.750 112.290 127.345 ;
        RECT 112.460 126.815 112.630 127.515 ;
        RECT 112.800 127.155 112.970 127.935 ;
        RECT 113.290 127.885 113.660 128.385 ;
        RECT 113.840 127.935 114.245 128.105 ;
        RECT 114.415 127.935 115.200 128.105 ;
        RECT 113.840 127.705 114.010 127.935 ;
        RECT 113.180 127.405 114.010 127.705 ;
        RECT 114.395 127.435 114.860 127.765 ;
        RECT 113.180 127.375 113.380 127.405 ;
        RECT 113.500 127.155 113.670 127.225 ;
        RECT 112.800 126.985 113.670 127.155 ;
        RECT 113.160 126.895 113.670 126.985 ;
        RECT 111.710 126.430 112.015 126.560 ;
        RECT 112.460 126.450 112.990 126.815 ;
        RECT 111.330 125.835 111.595 126.295 ;
        RECT 111.765 126.005 112.015 126.430 ;
        RECT 113.160 126.280 113.330 126.895 ;
        RECT 112.225 126.110 113.330 126.280 ;
        RECT 113.500 125.835 113.670 126.635 ;
        RECT 113.840 126.335 114.010 127.405 ;
        RECT 114.180 126.505 114.370 127.225 ;
        RECT 114.540 126.475 114.860 127.435 ;
        RECT 115.030 127.475 115.200 127.935 ;
        RECT 115.475 127.855 115.685 128.385 ;
        RECT 115.945 127.645 116.275 128.170 ;
        RECT 116.445 127.775 116.615 128.385 ;
        RECT 116.785 127.730 117.115 128.165 ;
        RECT 117.335 127.885 117.635 128.215 ;
        RECT 117.805 127.905 118.080 128.385 ;
        RECT 116.785 127.645 117.165 127.730 ;
        RECT 116.075 127.475 116.275 127.645 ;
        RECT 116.940 127.605 117.165 127.645 ;
        RECT 115.030 127.145 115.905 127.475 ;
        RECT 116.075 127.145 116.825 127.475 ;
        RECT 113.840 126.005 114.090 126.335 ;
        RECT 115.030 126.305 115.200 127.145 ;
        RECT 116.075 126.940 116.265 127.145 ;
        RECT 116.995 127.025 117.165 127.605 ;
        RECT 116.950 126.975 117.165 127.025 ;
        RECT 115.370 126.565 116.265 126.940 ;
        RECT 116.775 126.895 117.165 126.975 ;
        RECT 117.335 126.975 117.505 127.885 ;
        RECT 118.260 127.735 118.555 128.125 ;
        RECT 118.725 127.905 118.980 128.385 ;
        RECT 119.155 127.735 119.415 128.125 ;
        RECT 119.585 127.905 119.865 128.385 ;
        RECT 117.675 127.145 118.025 127.715 ;
        RECT 118.260 127.565 119.910 127.735 ;
        RECT 120.555 127.660 120.845 128.385 ;
        RECT 121.105 127.835 121.275 128.125 ;
        RECT 121.445 128.005 121.775 128.385 ;
        RECT 121.105 127.665 121.770 127.835 ;
        RECT 118.195 127.225 119.335 127.395 ;
        RECT 118.195 126.975 118.365 127.225 ;
        RECT 119.505 127.055 119.910 127.565 ;
        RECT 114.315 126.135 115.200 126.305 ;
        RECT 115.380 125.835 115.695 126.335 ;
        RECT 115.925 126.005 116.265 126.565 ;
        RECT 116.435 125.835 116.605 126.845 ;
        RECT 116.775 126.050 117.105 126.895 ;
        RECT 117.335 126.805 118.365 126.975 ;
        RECT 119.155 126.885 119.910 127.055 ;
        RECT 117.335 126.005 117.645 126.805 ;
        RECT 119.155 126.635 119.415 126.885 ;
        RECT 117.815 125.835 118.125 126.635 ;
        RECT 118.295 126.465 119.415 126.635 ;
        RECT 118.295 126.005 118.555 126.465 ;
        RECT 118.725 125.835 118.980 126.295 ;
        RECT 119.155 126.005 119.415 126.465 ;
        RECT 119.585 125.835 119.870 126.705 ;
        RECT 120.555 125.835 120.845 127.000 ;
        RECT 121.020 126.845 121.370 127.495 ;
        RECT 121.540 126.675 121.770 127.665 ;
        RECT 121.105 126.505 121.770 126.675 ;
        RECT 121.105 126.005 121.275 126.505 ;
        RECT 121.445 125.835 121.775 126.335 ;
        RECT 121.945 126.005 122.130 128.125 ;
        RECT 122.385 127.925 122.635 128.385 ;
        RECT 122.805 127.935 123.140 128.105 ;
        RECT 123.335 127.935 124.010 128.105 ;
        RECT 122.805 127.795 122.975 127.935 ;
        RECT 122.300 126.805 122.580 127.755 ;
        RECT 122.750 127.665 122.975 127.795 ;
        RECT 122.750 126.560 122.920 127.665 ;
        RECT 123.145 127.515 123.670 127.735 ;
        RECT 123.090 126.750 123.330 127.345 ;
        RECT 123.500 126.815 123.670 127.515 ;
        RECT 123.840 127.155 124.010 127.935 ;
        RECT 124.330 127.885 124.700 128.385 ;
        RECT 124.880 127.935 125.285 128.105 ;
        RECT 125.455 127.935 126.240 128.105 ;
        RECT 124.880 127.705 125.050 127.935 ;
        RECT 124.220 127.405 125.050 127.705 ;
        RECT 125.435 127.435 125.900 127.765 ;
        RECT 124.220 127.375 124.420 127.405 ;
        RECT 124.540 127.155 124.710 127.225 ;
        RECT 123.840 126.985 124.710 127.155 ;
        RECT 124.200 126.895 124.710 126.985 ;
        RECT 122.750 126.430 123.055 126.560 ;
        RECT 123.500 126.450 124.030 126.815 ;
        RECT 122.370 125.835 122.635 126.295 ;
        RECT 122.805 126.005 123.055 126.430 ;
        RECT 124.200 126.280 124.370 126.895 ;
        RECT 123.265 126.110 124.370 126.280 ;
        RECT 124.540 125.835 124.710 126.635 ;
        RECT 124.880 126.335 125.050 127.405 ;
        RECT 125.220 126.505 125.410 127.225 ;
        RECT 125.580 126.475 125.900 127.435 ;
        RECT 126.070 127.475 126.240 127.935 ;
        RECT 126.515 127.855 126.725 128.385 ;
        RECT 126.985 127.645 127.315 128.170 ;
        RECT 127.485 127.775 127.655 128.385 ;
        RECT 127.825 127.730 128.155 128.165 ;
        RECT 127.825 127.645 128.205 127.730 ;
        RECT 127.115 127.475 127.315 127.645 ;
        RECT 127.980 127.605 128.205 127.645 ;
        RECT 126.070 127.145 126.945 127.475 ;
        RECT 127.115 127.145 127.865 127.475 ;
        RECT 124.880 126.005 125.130 126.335 ;
        RECT 126.070 126.305 126.240 127.145 ;
        RECT 127.115 126.940 127.305 127.145 ;
        RECT 128.035 127.025 128.205 127.605 ;
        RECT 128.375 127.615 130.965 128.385 ;
        RECT 131.225 127.835 131.395 128.125 ;
        RECT 131.565 128.005 131.895 128.385 ;
        RECT 131.225 127.665 131.890 127.835 ;
        RECT 128.375 127.095 129.585 127.615 ;
        RECT 127.990 126.975 128.205 127.025 ;
        RECT 126.410 126.565 127.305 126.940 ;
        RECT 127.815 126.895 128.205 126.975 ;
        RECT 129.755 126.925 130.965 127.445 ;
        RECT 125.355 126.135 126.240 126.305 ;
        RECT 126.420 125.835 126.735 126.335 ;
        RECT 126.965 126.005 127.305 126.565 ;
        RECT 127.475 125.835 127.645 126.845 ;
        RECT 127.815 126.050 128.145 126.895 ;
        RECT 128.375 125.835 130.965 126.925 ;
        RECT 131.140 126.845 131.490 127.495 ;
        RECT 131.660 126.675 131.890 127.665 ;
        RECT 131.225 126.505 131.890 126.675 ;
        RECT 131.225 126.005 131.395 126.505 ;
        RECT 131.565 125.835 131.895 126.335 ;
        RECT 132.065 126.005 132.250 128.125 ;
        RECT 132.505 127.925 132.755 128.385 ;
        RECT 132.925 127.935 133.260 128.105 ;
        RECT 133.455 127.935 134.130 128.105 ;
        RECT 132.925 127.795 133.095 127.935 ;
        RECT 132.420 126.805 132.700 127.755 ;
        RECT 132.870 127.665 133.095 127.795 ;
        RECT 132.870 126.560 133.040 127.665 ;
        RECT 133.265 127.515 133.790 127.735 ;
        RECT 133.210 126.750 133.450 127.345 ;
        RECT 133.620 126.815 133.790 127.515 ;
        RECT 133.960 127.155 134.130 127.935 ;
        RECT 134.450 127.885 134.820 128.385 ;
        RECT 135.000 127.935 135.405 128.105 ;
        RECT 135.575 127.935 136.360 128.105 ;
        RECT 135.000 127.705 135.170 127.935 ;
        RECT 134.340 127.405 135.170 127.705 ;
        RECT 135.555 127.435 136.020 127.765 ;
        RECT 134.340 127.375 134.540 127.405 ;
        RECT 134.660 127.155 134.830 127.225 ;
        RECT 133.960 126.985 134.830 127.155 ;
        RECT 134.320 126.895 134.830 126.985 ;
        RECT 132.870 126.430 133.175 126.560 ;
        RECT 133.620 126.450 134.150 126.815 ;
        RECT 132.490 125.835 132.755 126.295 ;
        RECT 132.925 126.005 133.175 126.430 ;
        RECT 134.320 126.280 134.490 126.895 ;
        RECT 133.385 126.110 134.490 126.280 ;
        RECT 134.660 125.835 134.830 126.635 ;
        RECT 135.000 126.335 135.170 127.405 ;
        RECT 135.340 126.505 135.530 127.225 ;
        RECT 135.700 126.475 136.020 127.435 ;
        RECT 136.190 127.475 136.360 127.935 ;
        RECT 136.635 127.855 136.845 128.385 ;
        RECT 137.105 127.645 137.435 128.170 ;
        RECT 137.605 127.775 137.775 128.385 ;
        RECT 137.945 127.730 138.275 128.165 ;
        RECT 137.945 127.645 138.325 127.730 ;
        RECT 137.235 127.475 137.435 127.645 ;
        RECT 138.100 127.605 138.325 127.645 ;
        RECT 136.190 127.145 137.065 127.475 ;
        RECT 137.235 127.145 137.985 127.475 ;
        RECT 135.000 126.005 135.250 126.335 ;
        RECT 136.190 126.305 136.360 127.145 ;
        RECT 137.235 126.940 137.425 127.145 ;
        RECT 138.155 127.025 138.325 127.605 ;
        RECT 138.495 127.635 139.705 128.385 ;
        RECT 139.965 127.835 140.135 128.215 ;
        RECT 140.350 128.005 140.680 128.385 ;
        RECT 139.965 127.665 140.680 127.835 ;
        RECT 138.495 127.095 139.015 127.635 ;
        RECT 138.110 126.975 138.325 127.025 ;
        RECT 136.530 126.565 137.425 126.940 ;
        RECT 137.935 126.895 138.325 126.975 ;
        RECT 139.185 126.925 139.705 127.465 ;
        RECT 139.875 127.115 140.230 127.485 ;
        RECT 140.510 127.475 140.680 127.665 ;
        RECT 140.850 127.640 141.105 128.215 ;
        RECT 140.510 127.145 140.765 127.475 ;
        RECT 140.510 126.935 140.680 127.145 ;
        RECT 135.475 126.135 136.360 126.305 ;
        RECT 136.540 125.835 136.855 126.335 ;
        RECT 137.085 126.005 137.425 126.565 ;
        RECT 137.595 125.835 137.765 126.845 ;
        RECT 137.935 126.050 138.265 126.895 ;
        RECT 138.495 125.835 139.705 126.925 ;
        RECT 139.965 126.765 140.680 126.935 ;
        RECT 140.935 126.910 141.105 127.640 ;
        RECT 141.280 127.545 141.540 128.385 ;
        RECT 141.715 127.635 142.925 128.385 ;
        RECT 139.965 126.005 140.135 126.765 ;
        RECT 140.350 125.835 140.680 126.595 ;
        RECT 140.850 126.005 141.105 126.910 ;
        RECT 141.280 125.835 141.540 126.985 ;
        RECT 141.715 126.925 142.235 127.465 ;
        RECT 142.405 127.095 142.925 127.635 ;
        RECT 141.715 125.835 142.925 126.925 ;
        RECT 17.430 125.665 143.010 125.835 ;
        RECT 17.515 124.575 18.725 125.665 ;
        RECT 18.895 124.575 21.485 125.665 ;
        RECT 22.205 124.995 22.375 125.495 ;
        RECT 22.545 125.165 22.875 125.665 ;
        RECT 22.205 124.825 22.870 124.995 ;
        RECT 17.515 123.865 18.035 124.405 ;
        RECT 18.205 124.035 18.725 124.575 ;
        RECT 18.895 123.885 20.105 124.405 ;
        RECT 20.275 124.055 21.485 124.575 ;
        RECT 22.120 124.005 22.470 124.655 ;
        RECT 17.515 123.115 18.725 123.865 ;
        RECT 18.895 123.115 21.485 123.885 ;
        RECT 22.640 123.835 22.870 124.825 ;
        RECT 22.205 123.665 22.870 123.835 ;
        RECT 22.205 123.375 22.375 123.665 ;
        RECT 22.545 123.115 22.875 123.495 ;
        RECT 23.045 123.375 23.230 125.495 ;
        RECT 23.470 125.205 23.735 125.665 ;
        RECT 23.905 125.070 24.155 125.495 ;
        RECT 24.365 125.220 25.470 125.390 ;
        RECT 23.850 124.940 24.155 125.070 ;
        RECT 23.400 123.745 23.680 124.695 ;
        RECT 23.850 123.835 24.020 124.940 ;
        RECT 24.190 124.155 24.430 124.750 ;
        RECT 24.600 124.685 25.130 125.050 ;
        RECT 24.600 123.985 24.770 124.685 ;
        RECT 25.300 124.605 25.470 125.220 ;
        RECT 25.640 124.865 25.810 125.665 ;
        RECT 25.980 125.165 26.230 125.495 ;
        RECT 26.455 125.195 27.340 125.365 ;
        RECT 25.300 124.515 25.810 124.605 ;
        RECT 23.850 123.705 24.075 123.835 ;
        RECT 24.245 123.765 24.770 123.985 ;
        RECT 24.940 124.345 25.810 124.515 ;
        RECT 23.485 123.115 23.735 123.575 ;
        RECT 23.905 123.565 24.075 123.705 ;
        RECT 24.940 123.565 25.110 124.345 ;
        RECT 25.640 124.275 25.810 124.345 ;
        RECT 25.320 124.095 25.520 124.125 ;
        RECT 25.980 124.095 26.150 125.165 ;
        RECT 26.320 124.275 26.510 124.995 ;
        RECT 25.320 123.795 26.150 124.095 ;
        RECT 26.680 124.065 27.000 125.025 ;
        RECT 23.905 123.395 24.240 123.565 ;
        RECT 24.435 123.395 25.110 123.565 ;
        RECT 25.430 123.115 25.800 123.615 ;
        RECT 25.980 123.565 26.150 123.795 ;
        RECT 26.535 123.735 27.000 124.065 ;
        RECT 27.170 124.355 27.340 125.195 ;
        RECT 27.520 125.165 27.835 125.665 ;
        RECT 28.065 124.935 28.405 125.495 ;
        RECT 27.510 124.560 28.405 124.935 ;
        RECT 28.575 124.655 28.745 125.665 ;
        RECT 28.215 124.355 28.405 124.560 ;
        RECT 28.915 124.605 29.245 125.450 ;
        RECT 28.915 124.525 29.305 124.605 ;
        RECT 29.090 124.475 29.305 124.525 ;
        RECT 30.395 124.500 30.685 125.665 ;
        RECT 30.855 125.110 31.460 125.665 ;
        RECT 31.635 125.155 32.115 125.495 ;
        RECT 32.285 125.120 32.540 125.665 ;
        RECT 30.855 125.010 31.470 125.110 ;
        RECT 31.285 124.985 31.470 125.010 ;
        RECT 27.170 124.025 28.045 124.355 ;
        RECT 28.215 124.025 28.965 124.355 ;
        RECT 27.170 123.565 27.340 124.025 ;
        RECT 28.215 123.855 28.415 124.025 ;
        RECT 29.135 123.895 29.305 124.475 ;
        RECT 30.855 124.390 31.115 124.840 ;
        RECT 31.285 124.740 31.615 124.985 ;
        RECT 31.785 124.665 32.540 124.915 ;
        RECT 32.710 124.795 32.985 125.495 ;
        RECT 31.770 124.630 32.540 124.665 ;
        RECT 31.755 124.620 32.540 124.630 ;
        RECT 31.750 124.605 32.645 124.620 ;
        RECT 31.730 124.590 32.645 124.605 ;
        RECT 31.710 124.580 32.645 124.590 ;
        RECT 31.685 124.570 32.645 124.580 ;
        RECT 31.615 124.540 32.645 124.570 ;
        RECT 31.595 124.510 32.645 124.540 ;
        RECT 31.575 124.480 32.645 124.510 ;
        RECT 31.545 124.455 32.645 124.480 ;
        RECT 31.510 124.420 32.645 124.455 ;
        RECT 31.480 124.415 32.645 124.420 ;
        RECT 31.480 124.410 31.870 124.415 ;
        RECT 31.480 124.400 31.845 124.410 ;
        RECT 31.480 124.395 31.830 124.400 ;
        RECT 31.480 124.390 31.815 124.395 ;
        RECT 30.855 124.385 31.815 124.390 ;
        RECT 30.855 124.375 31.805 124.385 ;
        RECT 30.855 124.370 31.795 124.375 ;
        RECT 30.855 124.360 31.785 124.370 ;
        RECT 30.855 124.350 31.780 124.360 ;
        RECT 30.855 124.345 31.775 124.350 ;
        RECT 30.855 124.330 31.765 124.345 ;
        RECT 30.855 124.315 31.760 124.330 ;
        RECT 30.855 124.290 31.750 124.315 ;
        RECT 30.855 124.220 31.745 124.290 ;
        RECT 29.080 123.855 29.305 123.895 ;
        RECT 25.980 123.395 26.385 123.565 ;
        RECT 26.555 123.395 27.340 123.565 ;
        RECT 27.615 123.115 27.825 123.645 ;
        RECT 28.085 123.330 28.415 123.855 ;
        RECT 28.925 123.770 29.305 123.855 ;
        RECT 28.585 123.115 28.755 123.725 ;
        RECT 28.925 123.335 29.255 123.770 ;
        RECT 30.395 123.115 30.685 123.840 ;
        RECT 30.855 123.665 31.405 124.050 ;
        RECT 31.575 123.495 31.745 124.220 ;
        RECT 30.855 123.325 31.745 123.495 ;
        RECT 31.915 123.820 32.245 124.245 ;
        RECT 32.415 124.020 32.645 124.415 ;
        RECT 31.915 123.335 32.135 123.820 ;
        RECT 32.815 123.765 32.985 124.795 ;
        RECT 33.165 124.695 33.495 125.480 ;
        RECT 33.165 124.525 33.845 124.695 ;
        RECT 34.025 124.525 34.355 125.665 ;
        RECT 35.455 124.815 35.835 125.495 ;
        RECT 36.425 124.815 36.595 125.665 ;
        RECT 36.765 124.985 37.095 125.495 ;
        RECT 37.265 125.155 37.435 125.665 ;
        RECT 37.605 124.985 38.005 125.495 ;
        RECT 36.765 124.815 38.005 124.985 ;
        RECT 33.155 124.105 33.505 124.355 ;
        RECT 33.675 123.925 33.845 124.525 ;
        RECT 34.015 124.105 34.365 124.355 ;
        RECT 32.305 123.115 32.555 123.655 ;
        RECT 32.725 123.285 32.985 123.765 ;
        RECT 33.175 123.115 33.415 123.925 ;
        RECT 33.585 123.285 33.915 123.925 ;
        RECT 34.085 123.115 34.355 123.925 ;
        RECT 35.455 123.855 35.625 124.815 ;
        RECT 35.795 124.475 37.100 124.645 ;
        RECT 38.185 124.565 38.505 125.495 ;
        RECT 38.765 124.995 38.935 125.495 ;
        RECT 39.105 125.165 39.435 125.665 ;
        RECT 38.765 124.825 39.430 124.995 ;
        RECT 35.795 124.025 36.040 124.475 ;
        RECT 36.210 124.105 36.760 124.305 ;
        RECT 36.930 124.275 37.100 124.475 ;
        RECT 37.875 124.395 38.505 124.565 ;
        RECT 36.930 124.105 37.305 124.275 ;
        RECT 37.475 123.855 37.705 124.355 ;
        RECT 35.455 123.685 37.705 123.855 ;
        RECT 35.505 123.115 35.835 123.505 ;
        RECT 36.005 123.365 36.175 123.685 ;
        RECT 37.875 123.515 38.045 124.395 ;
        RECT 38.680 124.005 39.030 124.655 ;
        RECT 36.345 123.115 36.675 123.505 ;
        RECT 37.090 123.345 38.045 123.515 ;
        RECT 38.215 123.115 38.505 123.950 ;
        RECT 39.200 123.835 39.430 124.825 ;
        RECT 38.765 123.665 39.430 123.835 ;
        RECT 38.765 123.375 38.935 123.665 ;
        RECT 39.105 123.115 39.435 123.495 ;
        RECT 39.605 123.375 39.790 125.495 ;
        RECT 40.030 125.205 40.295 125.665 ;
        RECT 40.465 125.070 40.715 125.495 ;
        RECT 40.925 125.220 42.030 125.390 ;
        RECT 40.410 124.940 40.715 125.070 ;
        RECT 39.960 123.745 40.240 124.695 ;
        RECT 40.410 123.835 40.580 124.940 ;
        RECT 40.750 124.155 40.990 124.750 ;
        RECT 41.160 124.685 41.690 125.050 ;
        RECT 41.160 123.985 41.330 124.685 ;
        RECT 41.860 124.605 42.030 125.220 ;
        RECT 42.200 124.865 42.370 125.665 ;
        RECT 42.540 125.165 42.790 125.495 ;
        RECT 43.015 125.195 43.900 125.365 ;
        RECT 41.860 124.515 42.370 124.605 ;
        RECT 40.410 123.705 40.635 123.835 ;
        RECT 40.805 123.765 41.330 123.985 ;
        RECT 41.500 124.345 42.370 124.515 ;
        RECT 40.045 123.115 40.295 123.575 ;
        RECT 40.465 123.565 40.635 123.705 ;
        RECT 41.500 123.565 41.670 124.345 ;
        RECT 42.200 124.275 42.370 124.345 ;
        RECT 41.880 124.095 42.080 124.125 ;
        RECT 42.540 124.095 42.710 125.165 ;
        RECT 42.880 124.275 43.070 124.995 ;
        RECT 41.880 123.795 42.710 124.095 ;
        RECT 43.240 124.065 43.560 125.025 ;
        RECT 40.465 123.395 40.800 123.565 ;
        RECT 40.995 123.395 41.670 123.565 ;
        RECT 41.990 123.115 42.360 123.615 ;
        RECT 42.540 123.565 42.710 123.795 ;
        RECT 43.095 123.735 43.560 124.065 ;
        RECT 43.730 124.355 43.900 125.195 ;
        RECT 44.080 125.165 44.395 125.665 ;
        RECT 44.625 124.935 44.965 125.495 ;
        RECT 44.070 124.560 44.965 124.935 ;
        RECT 45.135 124.655 45.305 125.665 ;
        RECT 44.775 124.355 44.965 124.560 ;
        RECT 45.475 124.605 45.805 125.450 ;
        RECT 46.045 125.055 46.375 125.485 ;
        RECT 46.555 125.225 46.750 125.665 ;
        RECT 46.920 125.055 47.250 125.485 ;
        RECT 46.045 124.885 47.250 125.055 ;
        RECT 45.475 124.525 45.865 124.605 ;
        RECT 46.045 124.555 46.940 124.885 ;
        RECT 47.420 124.715 47.695 125.485 ;
        RECT 47.875 125.110 48.480 125.665 ;
        RECT 48.655 125.155 49.135 125.495 ;
        RECT 49.305 125.120 49.560 125.665 ;
        RECT 47.875 125.010 48.490 125.110 ;
        RECT 48.305 124.985 48.490 125.010 ;
        RECT 45.650 124.475 45.865 124.525 ;
        RECT 43.730 124.025 44.605 124.355 ;
        RECT 44.775 124.025 45.525 124.355 ;
        RECT 43.730 123.565 43.900 124.025 ;
        RECT 44.775 123.855 44.975 124.025 ;
        RECT 45.695 123.895 45.865 124.475 ;
        RECT 47.110 124.525 47.695 124.715 ;
        RECT 46.050 124.025 46.345 124.355 ;
        RECT 46.525 124.025 46.940 124.355 ;
        RECT 45.640 123.855 45.865 123.895 ;
        RECT 42.540 123.395 42.945 123.565 ;
        RECT 43.115 123.395 43.900 123.565 ;
        RECT 44.175 123.115 44.385 123.645 ;
        RECT 44.645 123.330 44.975 123.855 ;
        RECT 45.485 123.770 45.865 123.855 ;
        RECT 45.145 123.115 45.315 123.725 ;
        RECT 45.485 123.335 45.815 123.770 ;
        RECT 46.045 123.115 46.345 123.845 ;
        RECT 46.525 123.405 46.755 124.025 ;
        RECT 47.110 123.855 47.285 124.525 ;
        RECT 47.875 124.390 48.135 124.840 ;
        RECT 48.305 124.740 48.635 124.985 ;
        RECT 48.805 124.665 49.560 124.915 ;
        RECT 49.730 124.795 50.005 125.495 ;
        RECT 50.175 125.110 50.780 125.665 ;
        RECT 50.955 125.155 51.435 125.495 ;
        RECT 51.605 125.120 51.860 125.665 ;
        RECT 50.175 125.010 50.790 125.110 ;
        RECT 50.605 124.985 50.790 125.010 ;
        RECT 48.790 124.630 49.560 124.665 ;
        RECT 48.775 124.620 49.560 124.630 ;
        RECT 48.770 124.605 49.665 124.620 ;
        RECT 48.750 124.590 49.665 124.605 ;
        RECT 48.730 124.580 49.665 124.590 ;
        RECT 48.705 124.570 49.665 124.580 ;
        RECT 48.635 124.540 49.665 124.570 ;
        RECT 48.615 124.510 49.665 124.540 ;
        RECT 48.595 124.480 49.665 124.510 ;
        RECT 48.565 124.455 49.665 124.480 ;
        RECT 48.530 124.420 49.665 124.455 ;
        RECT 48.500 124.415 49.665 124.420 ;
        RECT 48.500 124.410 48.890 124.415 ;
        RECT 48.500 124.400 48.865 124.410 ;
        RECT 48.500 124.395 48.850 124.400 ;
        RECT 48.500 124.390 48.835 124.395 ;
        RECT 47.875 124.385 48.835 124.390 ;
        RECT 47.875 124.375 48.825 124.385 ;
        RECT 47.875 124.370 48.815 124.375 ;
        RECT 47.875 124.360 48.805 124.370 ;
        RECT 46.955 123.675 47.285 123.855 ;
        RECT 47.455 123.705 47.695 124.355 ;
        RECT 47.875 124.350 48.800 124.360 ;
        RECT 47.875 124.345 48.795 124.350 ;
        RECT 47.875 124.330 48.785 124.345 ;
        RECT 47.875 124.315 48.780 124.330 ;
        RECT 47.875 124.290 48.770 124.315 ;
        RECT 47.875 124.220 48.765 124.290 ;
        RECT 46.955 123.295 47.180 123.675 ;
        RECT 47.875 123.665 48.425 124.050 ;
        RECT 47.350 123.115 47.680 123.505 ;
        RECT 48.595 123.495 48.765 124.220 ;
        RECT 47.875 123.325 48.765 123.495 ;
        RECT 48.935 123.820 49.265 124.245 ;
        RECT 49.435 124.020 49.665 124.415 ;
        RECT 48.935 123.335 49.155 123.820 ;
        RECT 49.835 123.765 50.005 124.795 ;
        RECT 50.175 124.390 50.435 124.840 ;
        RECT 50.605 124.740 50.935 124.985 ;
        RECT 51.105 124.665 51.860 124.915 ;
        RECT 52.030 124.795 52.305 125.495 ;
        RECT 51.090 124.630 51.860 124.665 ;
        RECT 51.075 124.620 51.860 124.630 ;
        RECT 51.070 124.605 51.965 124.620 ;
        RECT 51.050 124.590 51.965 124.605 ;
        RECT 51.030 124.580 51.965 124.590 ;
        RECT 51.005 124.570 51.965 124.580 ;
        RECT 50.935 124.540 51.965 124.570 ;
        RECT 50.915 124.510 51.965 124.540 ;
        RECT 50.895 124.480 51.965 124.510 ;
        RECT 50.865 124.455 51.965 124.480 ;
        RECT 50.830 124.420 51.965 124.455 ;
        RECT 50.800 124.415 51.965 124.420 ;
        RECT 50.800 124.410 51.190 124.415 ;
        RECT 50.800 124.400 51.165 124.410 ;
        RECT 50.800 124.395 51.150 124.400 ;
        RECT 50.800 124.390 51.135 124.395 ;
        RECT 50.175 124.385 51.135 124.390 ;
        RECT 50.175 124.375 51.125 124.385 ;
        RECT 50.175 124.370 51.115 124.375 ;
        RECT 50.175 124.360 51.105 124.370 ;
        RECT 50.175 124.350 51.100 124.360 ;
        RECT 50.175 124.345 51.095 124.350 ;
        RECT 50.175 124.330 51.085 124.345 ;
        RECT 50.175 124.315 51.080 124.330 ;
        RECT 50.175 124.290 51.070 124.315 ;
        RECT 50.175 124.220 51.065 124.290 ;
        RECT 49.325 123.115 49.575 123.655 ;
        RECT 49.745 123.285 50.005 123.765 ;
        RECT 50.175 123.665 50.725 124.050 ;
        RECT 50.895 123.495 51.065 124.220 ;
        RECT 50.175 123.325 51.065 123.495 ;
        RECT 51.235 123.820 51.565 124.245 ;
        RECT 51.735 124.020 51.965 124.415 ;
        RECT 51.235 123.335 51.455 123.820 ;
        RECT 52.135 123.765 52.305 124.795 ;
        RECT 52.485 124.695 52.815 125.480 ;
        RECT 52.485 124.525 53.165 124.695 ;
        RECT 53.345 124.525 53.675 125.665 ;
        RECT 53.855 125.110 54.460 125.665 ;
        RECT 54.635 125.155 55.115 125.495 ;
        RECT 55.285 125.120 55.540 125.665 ;
        RECT 53.855 125.010 54.470 125.110 ;
        RECT 54.285 124.985 54.470 125.010 ;
        RECT 52.475 124.105 52.825 124.355 ;
        RECT 52.995 123.925 53.165 124.525 ;
        RECT 53.855 124.390 54.115 124.840 ;
        RECT 54.285 124.740 54.615 124.985 ;
        RECT 54.785 124.665 55.540 124.915 ;
        RECT 55.710 124.795 55.985 125.495 ;
        RECT 54.770 124.630 55.540 124.665 ;
        RECT 54.755 124.620 55.540 124.630 ;
        RECT 54.750 124.605 55.645 124.620 ;
        RECT 54.730 124.590 55.645 124.605 ;
        RECT 54.710 124.580 55.645 124.590 ;
        RECT 54.685 124.570 55.645 124.580 ;
        RECT 54.615 124.540 55.645 124.570 ;
        RECT 54.595 124.510 55.645 124.540 ;
        RECT 54.575 124.480 55.645 124.510 ;
        RECT 54.545 124.455 55.645 124.480 ;
        RECT 54.510 124.420 55.645 124.455 ;
        RECT 54.480 124.415 55.645 124.420 ;
        RECT 54.480 124.410 54.870 124.415 ;
        RECT 54.480 124.400 54.845 124.410 ;
        RECT 54.480 124.395 54.830 124.400 ;
        RECT 54.480 124.390 54.815 124.395 ;
        RECT 53.855 124.385 54.815 124.390 ;
        RECT 53.855 124.375 54.805 124.385 ;
        RECT 53.855 124.370 54.795 124.375 ;
        RECT 53.855 124.360 54.785 124.370 ;
        RECT 53.335 124.105 53.685 124.355 ;
        RECT 53.855 124.350 54.780 124.360 ;
        RECT 53.855 124.345 54.775 124.350 ;
        RECT 53.855 124.330 54.765 124.345 ;
        RECT 53.855 124.315 54.760 124.330 ;
        RECT 53.855 124.290 54.750 124.315 ;
        RECT 53.855 124.220 54.745 124.290 ;
        RECT 51.625 123.115 51.875 123.655 ;
        RECT 52.045 123.285 52.305 123.765 ;
        RECT 52.495 123.115 52.735 123.925 ;
        RECT 52.905 123.285 53.235 123.925 ;
        RECT 53.405 123.115 53.675 123.925 ;
        RECT 53.855 123.665 54.405 124.050 ;
        RECT 54.575 123.495 54.745 124.220 ;
        RECT 53.855 123.325 54.745 123.495 ;
        RECT 54.915 123.820 55.245 124.245 ;
        RECT 55.415 124.020 55.645 124.415 ;
        RECT 54.915 123.795 55.165 123.820 ;
        RECT 54.915 123.335 55.135 123.795 ;
        RECT 55.815 123.765 55.985 124.795 ;
        RECT 56.155 124.500 56.445 125.665 ;
        RECT 56.615 125.230 61.960 125.665 ;
        RECT 62.135 125.230 67.480 125.665 ;
        RECT 55.305 123.115 55.555 123.655 ;
        RECT 55.725 123.285 55.985 123.765 ;
        RECT 56.155 123.115 56.445 123.840 ;
        RECT 58.200 123.660 58.540 124.490 ;
        RECT 60.020 123.980 60.370 125.230 ;
        RECT 63.720 123.660 64.060 124.490 ;
        RECT 65.540 123.980 65.890 125.230 ;
        RECT 67.655 124.575 71.165 125.665 ;
        RECT 67.655 123.885 69.305 124.405 ;
        RECT 69.475 124.055 71.165 124.575 ;
        RECT 71.830 124.875 72.365 125.495 ;
        RECT 56.615 123.115 61.960 123.660 ;
        RECT 62.135 123.115 67.480 123.660 ;
        RECT 67.655 123.115 71.165 123.885 ;
        RECT 71.830 123.855 72.145 124.875 ;
        RECT 72.535 124.865 72.865 125.665 ;
        RECT 73.350 124.695 73.740 124.870 ;
        RECT 72.315 124.525 73.740 124.695 ;
        RECT 74.280 124.695 74.670 124.870 ;
        RECT 75.155 124.865 75.485 125.665 ;
        RECT 75.655 124.875 76.190 125.495 ;
        RECT 74.280 124.525 75.705 124.695 ;
        RECT 72.315 124.025 72.485 124.525 ;
        RECT 71.830 123.285 72.445 123.855 ;
        RECT 72.735 123.795 73.000 124.355 ;
        RECT 73.170 123.625 73.340 124.525 ;
        RECT 73.510 123.795 73.865 124.355 ;
        RECT 74.155 123.795 74.510 124.355 ;
        RECT 74.680 123.625 74.850 124.525 ;
        RECT 75.020 123.795 75.285 124.355 ;
        RECT 75.535 124.025 75.705 124.525 ;
        RECT 75.875 123.855 76.190 124.875 ;
        RECT 72.615 123.115 72.830 123.625 ;
        RECT 73.060 123.295 73.340 123.625 ;
        RECT 73.520 123.115 73.760 123.625 ;
        RECT 74.260 123.115 74.500 123.625 ;
        RECT 74.680 123.295 74.960 123.625 ;
        RECT 75.190 123.115 75.405 123.625 ;
        RECT 75.575 123.285 76.190 123.855 ;
        RECT 76.395 124.945 76.855 125.495 ;
        RECT 77.045 124.945 77.375 125.665 ;
        RECT 76.395 123.575 76.645 124.945 ;
        RECT 77.575 124.775 77.875 125.325 ;
        RECT 78.045 124.995 78.325 125.665 ;
        RECT 76.935 124.605 77.875 124.775 ;
        RECT 76.935 124.355 77.105 124.605 ;
        RECT 78.245 124.355 78.510 124.715 ;
        RECT 78.695 124.575 81.285 125.665 ;
        RECT 76.815 124.025 77.105 124.355 ;
        RECT 77.275 124.105 77.615 124.355 ;
        RECT 77.835 124.105 78.510 124.355 ;
        RECT 76.935 123.935 77.105 124.025 ;
        RECT 76.935 123.745 78.325 123.935 ;
        RECT 76.395 123.285 76.955 123.575 ;
        RECT 77.125 123.115 77.375 123.575 ;
        RECT 77.995 123.385 78.325 123.745 ;
        RECT 78.695 123.885 79.905 124.405 ;
        RECT 80.075 124.055 81.285 124.575 ;
        RECT 81.915 124.500 82.205 125.665 ;
        RECT 82.835 124.525 83.095 125.665 ;
        RECT 83.335 125.155 84.950 125.485 ;
        RECT 83.345 124.355 83.515 124.915 ;
        RECT 83.775 124.815 84.950 124.985 ;
        RECT 85.120 124.865 85.400 125.665 ;
        RECT 83.775 124.525 84.105 124.815 ;
        RECT 84.780 124.695 84.950 124.815 ;
        RECT 84.275 124.355 84.520 124.645 ;
        RECT 84.780 124.525 85.440 124.695 ;
        RECT 85.610 124.525 85.885 125.495 ;
        RECT 86.055 125.110 86.660 125.665 ;
        RECT 86.835 125.155 87.315 125.495 ;
        RECT 87.485 125.120 87.740 125.665 ;
        RECT 86.055 125.010 86.670 125.110 ;
        RECT 86.485 124.985 86.670 125.010 ;
        RECT 85.270 124.355 85.440 124.525 ;
        RECT 82.840 124.105 83.175 124.355 ;
        RECT 83.345 124.025 84.060 124.355 ;
        RECT 84.275 124.025 85.100 124.355 ;
        RECT 85.270 124.025 85.545 124.355 ;
        RECT 83.345 123.935 83.595 124.025 ;
        RECT 78.695 123.115 81.285 123.885 ;
        RECT 81.915 123.115 82.205 123.840 ;
        RECT 82.835 123.115 83.095 123.935 ;
        RECT 83.265 123.515 83.595 123.935 ;
        RECT 85.270 123.855 85.440 124.025 ;
        RECT 83.775 123.685 85.440 123.855 ;
        RECT 85.715 123.790 85.885 124.525 ;
        RECT 86.055 124.390 86.315 124.840 ;
        RECT 86.485 124.740 86.815 124.985 ;
        RECT 86.985 124.665 87.740 124.915 ;
        RECT 87.910 124.795 88.185 125.495 ;
        RECT 88.445 124.995 88.615 125.495 ;
        RECT 88.785 125.165 89.115 125.665 ;
        RECT 88.445 124.825 89.110 124.995 ;
        RECT 86.970 124.630 87.740 124.665 ;
        RECT 86.955 124.620 87.740 124.630 ;
        RECT 86.950 124.605 87.845 124.620 ;
        RECT 86.930 124.590 87.845 124.605 ;
        RECT 86.910 124.580 87.845 124.590 ;
        RECT 86.885 124.570 87.845 124.580 ;
        RECT 86.815 124.540 87.845 124.570 ;
        RECT 86.795 124.510 87.845 124.540 ;
        RECT 86.775 124.480 87.845 124.510 ;
        RECT 86.745 124.455 87.845 124.480 ;
        RECT 86.710 124.420 87.845 124.455 ;
        RECT 86.680 124.415 87.845 124.420 ;
        RECT 86.680 124.410 87.070 124.415 ;
        RECT 86.680 124.400 87.045 124.410 ;
        RECT 86.680 124.395 87.030 124.400 ;
        RECT 86.680 124.390 87.015 124.395 ;
        RECT 86.055 124.385 87.015 124.390 ;
        RECT 86.055 124.375 87.005 124.385 ;
        RECT 86.055 124.370 86.995 124.375 ;
        RECT 86.055 124.360 86.985 124.370 ;
        RECT 86.055 124.350 86.980 124.360 ;
        RECT 86.055 124.345 86.975 124.350 ;
        RECT 86.055 124.330 86.965 124.345 ;
        RECT 86.055 124.315 86.960 124.330 ;
        RECT 86.055 124.290 86.950 124.315 ;
        RECT 86.055 124.220 86.945 124.290 ;
        RECT 83.775 123.285 84.035 123.685 ;
        RECT 84.205 123.115 84.535 123.515 ;
        RECT 84.705 123.335 84.875 123.685 ;
        RECT 85.045 123.115 85.420 123.515 ;
        RECT 85.610 123.445 85.885 123.790 ;
        RECT 86.055 123.665 86.605 124.050 ;
        RECT 86.775 123.495 86.945 124.220 ;
        RECT 86.055 123.325 86.945 123.495 ;
        RECT 87.115 123.820 87.445 124.245 ;
        RECT 87.615 124.020 87.845 124.415 ;
        RECT 87.115 123.335 87.335 123.820 ;
        RECT 88.015 123.765 88.185 124.795 ;
        RECT 88.360 124.005 88.710 124.655 ;
        RECT 88.880 123.835 89.110 124.825 ;
        RECT 87.505 123.115 87.755 123.655 ;
        RECT 87.925 123.285 88.185 123.765 ;
        RECT 88.445 123.665 89.110 123.835 ;
        RECT 88.445 123.375 88.615 123.665 ;
        RECT 88.785 123.115 89.115 123.495 ;
        RECT 89.285 123.375 89.470 125.495 ;
        RECT 89.710 125.205 89.975 125.665 ;
        RECT 90.145 125.070 90.395 125.495 ;
        RECT 90.605 125.220 91.710 125.390 ;
        RECT 90.090 124.940 90.395 125.070 ;
        RECT 89.640 123.745 89.920 124.695 ;
        RECT 90.090 123.835 90.260 124.940 ;
        RECT 90.430 124.155 90.670 124.750 ;
        RECT 90.840 124.685 91.370 125.050 ;
        RECT 90.840 123.985 91.010 124.685 ;
        RECT 91.540 124.605 91.710 125.220 ;
        RECT 91.880 124.865 92.050 125.665 ;
        RECT 92.220 125.165 92.470 125.495 ;
        RECT 92.695 125.195 93.580 125.365 ;
        RECT 91.540 124.515 92.050 124.605 ;
        RECT 90.090 123.705 90.315 123.835 ;
        RECT 90.485 123.765 91.010 123.985 ;
        RECT 91.180 124.345 92.050 124.515 ;
        RECT 89.725 123.115 89.975 123.575 ;
        RECT 90.145 123.565 90.315 123.705 ;
        RECT 91.180 123.565 91.350 124.345 ;
        RECT 91.880 124.275 92.050 124.345 ;
        RECT 91.560 124.095 91.760 124.125 ;
        RECT 92.220 124.095 92.390 125.165 ;
        RECT 92.560 124.275 92.750 124.995 ;
        RECT 91.560 123.795 92.390 124.095 ;
        RECT 92.920 124.065 93.240 125.025 ;
        RECT 90.145 123.395 90.480 123.565 ;
        RECT 90.675 123.395 91.350 123.565 ;
        RECT 91.670 123.115 92.040 123.615 ;
        RECT 92.220 123.565 92.390 123.795 ;
        RECT 92.775 123.735 93.240 124.065 ;
        RECT 93.410 124.355 93.580 125.195 ;
        RECT 93.760 125.165 94.075 125.665 ;
        RECT 94.305 124.935 94.645 125.495 ;
        RECT 93.750 124.560 94.645 124.935 ;
        RECT 94.815 124.655 94.985 125.665 ;
        RECT 94.455 124.355 94.645 124.560 ;
        RECT 95.155 124.605 95.485 125.450 ;
        RECT 95.655 124.750 95.825 125.665 ;
        RECT 95.155 124.525 95.545 124.605 ;
        RECT 96.175 124.575 97.845 125.665 ;
        RECT 98.565 124.995 98.735 125.495 ;
        RECT 98.905 125.165 99.235 125.665 ;
        RECT 98.565 124.825 99.230 124.995 ;
        RECT 95.330 124.475 95.545 124.525 ;
        RECT 93.410 124.025 94.285 124.355 ;
        RECT 94.455 124.025 95.205 124.355 ;
        RECT 93.410 123.565 93.580 124.025 ;
        RECT 94.455 123.855 94.655 124.025 ;
        RECT 95.375 123.895 95.545 124.475 ;
        RECT 95.320 123.855 95.545 123.895 ;
        RECT 92.220 123.395 92.625 123.565 ;
        RECT 92.795 123.395 93.580 123.565 ;
        RECT 93.855 123.115 94.065 123.645 ;
        RECT 94.325 123.330 94.655 123.855 ;
        RECT 95.165 123.770 95.545 123.855 ;
        RECT 96.175 123.885 96.925 124.405 ;
        RECT 97.095 124.055 97.845 124.575 ;
        RECT 98.480 124.005 98.830 124.655 ;
        RECT 94.825 123.115 94.995 123.725 ;
        RECT 95.165 123.335 95.495 123.770 ;
        RECT 95.665 123.115 95.835 123.630 ;
        RECT 96.175 123.115 97.845 123.885 ;
        RECT 99.000 123.835 99.230 124.825 ;
        RECT 98.565 123.665 99.230 123.835 ;
        RECT 98.565 123.375 98.735 123.665 ;
        RECT 98.905 123.115 99.235 123.495 ;
        RECT 99.405 123.375 99.590 125.495 ;
        RECT 99.830 125.205 100.095 125.665 ;
        RECT 100.265 125.070 100.515 125.495 ;
        RECT 100.725 125.220 101.830 125.390 ;
        RECT 100.210 124.940 100.515 125.070 ;
        RECT 99.760 123.745 100.040 124.695 ;
        RECT 100.210 123.835 100.380 124.940 ;
        RECT 100.550 124.155 100.790 124.750 ;
        RECT 100.960 124.685 101.490 125.050 ;
        RECT 100.960 123.985 101.130 124.685 ;
        RECT 101.660 124.605 101.830 125.220 ;
        RECT 102.000 124.865 102.170 125.665 ;
        RECT 102.340 125.165 102.590 125.495 ;
        RECT 102.815 125.195 103.700 125.365 ;
        RECT 101.660 124.515 102.170 124.605 ;
        RECT 100.210 123.705 100.435 123.835 ;
        RECT 100.605 123.765 101.130 123.985 ;
        RECT 101.300 124.345 102.170 124.515 ;
        RECT 99.845 123.115 100.095 123.575 ;
        RECT 100.265 123.565 100.435 123.705 ;
        RECT 101.300 123.565 101.470 124.345 ;
        RECT 102.000 124.275 102.170 124.345 ;
        RECT 101.680 124.095 101.880 124.125 ;
        RECT 102.340 124.095 102.510 125.165 ;
        RECT 102.680 124.275 102.870 124.995 ;
        RECT 101.680 123.795 102.510 124.095 ;
        RECT 103.040 124.065 103.360 125.025 ;
        RECT 100.265 123.395 100.600 123.565 ;
        RECT 100.795 123.395 101.470 123.565 ;
        RECT 101.790 123.115 102.160 123.615 ;
        RECT 102.340 123.565 102.510 123.795 ;
        RECT 102.895 123.735 103.360 124.065 ;
        RECT 103.530 124.355 103.700 125.195 ;
        RECT 103.880 125.165 104.195 125.665 ;
        RECT 104.425 124.935 104.765 125.495 ;
        RECT 103.870 124.560 104.765 124.935 ;
        RECT 104.935 124.655 105.105 125.665 ;
        RECT 104.575 124.355 104.765 124.560 ;
        RECT 105.275 124.605 105.605 125.450 ;
        RECT 105.275 124.525 105.665 124.605 ;
        RECT 105.835 124.575 107.505 125.665 ;
        RECT 105.450 124.475 105.665 124.525 ;
        RECT 103.530 124.025 104.405 124.355 ;
        RECT 104.575 124.025 105.325 124.355 ;
        RECT 103.530 123.565 103.700 124.025 ;
        RECT 104.575 123.855 104.775 124.025 ;
        RECT 105.495 123.895 105.665 124.475 ;
        RECT 105.440 123.855 105.665 123.895 ;
        RECT 102.340 123.395 102.745 123.565 ;
        RECT 102.915 123.395 103.700 123.565 ;
        RECT 103.975 123.115 104.185 123.645 ;
        RECT 104.445 123.330 104.775 123.855 ;
        RECT 105.285 123.770 105.665 123.855 ;
        RECT 105.835 123.885 106.585 124.405 ;
        RECT 106.755 124.055 107.505 124.575 ;
        RECT 107.675 124.500 107.965 125.665 ;
        RECT 108.135 124.525 108.520 125.495 ;
        RECT 108.690 125.205 109.015 125.665 ;
        RECT 109.535 125.035 109.815 125.495 ;
        RECT 108.690 124.815 109.815 125.035 ;
        RECT 104.945 123.115 105.115 123.725 ;
        RECT 105.285 123.335 105.615 123.770 ;
        RECT 105.835 123.115 107.505 123.885 ;
        RECT 108.135 123.855 108.415 124.525 ;
        RECT 108.690 124.355 109.140 124.815 ;
        RECT 110.005 124.645 110.405 125.495 ;
        RECT 110.805 125.205 111.075 125.665 ;
        RECT 111.245 125.035 111.530 125.495 ;
        RECT 108.585 124.025 109.140 124.355 ;
        RECT 109.310 124.085 110.405 124.645 ;
        RECT 108.690 123.915 109.140 124.025 ;
        RECT 107.675 123.115 107.965 123.840 ;
        RECT 108.135 123.285 108.520 123.855 ;
        RECT 108.690 123.745 109.815 123.915 ;
        RECT 108.690 123.115 109.015 123.575 ;
        RECT 109.535 123.285 109.815 123.745 ;
        RECT 110.005 123.285 110.405 124.085 ;
        RECT 110.575 124.815 111.530 125.035 ;
        RECT 110.575 123.915 110.785 124.815 ;
        RECT 110.955 124.085 111.645 124.645 ;
        RECT 111.815 124.525 112.155 125.495 ;
        RECT 112.325 124.525 112.495 125.665 ;
        RECT 112.765 124.865 113.015 125.665 ;
        RECT 113.660 124.695 113.990 125.495 ;
        RECT 114.290 124.865 114.620 125.665 ;
        RECT 114.790 124.695 115.120 125.495 ;
        RECT 112.685 124.525 115.120 124.695 ;
        RECT 115.500 124.715 115.765 125.485 ;
        RECT 115.935 124.945 116.265 125.665 ;
        RECT 116.455 125.125 116.715 125.485 ;
        RECT 116.885 125.295 117.215 125.665 ;
        RECT 117.385 125.125 117.645 125.485 ;
        RECT 116.455 124.895 117.645 125.125 ;
        RECT 118.215 124.715 118.505 125.485 ;
        RECT 111.815 123.915 111.990 124.525 ;
        RECT 112.685 124.275 112.855 124.525 ;
        RECT 112.160 124.105 112.855 124.275 ;
        RECT 113.030 124.105 113.450 124.305 ;
        RECT 113.620 124.105 113.950 124.305 ;
        RECT 114.120 124.105 114.450 124.305 ;
        RECT 110.575 123.745 111.530 123.915 ;
        RECT 110.805 123.115 111.075 123.575 ;
        RECT 111.245 123.285 111.530 123.745 ;
        RECT 111.815 123.285 112.155 123.915 ;
        RECT 112.325 123.115 112.575 123.915 ;
        RECT 112.765 123.765 113.990 123.935 ;
        RECT 112.765 123.285 113.095 123.765 ;
        RECT 113.265 123.115 113.490 123.575 ;
        RECT 113.660 123.285 113.990 123.765 ;
        RECT 114.620 123.895 114.790 124.525 ;
        RECT 114.975 124.105 115.325 124.355 ;
        RECT 114.620 123.285 115.120 123.895 ;
        RECT 115.500 123.295 115.835 124.715 ;
        RECT 116.010 124.535 118.505 124.715 ;
        RECT 118.715 124.575 120.385 125.665 ;
        RECT 116.010 123.845 116.235 124.535 ;
        RECT 116.435 124.025 116.715 124.355 ;
        RECT 116.895 124.025 117.470 124.355 ;
        RECT 117.650 124.025 118.085 124.355 ;
        RECT 118.265 124.025 118.535 124.355 ;
        RECT 118.715 123.885 119.465 124.405 ;
        RECT 119.635 124.055 120.385 124.575 ;
        RECT 120.555 124.525 120.895 125.495 ;
        RECT 121.065 124.525 121.235 125.665 ;
        RECT 121.505 124.865 121.755 125.665 ;
        RECT 122.400 124.695 122.730 125.495 ;
        RECT 123.030 124.865 123.360 125.665 ;
        RECT 123.530 124.695 123.860 125.495 ;
        RECT 121.425 124.525 123.860 124.695 ;
        RECT 124.270 124.875 124.805 125.495 ;
        RECT 120.555 123.915 120.730 124.525 ;
        RECT 121.425 124.275 121.595 124.525 ;
        RECT 120.900 124.105 121.595 124.275 ;
        RECT 121.770 124.105 122.190 124.305 ;
        RECT 122.360 124.105 122.690 124.305 ;
        RECT 122.860 124.105 123.190 124.305 ;
        RECT 116.010 123.655 118.495 123.845 ;
        RECT 116.015 123.115 116.760 123.485 ;
        RECT 117.325 123.295 117.580 123.655 ;
        RECT 117.760 123.115 118.090 123.485 ;
        RECT 118.270 123.295 118.495 123.655 ;
        RECT 118.715 123.115 120.385 123.885 ;
        RECT 120.555 123.285 120.895 123.915 ;
        RECT 121.065 123.115 121.315 123.915 ;
        RECT 121.505 123.765 122.730 123.935 ;
        RECT 121.505 123.285 121.835 123.765 ;
        RECT 122.005 123.115 122.230 123.575 ;
        RECT 122.400 123.285 122.730 123.765 ;
        RECT 123.360 123.895 123.530 124.525 ;
        RECT 123.715 124.105 124.065 124.355 ;
        RECT 123.360 123.285 123.860 123.895 ;
        RECT 124.270 123.855 124.585 124.875 ;
        RECT 124.975 124.865 125.305 125.665 ;
        RECT 125.790 124.695 126.180 124.870 ;
        RECT 124.755 124.525 126.180 124.695 ;
        RECT 126.535 124.575 129.125 125.665 ;
        RECT 124.755 124.025 124.925 124.525 ;
        RECT 124.270 123.285 124.885 123.855 ;
        RECT 125.175 123.795 125.440 124.355 ;
        RECT 125.610 123.625 125.780 124.525 ;
        RECT 125.950 123.795 126.305 124.355 ;
        RECT 126.535 123.885 127.745 124.405 ;
        RECT 127.915 124.055 129.125 124.575 ;
        RECT 129.960 124.695 130.290 125.495 ;
        RECT 130.460 124.865 130.790 125.665 ;
        RECT 131.090 124.695 131.420 125.495 ;
        RECT 132.065 124.865 132.315 125.665 ;
        RECT 129.960 124.525 132.395 124.695 ;
        RECT 132.585 124.525 132.755 125.665 ;
        RECT 132.925 124.525 133.265 125.495 ;
        RECT 129.755 124.105 130.105 124.355 ;
        RECT 130.290 123.895 130.460 124.525 ;
        RECT 130.630 124.105 130.960 124.305 ;
        RECT 131.130 124.105 131.460 124.305 ;
        RECT 131.630 124.105 132.050 124.305 ;
        RECT 132.225 124.275 132.395 124.525 ;
        RECT 133.035 124.475 133.265 124.525 ;
        RECT 133.435 124.500 133.725 125.665 ;
        RECT 133.930 124.875 134.465 125.495 ;
        RECT 132.225 124.105 132.920 124.275 ;
        RECT 125.055 123.115 125.270 123.625 ;
        RECT 125.500 123.295 125.780 123.625 ;
        RECT 125.960 123.115 126.200 123.625 ;
        RECT 126.535 123.115 129.125 123.885 ;
        RECT 129.960 123.285 130.460 123.895 ;
        RECT 131.090 123.765 132.315 123.935 ;
        RECT 133.090 123.915 133.265 124.475 ;
        RECT 131.090 123.285 131.420 123.765 ;
        RECT 131.590 123.115 131.815 123.575 ;
        RECT 131.985 123.285 132.315 123.765 ;
        RECT 132.505 123.115 132.755 123.915 ;
        RECT 132.925 123.285 133.265 123.915 ;
        RECT 133.930 123.855 134.245 124.875 ;
        RECT 134.635 124.865 134.965 125.665 ;
        RECT 136.230 124.875 136.765 125.495 ;
        RECT 135.450 124.695 135.840 124.870 ;
        RECT 134.415 124.525 135.840 124.695 ;
        RECT 134.415 124.025 134.585 124.525 ;
        RECT 133.435 123.115 133.725 123.840 ;
        RECT 133.930 123.285 134.545 123.855 ;
        RECT 134.835 123.795 135.100 124.355 ;
        RECT 135.270 123.625 135.440 124.525 ;
        RECT 135.610 123.795 135.965 124.355 ;
        RECT 136.230 123.855 136.545 124.875 ;
        RECT 136.935 124.865 137.265 125.665 ;
        RECT 137.750 124.695 138.140 124.870 ;
        RECT 136.715 124.525 138.140 124.695 ;
        RECT 138.495 124.575 139.705 125.665 ;
        RECT 136.715 124.025 136.885 124.525 ;
        RECT 134.715 123.115 134.930 123.625 ;
        RECT 135.160 123.295 135.440 123.625 ;
        RECT 135.620 123.115 135.860 123.625 ;
        RECT 136.230 123.285 136.845 123.855 ;
        RECT 137.135 123.795 137.400 124.355 ;
        RECT 137.570 123.625 137.740 124.525 ;
        RECT 137.910 123.795 138.265 124.355 ;
        RECT 138.495 123.865 139.015 124.405 ;
        RECT 139.185 124.035 139.705 124.575 ;
        RECT 139.965 124.735 140.135 125.495 ;
        RECT 140.350 124.905 140.680 125.665 ;
        RECT 139.965 124.565 140.680 124.735 ;
        RECT 140.850 124.590 141.105 125.495 ;
        RECT 139.875 124.015 140.230 124.385 ;
        RECT 140.510 124.355 140.680 124.565 ;
        RECT 140.510 124.025 140.765 124.355 ;
        RECT 137.015 123.115 137.230 123.625 ;
        RECT 137.460 123.295 137.740 123.625 ;
        RECT 137.920 123.115 138.160 123.625 ;
        RECT 138.495 123.115 139.705 123.865 ;
        RECT 140.510 123.835 140.680 124.025 ;
        RECT 140.935 123.860 141.105 124.590 ;
        RECT 141.280 124.515 141.540 125.665 ;
        RECT 141.715 124.575 142.925 125.665 ;
        RECT 141.715 124.035 142.235 124.575 ;
        RECT 139.965 123.665 140.680 123.835 ;
        RECT 139.965 123.285 140.135 123.665 ;
        RECT 140.350 123.115 140.680 123.495 ;
        RECT 140.850 123.285 141.105 123.860 ;
        RECT 141.280 123.115 141.540 123.955 ;
        RECT 142.405 123.865 142.925 124.405 ;
        RECT 141.715 123.115 142.925 123.865 ;
        RECT 17.430 122.945 143.010 123.115 ;
        RECT 17.515 122.195 18.725 122.945 ;
        RECT 18.895 122.400 24.240 122.945 ;
        RECT 17.515 121.655 18.035 122.195 ;
        RECT 18.205 121.485 18.725 122.025 ;
        RECT 20.480 121.570 20.820 122.400 ;
        RECT 24.415 122.175 26.085 122.945 ;
        RECT 26.305 122.290 26.635 122.725 ;
        RECT 26.805 122.335 26.975 122.945 ;
        RECT 26.255 122.205 26.635 122.290 ;
        RECT 27.145 122.205 27.475 122.730 ;
        RECT 27.735 122.415 27.945 122.945 ;
        RECT 28.220 122.495 29.005 122.665 ;
        RECT 29.175 122.495 29.580 122.665 ;
        RECT 17.515 120.395 18.725 121.485 ;
        RECT 22.300 120.830 22.650 122.080 ;
        RECT 24.415 121.655 25.165 122.175 ;
        RECT 26.255 122.165 26.480 122.205 ;
        RECT 25.335 121.485 26.085 122.005 ;
        RECT 18.895 120.395 24.240 120.830 ;
        RECT 24.415 120.395 26.085 121.485 ;
        RECT 26.255 121.585 26.425 122.165 ;
        RECT 27.145 122.035 27.345 122.205 ;
        RECT 28.220 122.035 28.390 122.495 ;
        RECT 26.595 121.705 27.345 122.035 ;
        RECT 27.515 121.705 28.390 122.035 ;
        RECT 26.255 121.535 26.470 121.585 ;
        RECT 26.255 121.455 26.645 121.535 ;
        RECT 26.315 120.610 26.645 121.455 ;
        RECT 27.155 121.500 27.345 121.705 ;
        RECT 26.815 120.395 26.985 121.405 ;
        RECT 27.155 121.125 28.050 121.500 ;
        RECT 27.155 120.565 27.495 121.125 ;
        RECT 27.725 120.395 28.040 120.895 ;
        RECT 28.220 120.865 28.390 121.705 ;
        RECT 28.560 121.995 29.025 122.325 ;
        RECT 29.410 122.265 29.580 122.495 ;
        RECT 29.760 122.445 30.130 122.945 ;
        RECT 30.450 122.495 31.125 122.665 ;
        RECT 31.320 122.495 31.655 122.665 ;
        RECT 28.560 121.035 28.880 121.995 ;
        RECT 29.410 121.965 30.240 122.265 ;
        RECT 29.050 121.065 29.240 121.785 ;
        RECT 29.410 120.895 29.580 121.965 ;
        RECT 30.040 121.935 30.240 121.965 ;
        RECT 29.750 121.715 29.920 121.785 ;
        RECT 30.450 121.715 30.620 122.495 ;
        RECT 31.485 122.355 31.655 122.495 ;
        RECT 31.825 122.485 32.075 122.945 ;
        RECT 29.750 121.545 30.620 121.715 ;
        RECT 30.790 122.075 31.315 122.295 ;
        RECT 31.485 122.225 31.710 122.355 ;
        RECT 29.750 121.455 30.260 121.545 ;
        RECT 28.220 120.695 29.105 120.865 ;
        RECT 29.330 120.565 29.580 120.895 ;
        RECT 29.750 120.395 29.920 121.195 ;
        RECT 30.090 120.840 30.260 121.455 ;
        RECT 30.790 121.375 30.960 122.075 ;
        RECT 30.430 121.010 30.960 121.375 ;
        RECT 31.130 121.310 31.370 121.905 ;
        RECT 31.540 121.120 31.710 122.225 ;
        RECT 31.880 121.365 32.160 122.315 ;
        RECT 31.405 120.990 31.710 121.120 ;
        RECT 30.090 120.670 31.195 120.840 ;
        RECT 31.405 120.565 31.655 120.990 ;
        RECT 31.825 120.395 32.090 120.855 ;
        RECT 32.330 120.565 32.515 122.685 ;
        RECT 32.685 122.565 33.015 122.945 ;
        RECT 33.185 122.395 33.355 122.685 ;
        RECT 33.615 122.400 38.960 122.945 ;
        RECT 32.690 122.225 33.355 122.395 ;
        RECT 32.690 121.235 32.920 122.225 ;
        RECT 33.090 121.405 33.440 122.055 ;
        RECT 35.200 121.570 35.540 122.400 ;
        RECT 39.135 122.295 39.395 122.775 ;
        RECT 39.565 122.405 39.815 122.945 ;
        RECT 32.690 121.065 33.355 121.235 ;
        RECT 32.685 120.395 33.015 120.895 ;
        RECT 33.185 120.565 33.355 121.065 ;
        RECT 37.020 120.830 37.370 122.080 ;
        RECT 39.135 121.265 39.305 122.295 ;
        RECT 39.985 122.265 40.205 122.725 ;
        RECT 39.955 122.240 40.205 122.265 ;
        RECT 39.475 121.645 39.705 122.040 ;
        RECT 39.875 121.815 40.205 122.240 ;
        RECT 40.375 122.565 41.265 122.735 ;
        RECT 40.375 121.840 40.545 122.565 ;
        RECT 40.715 122.010 41.265 122.395 ;
        RECT 41.435 122.175 43.105 122.945 ;
        RECT 43.275 122.220 43.565 122.945 ;
        RECT 43.735 122.195 44.945 122.945 ;
        RECT 45.115 122.205 45.580 122.750 ;
        RECT 40.375 121.770 41.265 121.840 ;
        RECT 40.370 121.745 41.265 121.770 ;
        RECT 40.360 121.730 41.265 121.745 ;
        RECT 40.355 121.715 41.265 121.730 ;
        RECT 40.345 121.710 41.265 121.715 ;
        RECT 40.340 121.700 41.265 121.710 ;
        RECT 40.335 121.690 41.265 121.700 ;
        RECT 40.325 121.685 41.265 121.690 ;
        RECT 40.315 121.675 41.265 121.685 ;
        RECT 40.305 121.670 41.265 121.675 ;
        RECT 40.305 121.665 40.640 121.670 ;
        RECT 40.290 121.660 40.640 121.665 ;
        RECT 40.275 121.650 40.640 121.660 ;
        RECT 40.250 121.645 40.640 121.650 ;
        RECT 39.475 121.640 40.640 121.645 ;
        RECT 39.475 121.605 40.610 121.640 ;
        RECT 39.475 121.580 40.575 121.605 ;
        RECT 39.475 121.550 40.545 121.580 ;
        RECT 39.475 121.520 40.525 121.550 ;
        RECT 39.475 121.490 40.505 121.520 ;
        RECT 39.475 121.480 40.435 121.490 ;
        RECT 39.475 121.470 40.410 121.480 ;
        RECT 39.475 121.455 40.390 121.470 ;
        RECT 39.475 121.440 40.370 121.455 ;
        RECT 39.580 121.430 40.365 121.440 ;
        RECT 39.580 121.395 40.350 121.430 ;
        RECT 33.615 120.395 38.960 120.830 ;
        RECT 39.135 120.565 39.410 121.265 ;
        RECT 39.580 121.145 40.335 121.395 ;
        RECT 40.505 121.075 40.835 121.320 ;
        RECT 41.005 121.220 41.265 121.670 ;
        RECT 41.435 121.655 42.185 122.175 ;
        RECT 42.355 121.485 43.105 122.005 ;
        RECT 43.735 121.655 44.255 122.195 ;
        RECT 40.650 121.050 40.835 121.075 ;
        RECT 40.650 120.950 41.265 121.050 ;
        RECT 39.580 120.395 39.835 120.940 ;
        RECT 40.005 120.565 40.485 120.905 ;
        RECT 40.660 120.395 41.265 120.950 ;
        RECT 41.435 120.395 43.105 121.485 ;
        RECT 43.275 120.395 43.565 121.560 ;
        RECT 44.425 121.485 44.945 122.025 ;
        RECT 43.735 120.395 44.945 121.485 ;
        RECT 45.115 121.245 45.285 122.205 ;
        RECT 46.085 122.125 46.255 122.945 ;
        RECT 46.425 122.295 46.755 122.775 ;
        RECT 46.925 122.555 47.275 122.945 ;
        RECT 47.445 122.375 47.675 122.775 ;
        RECT 47.165 122.295 47.675 122.375 ;
        RECT 46.425 122.205 47.675 122.295 ;
        RECT 47.845 122.205 48.165 122.685 ;
        RECT 46.425 122.125 47.335 122.205 ;
        RECT 45.455 121.585 45.700 122.035 ;
        RECT 45.960 121.755 46.655 121.955 ;
        RECT 46.825 121.785 47.425 121.955 ;
        RECT 46.825 121.585 46.995 121.785 ;
        RECT 47.655 121.615 47.825 122.035 ;
        RECT 45.455 121.415 46.995 121.585 ;
        RECT 47.165 121.445 47.825 121.615 ;
        RECT 47.165 121.245 47.335 121.445 ;
        RECT 47.995 121.275 48.165 122.205 ;
        RECT 48.335 122.195 49.545 122.945 ;
        RECT 49.765 122.290 50.095 122.725 ;
        RECT 50.265 122.335 50.435 122.945 ;
        RECT 49.715 122.205 50.095 122.290 ;
        RECT 50.605 122.205 50.935 122.730 ;
        RECT 51.195 122.415 51.405 122.945 ;
        RECT 51.680 122.495 52.465 122.665 ;
        RECT 52.635 122.495 53.040 122.665 ;
        RECT 48.335 121.655 48.855 122.195 ;
        RECT 49.715 122.165 49.940 122.205 ;
        RECT 49.025 121.485 49.545 122.025 ;
        RECT 45.115 121.075 47.335 121.245 ;
        RECT 47.505 121.075 48.165 121.275 ;
        RECT 45.115 120.395 45.415 120.905 ;
        RECT 45.585 120.565 45.915 121.075 ;
        RECT 47.505 120.905 47.675 121.075 ;
        RECT 46.085 120.395 46.715 120.905 ;
        RECT 47.295 120.735 47.675 120.905 ;
        RECT 47.845 120.395 48.145 120.905 ;
        RECT 48.335 120.395 49.545 121.485 ;
        RECT 49.715 121.585 49.885 122.165 ;
        RECT 50.605 122.035 50.805 122.205 ;
        RECT 51.680 122.035 51.850 122.495 ;
        RECT 50.055 121.705 50.805 122.035 ;
        RECT 50.975 121.705 51.850 122.035 ;
        RECT 49.715 121.535 49.930 121.585 ;
        RECT 49.715 121.455 50.105 121.535 ;
        RECT 49.775 120.610 50.105 121.455 ;
        RECT 50.615 121.500 50.805 121.705 ;
        RECT 50.275 120.395 50.445 121.405 ;
        RECT 50.615 121.125 51.510 121.500 ;
        RECT 50.615 120.565 50.955 121.125 ;
        RECT 51.185 120.395 51.500 120.895 ;
        RECT 51.680 120.865 51.850 121.705 ;
        RECT 52.020 121.995 52.485 122.325 ;
        RECT 52.870 122.265 53.040 122.495 ;
        RECT 53.220 122.445 53.590 122.945 ;
        RECT 53.910 122.495 54.585 122.665 ;
        RECT 54.780 122.495 55.115 122.665 ;
        RECT 52.020 121.035 52.340 121.995 ;
        RECT 52.870 121.965 53.700 122.265 ;
        RECT 52.510 121.065 52.700 121.785 ;
        RECT 52.870 120.895 53.040 121.965 ;
        RECT 53.500 121.935 53.700 121.965 ;
        RECT 53.210 121.715 53.380 121.785 ;
        RECT 53.910 121.715 54.080 122.495 ;
        RECT 54.945 122.355 55.115 122.495 ;
        RECT 55.285 122.485 55.535 122.945 ;
        RECT 53.210 121.545 54.080 121.715 ;
        RECT 54.250 122.075 54.775 122.295 ;
        RECT 54.945 122.225 55.170 122.355 ;
        RECT 53.210 121.455 53.720 121.545 ;
        RECT 51.680 120.695 52.565 120.865 ;
        RECT 52.790 120.565 53.040 120.895 ;
        RECT 53.210 120.395 53.380 121.195 ;
        RECT 53.550 120.840 53.720 121.455 ;
        RECT 54.250 121.375 54.420 122.075 ;
        RECT 53.890 121.010 54.420 121.375 ;
        RECT 54.590 121.310 54.830 121.905 ;
        RECT 55.000 121.120 55.170 122.225 ;
        RECT 55.340 121.365 55.620 122.315 ;
        RECT 54.865 120.990 55.170 121.120 ;
        RECT 53.550 120.670 54.655 120.840 ;
        RECT 54.865 120.565 55.115 120.990 ;
        RECT 55.285 120.395 55.550 120.855 ;
        RECT 55.790 120.565 55.975 122.685 ;
        RECT 56.145 122.565 56.475 122.945 ;
        RECT 56.645 122.395 56.815 122.685 ;
        RECT 57.075 122.400 62.420 122.945 ;
        RECT 63.115 122.485 63.360 122.945 ;
        RECT 56.150 122.225 56.815 122.395 ;
        RECT 56.150 121.235 56.380 122.225 ;
        RECT 56.550 121.405 56.900 122.055 ;
        RECT 58.660 121.570 59.000 122.400 ;
        RECT 56.150 121.065 56.815 121.235 ;
        RECT 56.145 120.395 56.475 120.895 ;
        RECT 56.645 120.565 56.815 121.065 ;
        RECT 60.480 120.830 60.830 122.080 ;
        RECT 63.055 121.705 63.370 122.315 ;
        RECT 63.540 121.955 63.790 122.765 ;
        RECT 63.960 122.420 64.220 122.945 ;
        RECT 64.390 122.295 64.650 122.750 ;
        RECT 64.820 122.465 65.080 122.945 ;
        RECT 65.250 122.295 65.510 122.750 ;
        RECT 65.680 122.465 65.940 122.945 ;
        RECT 66.110 122.295 66.370 122.750 ;
        RECT 66.540 122.465 66.800 122.945 ;
        RECT 66.970 122.295 67.230 122.750 ;
        RECT 67.400 122.465 67.700 122.945 ;
        RECT 64.390 122.125 67.700 122.295 ;
        RECT 69.035 122.220 69.325 122.945 ;
        RECT 69.505 122.135 69.775 122.945 ;
        RECT 69.945 122.135 70.275 122.775 ;
        RECT 70.445 122.135 70.685 122.945 ;
        RECT 70.875 122.195 72.085 122.945 ;
        RECT 63.540 121.705 66.560 121.955 ;
        RECT 57.075 120.395 62.420 120.830 ;
        RECT 63.065 120.395 63.360 121.505 ;
        RECT 63.540 120.570 63.790 121.705 ;
        RECT 66.730 121.535 67.700 122.125 ;
        RECT 69.495 121.705 69.845 121.955 ;
        RECT 63.960 120.395 64.220 121.505 ;
        RECT 64.390 121.295 67.700 121.535 ;
        RECT 64.390 120.570 64.650 121.295 ;
        RECT 64.820 120.395 65.080 121.125 ;
        RECT 65.250 120.570 65.510 121.295 ;
        RECT 65.680 120.395 65.940 121.125 ;
        RECT 66.110 120.570 66.370 121.295 ;
        RECT 66.540 120.395 66.800 121.125 ;
        RECT 66.970 120.570 67.230 121.295 ;
        RECT 67.400 120.395 67.695 121.125 ;
        RECT 69.035 120.395 69.325 121.560 ;
        RECT 70.015 121.535 70.185 122.135 ;
        RECT 70.355 121.705 70.705 121.955 ;
        RECT 70.875 121.655 71.395 122.195 ;
        RECT 72.255 122.145 72.950 122.775 ;
        RECT 73.155 122.145 73.465 122.945 ;
        RECT 74.095 122.145 74.405 122.945 ;
        RECT 74.610 122.145 75.305 122.775 ;
        RECT 75.475 122.400 80.820 122.945 ;
        RECT 69.505 120.395 69.835 121.535 ;
        RECT 70.015 121.365 70.695 121.535 ;
        RECT 71.565 121.485 72.085 122.025 ;
        RECT 72.275 121.705 72.610 121.955 ;
        RECT 72.780 121.545 72.950 122.145 ;
        RECT 73.120 121.705 73.455 121.975 ;
        RECT 74.105 121.705 74.440 121.975 ;
        RECT 74.610 121.545 74.780 122.145 ;
        RECT 74.950 121.705 75.285 121.955 ;
        RECT 77.060 121.570 77.400 122.400 ;
        RECT 80.995 122.175 82.665 122.945 ;
        RECT 70.365 120.580 70.695 121.365 ;
        RECT 70.875 120.395 72.085 121.485 ;
        RECT 72.255 120.395 72.515 121.535 ;
        RECT 72.685 120.565 73.015 121.545 ;
        RECT 73.185 120.395 73.465 121.535 ;
        RECT 74.095 120.395 74.375 121.535 ;
        RECT 74.545 120.565 74.875 121.545 ;
        RECT 75.045 120.395 75.305 121.535 ;
        RECT 78.880 120.830 79.230 122.080 ;
        RECT 80.995 121.655 81.745 122.175 ;
        RECT 83.335 122.125 83.565 122.945 ;
        RECT 83.735 122.145 84.065 122.775 ;
        RECT 81.915 121.485 82.665 122.005 ;
        RECT 83.315 121.705 83.645 121.955 ;
        RECT 83.815 121.545 84.065 122.145 ;
        RECT 84.235 122.125 84.445 122.945 ;
        RECT 84.675 122.125 84.935 122.945 ;
        RECT 85.105 122.125 85.435 122.545 ;
        RECT 85.615 122.375 85.875 122.775 ;
        RECT 86.045 122.545 86.375 122.945 ;
        RECT 86.545 122.375 86.715 122.725 ;
        RECT 86.885 122.545 87.260 122.945 ;
        RECT 85.615 122.205 87.280 122.375 ;
        RECT 87.450 122.270 87.725 122.615 ;
        RECT 85.185 122.035 85.435 122.125 ;
        RECT 87.110 122.035 87.280 122.205 ;
        RECT 84.680 121.705 85.015 121.955 ;
        RECT 85.185 121.705 85.900 122.035 ;
        RECT 86.115 121.705 86.940 122.035 ;
        RECT 87.110 121.705 87.385 122.035 ;
        RECT 75.475 120.395 80.820 120.830 ;
        RECT 80.995 120.395 82.665 121.485 ;
        RECT 83.335 120.395 83.565 121.535 ;
        RECT 83.735 120.565 84.065 121.545 ;
        RECT 84.235 120.395 84.445 121.535 ;
        RECT 84.675 120.395 84.935 121.535 ;
        RECT 85.185 121.145 85.355 121.705 ;
        RECT 85.615 121.245 85.945 121.535 ;
        RECT 86.115 121.415 86.360 121.705 ;
        RECT 87.110 121.535 87.280 121.705 ;
        RECT 87.555 121.535 87.725 122.270 ;
        RECT 86.620 121.365 87.280 121.535 ;
        RECT 86.620 121.245 86.790 121.365 ;
        RECT 85.615 121.075 86.790 121.245 ;
        RECT 85.175 120.575 86.790 120.905 ;
        RECT 86.960 120.395 87.240 121.195 ;
        RECT 87.450 120.565 87.725 121.535 ;
        RECT 88.820 122.205 89.075 122.775 ;
        RECT 89.245 122.545 89.575 122.945 ;
        RECT 90.000 122.410 90.530 122.775 ;
        RECT 90.000 122.375 90.175 122.410 ;
        RECT 89.245 122.205 90.175 122.375 ;
        RECT 88.820 121.535 88.990 122.205 ;
        RECT 89.245 122.035 89.415 122.205 ;
        RECT 89.160 121.705 89.415 122.035 ;
        RECT 89.640 121.705 89.835 122.035 ;
        RECT 88.820 120.565 89.155 121.535 ;
        RECT 89.325 120.395 89.495 121.535 ;
        RECT 89.665 120.735 89.835 121.705 ;
        RECT 90.005 121.075 90.175 122.205 ;
        RECT 90.345 121.415 90.515 122.215 ;
        RECT 90.720 121.925 90.995 122.775 ;
        RECT 90.715 121.755 90.995 121.925 ;
        RECT 90.720 121.615 90.995 121.755 ;
        RECT 91.165 121.415 91.355 122.775 ;
        RECT 91.535 122.410 92.045 122.945 ;
        RECT 92.265 122.135 92.510 122.740 ;
        RECT 92.955 122.175 94.625 122.945 ;
        RECT 94.795 122.220 95.085 122.945 ;
        RECT 95.255 122.400 100.600 122.945 ;
        RECT 91.555 121.965 92.785 122.135 ;
        RECT 90.345 121.245 91.355 121.415 ;
        RECT 91.525 121.400 92.275 121.590 ;
        RECT 90.005 120.905 91.130 121.075 ;
        RECT 91.525 120.735 91.695 121.400 ;
        RECT 92.445 121.155 92.785 121.965 ;
        RECT 92.955 121.655 93.705 122.175 ;
        RECT 93.875 121.485 94.625 122.005 ;
        RECT 96.840 121.570 97.180 122.400 ;
        RECT 101.700 122.205 101.955 122.775 ;
        RECT 102.125 122.545 102.455 122.945 ;
        RECT 102.880 122.410 103.410 122.775 ;
        RECT 102.880 122.375 103.055 122.410 ;
        RECT 102.125 122.205 103.055 122.375 ;
        RECT 89.665 120.565 91.695 120.735 ;
        RECT 91.865 120.395 92.035 121.155 ;
        RECT 92.270 120.745 92.785 121.155 ;
        RECT 92.955 120.395 94.625 121.485 ;
        RECT 94.795 120.395 95.085 121.560 ;
        RECT 98.660 120.830 99.010 122.080 ;
        RECT 101.700 121.535 101.870 122.205 ;
        RECT 102.125 122.035 102.295 122.205 ;
        RECT 102.040 121.705 102.295 122.035 ;
        RECT 102.520 121.705 102.715 122.035 ;
        RECT 95.255 120.395 100.600 120.830 ;
        RECT 101.700 120.565 102.035 121.535 ;
        RECT 102.205 120.395 102.375 121.535 ;
        RECT 102.545 120.735 102.715 121.705 ;
        RECT 102.885 121.075 103.055 122.205 ;
        RECT 103.225 121.415 103.395 122.215 ;
        RECT 103.600 121.925 103.875 122.775 ;
        RECT 103.595 121.755 103.875 121.925 ;
        RECT 103.600 121.615 103.875 121.755 ;
        RECT 104.045 121.415 104.235 122.775 ;
        RECT 104.415 122.410 104.925 122.945 ;
        RECT 105.145 122.135 105.390 122.740 ;
        RECT 105.835 122.400 111.180 122.945 ;
        RECT 111.355 122.400 116.700 122.945 ;
        RECT 104.435 121.965 105.665 122.135 ;
        RECT 103.225 121.245 104.235 121.415 ;
        RECT 104.405 121.400 105.155 121.590 ;
        RECT 102.885 120.905 104.010 121.075 ;
        RECT 104.405 120.735 104.575 121.400 ;
        RECT 105.325 121.155 105.665 121.965 ;
        RECT 107.420 121.570 107.760 122.400 ;
        RECT 102.545 120.565 104.575 120.735 ;
        RECT 104.745 120.395 104.915 121.155 ;
        RECT 105.150 120.745 105.665 121.155 ;
        RECT 109.240 120.830 109.590 122.080 ;
        RECT 112.940 121.570 113.280 122.400 ;
        RECT 116.875 122.145 117.215 122.775 ;
        RECT 117.385 122.145 117.635 122.945 ;
        RECT 117.825 122.295 118.155 122.775 ;
        RECT 118.325 122.485 118.550 122.945 ;
        RECT 118.720 122.295 119.050 122.775 ;
        RECT 114.760 120.830 115.110 122.080 ;
        RECT 116.875 121.535 117.050 122.145 ;
        RECT 117.825 122.125 119.050 122.295 ;
        RECT 119.680 122.165 120.180 122.775 ;
        RECT 120.555 122.220 120.845 122.945 ;
        RECT 121.050 122.205 121.665 122.775 ;
        RECT 121.835 122.435 122.050 122.945 ;
        RECT 122.280 122.435 122.560 122.765 ;
        RECT 122.740 122.435 122.980 122.945 ;
        RECT 117.220 121.785 117.915 121.955 ;
        RECT 117.745 121.535 117.915 121.785 ;
        RECT 118.090 121.755 118.510 121.955 ;
        RECT 118.680 121.755 119.010 121.955 ;
        RECT 119.180 121.755 119.510 121.955 ;
        RECT 119.680 121.535 119.850 122.165 ;
        RECT 120.035 121.705 120.385 121.955 ;
        RECT 105.835 120.395 111.180 120.830 ;
        RECT 111.355 120.395 116.700 120.830 ;
        RECT 116.875 120.565 117.215 121.535 ;
        RECT 117.385 120.395 117.555 121.535 ;
        RECT 117.745 121.365 120.180 121.535 ;
        RECT 117.825 120.395 118.075 121.195 ;
        RECT 118.720 120.565 119.050 121.365 ;
        RECT 119.350 120.395 119.680 121.195 ;
        RECT 119.850 120.565 120.180 121.365 ;
        RECT 120.555 120.395 120.845 121.560 ;
        RECT 121.050 121.185 121.365 122.205 ;
        RECT 121.535 121.535 121.705 122.035 ;
        RECT 121.955 121.705 122.220 122.265 ;
        RECT 122.390 121.535 122.560 122.435 ;
        RECT 123.315 122.400 128.660 122.945 ;
        RECT 122.730 121.705 123.085 122.265 ;
        RECT 124.900 121.570 125.240 122.400 ;
        RECT 129.040 122.165 129.540 122.775 ;
        RECT 121.535 121.365 122.960 121.535 ;
        RECT 121.050 120.565 121.585 121.185 ;
        RECT 121.755 120.395 122.085 121.195 ;
        RECT 122.570 121.190 122.960 121.365 ;
        RECT 126.720 120.830 127.070 122.080 ;
        RECT 128.835 121.705 129.185 121.955 ;
        RECT 129.370 121.535 129.540 122.165 ;
        RECT 130.170 122.295 130.500 122.775 ;
        RECT 130.670 122.485 130.895 122.945 ;
        RECT 131.065 122.295 131.395 122.775 ;
        RECT 130.170 122.125 131.395 122.295 ;
        RECT 131.585 122.145 131.835 122.945 ;
        RECT 132.005 122.145 132.345 122.775 ;
        RECT 132.605 122.395 132.775 122.685 ;
        RECT 132.945 122.565 133.275 122.945 ;
        RECT 132.605 122.225 133.270 122.395 ;
        RECT 132.115 122.095 132.345 122.145 ;
        RECT 129.710 121.755 130.040 121.955 ;
        RECT 130.210 121.755 130.540 121.955 ;
        RECT 130.710 121.755 131.130 121.955 ;
        RECT 131.305 121.785 132.000 121.955 ;
        RECT 131.305 121.535 131.475 121.785 ;
        RECT 132.170 121.535 132.345 122.095 ;
        RECT 129.040 121.365 131.475 121.535 ;
        RECT 123.315 120.395 128.660 120.830 ;
        RECT 129.040 120.565 129.370 121.365 ;
        RECT 129.540 120.395 129.870 121.195 ;
        RECT 130.170 120.565 130.500 121.365 ;
        RECT 131.145 120.395 131.395 121.195 ;
        RECT 131.665 120.395 131.835 121.535 ;
        RECT 132.005 120.565 132.345 121.535 ;
        RECT 132.520 121.405 132.870 122.055 ;
        RECT 133.040 121.235 133.270 122.225 ;
        RECT 132.605 121.065 133.270 121.235 ;
        RECT 132.605 120.565 132.775 121.065 ;
        RECT 132.945 120.395 133.275 120.895 ;
        RECT 133.445 120.565 133.630 122.685 ;
        RECT 133.885 122.485 134.135 122.945 ;
        RECT 134.305 122.495 134.640 122.665 ;
        RECT 134.835 122.495 135.510 122.665 ;
        RECT 134.305 122.355 134.475 122.495 ;
        RECT 133.800 121.365 134.080 122.315 ;
        RECT 134.250 122.225 134.475 122.355 ;
        RECT 134.250 121.120 134.420 122.225 ;
        RECT 134.645 122.075 135.170 122.295 ;
        RECT 134.590 121.310 134.830 121.905 ;
        RECT 135.000 121.375 135.170 122.075 ;
        RECT 135.340 121.715 135.510 122.495 ;
        RECT 135.830 122.445 136.200 122.945 ;
        RECT 136.380 122.495 136.785 122.665 ;
        RECT 136.955 122.495 137.740 122.665 ;
        RECT 136.380 122.265 136.550 122.495 ;
        RECT 135.720 121.965 136.550 122.265 ;
        RECT 136.935 121.995 137.400 122.325 ;
        RECT 135.720 121.935 135.920 121.965 ;
        RECT 136.040 121.715 136.210 121.785 ;
        RECT 135.340 121.545 136.210 121.715 ;
        RECT 135.700 121.455 136.210 121.545 ;
        RECT 134.250 120.990 134.555 121.120 ;
        RECT 135.000 121.010 135.530 121.375 ;
        RECT 133.870 120.395 134.135 120.855 ;
        RECT 134.305 120.565 134.555 120.990 ;
        RECT 135.700 120.840 135.870 121.455 ;
        RECT 134.765 120.670 135.870 120.840 ;
        RECT 136.040 120.395 136.210 121.195 ;
        RECT 136.380 120.895 136.550 121.965 ;
        RECT 136.720 121.065 136.910 121.785 ;
        RECT 137.080 121.035 137.400 121.995 ;
        RECT 137.570 122.035 137.740 122.495 ;
        RECT 138.015 122.415 138.225 122.945 ;
        RECT 138.485 122.205 138.815 122.730 ;
        RECT 138.985 122.335 139.155 122.945 ;
        RECT 139.325 122.290 139.655 122.725 ;
        RECT 139.965 122.395 140.135 122.775 ;
        RECT 140.350 122.565 140.680 122.945 ;
        RECT 139.325 122.205 139.705 122.290 ;
        RECT 139.965 122.225 140.680 122.395 ;
        RECT 138.615 122.035 138.815 122.205 ;
        RECT 139.480 122.165 139.705 122.205 ;
        RECT 137.570 121.705 138.445 122.035 ;
        RECT 138.615 121.705 139.365 122.035 ;
        RECT 136.380 120.565 136.630 120.895 ;
        RECT 137.570 120.865 137.740 121.705 ;
        RECT 138.615 121.500 138.805 121.705 ;
        RECT 139.535 121.585 139.705 122.165 ;
        RECT 139.875 121.675 140.230 122.045 ;
        RECT 140.510 122.035 140.680 122.225 ;
        RECT 140.850 122.200 141.105 122.775 ;
        RECT 140.510 121.705 140.765 122.035 ;
        RECT 139.490 121.535 139.705 121.585 ;
        RECT 137.910 121.125 138.805 121.500 ;
        RECT 139.315 121.455 139.705 121.535 ;
        RECT 140.510 121.495 140.680 121.705 ;
        RECT 136.855 120.695 137.740 120.865 ;
        RECT 137.920 120.395 138.235 120.895 ;
        RECT 138.465 120.565 138.805 121.125 ;
        RECT 138.975 120.395 139.145 121.405 ;
        RECT 139.315 120.610 139.645 121.455 ;
        RECT 139.965 121.325 140.680 121.495 ;
        RECT 140.935 121.470 141.105 122.200 ;
        RECT 141.280 122.105 141.540 122.945 ;
        RECT 141.715 122.195 142.925 122.945 ;
        RECT 139.965 120.565 140.135 121.325 ;
        RECT 140.350 120.395 140.680 121.155 ;
        RECT 140.850 120.565 141.105 121.470 ;
        RECT 141.280 120.395 141.540 121.545 ;
        RECT 141.715 121.485 142.235 122.025 ;
        RECT 142.405 121.655 142.925 122.195 ;
        RECT 141.715 120.395 142.925 121.485 ;
        RECT 17.430 120.225 143.010 120.395 ;
        RECT 17.515 119.135 18.725 120.225 ;
        RECT 18.895 119.790 24.240 120.225 ;
        RECT 17.515 118.425 18.035 118.965 ;
        RECT 18.205 118.595 18.725 119.135 ;
        RECT 17.515 117.675 18.725 118.425 ;
        RECT 20.480 118.220 20.820 119.050 ;
        RECT 22.300 118.540 22.650 119.790 ;
        RECT 24.415 119.135 27.005 120.225 ;
        RECT 24.415 118.445 25.625 118.965 ;
        RECT 25.795 118.615 27.005 119.135 ;
        RECT 27.765 119.055 28.095 120.225 ;
        RECT 28.295 118.885 28.625 120.055 ;
        RECT 28.825 119.055 29.155 120.225 ;
        RECT 29.355 118.885 29.715 120.055 ;
        RECT 29.885 119.085 30.215 120.225 ;
        RECT 30.395 119.060 30.685 120.225 ;
        RECT 31.105 119.495 31.400 120.225 ;
        RECT 31.570 119.325 31.830 120.050 ;
        RECT 32.000 119.495 32.260 120.225 ;
        RECT 32.430 119.325 32.690 120.050 ;
        RECT 32.860 119.495 33.120 120.225 ;
        RECT 33.290 119.325 33.550 120.050 ;
        RECT 33.720 119.495 33.980 120.225 ;
        RECT 34.150 119.325 34.410 120.050 ;
        RECT 31.100 119.085 34.410 119.325 ;
        RECT 34.580 119.115 34.840 120.225 ;
        RECT 28.295 118.605 29.715 118.885 ;
        RECT 18.895 117.675 24.240 118.220 ;
        RECT 24.415 117.675 27.005 118.445 ;
        RECT 28.305 117.675 28.635 118.365 ;
        RECT 29.355 118.270 29.715 118.605 ;
        RECT 29.885 118.335 30.225 118.915 ;
        RECT 31.100 118.495 32.070 119.085 ;
        RECT 35.010 118.915 35.260 120.050 ;
        RECT 35.440 119.115 35.735 120.225 ;
        RECT 35.915 119.790 41.260 120.225 ;
        RECT 41.435 119.790 46.780 120.225 ;
        RECT 46.955 119.790 52.300 120.225 ;
        RECT 32.240 118.665 35.260 118.915 ;
        RECT 29.095 117.845 29.715 118.270 ;
        RECT 29.885 117.675 30.215 118.165 ;
        RECT 30.395 117.675 30.685 118.400 ;
        RECT 31.100 118.325 34.410 118.495 ;
        RECT 31.100 117.675 31.400 118.155 ;
        RECT 31.570 117.870 31.830 118.325 ;
        RECT 32.000 117.675 32.260 118.155 ;
        RECT 32.430 117.870 32.690 118.325 ;
        RECT 32.860 117.675 33.120 118.155 ;
        RECT 33.290 117.870 33.550 118.325 ;
        RECT 33.720 117.675 33.980 118.155 ;
        RECT 34.150 117.870 34.410 118.325 ;
        RECT 34.580 117.675 34.840 118.200 ;
        RECT 35.010 117.855 35.260 118.665 ;
        RECT 35.430 118.305 35.745 118.915 ;
        RECT 37.500 118.220 37.840 119.050 ;
        RECT 39.320 118.540 39.670 119.790 ;
        RECT 43.020 118.220 43.360 119.050 ;
        RECT 44.840 118.540 45.190 119.790 ;
        RECT 48.540 118.220 48.880 119.050 ;
        RECT 50.360 118.540 50.710 119.790 ;
        RECT 52.475 119.135 55.985 120.225 ;
        RECT 52.475 118.445 54.125 118.965 ;
        RECT 54.295 118.615 55.985 119.135 ;
        RECT 56.155 119.060 56.445 120.225 ;
        RECT 56.615 119.135 60.125 120.225 ;
        RECT 56.615 118.445 58.265 118.965 ;
        RECT 58.435 118.615 60.125 119.135 ;
        RECT 60.305 119.255 60.635 120.040 ;
        RECT 60.305 119.085 60.985 119.255 ;
        RECT 61.165 119.085 61.495 120.225 ;
        RECT 61.675 119.135 62.885 120.225 ;
        RECT 60.295 118.665 60.645 118.915 ;
        RECT 60.815 118.485 60.985 119.085 ;
        RECT 61.155 118.665 61.505 118.915 ;
        RECT 35.440 117.675 35.685 118.135 ;
        RECT 35.915 117.675 41.260 118.220 ;
        RECT 41.435 117.675 46.780 118.220 ;
        RECT 46.955 117.675 52.300 118.220 ;
        RECT 52.475 117.675 55.985 118.445 ;
        RECT 56.155 117.675 56.445 118.400 ;
        RECT 56.615 117.675 60.125 118.445 ;
        RECT 60.315 117.675 60.555 118.485 ;
        RECT 60.725 117.845 61.055 118.485 ;
        RECT 61.225 117.675 61.495 118.485 ;
        RECT 61.675 118.425 62.195 118.965 ;
        RECT 62.365 118.595 62.885 119.135 ;
        RECT 63.065 119.205 63.395 120.055 ;
        RECT 63.565 119.375 63.735 120.225 ;
        RECT 63.905 119.205 64.235 120.055 ;
        RECT 64.405 119.375 64.575 120.225 ;
        RECT 64.745 119.205 65.075 120.055 ;
        RECT 65.245 119.425 65.415 120.225 ;
        RECT 65.585 119.205 65.915 120.055 ;
        RECT 66.085 119.425 66.255 120.225 ;
        RECT 66.425 119.205 66.755 120.055 ;
        RECT 66.925 119.425 67.095 120.225 ;
        RECT 67.265 119.205 67.595 120.055 ;
        RECT 67.765 119.425 67.935 120.225 ;
        RECT 68.105 119.205 68.435 120.055 ;
        RECT 68.605 119.425 68.775 120.225 ;
        RECT 68.945 119.205 69.275 120.055 ;
        RECT 69.445 119.425 69.615 120.225 ;
        RECT 69.785 119.205 70.115 120.055 ;
        RECT 70.285 119.425 70.455 120.225 ;
        RECT 70.625 119.205 70.955 120.055 ;
        RECT 71.125 119.425 71.295 120.225 ;
        RECT 71.465 119.205 71.795 120.055 ;
        RECT 71.965 119.425 72.135 120.225 ;
        RECT 72.305 119.205 72.635 120.055 ;
        RECT 72.805 119.425 72.975 120.225 ;
        RECT 73.145 119.205 73.475 120.055 ;
        RECT 73.645 119.425 73.815 120.225 ;
        RECT 63.065 119.035 64.575 119.205 ;
        RECT 64.745 119.035 67.095 119.205 ;
        RECT 67.265 119.035 73.925 119.205 ;
        RECT 74.095 119.135 75.305 120.225 ;
        RECT 64.405 118.865 64.575 119.035 ;
        RECT 66.920 118.865 67.095 119.035 ;
        RECT 63.060 118.665 64.235 118.865 ;
        RECT 64.405 118.665 66.715 118.865 ;
        RECT 66.920 118.665 73.480 118.865 ;
        RECT 64.405 118.495 64.575 118.665 ;
        RECT 66.920 118.495 67.095 118.665 ;
        RECT 73.650 118.495 73.925 119.035 ;
        RECT 61.675 117.675 62.885 118.425 ;
        RECT 63.065 118.325 64.575 118.495 ;
        RECT 64.745 118.325 67.095 118.495 ;
        RECT 67.265 118.325 73.925 118.495 ;
        RECT 74.095 118.425 74.615 118.965 ;
        RECT 74.785 118.595 75.305 119.135 ;
        RECT 75.475 119.085 75.860 120.055 ;
        RECT 76.030 119.765 76.355 120.225 ;
        RECT 76.875 119.595 77.155 120.055 ;
        RECT 76.030 119.375 77.155 119.595 ;
        RECT 63.065 117.850 63.395 118.325 ;
        RECT 63.565 117.675 63.735 118.155 ;
        RECT 63.905 117.850 64.235 118.325 ;
        RECT 64.405 117.675 64.575 118.155 ;
        RECT 64.745 117.850 65.075 118.325 ;
        RECT 65.245 117.675 65.415 118.155 ;
        RECT 65.585 117.850 65.915 118.325 ;
        RECT 66.085 117.675 66.255 118.155 ;
        RECT 66.425 117.850 66.755 118.325 ;
        RECT 66.925 117.675 67.095 118.155 ;
        RECT 67.265 117.850 67.595 118.325 ;
        RECT 67.265 117.845 67.515 117.850 ;
        RECT 67.765 117.675 67.935 118.155 ;
        RECT 68.105 117.850 68.435 118.325 ;
        RECT 68.185 117.845 68.355 117.850 ;
        RECT 68.605 117.675 68.775 118.155 ;
        RECT 68.945 117.850 69.275 118.325 ;
        RECT 69.025 117.845 69.195 117.850 ;
        RECT 69.445 117.675 69.615 118.155 ;
        RECT 69.785 117.850 70.115 118.325 ;
        RECT 70.285 117.675 70.455 118.155 ;
        RECT 70.625 117.850 70.955 118.325 ;
        RECT 71.125 117.675 71.295 118.155 ;
        RECT 71.465 117.850 71.795 118.325 ;
        RECT 71.965 117.675 72.135 118.155 ;
        RECT 72.305 117.850 72.635 118.325 ;
        RECT 72.805 117.675 72.975 118.155 ;
        RECT 73.145 117.850 73.475 118.325 ;
        RECT 73.645 117.675 73.815 118.155 ;
        RECT 74.095 117.675 75.305 118.425 ;
        RECT 75.475 118.415 75.755 119.085 ;
        RECT 76.030 118.915 76.480 119.375 ;
        RECT 77.345 119.205 77.745 120.055 ;
        RECT 78.145 119.765 78.415 120.225 ;
        RECT 78.585 119.595 78.870 120.055 ;
        RECT 75.925 118.585 76.480 118.915 ;
        RECT 76.650 118.645 77.745 119.205 ;
        RECT 76.030 118.475 76.480 118.585 ;
        RECT 75.475 117.845 75.860 118.415 ;
        RECT 76.030 118.305 77.155 118.475 ;
        RECT 76.030 117.675 76.355 118.135 ;
        RECT 76.875 117.845 77.155 118.305 ;
        RECT 77.345 117.845 77.745 118.645 ;
        RECT 77.915 119.375 78.870 119.595 ;
        RECT 77.915 118.475 78.125 119.375 ;
        RECT 79.155 119.355 79.430 120.055 ;
        RECT 79.600 119.680 79.855 120.225 ;
        RECT 80.025 119.715 80.505 120.055 ;
        RECT 80.680 119.670 81.285 120.225 ;
        RECT 80.670 119.570 81.285 119.670 ;
        RECT 80.670 119.545 80.855 119.570 ;
        RECT 78.295 118.645 78.985 119.205 ;
        RECT 77.915 118.305 78.870 118.475 ;
        RECT 78.145 117.675 78.415 118.135 ;
        RECT 78.585 117.845 78.870 118.305 ;
        RECT 79.155 118.325 79.325 119.355 ;
        RECT 79.600 119.225 80.355 119.475 ;
        RECT 80.525 119.300 80.855 119.545 ;
        RECT 79.600 119.190 80.370 119.225 ;
        RECT 79.600 119.180 80.385 119.190 ;
        RECT 79.495 119.165 80.390 119.180 ;
        RECT 79.495 119.150 80.410 119.165 ;
        RECT 79.495 119.140 80.430 119.150 ;
        RECT 79.495 119.130 80.455 119.140 ;
        RECT 79.495 119.100 80.525 119.130 ;
        RECT 79.495 119.070 80.545 119.100 ;
        RECT 79.495 119.040 80.565 119.070 ;
        RECT 79.495 119.015 80.595 119.040 ;
        RECT 79.495 118.980 80.630 119.015 ;
        RECT 79.495 118.975 80.660 118.980 ;
        RECT 79.495 118.580 79.725 118.975 ;
        RECT 80.270 118.970 80.660 118.975 ;
        RECT 80.295 118.960 80.660 118.970 ;
        RECT 80.310 118.955 80.660 118.960 ;
        RECT 80.325 118.950 80.660 118.955 ;
        RECT 81.025 118.950 81.285 119.400 ;
        RECT 81.915 119.060 82.205 120.225 ;
        RECT 82.375 119.715 83.565 120.005 ;
        RECT 82.395 119.375 83.565 119.545 ;
        RECT 83.735 119.425 84.015 120.225 ;
        RECT 82.395 119.085 82.720 119.375 ;
        RECT 83.395 119.255 83.565 119.375 ;
        RECT 80.325 118.945 81.285 118.950 ;
        RECT 80.335 118.935 81.285 118.945 ;
        RECT 80.345 118.930 81.285 118.935 ;
        RECT 80.355 118.920 81.285 118.930 ;
        RECT 80.360 118.910 81.285 118.920 ;
        RECT 82.890 118.915 83.085 119.205 ;
        RECT 83.395 119.085 84.055 119.255 ;
        RECT 84.225 119.085 84.500 120.055 ;
        RECT 85.135 119.085 85.395 120.225 ;
        RECT 85.635 119.715 87.250 120.045 ;
        RECT 83.885 118.915 84.055 119.085 ;
        RECT 80.365 118.905 81.285 118.910 ;
        RECT 80.375 118.890 81.285 118.905 ;
        RECT 80.380 118.875 81.285 118.890 ;
        RECT 80.390 118.850 81.285 118.875 ;
        RECT 79.895 118.380 80.225 118.805 ;
        RECT 79.975 118.355 80.225 118.380 ;
        RECT 79.155 117.845 79.415 118.325 ;
        RECT 79.585 117.675 79.835 118.215 ;
        RECT 80.005 117.895 80.225 118.355 ;
        RECT 80.395 118.780 81.285 118.850 ;
        RECT 80.395 118.055 80.565 118.780 ;
        RECT 80.735 118.225 81.285 118.610 ;
        RECT 82.375 118.585 82.720 118.915 ;
        RECT 82.890 118.585 83.715 118.915 ;
        RECT 83.885 118.585 84.160 118.915 ;
        RECT 83.885 118.415 84.055 118.585 ;
        RECT 80.395 117.885 81.285 118.055 ;
        RECT 81.915 117.675 82.205 118.400 ;
        RECT 82.390 118.245 84.055 118.415 ;
        RECT 84.330 118.350 84.500 119.085 ;
        RECT 85.645 118.915 85.815 119.475 ;
        RECT 86.075 119.375 87.250 119.545 ;
        RECT 87.420 119.425 87.700 120.225 ;
        RECT 86.075 119.085 86.405 119.375 ;
        RECT 87.080 119.255 87.250 119.375 ;
        RECT 86.575 118.915 86.820 119.205 ;
        RECT 87.080 119.085 87.740 119.255 ;
        RECT 87.910 119.085 88.185 120.055 ;
        RECT 87.570 118.915 87.740 119.085 ;
        RECT 85.140 118.665 85.475 118.915 ;
        RECT 85.645 118.585 86.360 118.915 ;
        RECT 86.575 118.585 87.400 118.915 ;
        RECT 87.570 118.585 87.845 118.915 ;
        RECT 85.645 118.495 85.895 118.585 ;
        RECT 82.390 117.895 82.645 118.245 ;
        RECT 82.815 117.675 83.145 118.075 ;
        RECT 83.315 117.895 83.485 118.245 ;
        RECT 83.655 117.675 84.035 118.075 ;
        RECT 84.225 118.005 84.500 118.350 ;
        RECT 85.135 117.675 85.395 118.495 ;
        RECT 85.565 118.075 85.895 118.495 ;
        RECT 87.570 118.415 87.740 118.585 ;
        RECT 86.075 118.245 87.740 118.415 ;
        RECT 88.015 118.350 88.185 119.085 ;
        RECT 86.075 117.845 86.335 118.245 ;
        RECT 86.505 117.675 86.835 118.075 ;
        RECT 87.005 117.895 87.175 118.245 ;
        RECT 87.345 117.675 87.720 118.075 ;
        RECT 87.910 118.005 88.185 118.350 ;
        RECT 88.820 119.085 89.155 120.055 ;
        RECT 89.325 119.085 89.495 120.225 ;
        RECT 89.665 119.885 91.695 120.055 ;
        RECT 88.820 118.415 88.990 119.085 ;
        RECT 89.665 118.915 89.835 119.885 ;
        RECT 89.160 118.585 89.415 118.915 ;
        RECT 89.640 118.585 89.835 118.915 ;
        RECT 90.005 119.545 91.130 119.715 ;
        RECT 89.245 118.415 89.415 118.585 ;
        RECT 90.005 118.415 90.175 119.545 ;
        RECT 88.820 117.845 89.075 118.415 ;
        RECT 89.245 118.245 90.175 118.415 ;
        RECT 90.345 119.205 91.355 119.375 ;
        RECT 90.345 118.405 90.515 119.205 ;
        RECT 90.720 118.525 90.995 119.005 ;
        RECT 90.715 118.355 90.995 118.525 ;
        RECT 90.000 118.210 90.175 118.245 ;
        RECT 89.245 117.675 89.575 118.075 ;
        RECT 90.000 117.845 90.530 118.210 ;
        RECT 90.720 117.845 90.995 118.355 ;
        RECT 91.165 117.845 91.355 119.205 ;
        RECT 91.525 119.220 91.695 119.885 ;
        RECT 91.865 119.465 92.035 120.225 ;
        RECT 92.270 119.465 92.785 119.875 ;
        RECT 92.955 119.790 98.300 120.225 ;
        RECT 91.525 119.030 92.275 119.220 ;
        RECT 92.445 118.655 92.785 119.465 ;
        RECT 91.555 118.485 92.785 118.655 ;
        RECT 91.535 117.675 92.045 118.210 ;
        RECT 92.265 117.880 92.510 118.485 ;
        RECT 94.540 118.220 94.880 119.050 ;
        RECT 96.360 118.540 96.710 119.790 ;
        RECT 98.475 119.135 99.685 120.225 ;
        RECT 99.945 119.555 100.115 120.055 ;
        RECT 100.285 119.725 100.615 120.225 ;
        RECT 99.945 119.385 100.610 119.555 ;
        RECT 98.475 118.425 98.995 118.965 ;
        RECT 99.165 118.595 99.685 119.135 ;
        RECT 99.860 118.565 100.210 119.215 ;
        RECT 92.955 117.675 98.300 118.220 ;
        RECT 98.475 117.675 99.685 118.425 ;
        RECT 100.380 118.395 100.610 119.385 ;
        RECT 99.945 118.225 100.610 118.395 ;
        RECT 99.945 117.935 100.115 118.225 ;
        RECT 100.285 117.675 100.615 118.055 ;
        RECT 100.785 117.935 100.970 120.055 ;
        RECT 101.210 119.765 101.475 120.225 ;
        RECT 101.645 119.630 101.895 120.055 ;
        RECT 102.105 119.780 103.210 119.950 ;
        RECT 101.590 119.500 101.895 119.630 ;
        RECT 101.140 118.305 101.420 119.255 ;
        RECT 101.590 118.395 101.760 119.500 ;
        RECT 101.930 118.715 102.170 119.310 ;
        RECT 102.340 119.245 102.870 119.610 ;
        RECT 102.340 118.545 102.510 119.245 ;
        RECT 103.040 119.165 103.210 119.780 ;
        RECT 103.380 119.425 103.550 120.225 ;
        RECT 103.720 119.725 103.970 120.055 ;
        RECT 104.195 119.755 105.080 119.925 ;
        RECT 103.040 119.075 103.550 119.165 ;
        RECT 101.590 118.265 101.815 118.395 ;
        RECT 101.985 118.325 102.510 118.545 ;
        RECT 102.680 118.905 103.550 119.075 ;
        RECT 101.225 117.675 101.475 118.135 ;
        RECT 101.645 118.125 101.815 118.265 ;
        RECT 102.680 118.125 102.850 118.905 ;
        RECT 103.380 118.835 103.550 118.905 ;
        RECT 103.060 118.655 103.260 118.685 ;
        RECT 103.720 118.655 103.890 119.725 ;
        RECT 104.060 118.835 104.250 119.555 ;
        RECT 103.060 118.355 103.890 118.655 ;
        RECT 104.420 118.625 104.740 119.585 ;
        RECT 101.645 117.955 101.980 118.125 ;
        RECT 102.175 117.955 102.850 118.125 ;
        RECT 103.170 117.675 103.540 118.175 ;
        RECT 103.720 118.125 103.890 118.355 ;
        RECT 104.275 118.295 104.740 118.625 ;
        RECT 104.910 118.915 105.080 119.755 ;
        RECT 105.260 119.725 105.575 120.225 ;
        RECT 105.805 119.495 106.145 120.055 ;
        RECT 105.250 119.120 106.145 119.495 ;
        RECT 106.315 119.215 106.485 120.225 ;
        RECT 105.955 118.915 106.145 119.120 ;
        RECT 106.655 119.165 106.985 120.010 ;
        RECT 106.655 119.085 107.045 119.165 ;
        RECT 106.830 119.035 107.045 119.085 ;
        RECT 107.675 119.060 107.965 120.225 ;
        RECT 108.140 119.085 108.475 120.055 ;
        RECT 108.645 119.085 108.815 120.225 ;
        RECT 108.985 119.885 111.015 120.055 ;
        RECT 104.910 118.585 105.785 118.915 ;
        RECT 105.955 118.585 106.705 118.915 ;
        RECT 104.910 118.125 105.080 118.585 ;
        RECT 105.955 118.415 106.155 118.585 ;
        RECT 106.875 118.455 107.045 119.035 ;
        RECT 106.820 118.415 107.045 118.455 ;
        RECT 103.720 117.955 104.125 118.125 ;
        RECT 104.295 117.955 105.080 118.125 ;
        RECT 105.355 117.675 105.565 118.205 ;
        RECT 105.825 117.890 106.155 118.415 ;
        RECT 106.665 118.330 107.045 118.415 ;
        RECT 108.140 118.415 108.310 119.085 ;
        RECT 108.985 118.915 109.155 119.885 ;
        RECT 108.480 118.585 108.735 118.915 ;
        RECT 108.960 118.585 109.155 118.915 ;
        RECT 109.325 119.545 110.450 119.715 ;
        RECT 108.565 118.415 108.735 118.585 ;
        RECT 109.325 118.415 109.495 119.545 ;
        RECT 106.325 117.675 106.495 118.285 ;
        RECT 106.665 117.895 106.995 118.330 ;
        RECT 107.675 117.675 107.965 118.400 ;
        RECT 108.140 117.845 108.395 118.415 ;
        RECT 108.565 118.245 109.495 118.415 ;
        RECT 109.665 119.205 110.675 119.375 ;
        RECT 109.665 118.405 109.835 119.205 ;
        RECT 110.040 118.525 110.315 119.005 ;
        RECT 110.035 118.355 110.315 118.525 ;
        RECT 109.320 118.210 109.495 118.245 ;
        RECT 108.565 117.675 108.895 118.075 ;
        RECT 109.320 117.845 109.850 118.210 ;
        RECT 110.040 117.845 110.315 118.355 ;
        RECT 110.485 117.845 110.675 119.205 ;
        RECT 110.845 119.220 111.015 119.885 ;
        RECT 111.185 119.465 111.355 120.225 ;
        RECT 111.590 119.465 112.105 119.875 ;
        RECT 110.845 119.030 111.595 119.220 ;
        RECT 111.765 118.655 112.105 119.465 ;
        RECT 110.875 118.485 112.105 118.655 ;
        RECT 112.275 119.085 112.660 120.055 ;
        RECT 112.830 119.765 113.155 120.225 ;
        RECT 113.675 119.595 113.955 120.055 ;
        RECT 112.830 119.375 113.955 119.595 ;
        RECT 110.855 117.675 111.365 118.210 ;
        RECT 111.585 117.880 111.830 118.485 ;
        RECT 112.275 118.415 112.555 119.085 ;
        RECT 112.830 118.915 113.280 119.375 ;
        RECT 114.145 119.205 114.545 120.055 ;
        RECT 114.945 119.765 115.215 120.225 ;
        RECT 115.385 119.595 115.670 120.055 ;
        RECT 112.725 118.585 113.280 118.915 ;
        RECT 113.450 118.645 114.545 119.205 ;
        RECT 112.830 118.475 113.280 118.585 ;
        RECT 112.275 117.845 112.660 118.415 ;
        RECT 112.830 118.305 113.955 118.475 ;
        RECT 112.830 117.675 113.155 118.135 ;
        RECT 113.675 117.845 113.955 118.305 ;
        RECT 114.145 117.845 114.545 118.645 ;
        RECT 114.715 119.375 115.670 119.595 ;
        RECT 116.505 119.555 116.675 120.055 ;
        RECT 116.845 119.725 117.175 120.225 ;
        RECT 116.505 119.385 117.170 119.555 ;
        RECT 114.715 118.475 114.925 119.375 ;
        RECT 115.095 118.645 115.785 119.205 ;
        RECT 116.420 118.565 116.770 119.215 ;
        RECT 114.715 118.305 115.670 118.475 ;
        RECT 116.940 118.395 117.170 119.385 ;
        RECT 114.945 117.675 115.215 118.135 ;
        RECT 115.385 117.845 115.670 118.305 ;
        RECT 116.505 118.225 117.170 118.395 ;
        RECT 116.505 117.935 116.675 118.225 ;
        RECT 116.845 117.675 117.175 118.055 ;
        RECT 117.345 117.935 117.530 120.055 ;
        RECT 117.770 119.765 118.035 120.225 ;
        RECT 118.205 119.630 118.455 120.055 ;
        RECT 118.665 119.780 119.770 119.950 ;
        RECT 118.150 119.500 118.455 119.630 ;
        RECT 117.700 118.305 117.980 119.255 ;
        RECT 118.150 118.395 118.320 119.500 ;
        RECT 118.490 118.715 118.730 119.310 ;
        RECT 118.900 119.245 119.430 119.610 ;
        RECT 118.900 118.545 119.070 119.245 ;
        RECT 119.600 119.165 119.770 119.780 ;
        RECT 119.940 119.425 120.110 120.225 ;
        RECT 120.280 119.725 120.530 120.055 ;
        RECT 120.755 119.755 121.640 119.925 ;
        RECT 119.600 119.075 120.110 119.165 ;
        RECT 118.150 118.265 118.375 118.395 ;
        RECT 118.545 118.325 119.070 118.545 ;
        RECT 119.240 118.905 120.110 119.075 ;
        RECT 117.785 117.675 118.035 118.135 ;
        RECT 118.205 118.125 118.375 118.265 ;
        RECT 119.240 118.125 119.410 118.905 ;
        RECT 119.940 118.835 120.110 118.905 ;
        RECT 119.620 118.655 119.820 118.685 ;
        RECT 120.280 118.655 120.450 119.725 ;
        RECT 120.620 118.835 120.810 119.555 ;
        RECT 119.620 118.355 120.450 118.655 ;
        RECT 120.980 118.625 121.300 119.585 ;
        RECT 118.205 117.955 118.540 118.125 ;
        RECT 118.735 117.955 119.410 118.125 ;
        RECT 119.730 117.675 120.100 118.175 ;
        RECT 120.280 118.125 120.450 118.355 ;
        RECT 120.835 118.295 121.300 118.625 ;
        RECT 121.470 118.915 121.640 119.755 ;
        RECT 121.820 119.725 122.135 120.225 ;
        RECT 122.365 119.495 122.705 120.055 ;
        RECT 121.810 119.120 122.705 119.495 ;
        RECT 122.875 119.215 123.045 120.225 ;
        RECT 122.515 118.915 122.705 119.120 ;
        RECT 123.215 119.165 123.545 120.010 ;
        RECT 123.775 119.790 129.120 120.225 ;
        RECT 123.215 119.085 123.605 119.165 ;
        RECT 123.390 119.035 123.605 119.085 ;
        RECT 121.470 118.585 122.345 118.915 ;
        RECT 122.515 118.585 123.265 118.915 ;
        RECT 121.470 118.125 121.640 118.585 ;
        RECT 122.515 118.415 122.715 118.585 ;
        RECT 123.435 118.455 123.605 119.035 ;
        RECT 123.380 118.415 123.605 118.455 ;
        RECT 120.280 117.955 120.685 118.125 ;
        RECT 120.855 117.955 121.640 118.125 ;
        RECT 121.915 117.675 122.125 118.205 ;
        RECT 122.385 117.890 122.715 118.415 ;
        RECT 123.225 118.330 123.605 118.415 ;
        RECT 122.885 117.675 123.055 118.285 ;
        RECT 123.225 117.895 123.555 118.330 ;
        RECT 125.360 118.220 125.700 119.050 ;
        RECT 127.180 118.540 127.530 119.790 ;
        RECT 129.295 119.135 132.805 120.225 ;
        RECT 129.295 118.445 130.945 118.965 ;
        RECT 131.115 118.615 132.805 119.135 ;
        RECT 133.435 119.060 133.725 120.225 ;
        RECT 133.895 119.375 134.155 120.055 ;
        RECT 134.325 119.445 134.575 120.225 ;
        RECT 134.825 119.675 135.075 120.055 ;
        RECT 135.245 119.845 135.600 120.225 ;
        RECT 136.605 119.835 136.940 120.055 ;
        RECT 136.205 119.675 136.435 119.715 ;
        RECT 134.825 119.475 136.435 119.675 ;
        RECT 134.825 119.465 135.660 119.475 ;
        RECT 136.250 119.385 136.435 119.475 ;
        RECT 123.775 117.675 129.120 118.220 ;
        RECT 129.295 117.675 132.805 118.445 ;
        RECT 133.435 117.675 133.725 118.400 ;
        RECT 133.895 118.175 134.065 119.375 ;
        RECT 135.765 119.275 136.095 119.305 ;
        RECT 134.295 119.215 136.095 119.275 ;
        RECT 136.685 119.215 136.940 119.835 ;
        RECT 134.235 119.105 136.940 119.215 ;
        RECT 138.125 119.295 138.295 120.055 ;
        RECT 138.510 119.465 138.840 120.225 ;
        RECT 138.125 119.125 138.840 119.295 ;
        RECT 139.010 119.150 139.265 120.055 ;
        RECT 134.235 119.070 134.435 119.105 ;
        RECT 134.235 118.495 134.405 119.070 ;
        RECT 135.765 119.045 136.940 119.105 ;
        RECT 134.635 118.630 135.045 118.935 ;
        RECT 135.215 118.665 135.545 118.875 ;
        RECT 134.235 118.375 134.505 118.495 ;
        RECT 134.235 118.330 135.080 118.375 ;
        RECT 134.325 118.205 135.080 118.330 ;
        RECT 135.335 118.265 135.545 118.665 ;
        RECT 135.790 118.665 136.265 118.875 ;
        RECT 136.455 118.665 136.945 118.865 ;
        RECT 135.790 118.265 136.010 118.665 ;
        RECT 138.035 118.575 138.390 118.945 ;
        RECT 138.670 118.915 138.840 119.125 ;
        RECT 138.670 118.585 138.925 118.915 ;
        RECT 133.895 117.845 134.155 118.175 ;
        RECT 134.910 118.055 135.080 118.205 ;
        RECT 134.325 117.675 134.655 118.035 ;
        RECT 134.910 117.845 136.210 118.055 ;
        RECT 136.485 117.675 136.940 118.440 ;
        RECT 138.670 118.395 138.840 118.585 ;
        RECT 139.095 118.420 139.265 119.150 ;
        RECT 139.440 119.075 139.700 120.225 ;
        RECT 139.965 119.295 140.135 120.055 ;
        RECT 140.350 119.465 140.680 120.225 ;
        RECT 139.965 119.125 140.680 119.295 ;
        RECT 140.850 119.150 141.105 120.055 ;
        RECT 139.875 118.575 140.230 118.945 ;
        RECT 140.510 118.915 140.680 119.125 ;
        RECT 140.510 118.585 140.765 118.915 ;
        RECT 138.125 118.225 138.840 118.395 ;
        RECT 138.125 117.845 138.295 118.225 ;
        RECT 138.510 117.675 138.840 118.055 ;
        RECT 139.010 117.845 139.265 118.420 ;
        RECT 139.440 117.675 139.700 118.515 ;
        RECT 140.510 118.395 140.680 118.585 ;
        RECT 140.935 118.420 141.105 119.150 ;
        RECT 141.280 119.075 141.540 120.225 ;
        RECT 141.715 119.135 142.925 120.225 ;
        RECT 141.715 118.595 142.235 119.135 ;
        RECT 139.965 118.225 140.680 118.395 ;
        RECT 139.965 117.845 140.135 118.225 ;
        RECT 140.350 117.675 140.680 118.055 ;
        RECT 140.850 117.845 141.105 118.420 ;
        RECT 141.280 117.675 141.540 118.515 ;
        RECT 142.405 118.425 142.925 118.965 ;
        RECT 141.715 117.675 142.925 118.425 ;
        RECT 17.430 117.505 143.010 117.675 ;
        RECT 17.515 116.755 18.725 117.505 ;
        RECT 18.895 116.960 24.240 117.505 ;
        RECT 17.515 116.215 18.035 116.755 ;
        RECT 18.205 116.045 18.725 116.585 ;
        RECT 20.480 116.130 20.820 116.960 ;
        RECT 24.415 116.735 27.005 117.505 ;
        RECT 27.635 116.855 27.895 117.335 ;
        RECT 28.065 116.965 28.315 117.505 ;
        RECT 17.515 114.955 18.725 116.045 ;
        RECT 22.300 115.390 22.650 116.640 ;
        RECT 24.415 116.215 25.625 116.735 ;
        RECT 25.795 116.045 27.005 116.565 ;
        RECT 18.895 114.955 24.240 115.390 ;
        RECT 24.415 114.955 27.005 116.045 ;
        RECT 27.635 115.825 27.805 116.855 ;
        RECT 28.485 116.825 28.705 117.285 ;
        RECT 28.455 116.800 28.705 116.825 ;
        RECT 27.975 116.205 28.205 116.600 ;
        RECT 28.375 116.375 28.705 116.800 ;
        RECT 28.875 117.125 29.765 117.295 ;
        RECT 28.875 116.400 29.045 117.125 ;
        RECT 29.215 116.570 29.765 116.955 ;
        RECT 29.935 116.735 31.605 117.505 ;
        RECT 32.245 116.855 32.575 117.330 ;
        RECT 32.745 117.025 32.915 117.505 ;
        RECT 33.085 116.855 33.415 117.330 ;
        RECT 33.585 117.025 33.755 117.505 ;
        RECT 33.925 116.855 34.255 117.330 ;
        RECT 34.425 117.025 34.595 117.505 ;
        RECT 34.765 116.855 35.095 117.330 ;
        RECT 35.265 117.025 35.435 117.505 ;
        RECT 35.605 116.855 35.935 117.330 ;
        RECT 36.105 117.025 36.275 117.505 ;
        RECT 36.445 117.330 36.695 117.335 ;
        RECT 36.445 116.855 36.775 117.330 ;
        RECT 36.945 117.025 37.115 117.505 ;
        RECT 37.365 117.330 37.535 117.335 ;
        RECT 37.285 116.855 37.615 117.330 ;
        RECT 37.785 117.025 37.955 117.505 ;
        RECT 38.205 117.330 38.375 117.335 ;
        RECT 38.125 116.855 38.455 117.330 ;
        RECT 38.625 117.025 38.795 117.505 ;
        RECT 38.965 116.855 39.295 117.330 ;
        RECT 39.465 117.025 39.635 117.505 ;
        RECT 39.805 116.855 40.135 117.330 ;
        RECT 40.305 117.025 40.475 117.505 ;
        RECT 40.645 116.855 40.975 117.330 ;
        RECT 41.145 117.025 41.315 117.505 ;
        RECT 41.485 116.855 41.815 117.330 ;
        RECT 41.985 117.025 42.155 117.505 ;
        RECT 42.325 116.855 42.655 117.330 ;
        RECT 42.825 117.025 42.995 117.505 ;
        RECT 28.875 116.330 29.765 116.400 ;
        RECT 28.870 116.305 29.765 116.330 ;
        RECT 28.860 116.290 29.765 116.305 ;
        RECT 28.855 116.275 29.765 116.290 ;
        RECT 28.845 116.270 29.765 116.275 ;
        RECT 28.840 116.260 29.765 116.270 ;
        RECT 28.835 116.250 29.765 116.260 ;
        RECT 28.825 116.245 29.765 116.250 ;
        RECT 28.815 116.235 29.765 116.245 ;
        RECT 28.805 116.230 29.765 116.235 ;
        RECT 28.805 116.225 29.140 116.230 ;
        RECT 28.790 116.220 29.140 116.225 ;
        RECT 28.775 116.210 29.140 116.220 ;
        RECT 28.750 116.205 29.140 116.210 ;
        RECT 27.975 116.200 29.140 116.205 ;
        RECT 27.975 116.165 29.110 116.200 ;
        RECT 27.975 116.140 29.075 116.165 ;
        RECT 27.975 116.110 29.045 116.140 ;
        RECT 27.975 116.080 29.025 116.110 ;
        RECT 27.975 116.050 29.005 116.080 ;
        RECT 27.975 116.040 28.935 116.050 ;
        RECT 27.975 116.030 28.910 116.040 ;
        RECT 27.975 116.015 28.890 116.030 ;
        RECT 27.975 116.000 28.870 116.015 ;
        RECT 28.080 115.990 28.865 116.000 ;
        RECT 28.080 115.955 28.850 115.990 ;
        RECT 27.635 115.125 27.910 115.825 ;
        RECT 28.080 115.705 28.835 115.955 ;
        RECT 29.005 115.635 29.335 115.880 ;
        RECT 29.505 115.780 29.765 116.230 ;
        RECT 29.935 116.215 30.685 116.735 ;
        RECT 32.245 116.685 33.755 116.855 ;
        RECT 33.925 116.685 36.275 116.855 ;
        RECT 36.445 116.685 43.105 116.855 ;
        RECT 43.275 116.780 43.565 117.505 ;
        RECT 43.735 116.960 49.080 117.505 ;
        RECT 49.255 116.960 54.600 117.505 ;
        RECT 30.855 116.045 31.605 116.565 ;
        RECT 33.585 116.515 33.755 116.685 ;
        RECT 36.100 116.515 36.275 116.685 ;
        RECT 32.240 116.315 33.415 116.515 ;
        RECT 33.585 116.315 35.895 116.515 ;
        RECT 36.100 116.315 42.660 116.515 ;
        RECT 33.585 116.145 33.755 116.315 ;
        RECT 36.100 116.145 36.275 116.315 ;
        RECT 42.830 116.145 43.105 116.685 ;
        RECT 29.150 115.610 29.335 115.635 ;
        RECT 29.150 115.510 29.765 115.610 ;
        RECT 28.080 114.955 28.335 115.500 ;
        RECT 28.505 115.125 28.985 115.465 ;
        RECT 29.160 114.955 29.765 115.510 ;
        RECT 29.935 114.955 31.605 116.045 ;
        RECT 32.245 115.975 33.755 116.145 ;
        RECT 33.925 115.975 36.275 116.145 ;
        RECT 36.445 115.975 43.105 116.145 ;
        RECT 45.320 116.130 45.660 116.960 ;
        RECT 32.245 115.125 32.575 115.975 ;
        RECT 32.745 114.955 32.915 115.805 ;
        RECT 33.085 115.125 33.415 115.975 ;
        RECT 33.585 114.955 33.755 115.805 ;
        RECT 33.925 115.125 34.255 115.975 ;
        RECT 34.425 114.955 34.595 115.755 ;
        RECT 34.765 115.125 35.095 115.975 ;
        RECT 35.265 114.955 35.435 115.755 ;
        RECT 35.605 115.125 35.935 115.975 ;
        RECT 36.105 114.955 36.275 115.755 ;
        RECT 36.445 115.125 36.775 115.975 ;
        RECT 36.945 114.955 37.115 115.755 ;
        RECT 37.285 115.125 37.615 115.975 ;
        RECT 37.785 114.955 37.955 115.755 ;
        RECT 38.125 115.125 38.455 115.975 ;
        RECT 38.625 114.955 38.795 115.755 ;
        RECT 38.965 115.125 39.295 115.975 ;
        RECT 39.465 114.955 39.635 115.755 ;
        RECT 39.805 115.125 40.135 115.975 ;
        RECT 40.305 114.955 40.475 115.755 ;
        RECT 40.645 115.125 40.975 115.975 ;
        RECT 41.145 114.955 41.315 115.755 ;
        RECT 41.485 115.125 41.815 115.975 ;
        RECT 41.985 114.955 42.155 115.755 ;
        RECT 42.325 115.125 42.655 115.975 ;
        RECT 42.825 114.955 42.995 115.755 ;
        RECT 43.275 114.955 43.565 116.120 ;
        RECT 47.140 115.390 47.490 116.640 ;
        RECT 50.840 116.130 51.180 116.960 ;
        RECT 54.775 116.735 57.365 117.505 ;
        RECT 58.110 116.875 58.395 117.335 ;
        RECT 58.565 117.045 58.835 117.505 ;
        RECT 52.660 115.390 53.010 116.640 ;
        RECT 54.775 116.215 55.985 116.735 ;
        RECT 58.110 116.705 59.065 116.875 ;
        RECT 56.155 116.045 57.365 116.565 ;
        RECT 43.735 114.955 49.080 115.390 ;
        RECT 49.255 114.955 54.600 115.390 ;
        RECT 54.775 114.955 57.365 116.045 ;
        RECT 57.995 115.975 58.685 116.535 ;
        RECT 58.855 115.805 59.065 116.705 ;
        RECT 58.110 115.585 59.065 115.805 ;
        RECT 59.235 116.535 59.635 117.335 ;
        RECT 59.825 116.875 60.105 117.335 ;
        RECT 60.625 117.045 60.950 117.505 ;
        RECT 59.825 116.705 60.950 116.875 ;
        RECT 61.120 116.765 61.505 117.335 ;
        RECT 61.765 116.955 61.935 117.245 ;
        RECT 62.105 117.125 62.435 117.505 ;
        RECT 61.765 116.785 62.430 116.955 ;
        RECT 60.500 116.595 60.950 116.705 ;
        RECT 59.235 115.975 60.330 116.535 ;
        RECT 60.500 116.265 61.055 116.595 ;
        RECT 58.110 115.125 58.395 115.585 ;
        RECT 58.565 114.955 58.835 115.415 ;
        RECT 59.235 115.125 59.635 115.975 ;
        RECT 60.500 115.805 60.950 116.265 ;
        RECT 61.225 116.095 61.505 116.765 ;
        RECT 59.825 115.585 60.950 115.805 ;
        RECT 59.825 115.125 60.105 115.585 ;
        RECT 60.625 114.955 60.950 115.415 ;
        RECT 61.120 115.125 61.505 116.095 ;
        RECT 61.680 115.965 62.030 116.615 ;
        RECT 62.200 115.795 62.430 116.785 ;
        RECT 61.765 115.625 62.430 115.795 ;
        RECT 61.765 115.125 61.935 115.625 ;
        RECT 62.105 114.955 62.435 115.455 ;
        RECT 62.605 115.125 62.790 117.245 ;
        RECT 63.045 117.045 63.295 117.505 ;
        RECT 63.465 117.055 63.800 117.225 ;
        RECT 63.995 117.055 64.670 117.225 ;
        RECT 63.465 116.915 63.635 117.055 ;
        RECT 62.960 115.925 63.240 116.875 ;
        RECT 63.410 116.785 63.635 116.915 ;
        RECT 63.410 115.680 63.580 116.785 ;
        RECT 63.805 116.635 64.330 116.855 ;
        RECT 63.750 115.870 63.990 116.465 ;
        RECT 64.160 115.935 64.330 116.635 ;
        RECT 64.500 116.275 64.670 117.055 ;
        RECT 64.990 117.005 65.360 117.505 ;
        RECT 65.540 117.055 65.945 117.225 ;
        RECT 66.115 117.055 66.900 117.225 ;
        RECT 65.540 116.825 65.710 117.055 ;
        RECT 64.880 116.525 65.710 116.825 ;
        RECT 66.095 116.555 66.560 116.885 ;
        RECT 64.880 116.495 65.080 116.525 ;
        RECT 65.200 116.275 65.370 116.345 ;
        RECT 64.500 116.105 65.370 116.275 ;
        RECT 64.860 116.015 65.370 116.105 ;
        RECT 63.410 115.550 63.715 115.680 ;
        RECT 64.160 115.570 64.690 115.935 ;
        RECT 63.030 114.955 63.295 115.415 ;
        RECT 63.465 115.125 63.715 115.550 ;
        RECT 64.860 115.400 65.030 116.015 ;
        RECT 63.925 115.230 65.030 115.400 ;
        RECT 65.200 114.955 65.370 115.755 ;
        RECT 65.540 115.455 65.710 116.525 ;
        RECT 65.880 115.625 66.070 116.345 ;
        RECT 66.240 115.595 66.560 116.555 ;
        RECT 66.730 116.595 66.900 117.055 ;
        RECT 67.175 116.975 67.385 117.505 ;
        RECT 67.645 116.765 67.975 117.290 ;
        RECT 68.145 116.895 68.315 117.505 ;
        RECT 68.485 116.850 68.815 117.285 ;
        RECT 68.485 116.765 68.865 116.850 ;
        RECT 69.035 116.780 69.325 117.505 ;
        RECT 69.585 116.955 69.755 117.245 ;
        RECT 69.925 117.125 70.255 117.505 ;
        RECT 69.585 116.785 70.250 116.955 ;
        RECT 67.775 116.595 67.975 116.765 ;
        RECT 68.640 116.725 68.865 116.765 ;
        RECT 66.730 116.265 67.605 116.595 ;
        RECT 67.775 116.265 68.525 116.595 ;
        RECT 65.540 115.125 65.790 115.455 ;
        RECT 66.730 115.425 66.900 116.265 ;
        RECT 67.775 116.060 67.965 116.265 ;
        RECT 68.695 116.145 68.865 116.725 ;
        RECT 68.650 116.095 68.865 116.145 ;
        RECT 67.070 115.685 67.965 116.060 ;
        RECT 68.475 116.015 68.865 116.095 ;
        RECT 66.015 115.255 66.900 115.425 ;
        RECT 67.080 114.955 67.395 115.455 ;
        RECT 67.625 115.125 67.965 115.685 ;
        RECT 68.135 114.955 68.305 115.965 ;
        RECT 68.475 115.170 68.805 116.015 ;
        RECT 69.035 114.955 69.325 116.120 ;
        RECT 69.500 115.965 69.850 116.615 ;
        RECT 70.020 115.795 70.250 116.785 ;
        RECT 69.585 115.625 70.250 115.795 ;
        RECT 69.585 115.125 69.755 115.625 ;
        RECT 69.925 114.955 70.255 115.455 ;
        RECT 70.425 115.125 70.610 117.245 ;
        RECT 70.865 117.045 71.115 117.505 ;
        RECT 71.285 117.055 71.620 117.225 ;
        RECT 71.815 117.055 72.490 117.225 ;
        RECT 71.285 116.915 71.455 117.055 ;
        RECT 70.780 115.925 71.060 116.875 ;
        RECT 71.230 116.785 71.455 116.915 ;
        RECT 71.230 115.680 71.400 116.785 ;
        RECT 71.625 116.635 72.150 116.855 ;
        RECT 71.570 115.870 71.810 116.465 ;
        RECT 71.980 115.935 72.150 116.635 ;
        RECT 72.320 116.275 72.490 117.055 ;
        RECT 72.810 117.005 73.180 117.505 ;
        RECT 73.360 117.055 73.765 117.225 ;
        RECT 73.935 117.055 74.720 117.225 ;
        RECT 73.360 116.825 73.530 117.055 ;
        RECT 72.700 116.525 73.530 116.825 ;
        RECT 73.915 116.555 74.380 116.885 ;
        RECT 72.700 116.495 72.900 116.525 ;
        RECT 73.020 116.275 73.190 116.345 ;
        RECT 72.320 116.105 73.190 116.275 ;
        RECT 72.680 116.015 73.190 116.105 ;
        RECT 71.230 115.550 71.535 115.680 ;
        RECT 71.980 115.570 72.510 115.935 ;
        RECT 70.850 114.955 71.115 115.415 ;
        RECT 71.285 115.125 71.535 115.550 ;
        RECT 72.680 115.400 72.850 116.015 ;
        RECT 71.745 115.230 72.850 115.400 ;
        RECT 73.020 114.955 73.190 115.755 ;
        RECT 73.360 115.455 73.530 116.525 ;
        RECT 73.700 115.625 73.890 116.345 ;
        RECT 74.060 115.595 74.380 116.555 ;
        RECT 74.550 116.595 74.720 117.055 ;
        RECT 74.995 116.975 75.205 117.505 ;
        RECT 75.465 116.765 75.795 117.290 ;
        RECT 75.965 116.895 76.135 117.505 ;
        RECT 76.305 116.850 76.635 117.285 ;
        RECT 76.970 116.875 77.255 117.335 ;
        RECT 77.425 117.045 77.695 117.505 ;
        RECT 76.305 116.765 76.685 116.850 ;
        RECT 75.595 116.595 75.795 116.765 ;
        RECT 76.460 116.725 76.685 116.765 ;
        RECT 74.550 116.265 75.425 116.595 ;
        RECT 75.595 116.265 76.345 116.595 ;
        RECT 73.360 115.125 73.610 115.455 ;
        RECT 74.550 115.425 74.720 116.265 ;
        RECT 75.595 116.060 75.785 116.265 ;
        RECT 76.515 116.145 76.685 116.725 ;
        RECT 76.970 116.705 77.925 116.875 ;
        RECT 76.470 116.095 76.685 116.145 ;
        RECT 74.890 115.685 75.785 116.060 ;
        RECT 76.295 116.015 76.685 116.095 ;
        RECT 73.835 115.255 74.720 115.425 ;
        RECT 74.900 114.955 75.215 115.455 ;
        RECT 75.445 115.125 75.785 115.685 ;
        RECT 75.955 114.955 76.125 115.965 ;
        RECT 76.295 115.170 76.625 116.015 ;
        RECT 76.855 115.975 77.545 116.535 ;
        RECT 77.715 115.805 77.925 116.705 ;
        RECT 76.970 115.585 77.925 115.805 ;
        RECT 78.095 116.535 78.495 117.335 ;
        RECT 78.685 116.875 78.965 117.335 ;
        RECT 79.485 117.045 79.810 117.505 ;
        RECT 78.685 116.705 79.810 116.875 ;
        RECT 79.980 116.765 80.365 117.335 ;
        RECT 79.360 116.595 79.810 116.705 ;
        RECT 78.095 115.975 79.190 116.535 ;
        RECT 79.360 116.265 79.915 116.595 ;
        RECT 76.970 115.125 77.255 115.585 ;
        RECT 77.425 114.955 77.695 115.415 ;
        RECT 78.095 115.125 78.495 115.975 ;
        RECT 79.360 115.805 79.810 116.265 ;
        RECT 80.085 116.095 80.365 116.765 ;
        RECT 80.535 116.735 82.205 117.505 ;
        RECT 82.380 116.765 82.635 117.335 ;
        RECT 82.805 117.105 83.135 117.505 ;
        RECT 83.560 116.970 84.090 117.335 ;
        RECT 83.560 116.935 83.735 116.970 ;
        RECT 82.805 116.765 83.735 116.935 ;
        RECT 84.280 116.825 84.555 117.335 ;
        RECT 80.535 116.215 81.285 116.735 ;
        RECT 78.685 115.585 79.810 115.805 ;
        RECT 78.685 115.125 78.965 115.585 ;
        RECT 79.485 114.955 79.810 115.415 ;
        RECT 79.980 115.125 80.365 116.095 ;
        RECT 81.455 116.045 82.205 116.565 ;
        RECT 80.535 114.955 82.205 116.045 ;
        RECT 82.380 116.095 82.550 116.765 ;
        RECT 82.805 116.595 82.975 116.765 ;
        RECT 82.720 116.265 82.975 116.595 ;
        RECT 83.200 116.265 83.395 116.595 ;
        RECT 82.380 115.125 82.715 116.095 ;
        RECT 82.885 114.955 83.055 116.095 ;
        RECT 83.225 115.295 83.395 116.265 ;
        RECT 83.565 115.635 83.735 116.765 ;
        RECT 83.905 115.975 84.075 116.775 ;
        RECT 84.275 116.655 84.555 116.825 ;
        RECT 84.280 116.175 84.555 116.655 ;
        RECT 84.725 115.975 84.915 117.335 ;
        RECT 85.095 116.970 85.605 117.505 ;
        RECT 85.825 116.695 86.070 117.300 ;
        RECT 87.065 116.955 87.235 117.245 ;
        RECT 87.405 117.125 87.735 117.505 ;
        RECT 87.065 116.785 87.730 116.955 ;
        RECT 85.115 116.525 86.345 116.695 ;
        RECT 83.905 115.805 84.915 115.975 ;
        RECT 85.085 115.960 85.835 116.150 ;
        RECT 83.565 115.465 84.690 115.635 ;
        RECT 85.085 115.295 85.255 115.960 ;
        RECT 86.005 115.715 86.345 116.525 ;
        RECT 86.980 115.965 87.330 116.615 ;
        RECT 87.500 115.795 87.730 116.785 ;
        RECT 83.225 115.125 85.255 115.295 ;
        RECT 85.425 114.955 85.595 115.715 ;
        RECT 85.830 115.305 86.345 115.715 ;
        RECT 87.065 115.625 87.730 115.795 ;
        RECT 87.065 115.125 87.235 115.625 ;
        RECT 87.405 114.955 87.735 115.455 ;
        RECT 87.905 115.125 88.090 117.245 ;
        RECT 88.345 117.045 88.595 117.505 ;
        RECT 88.765 117.055 89.100 117.225 ;
        RECT 89.295 117.055 89.970 117.225 ;
        RECT 88.765 116.915 88.935 117.055 ;
        RECT 88.260 115.925 88.540 116.875 ;
        RECT 88.710 116.785 88.935 116.915 ;
        RECT 88.710 115.680 88.880 116.785 ;
        RECT 89.105 116.635 89.630 116.855 ;
        RECT 89.050 115.870 89.290 116.465 ;
        RECT 89.460 115.935 89.630 116.635 ;
        RECT 89.800 116.275 89.970 117.055 ;
        RECT 90.290 117.005 90.660 117.505 ;
        RECT 90.840 117.055 91.245 117.225 ;
        RECT 91.415 117.055 92.200 117.225 ;
        RECT 90.840 116.825 91.010 117.055 ;
        RECT 90.180 116.525 91.010 116.825 ;
        RECT 91.395 116.555 91.860 116.885 ;
        RECT 90.180 116.495 90.380 116.525 ;
        RECT 90.500 116.275 90.670 116.345 ;
        RECT 89.800 116.105 90.670 116.275 ;
        RECT 90.160 116.015 90.670 116.105 ;
        RECT 88.710 115.550 89.015 115.680 ;
        RECT 89.460 115.570 89.990 115.935 ;
        RECT 88.330 114.955 88.595 115.415 ;
        RECT 88.765 115.125 89.015 115.550 ;
        RECT 90.160 115.400 90.330 116.015 ;
        RECT 89.225 115.230 90.330 115.400 ;
        RECT 90.500 114.955 90.670 115.755 ;
        RECT 90.840 115.455 91.010 116.525 ;
        RECT 91.180 115.625 91.370 116.345 ;
        RECT 91.540 115.595 91.860 116.555 ;
        RECT 92.030 116.595 92.200 117.055 ;
        RECT 92.475 116.975 92.685 117.505 ;
        RECT 92.945 116.765 93.275 117.290 ;
        RECT 93.445 116.895 93.615 117.505 ;
        RECT 93.785 116.850 94.115 117.285 ;
        RECT 94.285 116.990 94.455 117.505 ;
        RECT 93.785 116.765 94.165 116.850 ;
        RECT 94.795 116.780 95.085 117.505 ;
        RECT 93.075 116.595 93.275 116.765 ;
        RECT 93.940 116.725 94.165 116.765 ;
        RECT 92.030 116.265 92.905 116.595 ;
        RECT 93.075 116.265 93.825 116.595 ;
        RECT 90.840 115.125 91.090 115.455 ;
        RECT 92.030 115.425 92.200 116.265 ;
        RECT 93.075 116.060 93.265 116.265 ;
        RECT 93.995 116.145 94.165 116.725 ;
        RECT 93.950 116.095 94.165 116.145 ;
        RECT 95.260 116.765 95.515 117.335 ;
        RECT 95.685 117.105 96.015 117.505 ;
        RECT 96.440 116.970 96.970 117.335 ;
        RECT 96.440 116.935 96.615 116.970 ;
        RECT 95.685 116.765 96.615 116.935 ;
        RECT 92.370 115.685 93.265 116.060 ;
        RECT 93.775 116.015 94.165 116.095 ;
        RECT 91.315 115.255 92.200 115.425 ;
        RECT 92.380 114.955 92.695 115.455 ;
        RECT 92.925 115.125 93.265 115.685 ;
        RECT 93.435 114.955 93.605 115.965 ;
        RECT 93.775 115.170 94.105 116.015 ;
        RECT 94.275 114.955 94.445 115.870 ;
        RECT 94.795 114.955 95.085 116.120 ;
        RECT 95.260 116.095 95.430 116.765 ;
        RECT 95.685 116.595 95.855 116.765 ;
        RECT 95.600 116.265 95.855 116.595 ;
        RECT 96.080 116.265 96.275 116.595 ;
        RECT 95.260 115.125 95.595 116.095 ;
        RECT 95.765 114.955 95.935 116.095 ;
        RECT 96.105 115.295 96.275 116.265 ;
        RECT 96.445 115.635 96.615 116.765 ;
        RECT 96.785 115.975 96.955 116.775 ;
        RECT 97.160 116.485 97.435 117.335 ;
        RECT 97.155 116.315 97.435 116.485 ;
        RECT 97.160 116.175 97.435 116.315 ;
        RECT 97.605 115.975 97.795 117.335 ;
        RECT 97.975 116.970 98.485 117.505 ;
        RECT 98.705 116.695 98.950 117.300 ;
        RECT 99.945 116.955 100.115 117.245 ;
        RECT 100.285 117.125 100.615 117.505 ;
        RECT 99.945 116.785 100.610 116.955 ;
        RECT 97.995 116.525 99.225 116.695 ;
        RECT 96.785 115.805 97.795 115.975 ;
        RECT 97.965 115.960 98.715 116.150 ;
        RECT 96.445 115.465 97.570 115.635 ;
        RECT 97.965 115.295 98.135 115.960 ;
        RECT 98.885 115.715 99.225 116.525 ;
        RECT 99.860 115.965 100.210 116.615 ;
        RECT 100.380 115.795 100.610 116.785 ;
        RECT 96.105 115.125 98.135 115.295 ;
        RECT 98.305 114.955 98.475 115.715 ;
        RECT 98.710 115.305 99.225 115.715 ;
        RECT 99.945 115.625 100.610 115.795 ;
        RECT 99.945 115.125 100.115 115.625 ;
        RECT 100.285 114.955 100.615 115.455 ;
        RECT 100.785 115.125 100.970 117.245 ;
        RECT 101.225 117.045 101.475 117.505 ;
        RECT 101.645 117.055 101.980 117.225 ;
        RECT 102.175 117.055 102.850 117.225 ;
        RECT 101.645 116.915 101.815 117.055 ;
        RECT 101.140 115.925 101.420 116.875 ;
        RECT 101.590 116.785 101.815 116.915 ;
        RECT 101.590 115.680 101.760 116.785 ;
        RECT 101.985 116.635 102.510 116.855 ;
        RECT 101.930 115.870 102.170 116.465 ;
        RECT 102.340 115.935 102.510 116.635 ;
        RECT 102.680 116.275 102.850 117.055 ;
        RECT 103.170 117.005 103.540 117.505 ;
        RECT 103.720 117.055 104.125 117.225 ;
        RECT 104.295 117.055 105.080 117.225 ;
        RECT 103.720 116.825 103.890 117.055 ;
        RECT 103.060 116.525 103.890 116.825 ;
        RECT 104.275 116.555 104.740 116.885 ;
        RECT 103.060 116.495 103.260 116.525 ;
        RECT 103.380 116.275 103.550 116.345 ;
        RECT 102.680 116.105 103.550 116.275 ;
        RECT 103.040 116.015 103.550 116.105 ;
        RECT 101.590 115.550 101.895 115.680 ;
        RECT 102.340 115.570 102.870 115.935 ;
        RECT 101.210 114.955 101.475 115.415 ;
        RECT 101.645 115.125 101.895 115.550 ;
        RECT 103.040 115.400 103.210 116.015 ;
        RECT 102.105 115.230 103.210 115.400 ;
        RECT 103.380 114.955 103.550 115.755 ;
        RECT 103.720 115.455 103.890 116.525 ;
        RECT 104.060 115.625 104.250 116.345 ;
        RECT 104.420 115.595 104.740 116.555 ;
        RECT 104.910 116.595 105.080 117.055 ;
        RECT 105.355 116.975 105.565 117.505 ;
        RECT 105.825 116.765 106.155 117.290 ;
        RECT 106.325 116.895 106.495 117.505 ;
        RECT 106.665 116.850 106.995 117.285 ;
        RECT 107.265 117.035 107.555 117.505 ;
        RECT 107.725 116.865 108.055 117.335 ;
        RECT 108.225 117.035 108.935 117.505 ;
        RECT 109.105 116.865 109.435 117.335 ;
        RECT 109.605 117.035 109.775 117.505 ;
        RECT 109.945 116.865 110.275 117.335 ;
        RECT 106.665 116.765 107.045 116.850 ;
        RECT 105.955 116.595 106.155 116.765 ;
        RECT 106.820 116.725 107.045 116.765 ;
        RECT 104.910 116.265 105.785 116.595 ;
        RECT 105.955 116.265 106.705 116.595 ;
        RECT 103.720 115.125 103.970 115.455 ;
        RECT 104.910 115.425 105.080 116.265 ;
        RECT 105.955 116.060 106.145 116.265 ;
        RECT 106.875 116.145 107.045 116.725 ;
        RECT 106.830 116.095 107.045 116.145 ;
        RECT 105.250 115.685 106.145 116.060 ;
        RECT 106.655 116.015 107.045 116.095 ;
        RECT 107.215 116.685 110.275 116.865 ;
        RECT 110.445 116.685 110.720 117.505 ;
        RECT 110.895 116.960 116.240 117.505 ;
        RECT 107.215 116.135 107.675 116.685 ;
        RECT 107.845 116.305 108.435 116.515 ;
        RECT 108.625 116.305 109.675 116.515 ;
        RECT 109.845 116.305 110.675 116.515 ;
        RECT 104.195 115.255 105.080 115.425 ;
        RECT 105.260 114.955 105.575 115.455 ;
        RECT 105.805 115.125 106.145 115.685 ;
        RECT 106.315 114.955 106.485 115.965 ;
        RECT 106.655 115.170 106.985 116.015 ;
        RECT 107.215 115.965 107.975 116.135 ;
        RECT 108.170 115.965 108.435 116.305 ;
        RECT 108.725 115.965 110.660 116.135 ;
        RECT 112.480 116.130 112.820 116.960 ;
        RECT 116.415 116.735 119.925 117.505 ;
        RECT 120.555 116.780 120.845 117.505 ;
        RECT 121.565 116.955 121.735 117.335 ;
        RECT 121.950 117.125 122.280 117.505 ;
        RECT 121.565 116.785 122.280 116.955 ;
        RECT 107.345 115.295 107.595 115.795 ;
        RECT 107.765 115.465 107.975 115.965 ;
        RECT 108.185 115.295 108.395 115.795 ;
        RECT 108.725 115.465 108.975 115.965 ;
        RECT 109.145 115.295 109.395 115.795 ;
        RECT 107.345 115.125 109.395 115.295 ;
        RECT 109.565 115.125 109.815 115.965 ;
        RECT 109.985 114.955 110.235 115.795 ;
        RECT 110.405 115.125 110.660 115.965 ;
        RECT 114.300 115.390 114.650 116.640 ;
        RECT 116.415 116.215 118.065 116.735 ;
        RECT 118.235 116.045 119.925 116.565 ;
        RECT 121.475 116.235 121.830 116.605 ;
        RECT 122.110 116.595 122.280 116.785 ;
        RECT 122.450 116.760 122.705 117.335 ;
        RECT 122.110 116.265 122.365 116.595 ;
        RECT 110.895 114.955 116.240 115.390 ;
        RECT 116.415 114.955 119.925 116.045 ;
        RECT 120.555 114.955 120.845 116.120 ;
        RECT 122.110 116.055 122.280 116.265 ;
        RECT 121.565 115.885 122.280 116.055 ;
        RECT 122.535 116.030 122.705 116.760 ;
        RECT 122.880 116.665 123.140 117.505 ;
        RECT 123.315 116.735 126.825 117.505 ;
        RECT 123.315 116.215 124.965 116.735 ;
        RECT 127.660 116.725 128.160 117.335 ;
        RECT 121.565 115.125 121.735 115.885 ;
        RECT 121.950 114.955 122.280 115.715 ;
        RECT 122.450 115.125 122.705 116.030 ;
        RECT 122.880 114.955 123.140 116.105 ;
        RECT 125.135 116.045 126.825 116.565 ;
        RECT 127.455 116.265 127.805 116.515 ;
        RECT 127.990 116.095 128.160 116.725 ;
        RECT 128.790 116.855 129.120 117.335 ;
        RECT 129.290 117.045 129.515 117.505 ;
        RECT 129.685 116.855 130.015 117.335 ;
        RECT 128.790 116.685 130.015 116.855 ;
        RECT 130.205 116.705 130.455 117.505 ;
        RECT 130.625 116.705 130.965 117.335 ;
        RECT 131.225 116.955 131.395 117.245 ;
        RECT 131.565 117.125 131.895 117.505 ;
        RECT 131.225 116.785 131.890 116.955 ;
        RECT 130.735 116.655 130.965 116.705 ;
        RECT 128.330 116.315 128.660 116.515 ;
        RECT 128.830 116.315 129.160 116.515 ;
        RECT 129.330 116.315 129.750 116.515 ;
        RECT 129.925 116.345 130.620 116.515 ;
        RECT 129.925 116.095 130.095 116.345 ;
        RECT 130.790 116.095 130.965 116.655 ;
        RECT 123.315 114.955 126.825 116.045 ;
        RECT 127.660 115.925 130.095 116.095 ;
        RECT 127.660 115.125 127.990 115.925 ;
        RECT 128.160 114.955 128.490 115.755 ;
        RECT 128.790 115.125 129.120 115.925 ;
        RECT 129.765 114.955 130.015 115.755 ;
        RECT 130.285 114.955 130.455 116.095 ;
        RECT 130.625 115.125 130.965 116.095 ;
        RECT 131.140 115.965 131.490 116.615 ;
        RECT 131.660 115.795 131.890 116.785 ;
        RECT 131.225 115.625 131.890 115.795 ;
        RECT 131.225 115.125 131.395 115.625 ;
        RECT 131.565 114.955 131.895 115.455 ;
        RECT 132.065 115.125 132.250 117.245 ;
        RECT 132.505 117.045 132.755 117.505 ;
        RECT 132.925 117.055 133.260 117.225 ;
        RECT 133.455 117.055 134.130 117.225 ;
        RECT 132.925 116.915 133.095 117.055 ;
        RECT 132.420 115.925 132.700 116.875 ;
        RECT 132.870 116.785 133.095 116.915 ;
        RECT 132.870 115.680 133.040 116.785 ;
        RECT 133.265 116.635 133.790 116.855 ;
        RECT 133.210 115.870 133.450 116.465 ;
        RECT 133.620 115.935 133.790 116.635 ;
        RECT 133.960 116.275 134.130 117.055 ;
        RECT 134.450 117.005 134.820 117.505 ;
        RECT 135.000 117.055 135.405 117.225 ;
        RECT 135.575 117.055 136.360 117.225 ;
        RECT 135.000 116.825 135.170 117.055 ;
        RECT 134.340 116.525 135.170 116.825 ;
        RECT 135.555 116.555 136.020 116.885 ;
        RECT 134.340 116.495 134.540 116.525 ;
        RECT 134.660 116.275 134.830 116.345 ;
        RECT 133.960 116.105 134.830 116.275 ;
        RECT 134.320 116.015 134.830 116.105 ;
        RECT 132.870 115.550 133.175 115.680 ;
        RECT 133.620 115.570 134.150 115.935 ;
        RECT 132.490 114.955 132.755 115.415 ;
        RECT 132.925 115.125 133.175 115.550 ;
        RECT 134.320 115.400 134.490 116.015 ;
        RECT 133.385 115.230 134.490 115.400 ;
        RECT 134.660 114.955 134.830 115.755 ;
        RECT 135.000 115.455 135.170 116.525 ;
        RECT 135.340 115.625 135.530 116.345 ;
        RECT 135.700 115.595 136.020 116.555 ;
        RECT 136.190 116.595 136.360 117.055 ;
        RECT 136.635 116.975 136.845 117.505 ;
        RECT 137.105 116.765 137.435 117.290 ;
        RECT 137.605 116.895 137.775 117.505 ;
        RECT 137.945 116.850 138.275 117.285 ;
        RECT 137.945 116.765 138.325 116.850 ;
        RECT 137.235 116.595 137.435 116.765 ;
        RECT 138.100 116.725 138.325 116.765 ;
        RECT 136.190 116.265 137.065 116.595 ;
        RECT 137.235 116.265 137.985 116.595 ;
        RECT 135.000 115.125 135.250 115.455 ;
        RECT 136.190 115.425 136.360 116.265 ;
        RECT 137.235 116.060 137.425 116.265 ;
        RECT 138.155 116.145 138.325 116.725 ;
        RECT 138.495 116.735 141.085 117.505 ;
        RECT 141.715 116.755 142.925 117.505 ;
        RECT 138.495 116.215 139.705 116.735 ;
        RECT 138.110 116.095 138.325 116.145 ;
        RECT 136.530 115.685 137.425 116.060 ;
        RECT 137.935 116.015 138.325 116.095 ;
        RECT 139.875 116.045 141.085 116.565 ;
        RECT 135.475 115.255 136.360 115.425 ;
        RECT 136.540 114.955 136.855 115.455 ;
        RECT 137.085 115.125 137.425 115.685 ;
        RECT 137.595 114.955 137.765 115.965 ;
        RECT 137.935 115.170 138.265 116.015 ;
        RECT 138.495 114.955 141.085 116.045 ;
        RECT 141.715 116.045 142.235 116.585 ;
        RECT 142.405 116.215 142.925 116.755 ;
        RECT 141.715 114.955 142.925 116.045 ;
        RECT 17.430 114.785 143.010 114.955 ;
        RECT 17.515 113.695 18.725 114.785 ;
        RECT 18.895 113.695 20.105 114.785 ;
        RECT 20.335 113.725 20.665 114.570 ;
        RECT 20.835 113.775 21.005 114.785 ;
        RECT 21.175 114.055 21.515 114.615 ;
        RECT 21.745 114.285 22.060 114.785 ;
        RECT 22.240 114.315 23.125 114.485 ;
        RECT 17.515 112.985 18.035 113.525 ;
        RECT 18.205 113.155 18.725 113.695 ;
        RECT 18.895 112.985 19.415 113.525 ;
        RECT 19.585 113.155 20.105 113.695 ;
        RECT 20.275 113.645 20.665 113.725 ;
        RECT 21.175 113.680 22.070 114.055 ;
        RECT 20.275 113.595 20.490 113.645 ;
        RECT 20.275 113.015 20.445 113.595 ;
        RECT 21.175 113.475 21.365 113.680 ;
        RECT 22.240 113.475 22.410 114.315 ;
        RECT 23.350 114.285 23.600 114.615 ;
        RECT 20.615 113.145 21.365 113.475 ;
        RECT 21.535 113.145 22.410 113.475 ;
        RECT 17.515 112.235 18.725 112.985 ;
        RECT 18.895 112.235 20.105 112.985 ;
        RECT 20.275 112.975 20.500 113.015 ;
        RECT 21.165 112.975 21.365 113.145 ;
        RECT 20.275 112.890 20.655 112.975 ;
        RECT 20.325 112.455 20.655 112.890 ;
        RECT 20.825 112.235 20.995 112.845 ;
        RECT 21.165 112.450 21.495 112.975 ;
        RECT 21.755 112.235 21.965 112.765 ;
        RECT 22.240 112.685 22.410 113.145 ;
        RECT 22.580 113.185 22.900 114.145 ;
        RECT 23.070 113.395 23.260 114.115 ;
        RECT 23.430 113.215 23.600 114.285 ;
        RECT 23.770 113.985 23.940 114.785 ;
        RECT 24.110 114.340 25.215 114.510 ;
        RECT 24.110 113.725 24.280 114.340 ;
        RECT 25.425 114.190 25.675 114.615 ;
        RECT 25.845 114.325 26.110 114.785 ;
        RECT 24.450 113.805 24.980 114.170 ;
        RECT 25.425 114.060 25.730 114.190 ;
        RECT 23.770 113.635 24.280 113.725 ;
        RECT 23.770 113.465 24.640 113.635 ;
        RECT 23.770 113.395 23.940 113.465 ;
        RECT 24.060 113.215 24.260 113.245 ;
        RECT 22.580 112.855 23.045 113.185 ;
        RECT 23.430 112.915 24.260 113.215 ;
        RECT 23.430 112.685 23.600 112.915 ;
        RECT 22.240 112.515 23.025 112.685 ;
        RECT 23.195 112.515 23.600 112.685 ;
        RECT 23.780 112.235 24.150 112.735 ;
        RECT 24.470 112.685 24.640 113.465 ;
        RECT 24.810 113.105 24.980 113.805 ;
        RECT 25.150 113.275 25.390 113.870 ;
        RECT 24.810 112.885 25.335 113.105 ;
        RECT 25.560 112.955 25.730 114.060 ;
        RECT 25.505 112.825 25.730 112.955 ;
        RECT 25.900 112.865 26.180 113.815 ;
        RECT 25.505 112.685 25.675 112.825 ;
        RECT 24.470 112.515 25.145 112.685 ;
        RECT 25.340 112.515 25.675 112.685 ;
        RECT 25.845 112.235 26.095 112.695 ;
        RECT 26.350 112.495 26.535 114.615 ;
        RECT 26.705 114.285 27.035 114.785 ;
        RECT 27.205 114.115 27.375 114.615 ;
        RECT 26.710 113.945 27.375 114.115 ;
        RECT 26.710 112.955 26.940 113.945 ;
        RECT 27.655 113.895 27.915 114.605 ;
        RECT 28.085 114.075 28.415 114.785 ;
        RECT 28.585 113.895 28.815 114.605 ;
        RECT 27.110 113.125 27.460 113.775 ;
        RECT 27.655 113.655 28.815 113.895 ;
        RECT 28.995 113.875 29.265 114.605 ;
        RECT 29.445 114.055 29.785 114.785 ;
        RECT 28.995 113.655 29.765 113.875 ;
        RECT 27.645 113.145 27.945 113.475 ;
        RECT 28.125 113.165 28.650 113.475 ;
        RECT 28.830 113.165 29.295 113.475 ;
        RECT 26.710 112.785 27.375 112.955 ;
        RECT 26.705 112.235 27.035 112.615 ;
        RECT 27.205 112.495 27.375 112.785 ;
        RECT 27.655 112.235 27.945 112.965 ;
        RECT 28.125 112.525 28.355 113.165 ;
        RECT 29.475 112.985 29.765 113.655 ;
        RECT 28.535 112.785 29.765 112.985 ;
        RECT 28.535 112.415 28.845 112.785 ;
        RECT 29.025 112.235 29.695 112.605 ;
        RECT 29.955 112.415 30.215 114.605 ;
        RECT 30.395 113.620 30.685 114.785 ;
        RECT 30.855 113.695 32.065 114.785 ;
        RECT 30.855 112.985 31.375 113.525 ;
        RECT 31.545 113.155 32.065 113.695 ;
        RECT 32.245 113.675 32.540 114.785 ;
        RECT 32.720 113.475 32.970 114.610 ;
        RECT 33.140 113.675 33.400 114.785 ;
        RECT 33.570 113.885 33.830 114.610 ;
        RECT 34.000 114.055 34.260 114.785 ;
        RECT 34.430 113.885 34.690 114.610 ;
        RECT 34.860 114.055 35.120 114.785 ;
        RECT 35.290 113.885 35.550 114.610 ;
        RECT 35.720 114.055 35.980 114.785 ;
        RECT 36.150 113.885 36.410 114.610 ;
        RECT 36.580 114.055 36.875 114.785 ;
        RECT 37.295 114.355 37.635 114.615 ;
        RECT 33.570 113.645 36.880 113.885 ;
        RECT 30.395 112.235 30.685 112.960 ;
        RECT 30.855 112.235 32.065 112.985 ;
        RECT 32.235 112.865 32.550 113.475 ;
        RECT 32.720 113.225 35.740 113.475 ;
        RECT 32.295 112.235 32.540 112.695 ;
        RECT 32.720 112.415 32.970 113.225 ;
        RECT 35.910 113.055 36.880 113.645 ;
        RECT 33.570 112.885 36.880 113.055 ;
        RECT 37.295 112.955 37.555 114.355 ;
        RECT 37.805 113.985 38.135 114.785 ;
        RECT 38.600 113.815 38.850 114.615 ;
        RECT 39.035 114.065 39.365 114.785 ;
        RECT 39.585 113.815 39.835 114.615 ;
        RECT 40.005 114.405 40.340 114.785 ;
        RECT 37.745 113.645 39.935 113.815 ;
        RECT 37.745 113.475 38.060 113.645 ;
        RECT 37.730 113.225 38.060 113.475 ;
        RECT 33.140 112.235 33.400 112.760 ;
        RECT 33.570 112.430 33.830 112.885 ;
        RECT 34.000 112.235 34.260 112.715 ;
        RECT 34.430 112.430 34.690 112.885 ;
        RECT 34.860 112.235 35.120 112.715 ;
        RECT 35.290 112.430 35.550 112.885 ;
        RECT 35.720 112.235 35.980 112.715 ;
        RECT 36.150 112.430 36.410 112.885 ;
        RECT 36.580 112.235 36.880 112.715 ;
        RECT 37.295 112.445 37.635 112.955 ;
        RECT 37.805 112.235 38.075 113.035 ;
        RECT 38.255 112.505 38.535 113.475 ;
        RECT 38.715 112.505 39.015 113.475 ;
        RECT 39.195 112.510 39.545 113.475 ;
        RECT 39.765 112.735 39.935 113.645 ;
        RECT 40.105 112.915 40.345 114.225 ;
        RECT 40.605 114.165 40.775 114.595 ;
        RECT 40.945 114.335 41.275 114.785 ;
        RECT 40.605 113.935 41.280 114.165 ;
        RECT 40.575 112.915 40.875 113.765 ;
        RECT 41.045 113.285 41.280 113.935 ;
        RECT 41.450 113.625 41.735 114.570 ;
        RECT 41.915 114.315 42.600 114.785 ;
        RECT 41.910 113.795 42.605 114.105 ;
        RECT 42.780 113.730 43.085 114.515 ;
        RECT 41.450 113.475 42.310 113.625 ;
        RECT 41.450 113.455 42.735 113.475 ;
        RECT 41.045 112.955 41.580 113.285 ;
        RECT 41.750 113.095 42.735 113.455 ;
        RECT 41.045 112.805 41.265 112.955 ;
        RECT 39.765 112.405 40.260 112.735 ;
        RECT 40.520 112.235 40.855 112.740 ;
        RECT 41.025 112.430 41.265 112.805 ;
        RECT 41.750 112.760 41.920 113.095 ;
        RECT 42.910 112.925 43.085 113.730 ;
        RECT 41.545 112.565 41.920 112.760 ;
        RECT 41.545 112.420 41.715 112.565 ;
        RECT 42.280 112.235 42.675 112.730 ;
        RECT 42.845 112.405 43.085 112.925 ;
        RECT 43.275 113.180 43.555 114.615 ;
        RECT 43.725 114.010 44.435 114.785 ;
        RECT 44.605 113.840 44.935 114.615 ;
        RECT 43.785 113.625 44.935 113.840 ;
        RECT 43.275 112.405 43.615 113.180 ;
        RECT 43.785 113.055 44.070 113.625 ;
        RECT 44.255 113.225 44.725 113.455 ;
        RECT 45.130 113.425 45.345 114.540 ;
        RECT 45.525 114.065 45.855 114.785 ;
        RECT 46.530 113.985 46.780 114.785 ;
        RECT 46.950 114.155 47.280 114.615 ;
        RECT 47.450 114.325 47.665 114.785 ;
        RECT 48.335 114.350 53.680 114.785 ;
        RECT 46.950 113.985 48.120 114.155 ;
        RECT 46.040 113.815 46.320 113.975 ;
        RECT 45.635 113.425 45.865 113.765 ;
        RECT 46.040 113.645 47.375 113.815 ;
        RECT 47.205 113.475 47.375 113.645 ;
        RECT 44.895 113.245 45.345 113.425 ;
        RECT 44.895 113.225 45.225 113.245 ;
        RECT 45.535 113.225 45.865 113.425 ;
        RECT 46.040 113.225 46.390 113.465 ;
        RECT 46.560 113.225 47.035 113.465 ;
        RECT 47.205 113.225 47.580 113.475 ;
        RECT 47.205 113.055 47.375 113.225 ;
        RECT 43.785 112.865 44.495 113.055 ;
        RECT 44.195 112.725 44.495 112.865 ;
        RECT 44.685 112.865 45.865 113.055 ;
        RECT 44.685 112.785 45.015 112.865 ;
        RECT 44.195 112.715 44.510 112.725 ;
        RECT 44.195 112.705 44.520 112.715 ;
        RECT 44.195 112.700 44.530 112.705 ;
        RECT 43.785 112.235 43.955 112.695 ;
        RECT 44.195 112.690 44.535 112.700 ;
        RECT 44.195 112.685 44.540 112.690 ;
        RECT 44.195 112.675 44.545 112.685 ;
        RECT 44.195 112.670 44.550 112.675 ;
        RECT 44.195 112.405 44.555 112.670 ;
        RECT 45.185 112.235 45.355 112.695 ;
        RECT 45.525 112.405 45.865 112.865 ;
        RECT 46.040 112.885 47.375 113.055 ;
        RECT 46.040 112.675 46.310 112.885 ;
        RECT 47.750 112.695 48.120 113.985 ;
        RECT 49.920 112.780 50.260 113.610 ;
        RECT 51.740 113.100 52.090 114.350 ;
        RECT 53.855 113.695 55.525 114.785 ;
        RECT 53.855 113.005 54.605 113.525 ;
        RECT 54.775 113.175 55.525 113.695 ;
        RECT 56.155 113.620 56.445 114.785 ;
        RECT 56.625 114.175 56.955 114.605 ;
        RECT 57.135 114.345 57.330 114.785 ;
        RECT 57.500 114.175 57.830 114.605 ;
        RECT 56.625 114.005 57.830 114.175 ;
        RECT 56.625 113.675 57.520 114.005 ;
        RECT 58.000 113.835 58.275 114.605 ;
        RECT 58.545 114.115 58.715 114.615 ;
        RECT 58.885 114.285 59.215 114.785 ;
        RECT 58.545 113.945 59.210 114.115 ;
        RECT 57.690 113.645 58.275 113.835 ;
        RECT 56.630 113.145 56.925 113.475 ;
        RECT 57.105 113.145 57.520 113.475 ;
        RECT 46.530 112.235 46.860 112.695 ;
        RECT 47.370 112.405 48.120 112.695 ;
        RECT 48.335 112.235 53.680 112.780 ;
        RECT 53.855 112.235 55.525 113.005 ;
        RECT 56.155 112.235 56.445 112.960 ;
        RECT 56.625 112.235 56.925 112.965 ;
        RECT 57.105 112.525 57.335 113.145 ;
        RECT 57.690 112.975 57.865 113.645 ;
        RECT 57.535 112.795 57.865 112.975 ;
        RECT 58.035 112.825 58.275 113.475 ;
        RECT 58.460 113.125 58.810 113.775 ;
        RECT 58.980 112.955 59.210 113.945 ;
        RECT 57.535 112.415 57.760 112.795 ;
        RECT 58.545 112.785 59.210 112.955 ;
        RECT 57.930 112.235 58.260 112.625 ;
        RECT 58.545 112.495 58.715 112.785 ;
        RECT 58.885 112.235 59.215 112.615 ;
        RECT 59.385 112.495 59.570 114.615 ;
        RECT 59.810 114.325 60.075 114.785 ;
        RECT 60.245 114.190 60.495 114.615 ;
        RECT 60.705 114.340 61.810 114.510 ;
        RECT 60.190 114.060 60.495 114.190 ;
        RECT 59.740 112.865 60.020 113.815 ;
        RECT 60.190 112.955 60.360 114.060 ;
        RECT 60.530 113.275 60.770 113.870 ;
        RECT 60.940 113.805 61.470 114.170 ;
        RECT 60.940 113.105 61.110 113.805 ;
        RECT 61.640 113.725 61.810 114.340 ;
        RECT 61.980 113.985 62.150 114.785 ;
        RECT 62.320 114.285 62.570 114.615 ;
        RECT 62.795 114.315 63.680 114.485 ;
        RECT 61.640 113.635 62.150 113.725 ;
        RECT 60.190 112.825 60.415 112.955 ;
        RECT 60.585 112.885 61.110 113.105 ;
        RECT 61.280 113.465 62.150 113.635 ;
        RECT 59.825 112.235 60.075 112.695 ;
        RECT 60.245 112.685 60.415 112.825 ;
        RECT 61.280 112.685 61.450 113.465 ;
        RECT 61.980 113.395 62.150 113.465 ;
        RECT 61.660 113.215 61.860 113.245 ;
        RECT 62.320 113.215 62.490 114.285 ;
        RECT 62.660 113.395 62.850 114.115 ;
        RECT 61.660 112.915 62.490 113.215 ;
        RECT 63.020 113.185 63.340 114.145 ;
        RECT 60.245 112.515 60.580 112.685 ;
        RECT 60.775 112.515 61.450 112.685 ;
        RECT 61.770 112.235 62.140 112.735 ;
        RECT 62.320 112.685 62.490 112.915 ;
        RECT 62.875 112.855 63.340 113.185 ;
        RECT 63.510 113.475 63.680 114.315 ;
        RECT 63.860 114.285 64.175 114.785 ;
        RECT 64.405 114.055 64.745 114.615 ;
        RECT 63.850 113.680 64.745 114.055 ;
        RECT 64.915 113.775 65.085 114.785 ;
        RECT 64.555 113.475 64.745 113.680 ;
        RECT 65.255 113.725 65.585 114.570 ;
        RECT 65.255 113.645 65.645 113.725 ;
        RECT 65.825 113.675 66.120 114.785 ;
        RECT 65.430 113.595 65.645 113.645 ;
        RECT 63.510 113.145 64.385 113.475 ;
        RECT 64.555 113.145 65.305 113.475 ;
        RECT 63.510 112.685 63.680 113.145 ;
        RECT 64.555 112.975 64.755 113.145 ;
        RECT 65.475 113.015 65.645 113.595 ;
        RECT 66.300 113.475 66.550 114.610 ;
        RECT 66.720 113.675 66.980 114.785 ;
        RECT 67.150 113.885 67.410 114.610 ;
        RECT 67.580 114.055 67.840 114.785 ;
        RECT 68.010 113.885 68.270 114.610 ;
        RECT 68.440 114.055 68.700 114.785 ;
        RECT 68.870 113.885 69.130 114.610 ;
        RECT 69.300 114.055 69.560 114.785 ;
        RECT 69.730 113.885 69.990 114.610 ;
        RECT 70.160 114.055 70.455 114.785 ;
        RECT 70.960 114.165 71.135 114.615 ;
        RECT 71.305 114.345 71.635 114.785 ;
        RECT 71.940 114.195 72.110 114.615 ;
        RECT 72.345 114.375 73.015 114.785 ;
        RECT 73.230 114.195 73.400 114.615 ;
        RECT 73.600 114.375 73.930 114.785 ;
        RECT 70.960 113.995 71.590 114.165 ;
        RECT 67.150 113.645 70.460 113.885 ;
        RECT 65.420 112.975 65.645 113.015 ;
        RECT 62.320 112.515 62.725 112.685 ;
        RECT 62.895 112.515 63.680 112.685 ;
        RECT 63.955 112.235 64.165 112.765 ;
        RECT 64.425 112.450 64.755 112.975 ;
        RECT 65.265 112.890 65.645 112.975 ;
        RECT 64.925 112.235 65.095 112.845 ;
        RECT 65.265 112.455 65.595 112.890 ;
        RECT 65.815 112.865 66.130 113.475 ;
        RECT 66.300 113.225 69.320 113.475 ;
        RECT 65.875 112.235 66.120 112.695 ;
        RECT 66.300 112.415 66.550 113.225 ;
        RECT 69.490 113.055 70.460 113.645 ;
        RECT 70.875 113.145 71.240 113.825 ;
        RECT 71.420 113.475 71.590 113.995 ;
        RECT 71.940 114.025 73.955 114.195 ;
        RECT 71.420 113.145 71.770 113.475 ;
        RECT 67.150 112.885 70.460 113.055 ;
        RECT 71.420 112.975 71.590 113.145 ;
        RECT 66.720 112.235 66.980 112.760 ;
        RECT 67.150 112.430 67.410 112.885 ;
        RECT 67.580 112.235 67.840 112.715 ;
        RECT 68.010 112.430 68.270 112.885 ;
        RECT 68.440 112.235 68.700 112.715 ;
        RECT 68.870 112.430 69.130 112.885 ;
        RECT 69.300 112.235 69.560 112.715 ;
        RECT 69.730 112.430 69.990 112.885 ;
        RECT 70.960 112.805 71.590 112.975 ;
        RECT 70.160 112.235 70.460 112.715 ;
        RECT 70.960 112.405 71.135 112.805 ;
        RECT 71.940 112.735 72.110 114.025 ;
        RECT 71.305 112.235 71.635 112.615 ;
        RECT 71.880 112.405 72.110 112.735 ;
        RECT 72.310 112.570 72.590 113.845 ;
        RECT 72.815 113.765 73.085 113.845 ;
        RECT 72.775 113.595 73.085 113.765 ;
        RECT 72.815 112.570 73.085 113.595 ;
        RECT 73.275 112.815 73.615 113.845 ;
        RECT 73.785 113.475 73.955 114.025 ;
        RECT 74.125 113.645 74.385 114.615 ;
        RECT 73.785 113.145 74.045 113.475 ;
        RECT 74.215 112.955 74.385 113.645 ;
        RECT 73.545 112.235 73.875 112.615 ;
        RECT 74.045 112.490 74.385 112.955 ;
        RECT 74.555 113.645 74.940 114.615 ;
        RECT 75.110 114.325 75.435 114.785 ;
        RECT 75.955 114.155 76.235 114.615 ;
        RECT 75.110 113.935 76.235 114.155 ;
        RECT 74.555 112.975 74.835 113.645 ;
        RECT 75.110 113.475 75.560 113.935 ;
        RECT 76.425 113.765 76.825 114.615 ;
        RECT 77.225 114.325 77.495 114.785 ;
        RECT 77.665 114.155 77.950 114.615 ;
        RECT 78.235 114.275 79.430 114.565 ;
        RECT 75.005 113.145 75.560 113.475 ;
        RECT 75.730 113.205 76.825 113.765 ;
        RECT 75.110 113.035 75.560 113.145 ;
        RECT 74.045 112.445 74.380 112.490 ;
        RECT 74.555 112.405 74.940 112.975 ;
        RECT 75.110 112.865 76.235 113.035 ;
        RECT 75.110 112.235 75.435 112.695 ;
        RECT 75.955 112.405 76.235 112.865 ;
        RECT 76.425 112.405 76.825 113.205 ;
        RECT 76.995 113.935 77.950 114.155 ;
        RECT 78.255 113.935 79.420 114.105 ;
        RECT 79.600 113.985 79.880 114.785 ;
        RECT 76.995 113.035 77.205 113.935 ;
        RECT 77.375 113.205 78.065 113.765 ;
        RECT 78.255 113.645 78.585 113.935 ;
        RECT 79.250 113.815 79.420 113.935 ;
        RECT 78.755 113.475 78.980 113.765 ;
        RECT 79.250 113.645 79.920 113.815 ;
        RECT 80.090 113.645 80.365 114.615 ;
        RECT 79.750 113.475 79.920 113.645 ;
        RECT 78.235 113.145 78.585 113.475 ;
        RECT 78.755 113.145 79.580 113.475 ;
        RECT 79.750 113.145 80.025 113.475 ;
        RECT 76.995 112.865 77.950 113.035 ;
        RECT 79.750 112.975 79.920 113.145 ;
        RECT 77.225 112.235 77.495 112.695 ;
        RECT 77.665 112.405 77.950 112.865 ;
        RECT 78.255 112.805 79.920 112.975 ;
        RECT 80.195 112.910 80.365 113.645 ;
        RECT 80.535 113.580 80.825 114.785 ;
        RECT 81.915 113.620 82.205 114.785 ;
        RECT 82.375 113.645 82.635 114.785 ;
        RECT 82.805 113.635 83.135 114.615 ;
        RECT 83.305 113.645 83.585 114.785 ;
        RECT 83.755 113.695 87.265 114.785 ;
        RECT 87.985 114.115 88.155 114.615 ;
        RECT 88.325 114.285 88.655 114.785 ;
        RECT 87.985 113.945 88.650 114.115 ;
        RECT 82.395 113.225 82.730 113.475 ;
        RECT 82.900 113.085 83.070 113.635 ;
        RECT 83.240 113.205 83.575 113.475 ;
        RECT 78.255 112.455 78.510 112.805 ;
        RECT 78.680 112.235 79.010 112.635 ;
        RECT 79.180 112.455 79.350 112.805 ;
        RECT 79.520 112.235 79.900 112.635 ;
        RECT 80.090 112.565 80.365 112.910 ;
        RECT 80.535 112.235 80.825 113.065 ;
        RECT 82.895 113.035 83.070 113.085 ;
        RECT 81.915 112.235 82.205 112.960 ;
        RECT 82.375 112.405 83.070 113.035 ;
        RECT 83.275 112.235 83.585 113.035 ;
        RECT 83.755 113.005 85.405 113.525 ;
        RECT 85.575 113.175 87.265 113.695 ;
        RECT 87.900 113.125 88.250 113.775 ;
        RECT 83.755 112.235 87.265 113.005 ;
        RECT 88.420 112.955 88.650 113.945 ;
        RECT 87.985 112.785 88.650 112.955 ;
        RECT 87.985 112.495 88.155 112.785 ;
        RECT 88.325 112.235 88.655 112.615 ;
        RECT 88.825 112.495 89.010 114.615 ;
        RECT 89.250 114.325 89.515 114.785 ;
        RECT 89.685 114.190 89.935 114.615 ;
        RECT 90.145 114.340 91.250 114.510 ;
        RECT 89.630 114.060 89.935 114.190 ;
        RECT 89.180 112.865 89.460 113.815 ;
        RECT 89.630 112.955 89.800 114.060 ;
        RECT 89.970 113.275 90.210 113.870 ;
        RECT 90.380 113.805 90.910 114.170 ;
        RECT 90.380 113.105 90.550 113.805 ;
        RECT 91.080 113.725 91.250 114.340 ;
        RECT 91.420 113.985 91.590 114.785 ;
        RECT 91.760 114.285 92.010 114.615 ;
        RECT 92.235 114.315 93.120 114.485 ;
        RECT 91.080 113.635 91.590 113.725 ;
        RECT 89.630 112.825 89.855 112.955 ;
        RECT 90.025 112.885 90.550 113.105 ;
        RECT 90.720 113.465 91.590 113.635 ;
        RECT 89.265 112.235 89.515 112.695 ;
        RECT 89.685 112.685 89.855 112.825 ;
        RECT 90.720 112.685 90.890 113.465 ;
        RECT 91.420 113.395 91.590 113.465 ;
        RECT 91.100 113.215 91.300 113.245 ;
        RECT 91.760 113.215 91.930 114.285 ;
        RECT 92.100 113.395 92.290 114.115 ;
        RECT 91.100 112.915 91.930 113.215 ;
        RECT 92.460 113.185 92.780 114.145 ;
        RECT 89.685 112.515 90.020 112.685 ;
        RECT 90.215 112.515 90.890 112.685 ;
        RECT 91.210 112.235 91.580 112.735 ;
        RECT 91.760 112.685 91.930 112.915 ;
        RECT 92.315 112.855 92.780 113.185 ;
        RECT 92.950 113.475 93.120 114.315 ;
        RECT 93.300 114.285 93.615 114.785 ;
        RECT 93.845 114.055 94.185 114.615 ;
        RECT 93.290 113.680 94.185 114.055 ;
        RECT 94.355 113.775 94.525 114.785 ;
        RECT 93.995 113.475 94.185 113.680 ;
        RECT 94.695 113.725 95.025 114.570 ;
        RECT 95.195 113.870 95.365 114.785 ;
        RECT 95.715 114.350 101.060 114.785 ;
        RECT 94.695 113.645 95.085 113.725 ;
        RECT 94.870 113.595 95.085 113.645 ;
        RECT 92.950 113.145 93.825 113.475 ;
        RECT 93.995 113.145 94.745 113.475 ;
        RECT 92.950 112.685 93.120 113.145 ;
        RECT 93.995 112.975 94.195 113.145 ;
        RECT 94.915 113.015 95.085 113.595 ;
        RECT 94.860 112.975 95.085 113.015 ;
        RECT 91.760 112.515 92.165 112.685 ;
        RECT 92.335 112.515 93.120 112.685 ;
        RECT 93.395 112.235 93.605 112.765 ;
        RECT 93.865 112.450 94.195 112.975 ;
        RECT 94.705 112.890 95.085 112.975 ;
        RECT 94.365 112.235 94.535 112.845 ;
        RECT 94.705 112.455 95.035 112.890 ;
        RECT 97.300 112.780 97.640 113.610 ;
        RECT 99.120 113.100 99.470 114.350 ;
        RECT 101.235 113.695 104.745 114.785 ;
        RECT 101.235 113.005 102.885 113.525 ;
        RECT 103.055 113.175 104.745 113.695 ;
        RECT 105.895 113.645 106.105 114.785 ;
        RECT 106.275 113.635 106.605 114.615 ;
        RECT 106.775 113.645 107.005 114.785 ;
        RECT 95.205 112.235 95.375 112.750 ;
        RECT 95.715 112.235 101.060 112.780 ;
        RECT 101.235 112.235 104.745 113.005 ;
        RECT 105.895 112.235 106.105 113.055 ;
        RECT 106.275 113.035 106.525 113.635 ;
        RECT 107.675 113.620 107.965 114.785 ;
        RECT 108.135 114.280 108.765 114.785 ;
        RECT 108.150 113.745 108.405 114.110 ;
        RECT 108.575 114.105 108.765 114.280 ;
        RECT 108.945 114.275 109.420 114.615 ;
        RECT 108.575 113.915 108.905 114.105 ;
        RECT 109.130 113.745 109.380 114.040 ;
        RECT 109.605 113.940 109.820 114.785 ;
        RECT 110.020 113.945 110.295 114.615 ;
        RECT 108.150 113.575 109.940 113.745 ;
        RECT 110.125 113.595 110.295 113.945 ;
        RECT 110.465 113.775 110.725 114.785 ;
        RECT 110.895 113.695 113.485 114.785 ;
        RECT 106.695 113.225 107.025 113.475 ;
        RECT 106.275 112.405 106.605 113.035 ;
        RECT 106.775 112.235 107.005 113.055 ;
        RECT 107.675 112.235 107.965 112.960 ;
        RECT 108.135 112.915 108.520 113.395 ;
        RECT 108.690 112.720 108.945 113.575 ;
        RECT 108.155 112.455 108.945 112.720 ;
        RECT 109.115 112.900 109.525 113.395 ;
        RECT 109.710 113.145 109.940 113.575 ;
        RECT 110.110 113.075 110.725 113.595 ;
        RECT 109.115 112.455 109.345 112.900 ;
        RECT 110.110 112.865 110.280 113.075 ;
        RECT 110.895 113.005 112.105 113.525 ;
        RECT 112.275 113.175 113.485 113.695 ;
        RECT 113.655 113.645 113.995 114.615 ;
        RECT 114.165 113.645 114.335 114.785 ;
        RECT 114.605 113.985 114.855 114.785 ;
        RECT 115.500 113.815 115.830 114.615 ;
        RECT 116.130 113.985 116.460 114.785 ;
        RECT 116.630 113.815 116.960 114.615 ;
        RECT 117.425 114.115 117.595 114.615 ;
        RECT 117.765 114.285 118.095 114.785 ;
        RECT 117.425 113.945 118.090 114.115 ;
        RECT 114.525 113.645 116.960 113.815 ;
        RECT 113.655 113.085 113.830 113.645 ;
        RECT 114.525 113.395 114.695 113.645 ;
        RECT 114.000 113.225 114.695 113.395 ;
        RECT 114.870 113.225 115.290 113.425 ;
        RECT 115.460 113.225 115.790 113.425 ;
        RECT 115.960 113.225 116.290 113.425 ;
        RECT 113.655 113.035 113.885 113.085 ;
        RECT 109.525 112.235 109.855 112.730 ;
        RECT 110.030 112.405 110.280 112.865 ;
        RECT 110.450 112.235 110.725 112.895 ;
        RECT 110.895 112.235 113.485 113.005 ;
        RECT 113.655 112.405 113.995 113.035 ;
        RECT 114.165 112.235 114.415 113.035 ;
        RECT 114.605 112.885 115.830 113.055 ;
        RECT 114.605 112.405 114.935 112.885 ;
        RECT 115.105 112.235 115.330 112.695 ;
        RECT 115.500 112.405 115.830 112.885 ;
        RECT 116.460 113.015 116.630 113.645 ;
        RECT 116.815 113.225 117.165 113.475 ;
        RECT 117.340 113.125 117.690 113.775 ;
        RECT 116.460 112.405 116.960 113.015 ;
        RECT 117.860 112.955 118.090 113.945 ;
        RECT 117.425 112.785 118.090 112.955 ;
        RECT 117.425 112.495 117.595 112.785 ;
        RECT 117.765 112.235 118.095 112.615 ;
        RECT 118.265 112.495 118.450 114.615 ;
        RECT 118.690 114.325 118.955 114.785 ;
        RECT 119.125 114.190 119.375 114.615 ;
        RECT 119.585 114.340 120.690 114.510 ;
        RECT 119.070 114.060 119.375 114.190 ;
        RECT 118.620 112.865 118.900 113.815 ;
        RECT 119.070 112.955 119.240 114.060 ;
        RECT 119.410 113.275 119.650 113.870 ;
        RECT 119.820 113.805 120.350 114.170 ;
        RECT 119.820 113.105 119.990 113.805 ;
        RECT 120.520 113.725 120.690 114.340 ;
        RECT 120.860 113.985 121.030 114.785 ;
        RECT 121.200 114.285 121.450 114.615 ;
        RECT 121.675 114.315 122.560 114.485 ;
        RECT 120.520 113.635 121.030 113.725 ;
        RECT 119.070 112.825 119.295 112.955 ;
        RECT 119.465 112.885 119.990 113.105 ;
        RECT 120.160 113.465 121.030 113.635 ;
        RECT 118.705 112.235 118.955 112.695 ;
        RECT 119.125 112.685 119.295 112.825 ;
        RECT 120.160 112.685 120.330 113.465 ;
        RECT 120.860 113.395 121.030 113.465 ;
        RECT 120.540 113.215 120.740 113.245 ;
        RECT 121.200 113.215 121.370 114.285 ;
        RECT 121.540 113.395 121.730 114.115 ;
        RECT 120.540 112.915 121.370 113.215 ;
        RECT 121.900 113.185 122.220 114.145 ;
        RECT 119.125 112.515 119.460 112.685 ;
        RECT 119.655 112.515 120.330 112.685 ;
        RECT 120.650 112.235 121.020 112.735 ;
        RECT 121.200 112.685 121.370 112.915 ;
        RECT 121.755 112.855 122.220 113.185 ;
        RECT 122.390 113.475 122.560 114.315 ;
        RECT 122.740 114.285 123.055 114.785 ;
        RECT 123.285 114.055 123.625 114.615 ;
        RECT 122.730 113.680 123.625 114.055 ;
        RECT 123.795 113.775 123.965 114.785 ;
        RECT 123.435 113.475 123.625 113.680 ;
        RECT 124.135 113.725 124.465 114.570 ;
        RECT 124.730 113.995 125.265 114.615 ;
        RECT 124.135 113.645 124.525 113.725 ;
        RECT 124.310 113.595 124.525 113.645 ;
        RECT 122.390 113.145 123.265 113.475 ;
        RECT 123.435 113.145 124.185 113.475 ;
        RECT 122.390 112.685 122.560 113.145 ;
        RECT 123.435 112.975 123.635 113.145 ;
        RECT 124.355 113.015 124.525 113.595 ;
        RECT 124.300 112.975 124.525 113.015 ;
        RECT 121.200 112.515 121.605 112.685 ;
        RECT 121.775 112.515 122.560 112.685 ;
        RECT 122.835 112.235 123.045 112.765 ;
        RECT 123.305 112.450 123.635 112.975 ;
        RECT 124.145 112.890 124.525 112.975 ;
        RECT 124.730 112.975 125.045 113.995 ;
        RECT 125.435 113.985 125.765 114.785 ;
        RECT 126.995 114.350 132.340 114.785 ;
        RECT 126.250 113.815 126.640 113.990 ;
        RECT 125.215 113.645 126.640 113.815 ;
        RECT 125.215 113.145 125.385 113.645 ;
        RECT 123.805 112.235 123.975 112.845 ;
        RECT 124.145 112.455 124.475 112.890 ;
        RECT 124.730 112.405 125.345 112.975 ;
        RECT 125.635 112.915 125.900 113.475 ;
        RECT 126.070 112.745 126.240 113.645 ;
        RECT 126.410 112.915 126.765 113.475 ;
        RECT 128.580 112.780 128.920 113.610 ;
        RECT 130.400 113.100 130.750 114.350 ;
        RECT 133.435 113.620 133.725 114.785 ;
        RECT 134.080 113.815 134.470 113.990 ;
        RECT 134.955 113.985 135.285 114.785 ;
        RECT 135.455 113.995 135.990 114.615 ;
        RECT 134.080 113.645 135.505 113.815 ;
        RECT 125.515 112.235 125.730 112.745 ;
        RECT 125.960 112.415 126.240 112.745 ;
        RECT 126.420 112.235 126.660 112.745 ;
        RECT 126.995 112.235 132.340 112.780 ;
        RECT 133.435 112.235 133.725 112.960 ;
        RECT 133.955 112.915 134.310 113.475 ;
        RECT 134.480 112.745 134.650 113.645 ;
        RECT 134.820 112.915 135.085 113.475 ;
        RECT 135.335 113.145 135.505 113.645 ;
        RECT 135.675 112.975 135.990 113.995 ;
        RECT 134.060 112.235 134.300 112.745 ;
        RECT 134.480 112.415 134.760 112.745 ;
        RECT 134.990 112.235 135.205 112.745 ;
        RECT 135.375 112.405 135.990 112.975 ;
        RECT 136.230 113.995 136.765 114.615 ;
        RECT 136.230 112.975 136.545 113.995 ;
        RECT 136.935 113.985 137.265 114.785 ;
        RECT 137.750 113.815 138.140 113.990 ;
        RECT 136.715 113.645 138.140 113.815 ;
        RECT 138.495 113.695 139.705 114.785 ;
        RECT 136.715 113.145 136.885 113.645 ;
        RECT 136.230 112.405 136.845 112.975 ;
        RECT 137.135 112.915 137.400 113.475 ;
        RECT 137.570 112.745 137.740 113.645 ;
        RECT 137.910 112.915 138.265 113.475 ;
        RECT 138.495 112.985 139.015 113.525 ;
        RECT 139.185 113.155 139.705 113.695 ;
        RECT 139.965 113.855 140.135 114.615 ;
        RECT 140.350 114.025 140.680 114.785 ;
        RECT 139.965 113.685 140.680 113.855 ;
        RECT 140.850 113.710 141.105 114.615 ;
        RECT 139.875 113.135 140.230 113.505 ;
        RECT 140.510 113.475 140.680 113.685 ;
        RECT 140.510 113.145 140.765 113.475 ;
        RECT 137.015 112.235 137.230 112.745 ;
        RECT 137.460 112.415 137.740 112.745 ;
        RECT 137.920 112.235 138.160 112.745 ;
        RECT 138.495 112.235 139.705 112.985 ;
        RECT 140.510 112.955 140.680 113.145 ;
        RECT 140.935 112.980 141.105 113.710 ;
        RECT 141.280 113.635 141.540 114.785 ;
        RECT 141.715 113.695 142.925 114.785 ;
        RECT 141.715 113.155 142.235 113.695 ;
        RECT 139.965 112.785 140.680 112.955 ;
        RECT 139.965 112.405 140.135 112.785 ;
        RECT 140.350 112.235 140.680 112.615 ;
        RECT 140.850 112.405 141.105 112.980 ;
        RECT 141.280 112.235 141.540 113.075 ;
        RECT 142.405 112.985 142.925 113.525 ;
        RECT 141.715 112.235 142.925 112.985 ;
        RECT 17.430 112.065 143.010 112.235 ;
        RECT 17.515 111.315 18.725 112.065 ;
        RECT 17.515 110.775 18.035 111.315 ;
        RECT 18.895 111.295 20.565 112.065 ;
        RECT 20.770 111.325 21.385 111.895 ;
        RECT 21.555 111.555 21.770 112.065 ;
        RECT 22.000 111.555 22.280 111.885 ;
        RECT 22.460 111.555 22.700 112.065 ;
        RECT 18.205 110.605 18.725 111.145 ;
        RECT 18.895 110.775 19.645 111.295 ;
        RECT 19.815 110.605 20.565 111.125 ;
        RECT 17.515 109.515 18.725 110.605 ;
        RECT 18.895 109.515 20.565 110.605 ;
        RECT 20.770 110.305 21.085 111.325 ;
        RECT 21.255 110.655 21.425 111.155 ;
        RECT 21.675 110.825 21.940 111.385 ;
        RECT 22.110 110.655 22.280 111.555 ;
        RECT 22.450 110.825 22.805 111.385 ;
        RECT 23.035 111.245 23.295 112.065 ;
        RECT 23.465 111.245 23.795 111.665 ;
        RECT 23.975 111.580 24.765 111.845 ;
        RECT 23.545 111.155 23.795 111.245 ;
        RECT 21.255 110.485 22.680 110.655 ;
        RECT 20.770 109.685 21.305 110.305 ;
        RECT 21.475 109.515 21.805 110.315 ;
        RECT 22.290 110.310 22.680 110.485 ;
        RECT 23.035 110.195 23.375 111.075 ;
        RECT 23.545 110.905 24.340 111.155 ;
        RECT 23.035 109.515 23.295 110.025 ;
        RECT 23.545 109.685 23.715 110.905 ;
        RECT 24.510 110.725 24.765 111.580 ;
        RECT 24.935 111.425 25.135 111.845 ;
        RECT 25.325 111.605 25.655 112.065 ;
        RECT 24.935 110.905 25.345 111.425 ;
        RECT 25.825 111.415 26.085 111.895 ;
        RECT 25.515 110.725 25.745 111.155 ;
        RECT 23.955 110.555 25.745 110.725 ;
        RECT 23.955 110.190 24.205 110.555 ;
        RECT 24.375 110.195 24.705 110.385 ;
        RECT 24.925 110.260 25.640 110.555 ;
        RECT 25.915 110.385 26.085 111.415 ;
        RECT 26.345 111.515 26.515 111.805 ;
        RECT 26.685 111.685 27.015 112.065 ;
        RECT 26.345 111.345 27.010 111.515 ;
        RECT 26.260 110.525 26.610 111.175 ;
        RECT 24.375 110.020 24.570 110.195 ;
        RECT 23.955 109.515 24.570 110.020 ;
        RECT 24.740 109.685 25.215 110.025 ;
        RECT 25.385 109.515 25.600 110.060 ;
        RECT 25.810 109.685 26.085 110.385 ;
        RECT 26.780 110.355 27.010 111.345 ;
        RECT 26.345 110.185 27.010 110.355 ;
        RECT 26.345 109.685 26.515 110.185 ;
        RECT 26.685 109.515 27.015 110.015 ;
        RECT 27.185 109.685 27.370 111.805 ;
        RECT 27.625 111.605 27.875 112.065 ;
        RECT 28.045 111.615 28.380 111.785 ;
        RECT 28.575 111.615 29.250 111.785 ;
        RECT 28.045 111.475 28.215 111.615 ;
        RECT 27.540 110.485 27.820 111.435 ;
        RECT 27.990 111.345 28.215 111.475 ;
        RECT 27.990 110.240 28.160 111.345 ;
        RECT 28.385 111.195 28.910 111.415 ;
        RECT 28.330 110.430 28.570 111.025 ;
        RECT 28.740 110.495 28.910 111.195 ;
        RECT 29.080 110.835 29.250 111.615 ;
        RECT 29.570 111.565 29.940 112.065 ;
        RECT 30.120 111.615 30.525 111.785 ;
        RECT 30.695 111.615 31.480 111.785 ;
        RECT 30.120 111.385 30.290 111.615 ;
        RECT 29.460 111.085 30.290 111.385 ;
        RECT 30.675 111.115 31.140 111.445 ;
        RECT 29.460 111.055 29.660 111.085 ;
        RECT 29.780 110.835 29.950 110.905 ;
        RECT 29.080 110.665 29.950 110.835 ;
        RECT 29.440 110.575 29.950 110.665 ;
        RECT 27.990 110.110 28.295 110.240 ;
        RECT 28.740 110.130 29.270 110.495 ;
        RECT 27.610 109.515 27.875 109.975 ;
        RECT 28.045 109.685 28.295 110.110 ;
        RECT 29.440 109.960 29.610 110.575 ;
        RECT 28.505 109.790 29.610 109.960 ;
        RECT 29.780 109.515 29.950 110.315 ;
        RECT 30.120 110.015 30.290 111.085 ;
        RECT 30.460 110.185 30.650 110.905 ;
        RECT 30.820 110.155 31.140 111.115 ;
        RECT 31.310 111.155 31.480 111.615 ;
        RECT 31.755 111.535 31.965 112.065 ;
        RECT 32.225 111.325 32.555 111.850 ;
        RECT 32.725 111.455 32.895 112.065 ;
        RECT 33.065 111.410 33.395 111.845 ;
        RECT 33.780 111.555 34.020 112.065 ;
        RECT 34.200 111.555 34.480 111.885 ;
        RECT 34.710 111.555 34.925 112.065 ;
        RECT 33.065 111.325 33.445 111.410 ;
        RECT 32.355 111.155 32.555 111.325 ;
        RECT 33.220 111.285 33.445 111.325 ;
        RECT 31.310 110.825 32.185 111.155 ;
        RECT 32.355 110.825 33.105 111.155 ;
        RECT 30.120 109.685 30.370 110.015 ;
        RECT 31.310 109.985 31.480 110.825 ;
        RECT 32.355 110.620 32.545 110.825 ;
        RECT 33.275 110.705 33.445 111.285 ;
        RECT 33.675 110.825 34.030 111.385 ;
        RECT 33.230 110.655 33.445 110.705 ;
        RECT 34.200 110.655 34.370 111.555 ;
        RECT 34.540 110.825 34.805 111.385 ;
        RECT 35.095 111.325 35.710 111.895 ;
        RECT 36.005 111.515 36.175 111.805 ;
        RECT 36.345 111.685 36.675 112.065 ;
        RECT 36.005 111.345 36.670 111.515 ;
        RECT 35.055 110.655 35.225 111.155 ;
        RECT 31.650 110.245 32.545 110.620 ;
        RECT 33.055 110.575 33.445 110.655 ;
        RECT 30.595 109.815 31.480 109.985 ;
        RECT 31.660 109.515 31.975 110.015 ;
        RECT 32.205 109.685 32.545 110.245 ;
        RECT 32.715 109.515 32.885 110.525 ;
        RECT 33.055 109.730 33.385 110.575 ;
        RECT 33.800 110.485 35.225 110.655 ;
        RECT 33.800 110.310 34.190 110.485 ;
        RECT 34.675 109.515 35.005 110.315 ;
        RECT 35.395 110.305 35.710 111.325 ;
        RECT 35.920 110.525 36.270 111.175 ;
        RECT 36.440 110.355 36.670 111.345 ;
        RECT 35.175 109.685 35.710 110.305 ;
        RECT 36.005 110.185 36.670 110.355 ;
        RECT 36.005 109.685 36.175 110.185 ;
        RECT 36.345 109.515 36.675 110.015 ;
        RECT 36.845 109.685 37.030 111.805 ;
        RECT 37.285 111.605 37.535 112.065 ;
        RECT 37.705 111.615 38.040 111.785 ;
        RECT 38.235 111.615 38.910 111.785 ;
        RECT 37.705 111.475 37.875 111.615 ;
        RECT 37.200 110.485 37.480 111.435 ;
        RECT 37.650 111.345 37.875 111.475 ;
        RECT 37.650 110.240 37.820 111.345 ;
        RECT 38.045 111.195 38.570 111.415 ;
        RECT 37.990 110.430 38.230 111.025 ;
        RECT 38.400 110.495 38.570 111.195 ;
        RECT 38.740 110.835 38.910 111.615 ;
        RECT 39.230 111.565 39.600 112.065 ;
        RECT 39.780 111.615 40.185 111.785 ;
        RECT 40.355 111.615 41.140 111.785 ;
        RECT 39.780 111.385 39.950 111.615 ;
        RECT 39.120 111.085 39.950 111.385 ;
        RECT 40.335 111.115 40.800 111.445 ;
        RECT 39.120 111.055 39.320 111.085 ;
        RECT 39.440 110.835 39.610 110.905 ;
        RECT 38.740 110.665 39.610 110.835 ;
        RECT 39.100 110.575 39.610 110.665 ;
        RECT 37.650 110.110 37.955 110.240 ;
        RECT 38.400 110.130 38.930 110.495 ;
        RECT 37.270 109.515 37.535 109.975 ;
        RECT 37.705 109.685 37.955 110.110 ;
        RECT 39.100 109.960 39.270 110.575 ;
        RECT 38.165 109.790 39.270 109.960 ;
        RECT 39.440 109.515 39.610 110.315 ;
        RECT 39.780 110.015 39.950 111.085 ;
        RECT 40.120 110.185 40.310 110.905 ;
        RECT 40.480 110.155 40.800 111.115 ;
        RECT 40.970 111.155 41.140 111.615 ;
        RECT 41.415 111.535 41.625 112.065 ;
        RECT 41.885 111.325 42.215 111.850 ;
        RECT 42.385 111.455 42.555 112.065 ;
        RECT 42.725 111.410 43.055 111.845 ;
        RECT 42.725 111.325 43.105 111.410 ;
        RECT 43.275 111.340 43.565 112.065 ;
        RECT 42.015 111.155 42.215 111.325 ;
        RECT 42.880 111.285 43.105 111.325 ;
        RECT 40.970 110.825 41.845 111.155 ;
        RECT 42.015 110.825 42.765 111.155 ;
        RECT 39.780 109.685 40.030 110.015 ;
        RECT 40.970 109.985 41.140 110.825 ;
        RECT 42.015 110.620 42.205 110.825 ;
        RECT 42.935 110.705 43.105 111.285 ;
        RECT 42.890 110.655 43.105 110.705 ;
        RECT 43.735 111.120 44.075 111.895 ;
        RECT 44.245 111.605 44.415 112.065 ;
        RECT 44.655 111.630 45.015 111.895 ;
        RECT 44.655 111.625 45.010 111.630 ;
        RECT 44.655 111.615 45.005 111.625 ;
        RECT 44.655 111.610 45.000 111.615 ;
        RECT 44.655 111.600 44.995 111.610 ;
        RECT 45.645 111.605 45.815 112.065 ;
        RECT 44.655 111.595 44.990 111.600 ;
        RECT 44.655 111.585 44.980 111.595 ;
        RECT 44.655 111.575 44.970 111.585 ;
        RECT 44.655 111.435 44.955 111.575 ;
        RECT 44.245 111.245 44.955 111.435 ;
        RECT 45.145 111.435 45.475 111.515 ;
        RECT 45.985 111.435 46.325 111.895 ;
        RECT 45.145 111.245 46.325 111.435 ;
        RECT 46.695 111.435 47.025 111.795 ;
        RECT 47.645 111.605 47.895 112.065 ;
        RECT 48.065 111.605 48.625 111.895 ;
        RECT 46.695 111.245 48.085 111.435 ;
        RECT 41.310 110.245 42.205 110.620 ;
        RECT 42.715 110.575 43.105 110.655 ;
        RECT 40.255 109.815 41.140 109.985 ;
        RECT 41.320 109.515 41.635 110.015 ;
        RECT 41.865 109.685 42.205 110.245 ;
        RECT 42.375 109.515 42.545 110.525 ;
        RECT 42.715 109.730 43.045 110.575 ;
        RECT 43.275 109.515 43.565 110.680 ;
        RECT 43.735 109.685 44.015 111.120 ;
        RECT 44.245 110.675 44.530 111.245 ;
        RECT 47.915 111.155 48.085 111.245 ;
        RECT 44.715 110.845 45.185 111.075 ;
        RECT 45.355 111.055 45.685 111.075 ;
        RECT 45.355 110.875 45.805 111.055 ;
        RECT 45.995 110.875 46.325 111.075 ;
        RECT 44.245 110.460 45.395 110.675 ;
        RECT 44.185 109.515 44.895 110.290 ;
        RECT 45.065 109.685 45.395 110.460 ;
        RECT 45.590 109.760 45.805 110.875 ;
        RECT 46.095 110.535 46.325 110.875 ;
        RECT 46.510 110.825 47.185 111.075 ;
        RECT 47.405 110.825 47.745 111.075 ;
        RECT 47.915 110.825 48.205 111.155 ;
        RECT 46.510 110.465 46.775 110.825 ;
        RECT 47.915 110.575 48.085 110.825 ;
        RECT 47.145 110.405 48.085 110.575 ;
        RECT 45.985 109.515 46.315 110.235 ;
        RECT 46.695 109.515 46.975 110.185 ;
        RECT 47.145 109.855 47.445 110.405 ;
        RECT 48.375 110.235 48.625 111.605 ;
        RECT 48.795 111.295 50.465 112.065 ;
        RECT 51.105 111.335 51.405 112.065 ;
        RECT 48.795 110.775 49.545 111.295 ;
        RECT 51.585 111.155 51.815 111.775 ;
        RECT 52.015 111.505 52.240 111.885 ;
        RECT 52.410 111.675 52.740 112.065 ;
        RECT 53.025 111.515 53.195 111.805 ;
        RECT 53.365 111.685 53.695 112.065 ;
        RECT 52.015 111.325 52.345 111.505 ;
        RECT 49.715 110.605 50.465 111.125 ;
        RECT 51.110 110.825 51.405 111.155 ;
        RECT 51.585 110.825 52.000 111.155 ;
        RECT 52.170 110.655 52.345 111.325 ;
        RECT 52.515 110.825 52.755 111.475 ;
        RECT 53.025 111.345 53.690 111.515 ;
        RECT 47.645 109.515 47.975 110.235 ;
        RECT 48.165 109.685 48.625 110.235 ;
        RECT 48.795 109.515 50.465 110.605 ;
        RECT 51.105 110.295 52.000 110.625 ;
        RECT 52.170 110.465 52.755 110.655 ;
        RECT 52.940 110.525 53.290 111.175 ;
        RECT 51.105 110.125 52.310 110.295 ;
        RECT 51.105 109.695 51.435 110.125 ;
        RECT 51.615 109.515 51.810 109.955 ;
        RECT 51.980 109.695 52.310 110.125 ;
        RECT 52.480 109.695 52.755 110.465 ;
        RECT 53.460 110.355 53.690 111.345 ;
        RECT 53.025 110.185 53.690 110.355 ;
        RECT 53.025 109.685 53.195 110.185 ;
        RECT 53.365 109.515 53.695 110.015 ;
        RECT 53.865 109.685 54.050 111.805 ;
        RECT 54.305 111.605 54.555 112.065 ;
        RECT 54.725 111.615 55.060 111.785 ;
        RECT 55.255 111.615 55.930 111.785 ;
        RECT 54.725 111.475 54.895 111.615 ;
        RECT 54.220 110.485 54.500 111.435 ;
        RECT 54.670 111.345 54.895 111.475 ;
        RECT 54.670 110.240 54.840 111.345 ;
        RECT 55.065 111.195 55.590 111.415 ;
        RECT 55.010 110.430 55.250 111.025 ;
        RECT 55.420 110.495 55.590 111.195 ;
        RECT 55.760 110.835 55.930 111.615 ;
        RECT 56.250 111.565 56.620 112.065 ;
        RECT 56.800 111.615 57.205 111.785 ;
        RECT 57.375 111.615 58.160 111.785 ;
        RECT 56.800 111.385 56.970 111.615 ;
        RECT 56.140 111.085 56.970 111.385 ;
        RECT 57.355 111.115 57.820 111.445 ;
        RECT 56.140 111.055 56.340 111.085 ;
        RECT 56.460 110.835 56.630 110.905 ;
        RECT 55.760 110.665 56.630 110.835 ;
        RECT 56.120 110.575 56.630 110.665 ;
        RECT 54.670 110.110 54.975 110.240 ;
        RECT 55.420 110.130 55.950 110.495 ;
        RECT 54.290 109.515 54.555 109.975 ;
        RECT 54.725 109.685 54.975 110.110 ;
        RECT 56.120 109.960 56.290 110.575 ;
        RECT 55.185 109.790 56.290 109.960 ;
        RECT 56.460 109.515 56.630 110.315 ;
        RECT 56.800 110.015 56.970 111.085 ;
        RECT 57.140 110.185 57.330 110.905 ;
        RECT 57.500 110.155 57.820 111.115 ;
        RECT 57.990 111.155 58.160 111.615 ;
        RECT 58.435 111.535 58.645 112.065 ;
        RECT 58.905 111.325 59.235 111.850 ;
        RECT 59.405 111.455 59.575 112.065 ;
        RECT 59.745 111.410 60.075 111.845 ;
        RECT 60.355 111.605 60.600 112.065 ;
        RECT 59.745 111.325 60.125 111.410 ;
        RECT 59.035 111.155 59.235 111.325 ;
        RECT 59.900 111.285 60.125 111.325 ;
        RECT 57.990 110.825 58.865 111.155 ;
        RECT 59.035 110.825 59.785 111.155 ;
        RECT 56.800 109.685 57.050 110.015 ;
        RECT 57.990 109.985 58.160 110.825 ;
        RECT 59.035 110.620 59.225 110.825 ;
        RECT 59.955 110.705 60.125 111.285 ;
        RECT 60.295 110.825 60.610 111.435 ;
        RECT 60.780 111.075 61.030 111.885 ;
        RECT 61.200 111.540 61.460 112.065 ;
        RECT 61.630 111.415 61.890 111.870 ;
        RECT 62.060 111.585 62.320 112.065 ;
        RECT 62.490 111.415 62.750 111.870 ;
        RECT 62.920 111.585 63.180 112.065 ;
        RECT 63.350 111.415 63.610 111.870 ;
        RECT 63.780 111.585 64.040 112.065 ;
        RECT 64.210 111.415 64.470 111.870 ;
        RECT 64.640 111.585 64.940 112.065 ;
        RECT 65.470 111.435 65.755 111.895 ;
        RECT 65.925 111.605 66.195 112.065 ;
        RECT 61.630 111.245 64.940 111.415 ;
        RECT 65.470 111.265 66.425 111.435 ;
        RECT 60.780 110.825 63.800 111.075 ;
        RECT 59.910 110.655 60.125 110.705 ;
        RECT 58.330 110.245 59.225 110.620 ;
        RECT 59.735 110.575 60.125 110.655 ;
        RECT 57.275 109.815 58.160 109.985 ;
        RECT 58.340 109.515 58.655 110.015 ;
        RECT 58.885 109.685 59.225 110.245 ;
        RECT 59.395 109.515 59.565 110.525 ;
        RECT 59.735 109.730 60.065 110.575 ;
        RECT 60.305 109.515 60.600 110.625 ;
        RECT 60.780 109.690 61.030 110.825 ;
        RECT 63.970 110.655 64.940 111.245 ;
        RECT 61.200 109.515 61.460 110.625 ;
        RECT 61.630 110.415 64.940 110.655 ;
        RECT 65.355 110.535 66.045 111.095 ;
        RECT 61.630 109.690 61.890 110.415 ;
        RECT 62.060 109.515 62.320 110.245 ;
        RECT 62.490 109.690 62.750 110.415 ;
        RECT 62.920 109.515 63.180 110.245 ;
        RECT 63.350 109.690 63.610 110.415 ;
        RECT 63.780 109.515 64.040 110.245 ;
        RECT 64.210 109.690 64.470 110.415 ;
        RECT 66.215 110.365 66.425 111.265 ;
        RECT 64.640 109.515 64.935 110.245 ;
        RECT 65.470 110.145 66.425 110.365 ;
        RECT 66.595 111.095 66.995 111.895 ;
        RECT 67.185 111.435 67.465 111.895 ;
        RECT 67.985 111.605 68.310 112.065 ;
        RECT 67.185 111.265 68.310 111.435 ;
        RECT 68.480 111.325 68.865 111.895 ;
        RECT 69.035 111.340 69.325 112.065 ;
        RECT 69.585 111.515 69.755 111.805 ;
        RECT 69.925 111.685 70.255 112.065 ;
        RECT 69.585 111.345 70.250 111.515 ;
        RECT 67.860 111.155 68.310 111.265 ;
        RECT 66.595 110.535 67.690 111.095 ;
        RECT 67.860 110.825 68.415 111.155 ;
        RECT 65.470 109.685 65.755 110.145 ;
        RECT 65.925 109.515 66.195 109.975 ;
        RECT 66.595 109.685 66.995 110.535 ;
        RECT 67.860 110.365 68.310 110.825 ;
        RECT 68.585 110.655 68.865 111.325 ;
        RECT 67.185 110.145 68.310 110.365 ;
        RECT 67.185 109.685 67.465 110.145 ;
        RECT 67.985 109.515 68.310 109.975 ;
        RECT 68.480 109.685 68.865 110.655 ;
        RECT 69.035 109.515 69.325 110.680 ;
        RECT 69.500 110.525 69.850 111.175 ;
        RECT 70.020 110.355 70.250 111.345 ;
        RECT 69.585 110.185 70.250 110.355 ;
        RECT 69.585 109.685 69.755 110.185 ;
        RECT 69.925 109.515 70.255 110.015 ;
        RECT 70.425 109.685 70.610 111.805 ;
        RECT 70.865 111.605 71.115 112.065 ;
        RECT 71.285 111.615 71.620 111.785 ;
        RECT 71.815 111.615 72.490 111.785 ;
        RECT 71.285 111.475 71.455 111.615 ;
        RECT 70.780 110.485 71.060 111.435 ;
        RECT 71.230 111.345 71.455 111.475 ;
        RECT 71.230 110.240 71.400 111.345 ;
        RECT 71.625 111.195 72.150 111.415 ;
        RECT 71.570 110.430 71.810 111.025 ;
        RECT 71.980 110.495 72.150 111.195 ;
        RECT 72.320 110.835 72.490 111.615 ;
        RECT 72.810 111.565 73.180 112.065 ;
        RECT 73.360 111.615 73.765 111.785 ;
        RECT 73.935 111.615 74.720 111.785 ;
        RECT 73.360 111.385 73.530 111.615 ;
        RECT 72.700 111.085 73.530 111.385 ;
        RECT 73.915 111.115 74.380 111.445 ;
        RECT 72.700 111.055 72.900 111.085 ;
        RECT 73.020 110.835 73.190 110.905 ;
        RECT 72.320 110.665 73.190 110.835 ;
        RECT 72.680 110.575 73.190 110.665 ;
        RECT 71.230 110.110 71.535 110.240 ;
        RECT 71.980 110.130 72.510 110.495 ;
        RECT 70.850 109.515 71.115 109.975 ;
        RECT 71.285 109.685 71.535 110.110 ;
        RECT 72.680 109.960 72.850 110.575 ;
        RECT 71.745 109.790 72.850 109.960 ;
        RECT 73.020 109.515 73.190 110.315 ;
        RECT 73.360 110.015 73.530 111.085 ;
        RECT 73.700 110.185 73.890 110.905 ;
        RECT 74.060 110.155 74.380 111.115 ;
        RECT 74.550 111.155 74.720 111.615 ;
        RECT 74.995 111.535 75.205 112.065 ;
        RECT 75.465 111.325 75.795 111.850 ;
        RECT 75.965 111.455 76.135 112.065 ;
        RECT 76.305 111.410 76.635 111.845 ;
        RECT 76.305 111.325 76.685 111.410 ;
        RECT 75.595 111.155 75.795 111.325 ;
        RECT 76.460 111.285 76.685 111.325 ;
        RECT 74.550 110.825 75.425 111.155 ;
        RECT 75.595 110.825 76.345 111.155 ;
        RECT 73.360 109.685 73.610 110.015 ;
        RECT 74.550 109.985 74.720 110.825 ;
        RECT 75.595 110.620 75.785 110.825 ;
        RECT 76.515 110.705 76.685 111.285 ;
        RECT 76.470 110.655 76.685 110.705 ;
        RECT 74.890 110.245 75.785 110.620 ;
        RECT 76.295 110.575 76.685 110.655 ;
        RECT 76.890 111.325 77.505 111.895 ;
        RECT 77.675 111.555 77.890 112.065 ;
        RECT 78.120 111.555 78.400 111.885 ;
        RECT 78.580 111.555 78.820 112.065 ;
        RECT 73.835 109.815 74.720 109.985 ;
        RECT 74.900 109.515 75.215 110.015 ;
        RECT 75.445 109.685 75.785 110.245 ;
        RECT 75.955 109.515 76.125 110.525 ;
        RECT 76.295 109.730 76.625 110.575 ;
        RECT 76.890 110.305 77.205 111.325 ;
        RECT 77.375 110.655 77.545 111.155 ;
        RECT 77.795 110.825 78.060 111.385 ;
        RECT 78.230 110.655 78.400 111.555 ;
        RECT 79.160 111.535 79.450 111.885 ;
        RECT 79.645 111.705 79.975 112.065 ;
        RECT 80.145 111.535 80.375 111.840 ;
        RECT 78.570 110.825 78.925 111.385 ;
        RECT 79.160 111.365 80.375 111.535 ;
        RECT 80.565 111.195 80.735 111.760 ;
        RECT 81.085 111.515 81.255 111.805 ;
        RECT 81.425 111.685 81.755 112.065 ;
        RECT 81.085 111.345 81.750 111.515 ;
        RECT 79.220 111.045 79.480 111.155 ;
        RECT 79.215 110.875 79.480 111.045 ;
        RECT 79.220 110.825 79.480 110.875 ;
        RECT 79.660 110.825 80.045 111.155 ;
        RECT 80.215 111.025 80.735 111.195 ;
        RECT 77.375 110.485 78.800 110.655 ;
        RECT 76.890 109.685 77.425 110.305 ;
        RECT 77.595 109.515 77.925 110.315 ;
        RECT 78.410 110.310 78.800 110.485 ;
        RECT 79.160 109.515 79.480 110.655 ;
        RECT 79.660 109.775 79.855 110.825 ;
        RECT 80.215 110.645 80.385 111.025 ;
        RECT 80.035 110.365 80.385 110.645 ;
        RECT 80.575 110.495 80.820 110.855 ;
        RECT 81.000 110.525 81.350 111.175 ;
        RECT 80.035 109.685 80.365 110.365 ;
        RECT 81.520 110.355 81.750 111.345 ;
        RECT 80.565 109.515 80.820 110.315 ;
        RECT 81.085 110.185 81.750 110.355 ;
        RECT 81.085 109.685 81.255 110.185 ;
        RECT 81.425 109.515 81.755 110.015 ;
        RECT 81.925 109.685 82.110 111.805 ;
        RECT 82.365 111.605 82.615 112.065 ;
        RECT 82.785 111.615 83.120 111.785 ;
        RECT 83.315 111.615 83.990 111.785 ;
        RECT 82.785 111.475 82.955 111.615 ;
        RECT 82.280 110.485 82.560 111.435 ;
        RECT 82.730 111.345 82.955 111.475 ;
        RECT 82.730 110.240 82.900 111.345 ;
        RECT 83.125 111.195 83.650 111.415 ;
        RECT 83.070 110.430 83.310 111.025 ;
        RECT 83.480 110.495 83.650 111.195 ;
        RECT 83.820 110.835 83.990 111.615 ;
        RECT 84.310 111.565 84.680 112.065 ;
        RECT 84.860 111.615 85.265 111.785 ;
        RECT 85.435 111.615 86.220 111.785 ;
        RECT 84.860 111.385 85.030 111.615 ;
        RECT 84.200 111.085 85.030 111.385 ;
        RECT 85.415 111.115 85.880 111.445 ;
        RECT 84.200 111.055 84.400 111.085 ;
        RECT 84.520 110.835 84.690 110.905 ;
        RECT 83.820 110.665 84.690 110.835 ;
        RECT 84.180 110.575 84.690 110.665 ;
        RECT 82.730 110.110 83.035 110.240 ;
        RECT 83.480 110.130 84.010 110.495 ;
        RECT 82.350 109.515 82.615 109.975 ;
        RECT 82.785 109.685 83.035 110.110 ;
        RECT 84.180 109.960 84.350 110.575 ;
        RECT 83.245 109.790 84.350 109.960 ;
        RECT 84.520 109.515 84.690 110.315 ;
        RECT 84.860 110.015 85.030 111.085 ;
        RECT 85.200 110.185 85.390 110.905 ;
        RECT 85.560 110.155 85.880 111.115 ;
        RECT 86.050 111.155 86.220 111.615 ;
        RECT 86.495 111.535 86.705 112.065 ;
        RECT 86.965 111.325 87.295 111.850 ;
        RECT 87.465 111.455 87.635 112.065 ;
        RECT 87.805 111.410 88.135 111.845 ;
        RECT 88.305 111.550 88.475 112.065 ;
        RECT 87.805 111.325 88.185 111.410 ;
        RECT 87.095 111.155 87.295 111.325 ;
        RECT 87.960 111.285 88.185 111.325 ;
        RECT 86.050 110.825 86.925 111.155 ;
        RECT 87.095 110.825 87.845 111.155 ;
        RECT 84.860 109.685 85.110 110.015 ;
        RECT 86.050 109.985 86.220 110.825 ;
        RECT 87.095 110.620 87.285 110.825 ;
        RECT 88.015 110.705 88.185 111.285 ;
        RECT 88.815 111.295 91.405 112.065 ;
        RECT 91.575 111.565 91.875 111.895 ;
        RECT 92.045 111.585 92.320 112.065 ;
        RECT 88.815 110.775 90.025 111.295 ;
        RECT 87.970 110.655 88.185 110.705 ;
        RECT 86.390 110.245 87.285 110.620 ;
        RECT 87.795 110.575 88.185 110.655 ;
        RECT 90.195 110.605 91.405 111.125 ;
        RECT 85.335 109.815 86.220 109.985 ;
        RECT 86.400 109.515 86.715 110.015 ;
        RECT 86.945 109.685 87.285 110.245 ;
        RECT 87.455 109.515 87.625 110.525 ;
        RECT 87.795 109.730 88.125 110.575 ;
        RECT 88.295 109.515 88.465 110.430 ;
        RECT 88.815 109.515 91.405 110.605 ;
        RECT 91.575 110.655 91.745 111.565 ;
        RECT 92.500 111.415 92.795 111.805 ;
        RECT 92.965 111.585 93.220 112.065 ;
        RECT 93.395 111.415 93.655 111.805 ;
        RECT 93.825 111.585 94.105 112.065 ;
        RECT 91.915 110.825 92.265 111.395 ;
        RECT 92.500 111.245 94.150 111.415 ;
        RECT 94.795 111.340 95.085 112.065 ;
        RECT 95.315 111.605 95.560 112.065 ;
        RECT 92.435 110.905 93.575 111.075 ;
        RECT 92.435 110.655 92.605 110.905 ;
        RECT 93.745 110.735 94.150 111.245 ;
        RECT 95.255 110.825 95.570 111.435 ;
        RECT 95.740 111.075 95.990 111.885 ;
        RECT 96.160 111.540 96.420 112.065 ;
        RECT 96.590 111.415 96.850 111.870 ;
        RECT 97.020 111.585 97.280 112.065 ;
        RECT 97.450 111.415 97.710 111.870 ;
        RECT 97.880 111.585 98.140 112.065 ;
        RECT 98.310 111.415 98.570 111.870 ;
        RECT 98.740 111.585 99.000 112.065 ;
        RECT 99.170 111.415 99.430 111.870 ;
        RECT 99.600 111.585 99.900 112.065 ;
        RECT 96.590 111.245 99.900 111.415 ;
        RECT 100.355 111.245 100.585 112.065 ;
        RECT 100.755 111.265 101.085 111.895 ;
        RECT 95.740 110.825 98.760 111.075 ;
        RECT 91.575 110.485 92.605 110.655 ;
        RECT 93.395 110.565 94.150 110.735 ;
        RECT 91.575 109.685 91.885 110.485 ;
        RECT 93.395 110.315 93.655 110.565 ;
        RECT 92.055 109.515 92.365 110.315 ;
        RECT 92.535 110.145 93.655 110.315 ;
        RECT 92.535 109.685 92.795 110.145 ;
        RECT 92.965 109.515 93.220 109.975 ;
        RECT 93.395 109.685 93.655 110.145 ;
        RECT 93.825 109.515 94.110 110.385 ;
        RECT 94.795 109.515 95.085 110.680 ;
        RECT 95.265 109.515 95.560 110.625 ;
        RECT 95.740 109.690 95.990 110.825 ;
        RECT 98.930 110.655 99.900 111.245 ;
        RECT 100.335 110.825 100.665 111.075 ;
        RECT 100.835 110.665 101.085 111.265 ;
        RECT 101.255 111.245 101.465 112.065 ;
        RECT 101.695 111.315 102.905 112.065 ;
        RECT 103.075 111.405 103.350 112.065 ;
        RECT 103.520 111.435 103.770 111.895 ;
        RECT 103.945 111.570 104.275 112.065 ;
        RECT 101.695 110.775 102.215 111.315 ;
        RECT 103.520 111.225 103.690 111.435 ;
        RECT 104.455 111.400 104.685 111.845 ;
        RECT 96.160 109.515 96.420 110.625 ;
        RECT 96.590 110.415 99.900 110.655 ;
        RECT 96.590 109.690 96.850 110.415 ;
        RECT 97.020 109.515 97.280 110.245 ;
        RECT 97.450 109.690 97.710 110.415 ;
        RECT 97.880 109.515 98.140 110.245 ;
        RECT 98.310 109.690 98.570 110.415 ;
        RECT 98.740 109.515 99.000 110.245 ;
        RECT 99.170 109.690 99.430 110.415 ;
        RECT 99.600 109.515 99.895 110.245 ;
        RECT 100.355 109.515 100.585 110.655 ;
        RECT 100.755 109.685 101.085 110.665 ;
        RECT 101.255 109.515 101.465 110.655 ;
        RECT 102.385 110.605 102.905 111.145 ;
        RECT 103.075 110.705 103.690 111.225 ;
        RECT 103.860 110.725 104.090 111.155 ;
        RECT 104.275 110.905 104.685 111.400 ;
        RECT 104.855 111.580 105.645 111.845 ;
        RECT 104.855 110.725 105.110 111.580 ;
        RECT 105.835 111.425 106.125 111.895 ;
        RECT 106.325 111.595 106.495 112.065 ;
        RECT 106.665 111.425 106.995 111.895 ;
        RECT 107.165 111.595 107.335 112.065 ;
        RECT 107.505 111.425 107.835 111.895 ;
        RECT 108.005 111.595 108.175 112.065 ;
        RECT 108.345 111.425 108.675 111.895 ;
        RECT 108.845 111.595 109.015 112.065 ;
        RECT 109.185 111.425 109.515 111.895 ;
        RECT 109.685 111.595 109.855 112.065 ;
        RECT 110.025 111.425 110.355 111.895 ;
        RECT 110.525 111.595 110.695 112.065 ;
        RECT 110.865 111.425 111.195 111.895 ;
        RECT 105.280 110.905 105.665 111.385 ;
        RECT 105.835 111.245 111.195 111.425 ;
        RECT 111.365 111.245 111.640 112.065 ;
        RECT 111.815 111.565 112.075 111.895 ;
        RECT 112.285 111.585 112.560 112.065 ;
        RECT 101.695 109.515 102.905 110.605 ;
        RECT 103.075 109.515 103.335 110.525 ;
        RECT 103.505 110.365 103.675 110.705 ;
        RECT 103.860 110.555 105.650 110.725 ;
        RECT 103.505 110.355 103.765 110.365 ;
        RECT 103.505 109.685 103.780 110.355 ;
        RECT 103.980 109.515 104.195 110.360 ;
        RECT 104.420 110.260 104.670 110.555 ;
        RECT 104.895 110.195 105.225 110.385 ;
        RECT 104.380 109.685 104.855 110.025 ;
        RECT 105.035 110.020 105.225 110.195 ;
        RECT 105.395 110.190 105.650 110.555 ;
        RECT 105.835 110.365 106.125 111.245 ;
        RECT 106.315 110.865 106.735 111.075 ;
        RECT 106.965 110.875 107.875 111.075 ;
        RECT 106.565 110.705 106.735 110.865 ;
        RECT 108.045 110.865 109.635 111.075 ;
        RECT 109.905 110.865 111.640 111.075 ;
        RECT 108.045 110.705 108.215 110.865 ;
        RECT 106.565 110.535 108.215 110.705 ;
        RECT 108.385 110.525 109.475 110.695 ;
        RECT 105.835 110.195 108.215 110.365 ;
        RECT 105.035 109.515 105.665 110.020 ;
        RECT 105.835 109.685 106.115 110.195 ;
        RECT 107.125 110.185 108.215 110.195 ;
        RECT 107.125 110.025 107.375 110.185 ;
        RECT 107.965 110.025 108.215 110.185 ;
        RECT 106.285 109.685 106.535 110.025 ;
        RECT 106.705 109.855 106.955 110.015 ;
        RECT 107.545 109.855 107.795 110.015 ;
        RECT 108.385 109.855 108.635 110.525 ;
        RECT 106.705 109.685 108.635 109.855 ;
        RECT 108.805 110.065 109.055 110.355 ;
        RECT 109.225 110.235 109.475 110.525 ;
        RECT 109.645 110.525 111.580 110.695 ;
        RECT 109.645 110.065 109.895 110.525 ;
        RECT 108.805 109.685 109.895 110.065 ;
        RECT 110.065 109.515 110.315 110.355 ;
        RECT 110.485 109.685 110.735 110.525 ;
        RECT 110.905 109.515 111.155 110.355 ;
        RECT 111.325 109.685 111.580 110.525 ;
        RECT 111.815 110.655 111.985 111.565 ;
        RECT 112.770 111.495 112.975 111.895 ;
        RECT 113.145 111.665 113.480 112.065 ;
        RECT 112.155 110.825 112.515 111.405 ;
        RECT 112.770 111.325 113.455 111.495 ;
        RECT 112.695 110.655 112.945 111.155 ;
        RECT 111.815 110.485 112.945 110.655 ;
        RECT 111.815 109.715 112.085 110.485 ;
        RECT 113.115 110.295 113.455 111.325 ;
        RECT 113.655 111.295 117.165 112.065 ;
        RECT 118.365 111.685 119.535 111.895 ;
        RECT 118.365 111.665 118.695 111.685 ;
        RECT 113.655 110.775 115.305 111.295 ;
        RECT 118.255 111.245 119.115 111.495 ;
        RECT 119.285 111.435 119.535 111.685 ;
        RECT 119.705 111.605 119.875 112.065 ;
        RECT 120.045 111.435 120.385 111.895 ;
        RECT 119.285 111.265 120.385 111.435 ;
        RECT 120.555 111.340 120.845 112.065 ;
        RECT 121.015 111.565 121.275 111.895 ;
        RECT 121.445 111.705 121.775 112.065 ;
        RECT 122.030 111.685 123.330 111.895 ;
        RECT 115.475 110.605 117.165 111.125 ;
        RECT 112.255 109.515 112.585 110.295 ;
        RECT 112.790 110.120 113.455 110.295 ;
        RECT 112.790 109.715 112.975 110.120 ;
        RECT 113.145 109.515 113.480 109.940 ;
        RECT 113.655 109.515 117.165 110.605 ;
        RECT 118.255 110.655 118.535 111.245 ;
        RECT 118.705 110.825 119.455 111.075 ;
        RECT 119.625 110.825 120.385 111.075 ;
        RECT 118.255 110.485 119.955 110.655 ;
        RECT 118.360 109.515 118.615 110.315 ;
        RECT 118.785 109.685 119.115 110.485 ;
        RECT 119.285 109.515 119.455 110.315 ;
        RECT 119.625 109.685 119.955 110.485 ;
        RECT 120.125 109.515 120.385 110.655 ;
        RECT 120.555 109.515 120.845 110.680 ;
        RECT 121.015 110.365 121.185 111.565 ;
        RECT 122.030 111.535 122.200 111.685 ;
        RECT 121.445 111.410 122.200 111.535 ;
        RECT 121.355 111.365 122.200 111.410 ;
        RECT 121.355 111.245 121.625 111.365 ;
        RECT 121.355 110.670 121.525 111.245 ;
        RECT 121.755 110.805 122.165 111.110 ;
        RECT 122.455 111.075 122.665 111.475 ;
        RECT 122.335 110.865 122.665 111.075 ;
        RECT 122.910 111.075 123.130 111.475 ;
        RECT 123.605 111.300 124.060 112.065 ;
        RECT 124.235 111.565 124.535 111.895 ;
        RECT 124.705 111.585 124.980 112.065 ;
        RECT 122.910 110.865 123.385 111.075 ;
        RECT 123.575 110.875 124.065 111.075 ;
        RECT 121.355 110.635 121.555 110.670 ;
        RECT 122.885 110.635 124.060 110.695 ;
        RECT 121.355 110.525 124.060 110.635 ;
        RECT 121.415 110.465 123.215 110.525 ;
        RECT 122.885 110.435 123.215 110.465 ;
        RECT 121.015 109.685 121.275 110.365 ;
        RECT 121.445 109.515 121.695 110.295 ;
        RECT 121.945 110.265 122.780 110.275 ;
        RECT 123.370 110.265 123.555 110.355 ;
        RECT 121.945 110.065 123.555 110.265 ;
        RECT 121.945 109.685 122.195 110.065 ;
        RECT 123.325 110.025 123.555 110.065 ;
        RECT 123.805 109.905 124.060 110.525 ;
        RECT 122.365 109.515 122.720 109.895 ;
        RECT 123.725 109.685 124.060 109.905 ;
        RECT 124.235 110.655 124.405 111.565 ;
        RECT 125.160 111.415 125.455 111.805 ;
        RECT 125.625 111.585 125.880 112.065 ;
        RECT 126.055 111.415 126.315 111.805 ;
        RECT 126.485 111.585 126.765 112.065 ;
        RECT 124.575 110.825 124.925 111.395 ;
        RECT 125.160 111.245 126.810 111.415 ;
        RECT 127.660 111.285 128.160 111.895 ;
        RECT 125.095 110.905 126.235 111.075 ;
        RECT 125.095 110.655 125.265 110.905 ;
        RECT 126.405 110.735 126.810 111.245 ;
        RECT 127.455 110.825 127.805 111.075 ;
        RECT 124.235 110.485 125.265 110.655 ;
        RECT 126.055 110.565 126.810 110.735 ;
        RECT 127.990 110.655 128.160 111.285 ;
        RECT 128.790 111.415 129.120 111.895 ;
        RECT 129.290 111.605 129.515 112.065 ;
        RECT 129.685 111.415 130.015 111.895 ;
        RECT 128.790 111.245 130.015 111.415 ;
        RECT 130.205 111.265 130.455 112.065 ;
        RECT 130.625 111.265 130.965 111.895 ;
        RECT 131.225 111.515 131.395 111.805 ;
        RECT 131.565 111.685 131.895 112.065 ;
        RECT 131.225 111.345 131.890 111.515 ;
        RECT 128.330 110.875 128.660 111.075 ;
        RECT 128.830 110.875 129.160 111.075 ;
        RECT 129.330 110.875 129.750 111.075 ;
        RECT 129.925 110.905 130.620 111.075 ;
        RECT 129.925 110.655 130.095 110.905 ;
        RECT 130.790 110.655 130.965 111.265 ;
        RECT 124.235 109.685 124.545 110.485 ;
        RECT 126.055 110.315 126.315 110.565 ;
        RECT 127.660 110.485 130.095 110.655 ;
        RECT 124.715 109.515 125.025 110.315 ;
        RECT 125.195 110.145 126.315 110.315 ;
        RECT 125.195 109.685 125.455 110.145 ;
        RECT 125.625 109.515 125.880 109.975 ;
        RECT 126.055 109.685 126.315 110.145 ;
        RECT 126.485 109.515 126.770 110.385 ;
        RECT 127.660 109.685 127.990 110.485 ;
        RECT 128.160 109.515 128.490 110.315 ;
        RECT 128.790 109.685 129.120 110.485 ;
        RECT 129.765 109.515 130.015 110.315 ;
        RECT 130.285 109.515 130.455 110.655 ;
        RECT 130.625 109.685 130.965 110.655 ;
        RECT 131.140 110.525 131.490 111.175 ;
        RECT 131.660 110.355 131.890 111.345 ;
        RECT 131.225 110.185 131.890 110.355 ;
        RECT 131.225 109.685 131.395 110.185 ;
        RECT 131.565 109.515 131.895 110.015 ;
        RECT 132.065 109.685 132.250 111.805 ;
        RECT 132.505 111.605 132.755 112.065 ;
        RECT 132.925 111.615 133.260 111.785 ;
        RECT 133.455 111.615 134.130 111.785 ;
        RECT 132.925 111.475 133.095 111.615 ;
        RECT 132.420 110.485 132.700 111.435 ;
        RECT 132.870 111.345 133.095 111.475 ;
        RECT 132.870 110.240 133.040 111.345 ;
        RECT 133.265 111.195 133.790 111.415 ;
        RECT 133.210 110.430 133.450 111.025 ;
        RECT 133.620 110.495 133.790 111.195 ;
        RECT 133.960 110.835 134.130 111.615 ;
        RECT 134.450 111.565 134.820 112.065 ;
        RECT 135.000 111.615 135.405 111.785 ;
        RECT 135.575 111.615 136.360 111.785 ;
        RECT 135.000 111.385 135.170 111.615 ;
        RECT 134.340 111.085 135.170 111.385 ;
        RECT 135.555 111.115 136.020 111.445 ;
        RECT 134.340 111.055 134.540 111.085 ;
        RECT 134.660 110.835 134.830 110.905 ;
        RECT 133.960 110.665 134.830 110.835 ;
        RECT 134.320 110.575 134.830 110.665 ;
        RECT 132.870 110.110 133.175 110.240 ;
        RECT 133.620 110.130 134.150 110.495 ;
        RECT 132.490 109.515 132.755 109.975 ;
        RECT 132.925 109.685 133.175 110.110 ;
        RECT 134.320 109.960 134.490 110.575 ;
        RECT 133.385 109.790 134.490 109.960 ;
        RECT 134.660 109.515 134.830 110.315 ;
        RECT 135.000 110.015 135.170 111.085 ;
        RECT 135.340 110.185 135.530 110.905 ;
        RECT 135.700 110.155 136.020 111.115 ;
        RECT 136.190 111.155 136.360 111.615 ;
        RECT 136.635 111.535 136.845 112.065 ;
        RECT 137.105 111.325 137.435 111.850 ;
        RECT 137.605 111.455 137.775 112.065 ;
        RECT 137.945 111.410 138.275 111.845 ;
        RECT 138.660 111.555 138.900 112.065 ;
        RECT 139.080 111.555 139.360 111.885 ;
        RECT 139.590 111.555 139.805 112.065 ;
        RECT 137.945 111.325 138.325 111.410 ;
        RECT 137.235 111.155 137.435 111.325 ;
        RECT 138.100 111.285 138.325 111.325 ;
        RECT 136.190 110.825 137.065 111.155 ;
        RECT 137.235 110.825 137.985 111.155 ;
        RECT 135.000 109.685 135.250 110.015 ;
        RECT 136.190 109.985 136.360 110.825 ;
        RECT 137.235 110.620 137.425 110.825 ;
        RECT 138.155 110.705 138.325 111.285 ;
        RECT 138.555 110.825 138.910 111.385 ;
        RECT 138.110 110.655 138.325 110.705 ;
        RECT 139.080 110.655 139.250 111.555 ;
        RECT 139.420 110.825 139.685 111.385 ;
        RECT 139.975 111.325 140.590 111.895 ;
        RECT 139.935 110.655 140.105 111.155 ;
        RECT 136.530 110.245 137.425 110.620 ;
        RECT 137.935 110.575 138.325 110.655 ;
        RECT 135.475 109.815 136.360 109.985 ;
        RECT 136.540 109.515 136.855 110.015 ;
        RECT 137.085 109.685 137.425 110.245 ;
        RECT 137.595 109.515 137.765 110.525 ;
        RECT 137.935 109.730 138.265 110.575 ;
        RECT 138.680 110.485 140.105 110.655 ;
        RECT 138.680 110.310 139.070 110.485 ;
        RECT 139.555 109.515 139.885 110.315 ;
        RECT 140.275 110.305 140.590 111.325 ;
        RECT 141.715 111.315 142.925 112.065 ;
        RECT 140.055 109.685 140.590 110.305 ;
        RECT 141.715 110.605 142.235 111.145 ;
        RECT 142.405 110.775 142.925 111.315 ;
        RECT 141.715 109.515 142.925 110.605 ;
        RECT 17.430 109.345 143.010 109.515 ;
        RECT 17.515 108.255 18.725 109.345 ;
        RECT 18.895 108.255 22.405 109.345 ;
        RECT 17.515 107.545 18.035 108.085 ;
        RECT 18.205 107.715 18.725 108.255 ;
        RECT 18.895 107.565 20.545 108.085 ;
        RECT 20.715 107.735 22.405 108.255 ;
        RECT 23.035 108.475 23.310 109.175 ;
        RECT 23.520 108.800 23.735 109.345 ;
        RECT 23.905 108.835 24.380 109.175 ;
        RECT 24.550 108.840 25.165 109.345 ;
        RECT 24.550 108.665 24.745 108.840 ;
        RECT 17.515 106.795 18.725 107.545 ;
        RECT 18.895 106.795 22.405 107.565 ;
        RECT 23.035 107.445 23.205 108.475 ;
        RECT 23.480 108.305 24.195 108.600 ;
        RECT 24.415 108.475 24.745 108.665 ;
        RECT 24.915 108.305 25.165 108.670 ;
        RECT 23.375 108.135 25.165 108.305 ;
        RECT 23.375 107.705 23.605 108.135 ;
        RECT 23.035 106.965 23.295 107.445 ;
        RECT 23.775 107.435 24.185 107.955 ;
        RECT 23.465 106.795 23.795 107.255 ;
        RECT 23.985 107.015 24.185 107.435 ;
        RECT 24.355 107.280 24.610 108.135 ;
        RECT 25.405 107.955 25.575 109.175 ;
        RECT 25.825 108.835 26.085 109.345 ;
        RECT 24.780 107.705 25.575 107.955 ;
        RECT 25.745 107.785 26.085 108.665 ;
        RECT 26.255 108.205 26.535 109.345 ;
        RECT 26.705 108.195 27.035 109.175 ;
        RECT 27.205 108.205 27.465 109.345 ;
        RECT 26.265 107.765 26.600 108.035 ;
        RECT 25.325 107.615 25.575 107.705 ;
        RECT 24.355 107.015 25.145 107.280 ;
        RECT 25.325 107.195 25.655 107.615 ;
        RECT 25.825 106.795 26.085 107.615 ;
        RECT 26.770 107.595 26.940 108.195 ;
        RECT 27.110 107.785 27.445 108.035 ;
        RECT 26.255 106.795 26.565 107.595 ;
        RECT 26.770 106.965 27.465 107.595 ;
        RECT 27.645 106.975 27.905 109.165 ;
        RECT 28.075 108.615 28.415 109.345 ;
        RECT 28.595 108.435 28.865 109.165 ;
        RECT 28.095 108.215 28.865 108.435 ;
        RECT 29.045 108.455 29.275 109.165 ;
        RECT 29.445 108.635 29.775 109.345 ;
        RECT 29.945 108.455 30.205 109.165 ;
        RECT 29.045 108.215 30.205 108.455 ;
        RECT 28.095 107.545 28.385 108.215 ;
        RECT 30.395 108.180 30.685 109.345 ;
        RECT 30.865 108.545 31.195 109.345 ;
        RECT 31.375 109.005 32.805 109.175 ;
        RECT 31.375 108.375 31.625 109.005 ;
        RECT 30.855 108.205 31.625 108.375 ;
        RECT 28.565 107.725 29.030 108.035 ;
        RECT 29.210 107.725 29.735 108.035 ;
        RECT 28.095 107.345 29.325 107.545 ;
        RECT 28.165 106.795 28.835 107.165 ;
        RECT 29.015 106.975 29.325 107.345 ;
        RECT 29.505 107.085 29.735 107.725 ;
        RECT 29.915 107.705 30.215 108.035 ;
        RECT 30.855 107.535 31.025 108.205 ;
        RECT 31.195 107.705 31.600 108.035 ;
        RECT 31.815 107.705 32.065 108.835 ;
        RECT 32.265 108.035 32.465 108.835 ;
        RECT 32.635 108.325 32.805 109.005 ;
        RECT 32.975 108.495 33.290 109.345 ;
        RECT 33.465 108.545 33.905 109.175 ;
        RECT 32.635 108.155 33.425 108.325 ;
        RECT 32.265 107.705 32.510 108.035 ;
        RECT 32.695 107.705 33.085 107.985 ;
        RECT 33.255 107.705 33.425 108.155 ;
        RECT 33.595 107.535 33.905 108.545 ;
        RECT 34.075 108.255 35.745 109.345 ;
        RECT 29.915 106.795 30.205 107.525 ;
        RECT 30.395 106.795 30.685 107.520 ;
        RECT 30.855 106.965 31.345 107.535 ;
        RECT 31.515 107.365 32.675 107.535 ;
        RECT 31.515 106.965 31.745 107.365 ;
        RECT 31.915 106.795 32.335 107.195 ;
        RECT 32.505 106.965 32.675 107.365 ;
        RECT 32.845 106.795 33.295 107.535 ;
        RECT 33.465 106.975 33.905 107.535 ;
        RECT 34.075 107.565 34.825 108.085 ;
        RECT 34.995 107.735 35.745 108.255 ;
        RECT 36.070 108.335 36.370 109.175 ;
        RECT 36.565 108.505 36.815 109.345 ;
        RECT 37.405 108.755 38.210 109.175 ;
        RECT 36.985 108.585 38.550 108.755 ;
        RECT 36.985 108.335 37.155 108.585 ;
        RECT 36.070 108.165 37.155 108.335 ;
        RECT 35.915 107.705 36.245 107.995 ;
        RECT 34.075 106.795 35.745 107.565 ;
        RECT 36.415 107.535 36.585 108.165 ;
        RECT 37.325 108.035 37.645 108.415 ;
        RECT 37.835 108.325 38.210 108.415 ;
        RECT 37.815 108.155 38.210 108.325 ;
        RECT 38.380 108.335 38.550 108.585 ;
        RECT 38.720 108.505 39.050 109.345 ;
        RECT 39.220 108.585 39.885 109.175 ;
        RECT 38.380 108.165 39.300 108.335 ;
        RECT 36.755 107.785 37.085 107.995 ;
        RECT 37.265 107.785 37.645 108.035 ;
        RECT 37.835 107.995 38.210 108.155 ;
        RECT 39.130 107.995 39.300 108.165 ;
        RECT 37.835 107.785 38.320 107.995 ;
        RECT 38.510 107.785 38.960 107.995 ;
        RECT 39.130 107.785 39.465 107.995 ;
        RECT 39.635 107.615 39.885 108.585 ;
        RECT 36.075 107.355 36.585 107.535 ;
        RECT 36.990 107.445 38.690 107.615 ;
        RECT 36.990 107.355 37.375 107.445 ;
        RECT 36.075 106.965 36.405 107.355 ;
        RECT 36.575 107.015 37.760 107.185 ;
        RECT 38.020 106.795 38.190 107.265 ;
        RECT 38.360 106.980 38.690 107.445 ;
        RECT 38.860 106.795 39.030 107.615 ;
        RECT 39.200 106.975 39.885 107.615 ;
        RECT 40.055 108.475 40.330 109.175 ;
        RECT 40.540 108.800 40.755 109.345 ;
        RECT 40.925 108.835 41.400 109.175 ;
        RECT 41.570 108.840 42.185 109.345 ;
        RECT 41.570 108.665 41.765 108.840 ;
        RECT 40.055 107.445 40.225 108.475 ;
        RECT 40.500 108.305 41.215 108.600 ;
        RECT 41.435 108.475 41.765 108.665 ;
        RECT 41.935 108.305 42.185 108.670 ;
        RECT 40.395 108.135 42.185 108.305 ;
        RECT 40.395 107.705 40.625 108.135 ;
        RECT 40.055 106.965 40.315 107.445 ;
        RECT 40.795 107.435 41.205 107.955 ;
        RECT 40.485 106.795 40.815 107.255 ;
        RECT 41.005 107.015 41.205 107.435 ;
        RECT 41.375 107.280 41.630 108.135 ;
        RECT 42.425 107.955 42.595 109.175 ;
        RECT 42.845 108.835 43.105 109.345 ;
        RECT 41.800 107.705 42.595 107.955 ;
        RECT 42.765 107.785 43.105 108.665 ;
        RECT 43.275 108.255 44.485 109.345 ;
        RECT 42.345 107.615 42.595 107.705 ;
        RECT 41.375 107.015 42.165 107.280 ;
        RECT 42.345 107.195 42.675 107.615 ;
        RECT 42.845 106.795 43.105 107.615 ;
        RECT 43.275 107.545 43.795 108.085 ;
        RECT 43.965 107.715 44.485 108.255 ;
        RECT 44.745 108.335 44.915 109.175 ;
        RECT 45.085 109.005 46.255 109.175 ;
        RECT 45.085 108.505 45.415 109.005 ;
        RECT 45.925 108.965 46.255 109.005 ;
        RECT 46.445 108.925 46.800 109.345 ;
        RECT 45.585 108.745 45.815 108.835 ;
        RECT 46.970 108.745 47.220 109.175 ;
        RECT 45.585 108.505 47.220 108.745 ;
        RECT 47.390 108.585 47.720 109.345 ;
        RECT 47.890 108.505 48.145 109.175 ;
        RECT 44.745 108.165 47.805 108.335 ;
        RECT 44.660 107.785 45.010 107.995 ;
        RECT 45.180 107.785 45.625 107.985 ;
        RECT 45.795 107.785 46.270 107.985 ;
        RECT 43.275 106.795 44.485 107.545 ;
        RECT 44.745 107.445 45.810 107.615 ;
        RECT 44.745 106.965 44.915 107.445 ;
        RECT 45.085 106.795 45.415 107.275 ;
        RECT 45.640 107.215 45.810 107.445 ;
        RECT 45.990 107.385 46.270 107.785 ;
        RECT 46.540 107.785 46.870 107.985 ;
        RECT 47.040 107.815 47.415 107.985 ;
        RECT 47.040 107.785 47.405 107.815 ;
        RECT 46.540 107.385 46.825 107.785 ;
        RECT 47.635 107.615 47.805 108.165 ;
        RECT 47.005 107.445 47.805 107.615 ;
        RECT 47.005 107.215 47.175 107.445 ;
        RECT 47.975 107.375 48.145 108.505 ;
        RECT 47.960 107.305 48.145 107.375 ;
        RECT 47.935 107.295 48.145 107.305 ;
        RECT 45.640 106.965 47.175 107.215 ;
        RECT 47.345 106.795 47.675 107.275 ;
        RECT 47.890 106.965 48.145 107.295 ;
        RECT 49.255 108.475 49.530 109.175 ;
        RECT 49.740 108.800 49.955 109.345 ;
        RECT 50.125 108.835 50.600 109.175 ;
        RECT 50.770 108.840 51.385 109.345 ;
        RECT 50.770 108.665 50.965 108.840 ;
        RECT 49.255 107.445 49.425 108.475 ;
        RECT 49.700 108.305 50.415 108.600 ;
        RECT 50.635 108.475 50.965 108.665 ;
        RECT 51.135 108.305 51.385 108.670 ;
        RECT 49.595 108.135 51.385 108.305 ;
        RECT 49.595 107.705 49.825 108.135 ;
        RECT 49.255 106.965 49.515 107.445 ;
        RECT 49.995 107.435 50.405 107.955 ;
        RECT 49.685 106.795 50.015 107.255 ;
        RECT 50.205 107.015 50.405 107.435 ;
        RECT 50.575 107.280 50.830 108.135 ;
        RECT 51.625 107.955 51.795 109.175 ;
        RECT 52.045 108.835 52.305 109.345 ;
        RECT 52.590 108.715 52.875 109.175 ;
        RECT 53.045 108.885 53.315 109.345 ;
        RECT 51.000 107.705 51.795 107.955 ;
        RECT 51.965 107.785 52.305 108.665 ;
        RECT 52.590 108.495 53.545 108.715 ;
        RECT 52.475 107.765 53.165 108.325 ;
        RECT 51.545 107.615 51.795 107.705 ;
        RECT 50.575 107.015 51.365 107.280 ;
        RECT 51.545 107.195 51.875 107.615 ;
        RECT 52.045 106.795 52.305 107.615 ;
        RECT 53.335 107.595 53.545 108.495 ;
        RECT 52.590 107.425 53.545 107.595 ;
        RECT 53.715 108.325 54.115 109.175 ;
        RECT 54.305 108.715 54.585 109.175 ;
        RECT 55.105 108.885 55.430 109.345 ;
        RECT 54.305 108.495 55.430 108.715 ;
        RECT 53.715 107.765 54.810 108.325 ;
        RECT 54.980 108.035 55.430 108.495 ;
        RECT 55.600 108.205 55.985 109.175 ;
        RECT 52.590 106.965 52.875 107.425 ;
        RECT 53.045 106.795 53.315 107.255 ;
        RECT 53.715 106.965 54.115 107.765 ;
        RECT 54.980 107.705 55.535 108.035 ;
        RECT 54.980 107.595 55.430 107.705 ;
        RECT 54.305 107.425 55.430 107.595 ;
        RECT 55.705 107.535 55.985 108.205 ;
        RECT 56.155 108.180 56.445 109.345 ;
        RECT 56.675 108.285 57.005 109.130 ;
        RECT 57.175 108.335 57.345 109.345 ;
        RECT 57.515 108.615 57.855 109.175 ;
        RECT 58.085 108.845 58.400 109.345 ;
        RECT 58.580 108.875 59.465 109.045 ;
        RECT 56.615 108.205 57.005 108.285 ;
        RECT 57.515 108.240 58.410 108.615 ;
        RECT 54.305 106.965 54.585 107.425 ;
        RECT 55.105 106.795 55.430 107.255 ;
        RECT 55.600 106.965 55.985 107.535 ;
        RECT 56.615 108.155 56.830 108.205 ;
        RECT 56.615 107.575 56.785 108.155 ;
        RECT 57.515 108.035 57.705 108.240 ;
        RECT 58.580 108.035 58.750 108.875 ;
        RECT 59.690 108.845 59.940 109.175 ;
        RECT 56.955 107.705 57.705 108.035 ;
        RECT 57.875 107.705 58.750 108.035 ;
        RECT 56.615 107.535 56.840 107.575 ;
        RECT 57.505 107.535 57.705 107.705 ;
        RECT 56.155 106.795 56.445 107.520 ;
        RECT 56.615 107.450 56.995 107.535 ;
        RECT 56.665 107.015 56.995 107.450 ;
        RECT 57.165 106.795 57.335 107.405 ;
        RECT 57.505 107.010 57.835 107.535 ;
        RECT 58.095 106.795 58.305 107.325 ;
        RECT 58.580 107.245 58.750 107.705 ;
        RECT 58.920 107.745 59.240 108.705 ;
        RECT 59.410 107.955 59.600 108.675 ;
        RECT 59.770 107.775 59.940 108.845 ;
        RECT 60.110 108.545 60.280 109.345 ;
        RECT 60.450 108.900 61.555 109.070 ;
        RECT 60.450 108.285 60.620 108.900 ;
        RECT 61.765 108.750 62.015 109.175 ;
        RECT 62.185 108.885 62.450 109.345 ;
        RECT 60.790 108.365 61.320 108.730 ;
        RECT 61.765 108.620 62.070 108.750 ;
        RECT 60.110 108.195 60.620 108.285 ;
        RECT 60.110 108.025 60.980 108.195 ;
        RECT 60.110 107.955 60.280 108.025 ;
        RECT 60.400 107.775 60.600 107.805 ;
        RECT 58.920 107.415 59.385 107.745 ;
        RECT 59.770 107.475 60.600 107.775 ;
        RECT 59.770 107.245 59.940 107.475 ;
        RECT 58.580 107.075 59.365 107.245 ;
        RECT 59.535 107.075 59.940 107.245 ;
        RECT 60.120 106.795 60.490 107.295 ;
        RECT 60.810 107.245 60.980 108.025 ;
        RECT 61.150 107.665 61.320 108.365 ;
        RECT 61.490 107.835 61.730 108.430 ;
        RECT 61.150 107.445 61.675 107.665 ;
        RECT 61.900 107.515 62.070 108.620 ;
        RECT 61.845 107.385 62.070 107.515 ;
        RECT 62.240 107.425 62.520 108.375 ;
        RECT 61.845 107.245 62.015 107.385 ;
        RECT 60.810 107.075 61.485 107.245 ;
        RECT 61.680 107.075 62.015 107.245 ;
        RECT 62.185 106.795 62.435 107.255 ;
        RECT 62.690 107.055 62.875 109.175 ;
        RECT 63.045 108.845 63.375 109.345 ;
        RECT 63.545 108.675 63.715 109.175 ;
        RECT 63.050 108.505 63.715 108.675 ;
        RECT 63.050 107.515 63.280 108.505 ;
        RECT 63.450 107.685 63.800 108.335 ;
        RECT 63.975 108.255 65.185 109.345 ;
        RECT 63.975 107.545 64.495 108.085 ;
        RECT 64.665 107.715 65.185 108.255 ;
        RECT 65.355 107.740 65.635 109.175 ;
        RECT 65.805 108.570 66.515 109.345 ;
        RECT 66.685 108.400 67.015 109.175 ;
        RECT 65.865 108.185 67.015 108.400 ;
        RECT 63.050 107.345 63.715 107.515 ;
        RECT 63.045 106.795 63.375 107.175 ;
        RECT 63.545 107.055 63.715 107.345 ;
        RECT 63.975 106.795 65.185 107.545 ;
        RECT 65.355 106.965 65.695 107.740 ;
        RECT 65.865 107.615 66.150 108.185 ;
        RECT 66.335 107.785 66.805 108.015 ;
        RECT 67.210 107.985 67.425 109.100 ;
        RECT 67.605 108.625 67.935 109.345 ;
        RECT 67.715 107.985 67.945 108.325 ;
        RECT 68.115 108.255 69.325 109.345 ;
        RECT 66.975 107.805 67.425 107.985 ;
        RECT 66.975 107.785 67.305 107.805 ;
        RECT 67.615 107.785 67.945 107.985 ;
        RECT 65.865 107.425 66.575 107.615 ;
        RECT 66.275 107.285 66.575 107.425 ;
        RECT 66.765 107.425 67.945 107.615 ;
        RECT 66.765 107.345 67.095 107.425 ;
        RECT 66.275 107.275 66.590 107.285 ;
        RECT 66.275 107.265 66.600 107.275 ;
        RECT 66.275 107.260 66.610 107.265 ;
        RECT 65.865 106.795 66.035 107.255 ;
        RECT 66.275 107.250 66.615 107.260 ;
        RECT 66.275 107.245 66.620 107.250 ;
        RECT 66.275 107.235 66.625 107.245 ;
        RECT 66.275 107.230 66.630 107.235 ;
        RECT 66.275 106.965 66.635 107.230 ;
        RECT 67.265 106.795 67.435 107.255 ;
        RECT 67.605 106.965 67.945 107.425 ;
        RECT 68.115 107.545 68.635 108.085 ;
        RECT 68.805 107.715 69.325 108.255 ;
        RECT 69.500 108.205 69.775 109.175 ;
        RECT 69.985 108.545 70.265 109.345 ;
        RECT 70.435 108.835 71.625 109.125 ;
        RECT 70.435 108.495 71.605 108.665 ;
        RECT 70.435 108.375 70.605 108.495 ;
        RECT 69.945 108.205 70.605 108.375 ;
        RECT 68.115 106.795 69.325 107.545 ;
        RECT 69.500 107.470 69.670 108.205 ;
        RECT 69.945 108.035 70.115 108.205 ;
        RECT 70.915 108.035 71.110 108.325 ;
        RECT 71.280 108.205 71.605 108.495 ;
        RECT 71.795 108.475 72.070 109.175 ;
        RECT 72.240 108.800 72.495 109.345 ;
        RECT 72.665 108.835 73.145 109.175 ;
        RECT 73.320 108.790 73.925 109.345 ;
        RECT 73.310 108.690 73.925 108.790 ;
        RECT 73.310 108.665 73.495 108.690 ;
        RECT 69.840 107.705 70.115 108.035 ;
        RECT 70.285 107.705 71.110 108.035 ;
        RECT 71.280 107.705 71.625 108.035 ;
        RECT 69.945 107.535 70.115 107.705 ;
        RECT 69.500 107.125 69.775 107.470 ;
        RECT 69.945 107.365 71.610 107.535 ;
        RECT 69.965 106.795 70.345 107.195 ;
        RECT 70.515 107.015 70.685 107.365 ;
        RECT 70.855 106.795 71.185 107.195 ;
        RECT 71.355 107.015 71.610 107.365 ;
        RECT 71.795 107.445 71.965 108.475 ;
        RECT 72.240 108.345 72.995 108.595 ;
        RECT 73.165 108.420 73.495 108.665 ;
        RECT 72.240 108.310 73.010 108.345 ;
        RECT 72.240 108.300 73.025 108.310 ;
        RECT 72.135 108.285 73.030 108.300 ;
        RECT 72.135 108.270 73.050 108.285 ;
        RECT 72.135 108.260 73.070 108.270 ;
        RECT 72.135 108.250 73.095 108.260 ;
        RECT 72.135 108.220 73.165 108.250 ;
        RECT 72.135 108.190 73.185 108.220 ;
        RECT 72.135 108.160 73.205 108.190 ;
        RECT 72.135 108.135 73.235 108.160 ;
        RECT 72.135 108.100 73.270 108.135 ;
        RECT 72.135 108.095 73.300 108.100 ;
        RECT 72.135 107.700 72.365 108.095 ;
        RECT 72.910 108.090 73.300 108.095 ;
        RECT 72.935 108.080 73.300 108.090 ;
        RECT 72.950 108.075 73.300 108.080 ;
        RECT 72.965 108.070 73.300 108.075 ;
        RECT 73.665 108.070 73.925 108.520 ;
        RECT 72.965 108.065 73.925 108.070 ;
        RECT 72.975 108.055 73.925 108.065 ;
        RECT 72.985 108.050 73.925 108.055 ;
        RECT 72.995 108.040 73.925 108.050 ;
        RECT 73.000 108.030 73.925 108.040 ;
        RECT 73.005 108.025 73.925 108.030 ;
        RECT 73.015 108.010 73.925 108.025 ;
        RECT 73.020 107.995 73.925 108.010 ;
        RECT 73.030 107.970 73.925 107.995 ;
        RECT 72.535 107.500 72.865 107.925 ;
        RECT 72.615 107.475 72.865 107.500 ;
        RECT 71.795 106.965 72.055 107.445 ;
        RECT 72.225 106.795 72.475 107.335 ;
        RECT 72.645 107.015 72.865 107.475 ;
        RECT 73.035 107.900 73.925 107.970 ;
        RECT 74.095 108.205 74.480 109.175 ;
        RECT 74.650 108.885 74.975 109.345 ;
        RECT 75.495 108.715 75.775 109.175 ;
        RECT 74.650 108.495 75.775 108.715 ;
        RECT 73.035 107.175 73.205 107.900 ;
        RECT 73.375 107.345 73.925 107.730 ;
        RECT 74.095 107.535 74.375 108.205 ;
        RECT 74.650 108.035 75.100 108.495 ;
        RECT 75.965 108.325 76.365 109.175 ;
        RECT 76.765 108.885 77.035 109.345 ;
        RECT 77.205 108.715 77.490 109.175 ;
        RECT 74.545 107.705 75.100 108.035 ;
        RECT 75.270 107.765 76.365 108.325 ;
        RECT 74.650 107.595 75.100 107.705 ;
        RECT 73.035 107.005 73.925 107.175 ;
        RECT 74.095 106.965 74.480 107.535 ;
        RECT 74.650 107.425 75.775 107.595 ;
        RECT 74.650 106.795 74.975 107.255 ;
        RECT 75.495 106.965 75.775 107.425 ;
        RECT 75.965 106.965 76.365 107.765 ;
        RECT 76.535 108.495 77.490 108.715 ;
        RECT 77.775 108.585 78.290 108.995 ;
        RECT 78.525 108.585 78.695 109.345 ;
        RECT 78.865 109.005 80.895 109.175 ;
        RECT 76.535 107.595 76.745 108.495 ;
        RECT 76.915 107.765 77.605 108.325 ;
        RECT 77.775 107.775 78.115 108.585 ;
        RECT 78.865 108.340 79.035 109.005 ;
        RECT 79.430 108.665 80.555 108.835 ;
        RECT 78.285 108.150 79.035 108.340 ;
        RECT 79.205 108.325 80.215 108.495 ;
        RECT 77.775 107.605 79.005 107.775 ;
        RECT 76.535 107.425 77.490 107.595 ;
        RECT 76.765 106.795 77.035 107.255 ;
        RECT 77.205 106.965 77.490 107.425 ;
        RECT 78.050 107.000 78.295 107.605 ;
        RECT 78.515 106.795 79.025 107.330 ;
        RECT 79.205 106.965 79.395 108.325 ;
        RECT 79.565 107.305 79.840 108.125 ;
        RECT 80.045 107.525 80.215 108.325 ;
        RECT 80.385 107.535 80.555 108.665 ;
        RECT 80.725 108.035 80.895 109.005 ;
        RECT 81.065 108.205 81.235 109.345 ;
        RECT 81.405 108.205 81.740 109.175 ;
        RECT 80.725 107.705 80.920 108.035 ;
        RECT 81.145 107.705 81.400 108.035 ;
        RECT 81.145 107.535 81.315 107.705 ;
        RECT 81.570 107.535 81.740 108.205 ;
        RECT 81.915 108.180 82.205 109.345 ;
        RECT 82.465 108.675 82.635 109.175 ;
        RECT 82.805 108.845 83.135 109.345 ;
        RECT 82.465 108.505 83.130 108.675 ;
        RECT 82.380 107.685 82.730 108.335 ;
        RECT 80.385 107.365 81.315 107.535 ;
        RECT 80.385 107.330 80.560 107.365 ;
        RECT 79.565 107.135 79.845 107.305 ;
        RECT 79.565 106.965 79.840 107.135 ;
        RECT 80.030 106.965 80.560 107.330 ;
        RECT 80.985 106.795 81.315 107.195 ;
        RECT 81.485 106.965 81.740 107.535 ;
        RECT 81.915 106.795 82.205 107.520 ;
        RECT 82.900 107.515 83.130 108.505 ;
        RECT 82.465 107.345 83.130 107.515 ;
        RECT 82.465 107.055 82.635 107.345 ;
        RECT 82.805 106.795 83.135 107.175 ;
        RECT 83.305 107.055 83.490 109.175 ;
        RECT 83.730 108.885 83.995 109.345 ;
        RECT 84.165 108.750 84.415 109.175 ;
        RECT 84.625 108.900 85.730 109.070 ;
        RECT 84.110 108.620 84.415 108.750 ;
        RECT 83.660 107.425 83.940 108.375 ;
        RECT 84.110 107.515 84.280 108.620 ;
        RECT 84.450 107.835 84.690 108.430 ;
        RECT 84.860 108.365 85.390 108.730 ;
        RECT 84.860 107.665 85.030 108.365 ;
        RECT 85.560 108.285 85.730 108.900 ;
        RECT 85.900 108.545 86.070 109.345 ;
        RECT 86.240 108.845 86.490 109.175 ;
        RECT 86.715 108.875 87.600 109.045 ;
        RECT 85.560 108.195 86.070 108.285 ;
        RECT 84.110 107.385 84.335 107.515 ;
        RECT 84.505 107.445 85.030 107.665 ;
        RECT 85.200 108.025 86.070 108.195 ;
        RECT 83.745 106.795 83.995 107.255 ;
        RECT 84.165 107.245 84.335 107.385 ;
        RECT 85.200 107.245 85.370 108.025 ;
        RECT 85.900 107.955 86.070 108.025 ;
        RECT 85.580 107.775 85.780 107.805 ;
        RECT 86.240 107.775 86.410 108.845 ;
        RECT 86.580 107.955 86.770 108.675 ;
        RECT 85.580 107.475 86.410 107.775 ;
        RECT 86.940 107.745 87.260 108.705 ;
        RECT 84.165 107.075 84.500 107.245 ;
        RECT 84.695 107.075 85.370 107.245 ;
        RECT 85.690 106.795 86.060 107.295 ;
        RECT 86.240 107.245 86.410 107.475 ;
        RECT 86.795 107.415 87.260 107.745 ;
        RECT 87.430 108.035 87.600 108.875 ;
        RECT 87.780 108.845 88.095 109.345 ;
        RECT 88.325 108.615 88.665 109.175 ;
        RECT 87.770 108.240 88.665 108.615 ;
        RECT 88.835 108.335 89.005 109.345 ;
        RECT 88.475 108.035 88.665 108.240 ;
        RECT 89.175 108.285 89.505 109.130 ;
        RECT 89.675 108.430 89.845 109.345 ;
        RECT 90.710 108.475 90.995 109.345 ;
        RECT 91.165 108.715 91.425 109.175 ;
        RECT 91.600 108.885 91.855 109.345 ;
        RECT 92.025 108.715 92.285 109.175 ;
        RECT 91.165 108.545 92.285 108.715 ;
        RECT 92.455 108.545 92.765 109.345 ;
        RECT 91.165 108.295 91.425 108.545 ;
        RECT 92.935 108.375 93.245 109.175 ;
        RECT 89.175 108.205 89.565 108.285 ;
        RECT 89.350 108.155 89.565 108.205 ;
        RECT 87.430 107.705 88.305 108.035 ;
        RECT 88.475 107.705 89.225 108.035 ;
        RECT 87.430 107.245 87.600 107.705 ;
        RECT 88.475 107.535 88.675 107.705 ;
        RECT 89.395 107.575 89.565 108.155 ;
        RECT 89.340 107.535 89.565 107.575 ;
        RECT 86.240 107.075 86.645 107.245 ;
        RECT 86.815 107.075 87.600 107.245 ;
        RECT 87.875 106.795 88.085 107.325 ;
        RECT 88.345 107.010 88.675 107.535 ;
        RECT 89.185 107.450 89.565 107.535 ;
        RECT 90.670 108.125 91.425 108.295 ;
        RECT 92.215 108.205 93.245 108.375 ;
        RECT 93.415 108.255 96.925 109.345 ;
        RECT 97.095 108.255 98.305 109.345 ;
        RECT 98.580 108.885 98.750 109.345 ;
        RECT 98.920 108.715 99.250 109.175 ;
        RECT 90.670 107.615 91.075 108.125 ;
        RECT 92.215 107.955 92.385 108.205 ;
        RECT 91.245 107.785 92.385 107.955 ;
        RECT 88.845 106.795 89.015 107.405 ;
        RECT 89.185 107.015 89.515 107.450 ;
        RECT 90.670 107.445 92.320 107.615 ;
        RECT 92.555 107.465 92.905 108.035 ;
        RECT 89.685 106.795 89.855 107.310 ;
        RECT 90.715 106.795 90.995 107.275 ;
        RECT 91.165 107.055 91.425 107.445 ;
        RECT 91.600 106.795 91.855 107.275 ;
        RECT 92.025 107.055 92.320 107.445 ;
        RECT 93.075 107.295 93.245 108.205 ;
        RECT 92.500 106.795 92.775 107.275 ;
        RECT 92.945 106.965 93.245 107.295 ;
        RECT 93.415 107.565 95.065 108.085 ;
        RECT 95.235 107.735 96.925 108.255 ;
        RECT 93.415 106.795 96.925 107.565 ;
        RECT 97.095 107.545 97.615 108.085 ;
        RECT 97.785 107.715 98.305 108.255 ;
        RECT 98.475 108.545 99.250 108.715 ;
        RECT 99.420 108.545 99.590 109.345 ;
        RECT 97.095 106.795 98.305 107.545 ;
        RECT 98.475 107.535 98.905 108.545 ;
        RECT 100.175 108.375 100.535 108.550 ;
        RECT 99.075 108.205 100.535 108.375 ;
        RECT 100.780 108.375 101.055 109.175 ;
        RECT 101.225 108.545 101.555 109.345 ;
        RECT 101.725 109.005 102.865 109.175 ;
        RECT 101.725 108.375 101.895 109.005 ;
        RECT 99.075 107.705 99.245 108.205 ;
        RECT 98.475 107.365 99.170 107.535 ;
        RECT 99.415 107.475 99.825 108.035 ;
        RECT 98.500 106.795 98.830 107.195 ;
        RECT 99.000 107.095 99.170 107.365 ;
        RECT 99.995 107.305 100.175 108.205 ;
        RECT 100.780 108.165 101.895 108.375 ;
        RECT 102.065 108.375 102.395 108.835 ;
        RECT 102.565 108.545 102.865 109.005 ;
        RECT 102.065 108.155 102.825 108.375 ;
        RECT 103.115 108.205 103.345 109.345 ;
        RECT 103.515 108.195 103.845 109.175 ;
        RECT 104.015 108.205 104.225 109.345 ;
        RECT 105.575 108.675 105.855 109.345 ;
        RECT 106.025 108.455 106.325 109.005 ;
        RECT 106.525 108.625 106.855 109.345 ;
        RECT 107.045 108.625 107.505 109.175 ;
        RECT 100.345 107.645 100.540 108.035 ;
        RECT 100.780 107.785 101.500 107.985 ;
        RECT 101.670 107.785 102.440 107.985 ;
        RECT 100.345 107.475 100.545 107.645 ;
        RECT 102.610 107.615 102.825 108.155 ;
        RECT 103.095 107.785 103.425 108.035 ;
        RECT 99.340 106.795 99.655 107.305 ;
        RECT 99.885 106.965 100.175 107.305 ;
        RECT 100.345 106.795 100.585 107.305 ;
        RECT 100.780 106.795 101.055 107.615 ;
        RECT 101.225 107.445 102.825 107.615 ;
        RECT 101.225 107.435 102.395 107.445 ;
        RECT 101.225 106.965 101.555 107.435 ;
        RECT 101.725 106.795 101.895 107.265 ;
        RECT 102.065 106.965 102.395 107.435 ;
        RECT 102.565 106.795 102.855 107.265 ;
        RECT 103.115 106.795 103.345 107.615 ;
        RECT 103.595 107.595 103.845 108.195 ;
        RECT 105.390 108.035 105.655 108.395 ;
        RECT 106.025 108.285 106.965 108.455 ;
        RECT 106.795 108.035 106.965 108.285 ;
        RECT 105.390 107.785 106.065 108.035 ;
        RECT 106.285 107.785 106.625 108.035 ;
        RECT 106.795 107.705 107.085 108.035 ;
        RECT 106.795 107.615 106.965 107.705 ;
        RECT 103.515 106.965 103.845 107.595 ;
        RECT 104.015 106.795 104.225 107.615 ;
        RECT 105.575 107.425 106.965 107.615 ;
        RECT 105.575 107.065 105.905 107.425 ;
        RECT 107.255 107.255 107.505 108.625 ;
        RECT 107.675 108.180 107.965 109.345 ;
        RECT 108.135 108.205 108.395 109.345 ;
        RECT 108.565 108.375 108.895 109.175 ;
        RECT 109.065 108.545 109.235 109.345 ;
        RECT 109.405 108.375 109.735 109.175 ;
        RECT 109.905 108.545 110.160 109.345 ;
        RECT 108.565 108.205 110.265 108.375 ;
        RECT 110.435 108.255 113.945 109.345 ;
        RECT 114.115 108.255 115.325 109.345 ;
        RECT 115.585 108.675 115.755 109.175 ;
        RECT 115.925 108.845 116.255 109.345 ;
        RECT 115.585 108.505 116.250 108.675 ;
        RECT 108.135 107.785 108.895 108.035 ;
        RECT 109.065 107.785 109.815 108.035 ;
        RECT 109.985 107.615 110.265 108.205 ;
        RECT 106.525 106.795 106.775 107.255 ;
        RECT 106.945 106.965 107.505 107.255 ;
        RECT 107.675 106.795 107.965 107.520 ;
        RECT 108.135 107.425 109.235 107.595 ;
        RECT 108.135 106.965 108.475 107.425 ;
        RECT 108.645 106.795 108.815 107.255 ;
        RECT 108.985 107.175 109.235 107.425 ;
        RECT 109.405 107.365 110.265 107.615 ;
        RECT 110.435 107.565 112.085 108.085 ;
        RECT 112.255 107.735 113.945 108.255 ;
        RECT 109.825 107.175 110.155 107.195 ;
        RECT 108.985 106.965 110.155 107.175 ;
        RECT 110.435 106.795 113.945 107.565 ;
        RECT 114.115 107.545 114.635 108.085 ;
        RECT 114.805 107.715 115.325 108.255 ;
        RECT 115.500 107.685 115.850 108.335 ;
        RECT 114.115 106.795 115.325 107.545 ;
        RECT 116.020 107.515 116.250 108.505 ;
        RECT 115.585 107.345 116.250 107.515 ;
        RECT 115.585 107.055 115.755 107.345 ;
        RECT 115.925 106.795 116.255 107.175 ;
        RECT 116.425 107.055 116.610 109.175 ;
        RECT 116.850 108.885 117.115 109.345 ;
        RECT 117.285 108.750 117.535 109.175 ;
        RECT 117.745 108.900 118.850 109.070 ;
        RECT 117.230 108.620 117.535 108.750 ;
        RECT 116.780 107.425 117.060 108.375 ;
        RECT 117.230 107.515 117.400 108.620 ;
        RECT 117.570 107.835 117.810 108.430 ;
        RECT 117.980 108.365 118.510 108.730 ;
        RECT 117.980 107.665 118.150 108.365 ;
        RECT 118.680 108.285 118.850 108.900 ;
        RECT 119.020 108.545 119.190 109.345 ;
        RECT 119.360 108.845 119.610 109.175 ;
        RECT 119.835 108.875 120.720 109.045 ;
        RECT 118.680 108.195 119.190 108.285 ;
        RECT 117.230 107.385 117.455 107.515 ;
        RECT 117.625 107.445 118.150 107.665 ;
        RECT 118.320 108.025 119.190 108.195 ;
        RECT 116.865 106.795 117.115 107.255 ;
        RECT 117.285 107.245 117.455 107.385 ;
        RECT 118.320 107.245 118.490 108.025 ;
        RECT 119.020 107.955 119.190 108.025 ;
        RECT 118.700 107.775 118.900 107.805 ;
        RECT 119.360 107.775 119.530 108.845 ;
        RECT 119.700 107.955 119.890 108.675 ;
        RECT 118.700 107.475 119.530 107.775 ;
        RECT 120.060 107.745 120.380 108.705 ;
        RECT 117.285 107.075 117.620 107.245 ;
        RECT 117.815 107.075 118.490 107.245 ;
        RECT 118.810 106.795 119.180 107.295 ;
        RECT 119.360 107.245 119.530 107.475 ;
        RECT 119.915 107.415 120.380 107.745 ;
        RECT 120.550 108.035 120.720 108.875 ;
        RECT 120.900 108.845 121.215 109.345 ;
        RECT 121.445 108.615 121.785 109.175 ;
        RECT 120.890 108.240 121.785 108.615 ;
        RECT 121.955 108.335 122.125 109.345 ;
        RECT 121.595 108.035 121.785 108.240 ;
        RECT 122.295 108.285 122.625 109.130 ;
        RECT 122.295 108.205 122.685 108.285 ;
        RECT 122.865 108.235 123.160 109.345 ;
        RECT 122.470 108.155 122.685 108.205 ;
        RECT 120.550 107.705 121.425 108.035 ;
        RECT 121.595 107.705 122.345 108.035 ;
        RECT 120.550 107.245 120.720 107.705 ;
        RECT 121.595 107.535 121.795 107.705 ;
        RECT 122.515 107.575 122.685 108.155 ;
        RECT 123.340 108.035 123.590 109.170 ;
        RECT 123.760 108.235 124.020 109.345 ;
        RECT 124.190 108.445 124.450 109.170 ;
        RECT 124.620 108.615 124.880 109.345 ;
        RECT 125.050 108.445 125.310 109.170 ;
        RECT 125.480 108.615 125.740 109.345 ;
        RECT 125.910 108.445 126.170 109.170 ;
        RECT 126.340 108.615 126.600 109.345 ;
        RECT 126.770 108.445 127.030 109.170 ;
        RECT 127.200 108.615 127.495 109.345 ;
        RECT 124.190 108.205 127.500 108.445 ;
        RECT 128.120 108.375 128.450 109.175 ;
        RECT 128.620 108.545 128.950 109.345 ;
        RECT 129.250 108.375 129.580 109.175 ;
        RECT 130.225 108.545 130.475 109.345 ;
        RECT 128.120 108.205 130.555 108.375 ;
        RECT 130.745 108.205 130.915 109.345 ;
        RECT 131.085 108.205 131.425 109.175 ;
        RECT 131.595 108.255 133.265 109.345 ;
        RECT 122.460 107.535 122.685 107.575 ;
        RECT 119.360 107.075 119.765 107.245 ;
        RECT 119.935 107.075 120.720 107.245 ;
        RECT 120.995 106.795 121.205 107.325 ;
        RECT 121.465 107.010 121.795 107.535 ;
        RECT 122.305 107.450 122.685 107.535 ;
        RECT 121.965 106.795 122.135 107.405 ;
        RECT 122.305 107.015 122.635 107.450 ;
        RECT 122.855 107.425 123.170 108.035 ;
        RECT 123.340 107.785 126.360 108.035 ;
        RECT 122.915 106.795 123.160 107.255 ;
        RECT 123.340 106.975 123.590 107.785 ;
        RECT 126.530 107.615 127.500 108.205 ;
        RECT 127.915 107.785 128.265 108.035 ;
        RECT 124.190 107.445 127.500 107.615 ;
        RECT 128.450 107.575 128.620 108.205 ;
        RECT 128.790 107.785 129.120 107.985 ;
        RECT 129.290 107.785 129.620 107.985 ;
        RECT 129.790 107.785 130.210 107.985 ;
        RECT 130.385 107.955 130.555 108.205 ;
        RECT 130.385 107.785 131.080 107.955 ;
        RECT 123.760 106.795 124.020 107.320 ;
        RECT 124.190 106.990 124.450 107.445 ;
        RECT 124.620 106.795 124.880 107.275 ;
        RECT 125.050 106.990 125.310 107.445 ;
        RECT 125.480 106.795 125.740 107.275 ;
        RECT 125.910 106.990 126.170 107.445 ;
        RECT 126.340 106.795 126.600 107.275 ;
        RECT 126.770 106.990 127.030 107.445 ;
        RECT 127.200 106.795 127.500 107.275 ;
        RECT 128.120 106.965 128.620 107.575 ;
        RECT 129.250 107.445 130.475 107.615 ;
        RECT 131.250 107.595 131.425 108.205 ;
        RECT 129.250 106.965 129.580 107.445 ;
        RECT 129.750 106.795 129.975 107.255 ;
        RECT 130.145 106.965 130.475 107.445 ;
        RECT 130.665 106.795 130.915 107.595 ;
        RECT 131.085 106.965 131.425 107.595 ;
        RECT 131.595 107.565 132.345 108.085 ;
        RECT 132.515 107.735 133.265 108.255 ;
        RECT 133.435 108.180 133.725 109.345 ;
        RECT 133.985 108.675 134.155 109.175 ;
        RECT 134.325 108.845 134.655 109.345 ;
        RECT 133.985 108.505 134.650 108.675 ;
        RECT 133.900 107.685 134.250 108.335 ;
        RECT 131.595 106.795 133.265 107.565 ;
        RECT 133.435 106.795 133.725 107.520 ;
        RECT 134.420 107.515 134.650 108.505 ;
        RECT 133.985 107.345 134.650 107.515 ;
        RECT 133.985 107.055 134.155 107.345 ;
        RECT 134.325 106.795 134.655 107.175 ;
        RECT 134.825 107.055 135.010 109.175 ;
        RECT 135.250 108.885 135.515 109.345 ;
        RECT 135.685 108.750 135.935 109.175 ;
        RECT 136.145 108.900 137.250 109.070 ;
        RECT 135.630 108.620 135.935 108.750 ;
        RECT 135.180 107.425 135.460 108.375 ;
        RECT 135.630 107.515 135.800 108.620 ;
        RECT 135.970 107.835 136.210 108.430 ;
        RECT 136.380 108.365 136.910 108.730 ;
        RECT 136.380 107.665 136.550 108.365 ;
        RECT 137.080 108.285 137.250 108.900 ;
        RECT 137.420 108.545 137.590 109.345 ;
        RECT 137.760 108.845 138.010 109.175 ;
        RECT 138.235 108.875 139.120 109.045 ;
        RECT 137.080 108.195 137.590 108.285 ;
        RECT 135.630 107.385 135.855 107.515 ;
        RECT 136.025 107.445 136.550 107.665 ;
        RECT 136.720 108.025 137.590 108.195 ;
        RECT 135.265 106.795 135.515 107.255 ;
        RECT 135.685 107.245 135.855 107.385 ;
        RECT 136.720 107.245 136.890 108.025 ;
        RECT 137.420 107.955 137.590 108.025 ;
        RECT 137.100 107.775 137.300 107.805 ;
        RECT 137.760 107.775 137.930 108.845 ;
        RECT 138.100 107.955 138.290 108.675 ;
        RECT 137.100 107.475 137.930 107.775 ;
        RECT 138.460 107.745 138.780 108.705 ;
        RECT 135.685 107.075 136.020 107.245 ;
        RECT 136.215 107.075 136.890 107.245 ;
        RECT 137.210 106.795 137.580 107.295 ;
        RECT 137.760 107.245 137.930 107.475 ;
        RECT 138.315 107.415 138.780 107.745 ;
        RECT 138.950 108.035 139.120 108.875 ;
        RECT 139.300 108.845 139.615 109.345 ;
        RECT 139.845 108.615 140.185 109.175 ;
        RECT 139.290 108.240 140.185 108.615 ;
        RECT 140.355 108.335 140.525 109.345 ;
        RECT 139.995 108.035 140.185 108.240 ;
        RECT 140.695 108.285 141.025 109.130 ;
        RECT 140.695 108.205 141.085 108.285 ;
        RECT 140.870 108.155 141.085 108.205 ;
        RECT 138.950 107.705 139.825 108.035 ;
        RECT 139.995 107.705 140.745 108.035 ;
        RECT 138.950 107.245 139.120 107.705 ;
        RECT 139.995 107.535 140.195 107.705 ;
        RECT 140.915 107.575 141.085 108.155 ;
        RECT 141.715 108.255 142.925 109.345 ;
        RECT 141.715 107.715 142.235 108.255 ;
        RECT 140.860 107.535 141.085 107.575 ;
        RECT 142.405 107.545 142.925 108.085 ;
        RECT 137.760 107.075 138.165 107.245 ;
        RECT 138.335 107.075 139.120 107.245 ;
        RECT 139.395 106.795 139.605 107.325 ;
        RECT 139.865 107.010 140.195 107.535 ;
        RECT 140.705 107.450 141.085 107.535 ;
        RECT 140.365 106.795 140.535 107.405 ;
        RECT 140.705 107.015 141.035 107.450 ;
        RECT 141.715 106.795 142.925 107.545 ;
        RECT 17.430 106.625 143.010 106.795 ;
        RECT 17.515 105.875 18.725 106.625 ;
        RECT 17.515 105.335 18.035 105.875 ;
        RECT 18.895 105.855 21.485 106.625 ;
        RECT 22.205 106.075 22.375 106.365 ;
        RECT 22.545 106.245 22.875 106.625 ;
        RECT 22.205 105.905 22.870 106.075 ;
        RECT 18.205 105.165 18.725 105.705 ;
        RECT 18.895 105.335 20.105 105.855 ;
        RECT 20.275 105.165 21.485 105.685 ;
        RECT 17.515 104.075 18.725 105.165 ;
        RECT 18.895 104.075 21.485 105.165 ;
        RECT 22.120 105.085 22.470 105.735 ;
        RECT 22.640 104.915 22.870 105.905 ;
        RECT 22.205 104.745 22.870 104.915 ;
        RECT 22.205 104.245 22.375 104.745 ;
        RECT 22.545 104.075 22.875 104.575 ;
        RECT 23.045 104.245 23.230 106.365 ;
        RECT 23.485 106.165 23.735 106.625 ;
        RECT 23.905 106.175 24.240 106.345 ;
        RECT 24.435 106.175 25.110 106.345 ;
        RECT 23.905 106.035 24.075 106.175 ;
        RECT 23.400 105.045 23.680 105.995 ;
        RECT 23.850 105.905 24.075 106.035 ;
        RECT 23.850 104.800 24.020 105.905 ;
        RECT 24.245 105.755 24.770 105.975 ;
        RECT 24.190 104.990 24.430 105.585 ;
        RECT 24.600 105.055 24.770 105.755 ;
        RECT 24.940 105.395 25.110 106.175 ;
        RECT 25.430 106.125 25.800 106.625 ;
        RECT 25.980 106.175 26.385 106.345 ;
        RECT 26.555 106.175 27.340 106.345 ;
        RECT 25.980 105.945 26.150 106.175 ;
        RECT 25.320 105.645 26.150 105.945 ;
        RECT 26.535 105.675 27.000 106.005 ;
        RECT 25.320 105.615 25.520 105.645 ;
        RECT 25.640 105.395 25.810 105.465 ;
        RECT 24.940 105.225 25.810 105.395 ;
        RECT 25.300 105.135 25.810 105.225 ;
        RECT 23.850 104.670 24.155 104.800 ;
        RECT 24.600 104.690 25.130 105.055 ;
        RECT 23.470 104.075 23.735 104.535 ;
        RECT 23.905 104.245 24.155 104.670 ;
        RECT 25.300 104.520 25.470 105.135 ;
        RECT 24.365 104.350 25.470 104.520 ;
        RECT 25.640 104.075 25.810 104.875 ;
        RECT 25.980 104.575 26.150 105.645 ;
        RECT 26.320 104.745 26.510 105.465 ;
        RECT 26.680 104.715 27.000 105.675 ;
        RECT 27.170 105.715 27.340 106.175 ;
        RECT 27.615 106.095 27.825 106.625 ;
        RECT 28.085 105.885 28.415 106.410 ;
        RECT 28.585 106.015 28.755 106.625 ;
        RECT 28.925 105.970 29.255 106.405 ;
        RECT 28.925 105.885 29.305 105.970 ;
        RECT 28.215 105.715 28.415 105.885 ;
        RECT 29.080 105.845 29.305 105.885 ;
        RECT 27.170 105.385 28.045 105.715 ;
        RECT 28.215 105.385 28.965 105.715 ;
        RECT 25.980 104.245 26.230 104.575 ;
        RECT 27.170 104.545 27.340 105.385 ;
        RECT 28.215 105.180 28.405 105.385 ;
        RECT 29.135 105.265 29.305 105.845 ;
        RECT 29.475 105.855 31.145 106.625 ;
        RECT 31.315 105.975 31.575 106.455 ;
        RECT 31.745 106.085 31.995 106.625 ;
        RECT 29.475 105.335 30.225 105.855 ;
        RECT 29.090 105.215 29.305 105.265 ;
        RECT 27.510 104.805 28.405 105.180 ;
        RECT 28.915 105.135 29.305 105.215 ;
        RECT 30.395 105.165 31.145 105.685 ;
        RECT 26.455 104.375 27.340 104.545 ;
        RECT 27.520 104.075 27.835 104.575 ;
        RECT 28.065 104.245 28.405 104.805 ;
        RECT 28.575 104.075 28.745 105.085 ;
        RECT 28.915 104.290 29.245 105.135 ;
        RECT 29.475 104.075 31.145 105.165 ;
        RECT 31.315 104.945 31.485 105.975 ;
        RECT 32.165 105.945 32.385 106.405 ;
        RECT 32.135 105.920 32.385 105.945 ;
        RECT 31.655 105.325 31.885 105.720 ;
        RECT 32.055 105.495 32.385 105.920 ;
        RECT 32.555 106.245 33.445 106.415 ;
        RECT 32.555 105.520 32.725 106.245 ;
        RECT 33.615 106.165 34.175 106.455 ;
        RECT 34.345 106.165 34.595 106.625 ;
        RECT 32.895 105.690 33.445 106.075 ;
        RECT 32.555 105.450 33.445 105.520 ;
        RECT 32.550 105.425 33.445 105.450 ;
        RECT 32.540 105.410 33.445 105.425 ;
        RECT 32.535 105.395 33.445 105.410 ;
        RECT 32.525 105.390 33.445 105.395 ;
        RECT 32.520 105.380 33.445 105.390 ;
        RECT 32.515 105.370 33.445 105.380 ;
        RECT 32.505 105.365 33.445 105.370 ;
        RECT 32.495 105.355 33.445 105.365 ;
        RECT 32.485 105.350 33.445 105.355 ;
        RECT 32.485 105.345 32.820 105.350 ;
        RECT 32.470 105.340 32.820 105.345 ;
        RECT 32.455 105.330 32.820 105.340 ;
        RECT 32.430 105.325 32.820 105.330 ;
        RECT 31.655 105.320 32.820 105.325 ;
        RECT 31.655 105.285 32.790 105.320 ;
        RECT 31.655 105.260 32.755 105.285 ;
        RECT 31.655 105.230 32.725 105.260 ;
        RECT 31.655 105.200 32.705 105.230 ;
        RECT 31.655 105.170 32.685 105.200 ;
        RECT 31.655 105.160 32.615 105.170 ;
        RECT 31.655 105.150 32.590 105.160 ;
        RECT 31.655 105.135 32.570 105.150 ;
        RECT 31.655 105.120 32.550 105.135 ;
        RECT 31.760 105.110 32.545 105.120 ;
        RECT 31.760 105.075 32.530 105.110 ;
        RECT 31.315 104.245 31.590 104.945 ;
        RECT 31.760 104.825 32.515 105.075 ;
        RECT 32.685 104.755 33.015 105.000 ;
        RECT 33.185 104.900 33.445 105.350 ;
        RECT 32.830 104.730 33.015 104.755 ;
        RECT 33.615 104.795 33.865 106.165 ;
        RECT 35.215 105.995 35.545 106.355 ;
        RECT 35.915 106.080 41.260 106.625 ;
        RECT 34.155 105.805 35.545 105.995 ;
        RECT 34.155 105.715 34.325 105.805 ;
        RECT 34.035 105.385 34.325 105.715 ;
        RECT 34.495 105.385 34.835 105.635 ;
        RECT 35.055 105.385 35.730 105.635 ;
        RECT 34.155 105.135 34.325 105.385 ;
        RECT 34.155 104.965 35.095 105.135 ;
        RECT 35.465 105.025 35.730 105.385 ;
        RECT 37.500 105.250 37.840 106.080 ;
        RECT 41.435 105.855 43.105 106.625 ;
        RECT 43.275 105.900 43.565 106.625 ;
        RECT 43.735 105.855 45.405 106.625 ;
        RECT 46.210 105.975 46.540 106.455 ;
        RECT 46.710 106.145 46.960 106.625 ;
        RECT 47.130 105.975 47.460 106.455 ;
        RECT 47.630 106.145 47.880 106.625 ;
        RECT 48.050 106.145 48.380 106.455 ;
        RECT 48.050 105.975 48.220 106.145 ;
        RECT 48.745 105.975 49.085 106.455 ;
        RECT 32.830 104.630 33.445 104.730 ;
        RECT 31.760 104.075 32.015 104.620 ;
        RECT 32.185 104.245 32.665 104.585 ;
        RECT 32.840 104.075 33.445 104.630 ;
        RECT 33.615 104.245 34.075 104.795 ;
        RECT 34.265 104.075 34.595 104.795 ;
        RECT 34.795 104.415 35.095 104.965 ;
        RECT 35.265 104.075 35.545 104.745 ;
        RECT 39.320 104.510 39.670 105.760 ;
        RECT 41.435 105.335 42.185 105.855 ;
        RECT 42.355 105.165 43.105 105.685 ;
        RECT 43.735 105.335 44.485 105.855 ;
        RECT 46.210 105.805 48.220 105.975 ;
        RECT 48.390 105.805 49.085 105.975 ;
        RECT 35.915 104.075 41.260 104.510 ;
        RECT 41.435 104.075 43.105 105.165 ;
        RECT 43.275 104.075 43.565 105.240 ;
        RECT 44.655 105.165 45.405 105.685 ;
        RECT 46.090 105.385 46.670 105.635 ;
        RECT 46.840 105.295 47.170 105.635 ;
        RECT 47.340 105.465 47.670 105.635 ;
        RECT 43.735 104.075 45.405 105.165 ;
        RECT 46.210 104.075 46.540 105.215 ;
        RECT 46.840 104.355 47.180 105.295 ;
        RECT 47.350 104.355 47.670 105.465 ;
        RECT 47.850 105.465 48.180 105.635 ;
        RECT 47.850 104.355 48.155 105.465 ;
        RECT 48.390 105.225 48.560 105.805 ;
        RECT 48.730 105.435 49.065 105.635 ;
        RECT 48.325 104.245 48.655 105.225 ;
        RECT 48.825 104.075 49.085 105.265 ;
        RECT 49.265 104.255 49.525 106.445 ;
        RECT 49.785 106.255 50.455 106.625 ;
        RECT 50.635 106.075 50.945 106.445 ;
        RECT 49.715 105.875 50.945 106.075 ;
        RECT 49.715 105.205 50.005 105.875 ;
        RECT 51.125 105.695 51.355 106.335 ;
        RECT 51.535 105.895 51.825 106.625 ;
        RECT 52.015 105.950 52.290 106.295 ;
        RECT 52.480 106.225 52.860 106.625 ;
        RECT 53.030 106.055 53.200 106.405 ;
        RECT 53.370 106.225 53.700 106.625 ;
        RECT 53.875 106.055 54.045 106.405 ;
        RECT 54.245 106.125 54.575 106.625 ;
        RECT 50.185 105.385 50.650 105.695 ;
        RECT 50.830 105.385 51.355 105.695 ;
        RECT 51.535 105.385 51.835 105.715 ;
        RECT 52.015 105.215 52.185 105.950 ;
        RECT 52.460 105.885 54.045 106.055 ;
        RECT 52.460 105.715 52.630 105.885 ;
        RECT 54.770 105.715 55.015 106.405 ;
        RECT 55.185 106.125 55.525 106.625 ;
        RECT 55.860 106.115 56.100 106.625 ;
        RECT 56.280 106.115 56.560 106.445 ;
        RECT 56.790 106.115 57.005 106.625 ;
        RECT 52.355 105.385 52.630 105.715 ;
        RECT 52.800 105.385 53.180 105.715 ;
        RECT 52.460 105.215 52.630 105.385 ;
        RECT 49.715 104.985 50.485 105.205 ;
        RECT 49.695 104.075 50.035 104.805 ;
        RECT 50.215 104.255 50.485 104.985 ;
        RECT 50.665 104.965 51.825 105.205 ;
        RECT 50.665 104.255 50.895 104.965 ;
        RECT 51.065 104.075 51.395 104.785 ;
        RECT 51.565 104.255 51.825 104.965 ;
        RECT 52.015 104.245 52.290 105.215 ;
        RECT 52.460 105.045 53.120 105.215 ;
        RECT 53.350 105.095 54.090 105.715 ;
        RECT 54.360 105.385 55.015 105.715 ;
        RECT 55.185 105.385 55.525 105.955 ;
        RECT 55.755 105.385 56.110 105.945 ;
        RECT 52.950 104.925 53.120 105.045 ;
        RECT 54.260 104.925 54.580 105.215 ;
        RECT 52.500 104.075 52.780 104.875 ;
        RECT 52.950 104.755 54.580 104.925 ;
        RECT 54.775 104.790 55.015 105.385 ;
        RECT 56.280 105.215 56.450 106.115 ;
        RECT 56.620 105.385 56.885 105.945 ;
        RECT 57.175 105.885 57.790 106.455 ;
        RECT 57.995 106.080 63.340 106.625 ;
        RECT 63.980 106.095 64.270 106.445 ;
        RECT 64.465 106.265 64.795 106.625 ;
        RECT 64.965 106.095 65.195 106.400 ;
        RECT 57.135 105.215 57.305 105.715 ;
        RECT 52.950 104.415 55.005 104.585 ;
        RECT 52.950 104.295 55.000 104.415 ;
        RECT 55.185 104.075 55.525 105.150 ;
        RECT 55.880 105.045 57.305 105.215 ;
        RECT 55.880 104.870 56.270 105.045 ;
        RECT 56.755 104.075 57.085 104.875 ;
        RECT 57.475 104.865 57.790 105.885 ;
        RECT 59.580 105.250 59.920 106.080 ;
        RECT 63.980 105.925 65.195 106.095 ;
        RECT 65.385 106.285 65.555 106.320 ;
        RECT 65.385 106.115 65.585 106.285 ;
        RECT 57.255 104.245 57.790 104.865 ;
        RECT 61.400 104.510 61.750 105.760 ;
        RECT 65.385 105.755 65.555 106.115 ;
        RECT 64.040 105.605 64.300 105.715 ;
        RECT 64.035 105.435 64.300 105.605 ;
        RECT 64.040 105.385 64.300 105.435 ;
        RECT 64.480 105.385 64.865 105.715 ;
        RECT 65.035 105.585 65.555 105.755 ;
        RECT 65.815 105.885 66.280 106.430 ;
        RECT 57.995 104.075 63.340 104.510 ;
        RECT 63.980 104.075 64.300 105.215 ;
        RECT 64.480 104.335 64.675 105.385 ;
        RECT 65.035 105.205 65.205 105.585 ;
        RECT 64.855 104.925 65.205 105.205 ;
        RECT 65.395 105.055 65.640 105.415 ;
        RECT 65.815 104.925 65.985 105.885 ;
        RECT 66.785 105.805 66.955 106.625 ;
        RECT 67.125 105.975 67.455 106.455 ;
        RECT 67.625 106.235 67.975 106.625 ;
        RECT 68.145 106.055 68.375 106.455 ;
        RECT 67.865 105.975 68.375 106.055 ;
        RECT 67.125 105.885 68.375 105.975 ;
        RECT 68.545 105.885 68.865 106.365 ;
        RECT 69.035 105.900 69.325 106.625 ;
        RECT 67.125 105.805 68.035 105.885 ;
        RECT 66.155 105.265 66.400 105.715 ;
        RECT 66.660 105.435 67.355 105.635 ;
        RECT 67.525 105.465 68.125 105.635 ;
        RECT 67.525 105.265 67.695 105.465 ;
        RECT 68.355 105.295 68.525 105.715 ;
        RECT 66.155 105.095 67.695 105.265 ;
        RECT 67.865 105.125 68.525 105.295 ;
        RECT 67.865 104.925 68.035 105.125 ;
        RECT 68.695 104.955 68.865 105.885 ;
        RECT 69.495 105.825 70.190 106.455 ;
        RECT 70.395 105.825 70.705 106.625 ;
        RECT 70.925 106.105 71.180 106.405 ;
        RECT 71.350 106.225 71.680 106.625 ;
        RECT 70.875 106.055 71.180 106.105 ;
        RECT 71.850 106.055 72.020 106.405 ;
        RECT 72.320 106.145 72.490 106.625 ;
        RECT 72.725 106.115 73.075 106.445 ;
        RECT 73.245 106.145 73.415 106.625 ;
        RECT 70.875 105.975 72.020 106.055 ;
        RECT 70.875 105.945 72.585 105.975 ;
        RECT 70.875 105.885 72.735 105.945 ;
        RECT 69.515 105.385 69.850 105.635 ;
        RECT 64.855 104.245 65.185 104.925 ;
        RECT 65.385 104.075 65.640 104.875 ;
        RECT 65.815 104.755 68.035 104.925 ;
        RECT 68.205 104.755 68.865 104.955 ;
        RECT 65.815 104.075 66.115 104.585 ;
        RECT 66.285 104.245 66.615 104.755 ;
        RECT 68.205 104.585 68.375 104.755 ;
        RECT 66.785 104.075 67.415 104.585 ;
        RECT 67.995 104.415 68.375 104.585 ;
        RECT 68.545 104.075 68.845 104.585 ;
        RECT 69.035 104.075 69.325 105.240 ;
        RECT 70.020 105.225 70.190 105.825 ;
        RECT 70.360 105.385 70.695 105.655 ;
        RECT 69.495 104.075 69.755 105.215 ;
        RECT 69.925 104.245 70.255 105.225 ;
        RECT 70.875 105.215 71.045 105.885 ;
        RECT 71.850 105.805 72.735 105.885 ;
        RECT 72.415 105.775 72.735 105.805 ;
        RECT 71.220 105.385 71.520 105.715 ;
        RECT 70.425 104.075 70.705 105.215 ;
        RECT 70.875 104.785 71.180 105.215 ;
        RECT 71.350 104.925 71.520 105.385 ;
        RECT 71.780 105.095 72.315 105.635 ;
        RECT 72.565 105.385 72.735 105.775 ;
        RECT 72.905 105.215 73.075 106.115 ;
        RECT 73.665 105.975 73.925 106.420 ;
        RECT 72.680 105.010 73.075 105.215 ;
        RECT 73.245 105.805 73.925 105.975 ;
        RECT 71.350 104.840 72.460 104.925 ;
        RECT 73.245 104.900 73.415 105.805 ;
        RECT 74.185 105.755 74.355 106.320 ;
        RECT 74.545 106.095 74.775 106.400 ;
        RECT 74.945 106.265 75.275 106.625 ;
        RECT 75.470 106.095 75.760 106.445 ;
        RECT 74.545 105.925 75.760 106.095 ;
        RECT 75.935 106.080 81.280 106.625 ;
        RECT 81.455 106.080 86.800 106.625 ;
        RECT 73.585 105.070 73.925 105.635 ;
        RECT 74.185 105.585 74.705 105.755 ;
        RECT 74.100 105.055 74.345 105.415 ;
        RECT 74.535 105.205 74.705 105.585 ;
        RECT 74.875 105.385 75.260 105.715 ;
        RECT 75.440 105.605 75.700 105.715 ;
        RECT 75.440 105.435 75.705 105.605 ;
        RECT 75.440 105.385 75.700 105.435 ;
        RECT 74.535 104.925 74.885 105.205 ;
        RECT 73.245 104.840 73.925 104.900 ;
        RECT 71.350 104.755 73.925 104.840 ;
        RECT 72.290 104.670 73.925 104.755 ;
        RECT 70.875 104.345 72.075 104.585 ;
        RECT 72.255 104.075 72.585 104.500 ;
        RECT 73.100 104.075 73.460 104.500 ;
        RECT 73.665 104.490 73.925 104.670 ;
        RECT 74.100 104.075 74.355 104.875 ;
        RECT 74.555 104.245 74.885 104.925 ;
        RECT 75.065 104.335 75.260 105.385 ;
        RECT 77.520 105.250 77.860 106.080 ;
        RECT 75.440 104.075 75.760 105.215 ;
        RECT 79.340 104.510 79.690 105.760 ;
        RECT 83.040 105.250 83.380 106.080 ;
        RECT 87.525 106.075 87.695 106.365 ;
        RECT 87.865 106.245 88.195 106.625 ;
        RECT 87.525 105.905 88.190 106.075 ;
        RECT 84.860 104.510 85.210 105.760 ;
        RECT 87.440 105.085 87.790 105.735 ;
        RECT 87.960 104.915 88.190 105.905 ;
        RECT 87.525 104.745 88.190 104.915 ;
        RECT 75.935 104.075 81.280 104.510 ;
        RECT 81.455 104.075 86.800 104.510 ;
        RECT 87.525 104.245 87.695 104.745 ;
        RECT 87.865 104.075 88.195 104.575 ;
        RECT 88.365 104.245 88.550 106.365 ;
        RECT 88.805 106.165 89.055 106.625 ;
        RECT 89.225 106.175 89.560 106.345 ;
        RECT 89.755 106.175 90.430 106.345 ;
        RECT 89.225 106.035 89.395 106.175 ;
        RECT 88.720 105.045 89.000 105.995 ;
        RECT 89.170 105.905 89.395 106.035 ;
        RECT 89.170 104.800 89.340 105.905 ;
        RECT 89.565 105.755 90.090 105.975 ;
        RECT 89.510 104.990 89.750 105.585 ;
        RECT 89.920 105.055 90.090 105.755 ;
        RECT 90.260 105.395 90.430 106.175 ;
        RECT 90.750 106.125 91.120 106.625 ;
        RECT 91.300 106.175 91.705 106.345 ;
        RECT 91.875 106.175 92.660 106.345 ;
        RECT 91.300 105.945 91.470 106.175 ;
        RECT 90.640 105.645 91.470 105.945 ;
        RECT 91.855 105.675 92.320 106.005 ;
        RECT 90.640 105.615 90.840 105.645 ;
        RECT 90.960 105.395 91.130 105.465 ;
        RECT 90.260 105.225 91.130 105.395 ;
        RECT 90.620 105.135 91.130 105.225 ;
        RECT 89.170 104.670 89.475 104.800 ;
        RECT 89.920 104.690 90.450 105.055 ;
        RECT 88.790 104.075 89.055 104.535 ;
        RECT 89.225 104.245 89.475 104.670 ;
        RECT 90.620 104.520 90.790 105.135 ;
        RECT 89.685 104.350 90.790 104.520 ;
        RECT 90.960 104.075 91.130 104.875 ;
        RECT 91.300 104.575 91.470 105.645 ;
        RECT 91.640 104.745 91.830 105.465 ;
        RECT 92.000 104.715 92.320 105.675 ;
        RECT 92.490 105.715 92.660 106.175 ;
        RECT 92.935 106.095 93.145 106.625 ;
        RECT 93.405 105.885 93.735 106.410 ;
        RECT 93.905 106.015 94.075 106.625 ;
        RECT 94.245 105.970 94.575 106.405 ;
        RECT 94.245 105.885 94.625 105.970 ;
        RECT 94.795 105.900 95.085 106.625 ;
        RECT 93.535 105.715 93.735 105.885 ;
        RECT 94.400 105.845 94.625 105.885 ;
        RECT 92.490 105.385 93.365 105.715 ;
        RECT 93.535 105.385 94.285 105.715 ;
        RECT 91.300 104.245 91.550 104.575 ;
        RECT 92.490 104.545 92.660 105.385 ;
        RECT 93.535 105.180 93.725 105.385 ;
        RECT 94.455 105.265 94.625 105.845 ;
        RECT 94.410 105.215 94.625 105.265 ;
        RECT 92.830 104.805 93.725 105.180 ;
        RECT 94.235 105.135 94.625 105.215 ;
        RECT 91.775 104.375 92.660 104.545 ;
        RECT 92.840 104.075 93.155 104.575 ;
        RECT 93.385 104.245 93.725 104.805 ;
        RECT 93.895 104.075 94.065 105.085 ;
        RECT 94.235 104.290 94.565 105.135 ;
        RECT 94.795 104.075 95.085 105.240 ;
        RECT 95.260 105.025 95.595 106.445 ;
        RECT 95.775 106.255 96.520 106.625 ;
        RECT 97.085 106.085 97.340 106.445 ;
        RECT 97.520 106.255 97.850 106.625 ;
        RECT 98.030 106.085 98.255 106.445 ;
        RECT 95.770 105.895 98.255 106.085 ;
        RECT 98.475 106.080 103.820 106.625 ;
        RECT 95.770 105.205 95.995 105.895 ;
        RECT 96.195 105.385 96.475 105.715 ;
        RECT 96.655 105.385 97.230 105.715 ;
        RECT 97.410 105.385 97.845 105.715 ;
        RECT 98.025 105.385 98.295 105.715 ;
        RECT 100.060 105.250 100.400 106.080 ;
        RECT 103.995 105.855 105.665 106.625 ;
        RECT 95.770 105.025 98.265 105.205 ;
        RECT 95.260 104.255 95.525 105.025 ;
        RECT 95.695 104.075 96.025 104.795 ;
        RECT 96.215 104.615 97.405 104.845 ;
        RECT 96.215 104.255 96.475 104.615 ;
        RECT 96.645 104.075 96.975 104.445 ;
        RECT 97.145 104.255 97.405 104.615 ;
        RECT 97.975 104.255 98.265 105.025 ;
        RECT 101.880 104.510 102.230 105.760 ;
        RECT 103.995 105.335 104.745 105.855 ;
        RECT 106.295 105.825 106.635 106.455 ;
        RECT 106.805 105.825 107.055 106.625 ;
        RECT 107.245 105.975 107.575 106.455 ;
        RECT 107.745 106.165 107.970 106.625 ;
        RECT 108.140 105.975 108.470 106.455 ;
        RECT 104.915 105.165 105.665 105.685 ;
        RECT 98.475 104.075 103.820 104.510 ;
        RECT 103.995 104.075 105.665 105.165 ;
        RECT 106.295 105.215 106.470 105.825 ;
        RECT 107.245 105.805 108.470 105.975 ;
        RECT 109.100 105.845 109.600 106.455 ;
        RECT 110.010 105.885 110.625 106.455 ;
        RECT 110.795 106.115 111.010 106.625 ;
        RECT 111.240 106.115 111.520 106.445 ;
        RECT 111.700 106.115 111.940 106.625 ;
        RECT 106.640 105.465 107.335 105.635 ;
        RECT 107.165 105.215 107.335 105.465 ;
        RECT 107.510 105.435 107.930 105.635 ;
        RECT 108.100 105.435 108.430 105.635 ;
        RECT 108.600 105.435 108.930 105.635 ;
        RECT 109.100 105.215 109.270 105.845 ;
        RECT 109.455 105.385 109.805 105.635 ;
        RECT 106.295 104.245 106.635 105.215 ;
        RECT 106.805 104.075 106.975 105.215 ;
        RECT 107.165 105.045 109.600 105.215 ;
        RECT 107.245 104.075 107.495 104.875 ;
        RECT 108.140 104.245 108.470 105.045 ;
        RECT 108.770 104.075 109.100 104.875 ;
        RECT 109.270 104.245 109.600 105.045 ;
        RECT 110.010 104.865 110.325 105.885 ;
        RECT 110.495 105.215 110.665 105.715 ;
        RECT 110.915 105.385 111.180 105.945 ;
        RECT 111.350 105.215 111.520 106.115 ;
        RECT 111.690 105.385 112.045 105.945 ;
        RECT 112.275 105.875 113.485 106.625 ;
        RECT 113.820 106.115 114.060 106.625 ;
        RECT 114.240 106.115 114.520 106.445 ;
        RECT 114.750 106.115 114.965 106.625 ;
        RECT 112.275 105.335 112.795 105.875 ;
        RECT 110.495 105.045 111.920 105.215 ;
        RECT 112.965 105.165 113.485 105.705 ;
        RECT 113.715 105.385 114.070 105.945 ;
        RECT 114.240 105.215 114.410 106.115 ;
        RECT 114.580 105.385 114.845 105.945 ;
        RECT 115.135 105.885 115.750 106.455 ;
        RECT 115.095 105.215 115.265 105.715 ;
        RECT 110.010 104.245 110.545 104.865 ;
        RECT 110.715 104.075 111.045 104.875 ;
        RECT 111.530 104.870 111.920 105.045 ;
        RECT 112.275 104.075 113.485 105.165 ;
        RECT 113.840 105.045 115.265 105.215 ;
        RECT 113.840 104.870 114.230 105.045 ;
        RECT 114.715 104.075 115.045 104.875 ;
        RECT 115.435 104.865 115.750 105.885 ;
        RECT 115.215 104.245 115.750 104.865 ;
        RECT 115.955 105.825 116.295 106.455 ;
        RECT 116.465 105.825 116.715 106.625 ;
        RECT 116.905 105.975 117.235 106.455 ;
        RECT 117.405 106.165 117.630 106.625 ;
        RECT 117.800 105.975 118.130 106.455 ;
        RECT 115.955 105.215 116.130 105.825 ;
        RECT 116.905 105.805 118.130 105.975 ;
        RECT 118.760 105.845 119.260 106.455 ;
        RECT 120.555 105.900 120.845 106.625 ;
        RECT 121.075 106.165 121.320 106.625 ;
        RECT 116.300 105.465 116.995 105.635 ;
        RECT 116.825 105.215 116.995 105.465 ;
        RECT 117.170 105.435 117.590 105.635 ;
        RECT 117.760 105.435 118.090 105.635 ;
        RECT 118.260 105.435 118.590 105.635 ;
        RECT 118.760 105.215 118.930 105.845 ;
        RECT 119.115 105.385 119.465 105.635 ;
        RECT 121.015 105.385 121.330 105.995 ;
        RECT 121.500 105.635 121.750 106.445 ;
        RECT 121.920 106.100 122.180 106.625 ;
        RECT 122.350 105.975 122.610 106.430 ;
        RECT 122.780 106.145 123.040 106.625 ;
        RECT 123.210 105.975 123.470 106.430 ;
        RECT 123.640 106.145 123.900 106.625 ;
        RECT 124.070 105.975 124.330 106.430 ;
        RECT 124.500 106.145 124.760 106.625 ;
        RECT 124.930 105.975 125.190 106.430 ;
        RECT 125.360 106.145 125.660 106.625 ;
        RECT 122.350 105.805 125.660 105.975 ;
        RECT 121.500 105.385 124.520 105.635 ;
        RECT 115.955 104.245 116.295 105.215 ;
        RECT 116.465 104.075 116.635 105.215 ;
        RECT 116.825 105.045 119.260 105.215 ;
        RECT 116.905 104.075 117.155 104.875 ;
        RECT 117.800 104.245 118.130 105.045 ;
        RECT 118.430 104.075 118.760 104.875 ;
        RECT 118.930 104.245 119.260 105.045 ;
        RECT 120.555 104.075 120.845 105.240 ;
        RECT 121.025 104.075 121.320 105.185 ;
        RECT 121.500 104.250 121.750 105.385 ;
        RECT 124.690 105.215 125.660 105.805 ;
        RECT 126.075 105.855 127.745 106.625 ;
        RECT 126.075 105.335 126.825 105.855 ;
        RECT 128.120 105.845 128.620 106.455 ;
        RECT 121.920 104.075 122.180 105.185 ;
        RECT 122.350 104.975 125.660 105.215 ;
        RECT 126.995 105.165 127.745 105.685 ;
        RECT 127.915 105.385 128.265 105.635 ;
        RECT 128.450 105.215 128.620 105.845 ;
        RECT 129.250 105.975 129.580 106.455 ;
        RECT 129.750 106.165 129.975 106.625 ;
        RECT 130.145 105.975 130.475 106.455 ;
        RECT 129.250 105.805 130.475 105.975 ;
        RECT 130.665 105.825 130.915 106.625 ;
        RECT 131.085 105.825 131.425 106.455 ;
        RECT 131.685 106.075 131.855 106.365 ;
        RECT 132.025 106.245 132.355 106.625 ;
        RECT 131.685 105.905 132.350 106.075 ;
        RECT 128.790 105.435 129.120 105.635 ;
        RECT 129.290 105.435 129.620 105.635 ;
        RECT 129.790 105.435 130.210 105.635 ;
        RECT 130.385 105.465 131.080 105.635 ;
        RECT 130.385 105.215 130.555 105.465 ;
        RECT 131.250 105.265 131.425 105.825 ;
        RECT 131.195 105.215 131.425 105.265 ;
        RECT 122.350 104.250 122.610 104.975 ;
        RECT 122.780 104.075 123.040 104.805 ;
        RECT 123.210 104.250 123.470 104.975 ;
        RECT 123.640 104.075 123.900 104.805 ;
        RECT 124.070 104.250 124.330 104.975 ;
        RECT 124.500 104.075 124.760 104.805 ;
        RECT 124.930 104.250 125.190 104.975 ;
        RECT 125.360 104.075 125.655 104.805 ;
        RECT 126.075 104.075 127.745 105.165 ;
        RECT 128.120 105.045 130.555 105.215 ;
        RECT 128.120 104.245 128.450 105.045 ;
        RECT 128.620 104.075 128.950 104.875 ;
        RECT 129.250 104.245 129.580 105.045 ;
        RECT 130.225 104.075 130.475 104.875 ;
        RECT 130.745 104.075 130.915 105.215 ;
        RECT 131.085 104.245 131.425 105.215 ;
        RECT 131.600 105.085 131.950 105.735 ;
        RECT 132.120 104.915 132.350 105.905 ;
        RECT 131.685 104.745 132.350 104.915 ;
        RECT 131.685 104.245 131.855 104.745 ;
        RECT 132.025 104.075 132.355 104.575 ;
        RECT 132.525 104.245 132.710 106.365 ;
        RECT 132.965 106.165 133.215 106.625 ;
        RECT 133.385 106.175 133.720 106.345 ;
        RECT 133.915 106.175 134.590 106.345 ;
        RECT 133.385 106.035 133.555 106.175 ;
        RECT 132.880 105.045 133.160 105.995 ;
        RECT 133.330 105.905 133.555 106.035 ;
        RECT 133.330 104.800 133.500 105.905 ;
        RECT 133.725 105.755 134.250 105.975 ;
        RECT 133.670 104.990 133.910 105.585 ;
        RECT 134.080 105.055 134.250 105.755 ;
        RECT 134.420 105.395 134.590 106.175 ;
        RECT 134.910 106.125 135.280 106.625 ;
        RECT 135.460 106.175 135.865 106.345 ;
        RECT 136.035 106.175 136.820 106.345 ;
        RECT 135.460 105.945 135.630 106.175 ;
        RECT 134.800 105.645 135.630 105.945 ;
        RECT 136.015 105.675 136.480 106.005 ;
        RECT 134.800 105.615 135.000 105.645 ;
        RECT 135.120 105.395 135.290 105.465 ;
        RECT 134.420 105.225 135.290 105.395 ;
        RECT 134.780 105.135 135.290 105.225 ;
        RECT 133.330 104.670 133.635 104.800 ;
        RECT 134.080 104.690 134.610 105.055 ;
        RECT 132.950 104.075 133.215 104.535 ;
        RECT 133.385 104.245 133.635 104.670 ;
        RECT 134.780 104.520 134.950 105.135 ;
        RECT 133.845 104.350 134.950 104.520 ;
        RECT 135.120 104.075 135.290 104.875 ;
        RECT 135.460 104.575 135.630 105.645 ;
        RECT 135.800 104.745 135.990 105.465 ;
        RECT 136.160 104.715 136.480 105.675 ;
        RECT 136.650 105.715 136.820 106.175 ;
        RECT 137.095 106.095 137.305 106.625 ;
        RECT 137.565 105.885 137.895 106.410 ;
        RECT 138.065 106.015 138.235 106.625 ;
        RECT 138.405 105.970 138.735 106.405 ;
        RECT 139.965 106.075 140.135 106.455 ;
        RECT 140.350 106.245 140.680 106.625 ;
        RECT 138.405 105.885 138.785 105.970 ;
        RECT 139.965 105.905 140.680 106.075 ;
        RECT 137.695 105.715 137.895 105.885 ;
        RECT 138.560 105.845 138.785 105.885 ;
        RECT 136.650 105.385 137.525 105.715 ;
        RECT 137.695 105.385 138.445 105.715 ;
        RECT 135.460 104.245 135.710 104.575 ;
        RECT 136.650 104.545 136.820 105.385 ;
        RECT 137.695 105.180 137.885 105.385 ;
        RECT 138.615 105.265 138.785 105.845 ;
        RECT 139.875 105.355 140.230 105.725 ;
        RECT 140.510 105.715 140.680 105.905 ;
        RECT 140.850 105.880 141.105 106.455 ;
        RECT 140.510 105.385 140.765 105.715 ;
        RECT 138.570 105.215 138.785 105.265 ;
        RECT 136.990 104.805 137.885 105.180 ;
        RECT 138.395 105.135 138.785 105.215 ;
        RECT 140.510 105.175 140.680 105.385 ;
        RECT 135.935 104.375 136.820 104.545 ;
        RECT 137.000 104.075 137.315 104.575 ;
        RECT 137.545 104.245 137.885 104.805 ;
        RECT 138.055 104.075 138.225 105.085 ;
        RECT 138.395 104.290 138.725 105.135 ;
        RECT 139.965 105.005 140.680 105.175 ;
        RECT 140.935 105.150 141.105 105.880 ;
        RECT 141.280 105.785 141.540 106.625 ;
        RECT 141.715 105.875 142.925 106.625 ;
        RECT 139.965 104.245 140.135 105.005 ;
        RECT 140.350 104.075 140.680 104.835 ;
        RECT 140.850 104.245 141.105 105.150 ;
        RECT 141.280 104.075 141.540 105.225 ;
        RECT 141.715 105.165 142.235 105.705 ;
        RECT 142.405 105.335 142.925 105.875 ;
        RECT 141.715 104.075 142.925 105.165 ;
        RECT 17.430 103.905 143.010 104.075 ;
        RECT 17.515 102.815 18.725 103.905 ;
        RECT 18.895 102.815 21.485 103.905 ;
        RECT 21.745 103.235 21.915 103.735 ;
        RECT 22.085 103.405 22.415 103.905 ;
        RECT 21.745 103.065 22.410 103.235 ;
        RECT 17.515 102.105 18.035 102.645 ;
        RECT 18.205 102.275 18.725 102.815 ;
        RECT 18.895 102.125 20.105 102.645 ;
        RECT 20.275 102.295 21.485 102.815 ;
        RECT 21.660 102.245 22.010 102.895 ;
        RECT 17.515 101.355 18.725 102.105 ;
        RECT 18.895 101.355 21.485 102.125 ;
        RECT 22.180 102.075 22.410 103.065 ;
        RECT 21.745 101.905 22.410 102.075 ;
        RECT 21.745 101.615 21.915 101.905 ;
        RECT 22.085 101.355 22.415 101.735 ;
        RECT 22.585 101.615 22.770 103.735 ;
        RECT 23.010 103.445 23.275 103.905 ;
        RECT 23.445 103.310 23.695 103.735 ;
        RECT 23.905 103.460 25.010 103.630 ;
        RECT 23.390 103.180 23.695 103.310 ;
        RECT 22.940 101.985 23.220 102.935 ;
        RECT 23.390 102.075 23.560 103.180 ;
        RECT 23.730 102.395 23.970 102.990 ;
        RECT 24.140 102.925 24.670 103.290 ;
        RECT 24.140 102.225 24.310 102.925 ;
        RECT 24.840 102.845 25.010 103.460 ;
        RECT 25.180 103.105 25.350 103.905 ;
        RECT 25.520 103.405 25.770 103.735 ;
        RECT 25.995 103.435 26.880 103.605 ;
        RECT 24.840 102.755 25.350 102.845 ;
        RECT 23.390 101.945 23.615 102.075 ;
        RECT 23.785 102.005 24.310 102.225 ;
        RECT 24.480 102.585 25.350 102.755 ;
        RECT 23.025 101.355 23.275 101.815 ;
        RECT 23.445 101.805 23.615 101.945 ;
        RECT 24.480 101.805 24.650 102.585 ;
        RECT 25.180 102.515 25.350 102.585 ;
        RECT 24.860 102.335 25.060 102.365 ;
        RECT 25.520 102.335 25.690 103.405 ;
        RECT 25.860 102.515 26.050 103.235 ;
        RECT 24.860 102.035 25.690 102.335 ;
        RECT 26.220 102.305 26.540 103.265 ;
        RECT 23.445 101.635 23.780 101.805 ;
        RECT 23.975 101.635 24.650 101.805 ;
        RECT 24.970 101.355 25.340 101.855 ;
        RECT 25.520 101.805 25.690 102.035 ;
        RECT 26.075 101.975 26.540 102.305 ;
        RECT 26.710 102.595 26.880 103.435 ;
        RECT 27.060 103.405 27.375 103.905 ;
        RECT 27.605 103.175 27.945 103.735 ;
        RECT 27.050 102.800 27.945 103.175 ;
        RECT 28.115 102.895 28.285 103.905 ;
        RECT 27.755 102.595 27.945 102.800 ;
        RECT 28.455 102.845 28.785 103.690 ;
        RECT 28.455 102.765 28.845 102.845 ;
        RECT 29.015 102.815 30.225 103.905 ;
        RECT 28.630 102.715 28.845 102.765 ;
        RECT 26.710 102.265 27.585 102.595 ;
        RECT 27.755 102.265 28.505 102.595 ;
        RECT 26.710 101.805 26.880 102.265 ;
        RECT 27.755 102.095 27.955 102.265 ;
        RECT 28.675 102.135 28.845 102.715 ;
        RECT 28.620 102.095 28.845 102.135 ;
        RECT 25.520 101.635 25.925 101.805 ;
        RECT 26.095 101.635 26.880 101.805 ;
        RECT 27.155 101.355 27.365 101.885 ;
        RECT 27.625 101.570 27.955 102.095 ;
        RECT 28.465 102.010 28.845 102.095 ;
        RECT 29.015 102.105 29.535 102.645 ;
        RECT 29.705 102.275 30.225 102.815 ;
        RECT 30.395 102.740 30.685 103.905 ;
        RECT 30.860 103.525 31.195 103.905 ;
        RECT 28.125 101.355 28.295 101.965 ;
        RECT 28.465 101.575 28.795 102.010 ;
        RECT 29.015 101.355 30.225 102.105 ;
        RECT 30.395 101.355 30.685 102.080 ;
        RECT 30.855 102.035 31.095 103.345 ;
        RECT 31.365 102.935 31.615 103.735 ;
        RECT 31.835 103.185 32.165 103.905 ;
        RECT 32.350 102.935 32.600 103.735 ;
        RECT 33.065 103.105 33.395 103.905 ;
        RECT 33.565 103.475 33.905 103.735 ;
        RECT 31.265 102.765 33.455 102.935 ;
        RECT 31.265 101.855 31.435 102.765 ;
        RECT 33.140 102.595 33.455 102.765 ;
        RECT 30.940 101.525 31.435 101.855 ;
        RECT 31.655 101.630 32.005 102.595 ;
        RECT 32.185 101.625 32.485 102.595 ;
        RECT 32.665 101.625 32.945 102.595 ;
        RECT 33.140 102.345 33.470 102.595 ;
        RECT 33.125 101.355 33.395 102.155 ;
        RECT 33.645 102.075 33.905 103.475 ;
        RECT 34.075 103.470 39.420 103.905 ;
        RECT 39.595 103.470 44.940 103.905 ;
        RECT 33.565 101.565 33.905 102.075 ;
        RECT 35.660 101.900 36.000 102.730 ;
        RECT 37.480 102.220 37.830 103.470 ;
        RECT 41.180 101.900 41.520 102.730 ;
        RECT 43.000 102.220 43.350 103.470 ;
        RECT 45.115 102.815 46.785 103.905 ;
        RECT 45.115 102.125 45.865 102.645 ;
        RECT 46.035 102.295 46.785 102.815 ;
        RECT 46.955 102.935 47.225 103.705 ;
        RECT 47.395 103.125 47.725 103.905 ;
        RECT 47.930 103.300 48.115 103.705 ;
        RECT 48.285 103.480 48.620 103.905 ;
        RECT 47.930 103.125 48.595 103.300 ;
        RECT 46.955 102.765 48.085 102.935 ;
        RECT 34.075 101.355 39.420 101.900 ;
        RECT 39.595 101.355 44.940 101.900 ;
        RECT 45.115 101.355 46.785 102.125 ;
        RECT 46.955 101.855 47.125 102.765 ;
        RECT 47.295 102.015 47.655 102.595 ;
        RECT 47.835 102.265 48.085 102.765 ;
        RECT 48.255 102.095 48.595 103.125 ;
        RECT 48.855 102.845 49.185 103.690 ;
        RECT 49.355 102.895 49.525 103.905 ;
        RECT 49.695 103.175 50.035 103.735 ;
        RECT 50.265 103.405 50.580 103.905 ;
        RECT 50.760 103.435 51.645 103.605 ;
        RECT 47.910 101.925 48.595 102.095 ;
        RECT 48.795 102.765 49.185 102.845 ;
        RECT 49.695 102.800 50.590 103.175 ;
        RECT 48.795 102.715 49.010 102.765 ;
        RECT 48.795 102.135 48.965 102.715 ;
        RECT 49.695 102.595 49.885 102.800 ;
        RECT 50.760 102.595 50.930 103.435 ;
        RECT 51.870 103.405 52.120 103.735 ;
        RECT 49.135 102.265 49.885 102.595 ;
        RECT 50.055 102.265 50.930 102.595 ;
        RECT 48.795 102.095 49.020 102.135 ;
        RECT 49.685 102.095 49.885 102.265 ;
        RECT 48.795 102.010 49.175 102.095 ;
        RECT 46.955 101.525 47.215 101.855 ;
        RECT 47.425 101.355 47.700 101.835 ;
        RECT 47.910 101.525 48.115 101.925 ;
        RECT 48.285 101.355 48.620 101.755 ;
        RECT 48.845 101.575 49.175 102.010 ;
        RECT 49.345 101.355 49.515 101.965 ;
        RECT 49.685 101.570 50.015 102.095 ;
        RECT 50.275 101.355 50.485 101.885 ;
        RECT 50.760 101.805 50.930 102.265 ;
        RECT 51.100 102.305 51.420 103.265 ;
        RECT 51.590 102.515 51.780 103.235 ;
        RECT 51.950 102.335 52.120 103.405 ;
        RECT 52.290 103.105 52.460 103.905 ;
        RECT 52.630 103.460 53.735 103.630 ;
        RECT 52.630 102.845 52.800 103.460 ;
        RECT 53.945 103.310 54.195 103.735 ;
        RECT 54.365 103.445 54.630 103.905 ;
        RECT 52.970 102.925 53.500 103.290 ;
        RECT 53.945 103.180 54.250 103.310 ;
        RECT 52.290 102.755 52.800 102.845 ;
        RECT 52.290 102.585 53.160 102.755 ;
        RECT 52.290 102.515 52.460 102.585 ;
        RECT 52.580 102.335 52.780 102.365 ;
        RECT 51.100 101.975 51.565 102.305 ;
        RECT 51.950 102.035 52.780 102.335 ;
        RECT 51.950 101.805 52.120 102.035 ;
        RECT 50.760 101.635 51.545 101.805 ;
        RECT 51.715 101.635 52.120 101.805 ;
        RECT 52.300 101.355 52.670 101.855 ;
        RECT 52.990 101.805 53.160 102.585 ;
        RECT 53.330 102.225 53.500 102.925 ;
        RECT 53.670 102.395 53.910 102.990 ;
        RECT 53.330 102.005 53.855 102.225 ;
        RECT 54.080 102.075 54.250 103.180 ;
        RECT 54.025 101.945 54.250 102.075 ;
        RECT 54.420 101.985 54.700 102.935 ;
        RECT 54.025 101.805 54.195 101.945 ;
        RECT 52.990 101.635 53.665 101.805 ;
        RECT 53.860 101.635 54.195 101.805 ;
        RECT 54.365 101.355 54.615 101.815 ;
        RECT 54.870 101.615 55.055 103.735 ;
        RECT 55.225 103.405 55.555 103.905 ;
        RECT 55.725 103.235 55.895 103.735 ;
        RECT 55.230 103.065 55.895 103.235 ;
        RECT 55.230 102.075 55.460 103.065 ;
        RECT 55.630 102.245 55.980 102.895 ;
        RECT 56.155 102.740 56.445 103.905 ;
        RECT 56.730 103.275 57.015 103.735 ;
        RECT 57.185 103.445 57.455 103.905 ;
        RECT 56.730 103.055 57.685 103.275 ;
        RECT 56.615 102.325 57.305 102.885 ;
        RECT 57.475 102.155 57.685 103.055 ;
        RECT 55.230 101.905 55.895 102.075 ;
        RECT 55.225 101.355 55.555 101.735 ;
        RECT 55.725 101.615 55.895 101.905 ;
        RECT 56.155 101.355 56.445 102.080 ;
        RECT 56.730 101.985 57.685 102.155 ;
        RECT 57.855 102.885 58.255 103.735 ;
        RECT 58.445 103.275 58.725 103.735 ;
        RECT 59.245 103.445 59.570 103.905 ;
        RECT 58.445 103.055 59.570 103.275 ;
        RECT 57.855 102.325 58.950 102.885 ;
        RECT 59.120 102.595 59.570 103.055 ;
        RECT 59.740 102.765 60.125 103.735 ;
        RECT 60.335 102.765 60.565 103.905 ;
        RECT 56.730 101.525 57.015 101.985 ;
        RECT 57.185 101.355 57.455 101.815 ;
        RECT 57.855 101.525 58.255 102.325 ;
        RECT 59.120 102.265 59.675 102.595 ;
        RECT 59.120 102.155 59.570 102.265 ;
        RECT 58.445 101.985 59.570 102.155 ;
        RECT 59.845 102.095 60.125 102.765 ;
        RECT 60.735 102.755 61.065 103.735 ;
        RECT 61.235 102.765 61.445 103.905 ;
        RECT 61.675 102.815 65.185 103.905 ;
        RECT 60.315 102.345 60.645 102.595 ;
        RECT 58.445 101.525 58.725 101.985 ;
        RECT 59.245 101.355 59.570 101.815 ;
        RECT 59.740 101.525 60.125 102.095 ;
        RECT 60.335 101.355 60.565 102.175 ;
        RECT 60.815 102.155 61.065 102.755 ;
        RECT 60.735 101.525 61.065 102.155 ;
        RECT 61.235 101.355 61.445 102.175 ;
        RECT 61.675 102.125 63.325 102.645 ;
        RECT 63.495 102.295 65.185 102.815 ;
        RECT 65.360 102.765 65.680 103.905 ;
        RECT 65.860 102.595 66.055 103.645 ;
        RECT 66.235 103.055 66.565 103.735 ;
        RECT 66.765 103.105 67.020 103.905 ;
        RECT 67.285 103.235 67.455 103.735 ;
        RECT 67.625 103.405 67.955 103.905 ;
        RECT 67.285 103.065 67.950 103.235 ;
        RECT 66.235 102.775 66.585 103.055 ;
        RECT 65.420 102.545 65.680 102.595 ;
        RECT 65.415 102.375 65.680 102.545 ;
        RECT 65.420 102.265 65.680 102.375 ;
        RECT 65.860 102.265 66.245 102.595 ;
        RECT 66.415 102.395 66.585 102.775 ;
        RECT 66.775 102.565 67.020 102.925 ;
        RECT 66.415 102.225 66.935 102.395 ;
        RECT 67.200 102.245 67.550 102.895 ;
        RECT 61.675 101.355 65.185 102.125 ;
        RECT 65.360 101.885 66.575 102.055 ;
        RECT 65.360 101.535 65.650 101.885 ;
        RECT 65.845 101.355 66.175 101.715 ;
        RECT 66.345 101.580 66.575 101.885 ;
        RECT 66.765 101.865 66.935 102.225 ;
        RECT 67.720 102.075 67.950 103.065 ;
        RECT 67.285 101.905 67.950 102.075 ;
        RECT 66.765 101.695 66.965 101.865 ;
        RECT 66.765 101.660 66.935 101.695 ;
        RECT 67.285 101.615 67.455 101.905 ;
        RECT 67.625 101.355 67.955 101.735 ;
        RECT 68.125 101.615 68.310 103.735 ;
        RECT 68.550 103.445 68.815 103.905 ;
        RECT 68.985 103.310 69.235 103.735 ;
        RECT 69.445 103.460 70.550 103.630 ;
        RECT 68.930 103.180 69.235 103.310 ;
        RECT 68.480 101.985 68.760 102.935 ;
        RECT 68.930 102.075 69.100 103.180 ;
        RECT 69.270 102.395 69.510 102.990 ;
        RECT 69.680 102.925 70.210 103.290 ;
        RECT 69.680 102.225 69.850 102.925 ;
        RECT 70.380 102.845 70.550 103.460 ;
        RECT 70.720 103.105 70.890 103.905 ;
        RECT 71.060 103.405 71.310 103.735 ;
        RECT 71.535 103.435 72.420 103.605 ;
        RECT 70.380 102.755 70.890 102.845 ;
        RECT 68.930 101.945 69.155 102.075 ;
        RECT 69.325 102.005 69.850 102.225 ;
        RECT 70.020 102.585 70.890 102.755 ;
        RECT 68.565 101.355 68.815 101.815 ;
        RECT 68.985 101.805 69.155 101.945 ;
        RECT 70.020 101.805 70.190 102.585 ;
        RECT 70.720 102.515 70.890 102.585 ;
        RECT 70.400 102.335 70.600 102.365 ;
        RECT 71.060 102.335 71.230 103.405 ;
        RECT 71.400 102.515 71.590 103.235 ;
        RECT 70.400 102.035 71.230 102.335 ;
        RECT 71.760 102.305 72.080 103.265 ;
        RECT 68.985 101.635 69.320 101.805 ;
        RECT 69.515 101.635 70.190 101.805 ;
        RECT 70.510 101.355 70.880 101.855 ;
        RECT 71.060 101.805 71.230 102.035 ;
        RECT 71.615 101.975 72.080 102.305 ;
        RECT 72.250 102.595 72.420 103.435 ;
        RECT 72.600 103.405 72.915 103.905 ;
        RECT 73.145 103.175 73.485 103.735 ;
        RECT 72.590 102.800 73.485 103.175 ;
        RECT 73.655 102.895 73.825 103.905 ;
        RECT 73.295 102.595 73.485 102.800 ;
        RECT 73.995 102.845 74.325 103.690 ;
        RECT 74.555 103.470 79.900 103.905 ;
        RECT 73.995 102.765 74.385 102.845 ;
        RECT 74.170 102.715 74.385 102.765 ;
        RECT 72.250 102.265 73.125 102.595 ;
        RECT 73.295 102.265 74.045 102.595 ;
        RECT 72.250 101.805 72.420 102.265 ;
        RECT 73.295 102.095 73.495 102.265 ;
        RECT 74.215 102.135 74.385 102.715 ;
        RECT 74.160 102.095 74.385 102.135 ;
        RECT 71.060 101.635 71.465 101.805 ;
        RECT 71.635 101.635 72.420 101.805 ;
        RECT 72.695 101.355 72.905 101.885 ;
        RECT 73.165 101.570 73.495 102.095 ;
        RECT 74.005 102.010 74.385 102.095 ;
        RECT 73.665 101.355 73.835 101.965 ;
        RECT 74.005 101.575 74.335 102.010 ;
        RECT 76.140 101.900 76.480 102.730 ;
        RECT 77.960 102.220 78.310 103.470 ;
        RECT 80.075 102.815 81.745 103.905 ;
        RECT 80.075 102.125 80.825 102.645 ;
        RECT 80.995 102.295 81.745 102.815 ;
        RECT 81.915 102.740 82.205 103.905 ;
        RECT 82.560 102.935 82.950 103.110 ;
        RECT 83.435 103.105 83.765 103.905 ;
        RECT 83.935 103.115 84.470 103.735 ;
        RECT 82.560 102.765 83.985 102.935 ;
        RECT 74.555 101.355 79.900 101.900 ;
        RECT 80.075 101.355 81.745 102.125 ;
        RECT 81.915 101.355 82.205 102.080 ;
        RECT 82.435 102.035 82.790 102.595 ;
        RECT 82.960 101.865 83.130 102.765 ;
        RECT 83.300 102.035 83.565 102.595 ;
        RECT 83.815 102.265 83.985 102.765 ;
        RECT 84.155 102.095 84.470 103.115 ;
        RECT 84.675 102.815 86.345 103.905 ;
        RECT 82.540 101.355 82.780 101.865 ;
        RECT 82.960 101.535 83.240 101.865 ;
        RECT 83.470 101.355 83.685 101.865 ;
        RECT 83.855 101.525 84.470 102.095 ;
        RECT 84.675 102.125 85.425 102.645 ;
        RECT 85.595 102.295 86.345 102.815 ;
        RECT 86.520 102.955 86.785 103.725 ;
        RECT 86.955 103.185 87.285 103.905 ;
        RECT 87.475 103.365 87.735 103.725 ;
        RECT 87.905 103.535 88.235 103.905 ;
        RECT 88.405 103.365 88.665 103.725 ;
        RECT 87.475 103.135 88.665 103.365 ;
        RECT 89.235 102.955 89.525 103.725 ;
        RECT 90.905 103.175 91.200 103.905 ;
        RECT 91.370 103.005 91.630 103.730 ;
        RECT 91.800 103.175 92.060 103.905 ;
        RECT 92.230 103.005 92.490 103.730 ;
        RECT 92.660 103.175 92.920 103.905 ;
        RECT 93.090 103.005 93.350 103.730 ;
        RECT 93.520 103.175 93.780 103.905 ;
        RECT 93.950 103.005 94.210 103.730 ;
        RECT 84.675 101.355 86.345 102.125 ;
        RECT 86.520 101.535 86.855 102.955 ;
        RECT 87.030 102.775 89.525 102.955 ;
        RECT 87.030 102.085 87.255 102.775 ;
        RECT 90.900 102.765 94.210 103.005 ;
        RECT 94.380 102.795 94.640 103.905 ;
        RECT 87.455 102.265 87.735 102.595 ;
        RECT 87.915 102.265 88.490 102.595 ;
        RECT 88.670 102.265 89.105 102.595 ;
        RECT 89.285 102.265 89.555 102.595 ;
        RECT 90.900 102.175 91.870 102.765 ;
        RECT 94.810 102.595 95.060 103.730 ;
        RECT 95.240 102.795 95.535 103.905 ;
        RECT 95.750 103.115 96.285 103.735 ;
        RECT 92.040 102.345 95.060 102.595 ;
        RECT 87.030 101.895 89.515 102.085 ;
        RECT 90.900 102.005 94.210 102.175 ;
        RECT 87.035 101.355 87.780 101.725 ;
        RECT 88.345 101.535 88.600 101.895 ;
        RECT 88.780 101.355 89.110 101.725 ;
        RECT 89.290 101.535 89.515 101.895 ;
        RECT 90.900 101.355 91.200 101.835 ;
        RECT 91.370 101.550 91.630 102.005 ;
        RECT 91.800 101.355 92.060 101.835 ;
        RECT 92.230 101.550 92.490 102.005 ;
        RECT 92.660 101.355 92.920 101.835 ;
        RECT 93.090 101.550 93.350 102.005 ;
        RECT 93.520 101.355 93.780 101.835 ;
        RECT 93.950 101.550 94.210 102.005 ;
        RECT 94.380 101.355 94.640 101.880 ;
        RECT 94.810 101.535 95.060 102.345 ;
        RECT 95.230 101.985 95.545 102.595 ;
        RECT 95.750 102.095 96.065 103.115 ;
        RECT 96.455 103.105 96.785 103.905 ;
        RECT 97.270 102.935 97.660 103.110 ;
        RECT 96.235 102.765 97.660 102.935 ;
        RECT 98.015 102.815 101.525 103.905 ;
        RECT 96.235 102.265 96.405 102.765 ;
        RECT 95.240 101.355 95.485 101.815 ;
        RECT 95.750 101.525 96.365 102.095 ;
        RECT 96.655 102.035 96.920 102.595 ;
        RECT 97.090 101.865 97.260 102.765 ;
        RECT 97.430 102.035 97.785 102.595 ;
        RECT 98.015 102.125 99.665 102.645 ;
        RECT 99.835 102.295 101.525 102.815 ;
        RECT 101.730 103.115 102.265 103.735 ;
        RECT 96.535 101.355 96.750 101.865 ;
        RECT 96.980 101.535 97.260 101.865 ;
        RECT 97.440 101.355 97.680 101.865 ;
        RECT 98.015 101.355 101.525 102.125 ;
        RECT 101.730 102.095 102.045 103.115 ;
        RECT 102.435 103.105 102.765 103.905 ;
        RECT 103.250 102.935 103.640 103.110 ;
        RECT 102.215 102.765 103.640 102.935 ;
        RECT 104.200 102.935 104.530 103.735 ;
        RECT 104.700 103.105 105.030 103.905 ;
        RECT 105.330 102.935 105.660 103.735 ;
        RECT 106.305 103.105 106.555 103.905 ;
        RECT 104.200 102.765 106.635 102.935 ;
        RECT 106.825 102.765 106.995 103.905 ;
        RECT 107.165 102.765 107.505 103.735 ;
        RECT 102.215 102.265 102.385 102.765 ;
        RECT 101.730 101.525 102.345 102.095 ;
        RECT 102.635 102.035 102.900 102.595 ;
        RECT 103.070 101.865 103.240 102.765 ;
        RECT 103.410 102.035 103.765 102.595 ;
        RECT 103.995 102.345 104.345 102.595 ;
        RECT 104.530 102.135 104.700 102.765 ;
        RECT 104.870 102.345 105.200 102.545 ;
        RECT 105.370 102.345 105.700 102.545 ;
        RECT 105.870 102.345 106.290 102.545 ;
        RECT 106.465 102.515 106.635 102.765 ;
        RECT 106.465 102.345 107.160 102.515 ;
        RECT 107.330 102.205 107.505 102.765 ;
        RECT 107.675 102.740 107.965 103.905 ;
        RECT 108.225 103.235 108.395 103.735 ;
        RECT 108.565 103.405 108.895 103.905 ;
        RECT 108.225 103.065 108.890 103.235 ;
        RECT 108.140 102.245 108.490 102.895 ;
        RECT 102.515 101.355 102.730 101.865 ;
        RECT 102.960 101.535 103.240 101.865 ;
        RECT 103.420 101.355 103.660 101.865 ;
        RECT 104.200 101.525 104.700 102.135 ;
        RECT 105.330 102.005 106.555 102.175 ;
        RECT 107.275 102.155 107.505 102.205 ;
        RECT 105.330 101.525 105.660 102.005 ;
        RECT 105.830 101.355 106.055 101.815 ;
        RECT 106.225 101.525 106.555 102.005 ;
        RECT 106.745 101.355 106.995 102.155 ;
        RECT 107.165 101.525 107.505 102.155 ;
        RECT 107.675 101.355 107.965 102.080 ;
        RECT 108.660 102.075 108.890 103.065 ;
        RECT 108.225 101.905 108.890 102.075 ;
        RECT 108.225 101.615 108.395 101.905 ;
        RECT 108.565 101.355 108.895 101.735 ;
        RECT 109.065 101.615 109.250 103.735 ;
        RECT 109.490 103.445 109.755 103.905 ;
        RECT 109.925 103.310 110.175 103.735 ;
        RECT 110.385 103.460 111.490 103.630 ;
        RECT 109.870 103.180 110.175 103.310 ;
        RECT 109.420 101.985 109.700 102.935 ;
        RECT 109.870 102.075 110.040 103.180 ;
        RECT 110.210 102.395 110.450 102.990 ;
        RECT 110.620 102.925 111.150 103.290 ;
        RECT 110.620 102.225 110.790 102.925 ;
        RECT 111.320 102.845 111.490 103.460 ;
        RECT 111.660 103.105 111.830 103.905 ;
        RECT 112.000 103.405 112.250 103.735 ;
        RECT 112.475 103.435 113.360 103.605 ;
        RECT 111.320 102.755 111.830 102.845 ;
        RECT 109.870 101.945 110.095 102.075 ;
        RECT 110.265 102.005 110.790 102.225 ;
        RECT 110.960 102.585 111.830 102.755 ;
        RECT 109.505 101.355 109.755 101.815 ;
        RECT 109.925 101.805 110.095 101.945 ;
        RECT 110.960 101.805 111.130 102.585 ;
        RECT 111.660 102.515 111.830 102.585 ;
        RECT 111.340 102.335 111.540 102.365 ;
        RECT 112.000 102.335 112.170 103.405 ;
        RECT 112.340 102.515 112.530 103.235 ;
        RECT 111.340 102.035 112.170 102.335 ;
        RECT 112.700 102.305 113.020 103.265 ;
        RECT 109.925 101.635 110.260 101.805 ;
        RECT 110.455 101.635 111.130 101.805 ;
        RECT 111.450 101.355 111.820 101.855 ;
        RECT 112.000 101.805 112.170 102.035 ;
        RECT 112.555 101.975 113.020 102.305 ;
        RECT 113.190 102.595 113.360 103.435 ;
        RECT 113.540 103.405 113.855 103.905 ;
        RECT 114.085 103.175 114.425 103.735 ;
        RECT 113.530 102.800 114.425 103.175 ;
        RECT 114.595 102.895 114.765 103.905 ;
        RECT 114.235 102.595 114.425 102.800 ;
        RECT 114.935 102.845 115.265 103.690 ;
        RECT 115.700 102.935 116.030 103.735 ;
        RECT 116.200 103.105 116.530 103.905 ;
        RECT 116.830 102.935 117.160 103.735 ;
        RECT 117.805 103.105 118.055 103.905 ;
        RECT 114.935 102.765 115.325 102.845 ;
        RECT 115.700 102.765 118.135 102.935 ;
        RECT 118.325 102.765 118.495 103.905 ;
        RECT 118.665 102.765 119.005 103.735 ;
        RECT 119.175 102.815 122.685 103.905 ;
        RECT 123.055 103.235 123.335 103.905 ;
        RECT 123.505 103.015 123.805 103.565 ;
        RECT 124.005 103.185 124.335 103.905 ;
        RECT 124.525 103.185 124.985 103.735 ;
        RECT 115.110 102.715 115.325 102.765 ;
        RECT 113.190 102.265 114.065 102.595 ;
        RECT 114.235 102.265 114.985 102.595 ;
        RECT 113.190 101.805 113.360 102.265 ;
        RECT 114.235 102.095 114.435 102.265 ;
        RECT 115.155 102.135 115.325 102.715 ;
        RECT 115.495 102.345 115.845 102.595 ;
        RECT 116.030 102.135 116.200 102.765 ;
        RECT 116.370 102.345 116.700 102.545 ;
        RECT 116.870 102.345 117.200 102.545 ;
        RECT 117.370 102.345 117.790 102.545 ;
        RECT 117.965 102.515 118.135 102.765 ;
        RECT 117.965 102.345 118.660 102.515 ;
        RECT 115.100 102.095 115.325 102.135 ;
        RECT 112.000 101.635 112.405 101.805 ;
        RECT 112.575 101.635 113.360 101.805 ;
        RECT 113.635 101.355 113.845 101.885 ;
        RECT 114.105 101.570 114.435 102.095 ;
        RECT 114.945 102.010 115.325 102.095 ;
        RECT 114.605 101.355 114.775 101.965 ;
        RECT 114.945 101.575 115.275 102.010 ;
        RECT 115.700 101.525 116.200 102.135 ;
        RECT 116.830 102.005 118.055 102.175 ;
        RECT 118.830 102.155 119.005 102.765 ;
        RECT 116.830 101.525 117.160 102.005 ;
        RECT 117.330 101.355 117.555 101.815 ;
        RECT 117.725 101.525 118.055 102.005 ;
        RECT 118.245 101.355 118.495 102.155 ;
        RECT 118.665 101.525 119.005 102.155 ;
        RECT 119.175 102.125 120.825 102.645 ;
        RECT 120.995 102.295 122.685 102.815 ;
        RECT 122.870 102.595 123.135 102.955 ;
        RECT 123.505 102.845 124.445 103.015 ;
        RECT 124.275 102.595 124.445 102.845 ;
        RECT 122.870 102.345 123.545 102.595 ;
        RECT 123.765 102.345 124.105 102.595 ;
        RECT 124.275 102.265 124.565 102.595 ;
        RECT 124.275 102.175 124.445 102.265 ;
        RECT 119.175 101.355 122.685 102.125 ;
        RECT 123.055 101.985 124.445 102.175 ;
        RECT 123.055 101.625 123.385 101.985 ;
        RECT 124.735 101.815 124.985 103.185 ;
        RECT 124.005 101.355 124.255 101.815 ;
        RECT 124.425 101.525 124.985 101.815 ;
        RECT 125.190 103.115 125.725 103.735 ;
        RECT 125.190 102.095 125.505 103.115 ;
        RECT 125.895 103.105 126.225 103.905 ;
        RECT 126.710 102.935 127.100 103.110 ;
        RECT 125.675 102.765 127.100 102.935 ;
        RECT 127.455 102.815 129.125 103.905 ;
        RECT 125.675 102.265 125.845 102.765 ;
        RECT 125.190 101.525 125.805 102.095 ;
        RECT 126.095 102.035 126.360 102.595 ;
        RECT 126.530 101.865 126.700 102.765 ;
        RECT 126.870 102.035 127.225 102.595 ;
        RECT 127.455 102.125 128.205 102.645 ;
        RECT 128.375 102.295 129.125 102.815 ;
        RECT 129.330 103.115 129.865 103.735 ;
        RECT 125.975 101.355 126.190 101.865 ;
        RECT 126.420 101.535 126.700 101.865 ;
        RECT 126.880 101.355 127.120 101.865 ;
        RECT 127.455 101.355 129.125 102.125 ;
        RECT 129.330 102.095 129.645 103.115 ;
        RECT 130.035 103.105 130.365 103.905 ;
        RECT 130.850 102.935 131.240 103.110 ;
        RECT 129.815 102.765 131.240 102.935 ;
        RECT 131.595 102.815 133.265 103.905 ;
        RECT 129.815 102.265 129.985 102.765 ;
        RECT 129.330 101.525 129.945 102.095 ;
        RECT 130.235 102.035 130.500 102.595 ;
        RECT 130.670 101.865 130.840 102.765 ;
        RECT 131.010 102.035 131.365 102.595 ;
        RECT 131.595 102.125 132.345 102.645 ;
        RECT 132.515 102.295 133.265 102.815 ;
        RECT 133.435 102.740 133.725 103.905 ;
        RECT 133.895 103.055 134.155 103.735 ;
        RECT 134.325 103.125 134.575 103.905 ;
        RECT 134.825 103.355 135.075 103.735 ;
        RECT 135.245 103.525 135.600 103.905 ;
        RECT 136.605 103.515 136.940 103.735 ;
        RECT 136.205 103.355 136.435 103.395 ;
        RECT 134.825 103.155 136.435 103.355 ;
        RECT 134.825 103.145 135.660 103.155 ;
        RECT 136.250 103.065 136.435 103.155 ;
        RECT 130.115 101.355 130.330 101.865 ;
        RECT 130.560 101.535 130.840 101.865 ;
        RECT 131.020 101.355 131.260 101.865 ;
        RECT 131.595 101.355 133.265 102.125 ;
        RECT 133.435 101.355 133.725 102.080 ;
        RECT 133.895 101.865 134.065 103.055 ;
        RECT 135.765 102.955 136.095 102.985 ;
        RECT 134.295 102.895 136.095 102.955 ;
        RECT 136.685 102.895 136.940 103.515 ;
        RECT 134.235 102.785 136.940 102.895 ;
        RECT 138.125 102.975 138.295 103.735 ;
        RECT 138.510 103.145 138.840 103.905 ;
        RECT 138.125 102.805 138.840 102.975 ;
        RECT 139.010 102.830 139.265 103.735 ;
        RECT 134.235 102.750 134.435 102.785 ;
        RECT 134.235 102.175 134.405 102.750 ;
        RECT 135.765 102.725 136.940 102.785 ;
        RECT 134.635 102.310 135.045 102.615 ;
        RECT 135.215 102.345 135.545 102.555 ;
        RECT 134.235 102.055 134.505 102.175 ;
        RECT 134.235 102.010 135.080 102.055 ;
        RECT 134.325 101.885 135.080 102.010 ;
        RECT 135.335 101.945 135.545 102.345 ;
        RECT 135.790 102.345 136.265 102.555 ;
        RECT 136.455 102.345 136.945 102.545 ;
        RECT 135.790 101.945 136.010 102.345 ;
        RECT 138.035 102.255 138.390 102.625 ;
        RECT 138.670 102.595 138.840 102.805 ;
        RECT 138.670 102.265 138.925 102.595 ;
        RECT 133.895 101.855 134.125 101.865 ;
        RECT 133.895 101.525 134.155 101.855 ;
        RECT 134.910 101.735 135.080 101.885 ;
        RECT 134.325 101.355 134.655 101.715 ;
        RECT 134.910 101.525 136.210 101.735 ;
        RECT 136.485 101.355 136.940 102.120 ;
        RECT 138.670 102.075 138.840 102.265 ;
        RECT 139.095 102.100 139.265 102.830 ;
        RECT 139.440 102.755 139.700 103.905 ;
        RECT 139.965 102.975 140.135 103.735 ;
        RECT 140.350 103.145 140.680 103.905 ;
        RECT 139.965 102.805 140.680 102.975 ;
        RECT 140.850 102.830 141.105 103.735 ;
        RECT 139.875 102.255 140.230 102.625 ;
        RECT 140.510 102.595 140.680 102.805 ;
        RECT 140.510 102.265 140.765 102.595 ;
        RECT 138.125 101.905 138.840 102.075 ;
        RECT 138.125 101.525 138.295 101.905 ;
        RECT 138.510 101.355 138.840 101.735 ;
        RECT 139.010 101.525 139.265 102.100 ;
        RECT 139.440 101.355 139.700 102.195 ;
        RECT 140.510 102.075 140.680 102.265 ;
        RECT 140.935 102.100 141.105 102.830 ;
        RECT 141.280 102.755 141.540 103.905 ;
        RECT 141.715 102.815 142.925 103.905 ;
        RECT 141.715 102.275 142.235 102.815 ;
        RECT 139.965 101.905 140.680 102.075 ;
        RECT 139.965 101.525 140.135 101.905 ;
        RECT 140.350 101.355 140.680 101.735 ;
        RECT 140.850 101.525 141.105 102.100 ;
        RECT 141.280 101.355 141.540 102.195 ;
        RECT 142.405 102.105 142.925 102.645 ;
        RECT 141.715 101.355 142.925 102.105 ;
        RECT 17.430 101.185 143.010 101.355 ;
        RECT 17.515 100.435 18.725 101.185 ;
        RECT 17.515 99.895 18.035 100.435 ;
        RECT 18.895 100.415 21.485 101.185 ;
        RECT 21.660 100.695 21.915 101.185 ;
        RECT 22.085 100.675 23.315 101.015 ;
        RECT 18.205 99.725 18.725 100.265 ;
        RECT 18.895 99.895 20.105 100.415 ;
        RECT 20.275 99.725 21.485 100.245 ;
        RECT 21.680 99.945 21.900 100.525 ;
        RECT 22.085 99.775 22.265 100.675 ;
        RECT 22.435 99.945 22.810 100.505 ;
        RECT 22.985 100.445 23.315 100.675 ;
        RECT 23.495 100.535 23.755 101.015 ;
        RECT 23.925 100.645 24.175 101.185 ;
        RECT 23.015 99.945 23.325 100.275 ;
        RECT 17.515 98.635 18.725 99.725 ;
        RECT 18.895 98.635 21.485 99.725 ;
        RECT 21.660 98.635 21.915 99.775 ;
        RECT 22.085 99.605 23.315 99.775 ;
        RECT 22.085 98.805 22.415 99.605 ;
        RECT 22.585 98.635 22.815 99.435 ;
        RECT 22.985 98.805 23.315 99.605 ;
        RECT 23.495 99.505 23.665 100.535 ;
        RECT 24.345 100.505 24.565 100.965 ;
        RECT 24.315 100.480 24.565 100.505 ;
        RECT 23.835 99.885 24.065 100.280 ;
        RECT 24.235 100.055 24.565 100.480 ;
        RECT 24.735 100.805 25.625 100.975 ;
        RECT 24.735 100.080 24.905 100.805 ;
        RECT 25.075 100.250 25.625 100.635 ;
        RECT 25.805 100.460 26.135 100.970 ;
        RECT 26.305 100.785 26.635 101.185 ;
        RECT 27.685 100.615 28.015 100.955 ;
        RECT 28.185 100.785 28.515 101.185 ;
        RECT 24.735 100.010 25.625 100.080 ;
        RECT 24.730 99.985 25.625 100.010 ;
        RECT 24.720 99.970 25.625 99.985 ;
        RECT 24.715 99.955 25.625 99.970 ;
        RECT 24.705 99.950 25.625 99.955 ;
        RECT 24.700 99.940 25.625 99.950 ;
        RECT 24.695 99.930 25.625 99.940 ;
        RECT 24.685 99.925 25.625 99.930 ;
        RECT 24.675 99.915 25.625 99.925 ;
        RECT 24.665 99.910 25.625 99.915 ;
        RECT 24.665 99.905 25.000 99.910 ;
        RECT 24.650 99.900 25.000 99.905 ;
        RECT 24.635 99.890 25.000 99.900 ;
        RECT 24.610 99.885 25.000 99.890 ;
        RECT 23.835 99.880 25.000 99.885 ;
        RECT 23.835 99.845 24.970 99.880 ;
        RECT 23.835 99.820 24.935 99.845 ;
        RECT 23.835 99.790 24.905 99.820 ;
        RECT 23.835 99.760 24.885 99.790 ;
        RECT 23.835 99.730 24.865 99.760 ;
        RECT 23.835 99.720 24.795 99.730 ;
        RECT 23.835 99.710 24.770 99.720 ;
        RECT 23.835 99.695 24.750 99.710 ;
        RECT 23.835 99.680 24.730 99.695 ;
        RECT 23.940 99.670 24.725 99.680 ;
        RECT 23.940 99.635 24.710 99.670 ;
        RECT 23.495 98.805 23.770 99.505 ;
        RECT 23.940 99.385 24.695 99.635 ;
        RECT 24.865 99.315 25.195 99.560 ;
        RECT 25.365 99.460 25.625 99.910 ;
        RECT 25.805 99.695 25.995 100.460 ;
        RECT 26.305 100.445 28.670 100.615 ;
        RECT 29.035 100.455 29.325 101.185 ;
        RECT 26.305 100.275 26.475 100.445 ;
        RECT 26.165 99.945 26.475 100.275 ;
        RECT 26.645 99.945 26.950 100.275 ;
        RECT 25.010 99.290 25.195 99.315 ;
        RECT 25.010 99.190 25.625 99.290 ;
        RECT 23.940 98.635 24.195 99.180 ;
        RECT 24.365 98.805 24.845 99.145 ;
        RECT 25.020 98.635 25.625 99.190 ;
        RECT 25.805 98.845 26.135 99.695 ;
        RECT 26.305 98.635 26.555 99.775 ;
        RECT 26.735 99.615 26.950 99.945 ;
        RECT 27.125 99.615 27.410 100.275 ;
        RECT 27.605 99.615 27.870 100.275 ;
        RECT 28.085 99.615 28.330 100.275 ;
        RECT 28.500 99.445 28.670 100.445 ;
        RECT 29.025 99.945 29.325 100.275 ;
        RECT 29.505 100.255 29.735 100.895 ;
        RECT 29.915 100.635 30.225 101.005 ;
        RECT 30.405 100.815 31.075 101.185 ;
        RECT 29.915 100.435 31.145 100.635 ;
        RECT 29.505 99.945 30.030 100.255 ;
        RECT 30.210 99.945 30.675 100.255 ;
        RECT 30.855 99.765 31.145 100.435 ;
        RECT 26.745 99.275 28.035 99.445 ;
        RECT 26.745 98.855 26.995 99.275 ;
        RECT 27.225 98.635 27.555 99.105 ;
        RECT 27.785 98.855 28.035 99.275 ;
        RECT 28.215 99.275 28.670 99.445 ;
        RECT 29.035 99.525 30.195 99.765 ;
        RECT 28.215 98.845 28.545 99.275 ;
        RECT 29.035 98.815 29.295 99.525 ;
        RECT 29.465 98.635 29.795 99.345 ;
        RECT 29.965 98.815 30.195 99.525 ;
        RECT 30.375 99.545 31.145 99.765 ;
        RECT 30.375 98.815 30.645 99.545 ;
        RECT 30.825 98.635 31.165 99.365 ;
        RECT 31.335 98.815 31.595 101.005 ;
        RECT 31.775 100.640 37.120 101.185 ;
        RECT 37.755 100.805 38.645 100.975 ;
        RECT 33.360 99.810 33.700 100.640 ;
        RECT 35.180 99.070 35.530 100.320 ;
        RECT 37.755 100.250 38.305 100.635 ;
        RECT 38.475 100.080 38.645 100.805 ;
        RECT 37.755 100.010 38.645 100.080 ;
        RECT 38.815 100.480 39.035 100.965 ;
        RECT 39.205 100.645 39.455 101.185 ;
        RECT 39.625 100.535 39.885 101.015 ;
        RECT 38.815 100.055 39.145 100.480 ;
        RECT 37.755 99.985 38.650 100.010 ;
        RECT 37.755 99.970 38.660 99.985 ;
        RECT 37.755 99.955 38.665 99.970 ;
        RECT 37.755 99.950 38.675 99.955 ;
        RECT 37.755 99.940 38.680 99.950 ;
        RECT 37.755 99.930 38.685 99.940 ;
        RECT 37.755 99.925 38.695 99.930 ;
        RECT 37.755 99.915 38.705 99.925 ;
        RECT 37.755 99.910 38.715 99.915 ;
        RECT 37.755 99.460 38.015 99.910 ;
        RECT 38.380 99.905 38.715 99.910 ;
        RECT 38.380 99.900 38.730 99.905 ;
        RECT 38.380 99.890 38.745 99.900 ;
        RECT 38.380 99.885 38.770 99.890 ;
        RECT 39.315 99.885 39.545 100.280 ;
        RECT 38.380 99.880 39.545 99.885 ;
        RECT 38.410 99.845 39.545 99.880 ;
        RECT 38.445 99.820 39.545 99.845 ;
        RECT 38.475 99.790 39.545 99.820 ;
        RECT 38.495 99.760 39.545 99.790 ;
        RECT 38.515 99.730 39.545 99.760 ;
        RECT 38.585 99.720 39.545 99.730 ;
        RECT 38.610 99.710 39.545 99.720 ;
        RECT 38.630 99.695 39.545 99.710 ;
        RECT 38.650 99.680 39.545 99.695 ;
        RECT 38.655 99.670 39.440 99.680 ;
        RECT 38.670 99.635 39.440 99.670 ;
        RECT 38.185 99.315 38.515 99.560 ;
        RECT 38.685 99.385 39.440 99.635 ;
        RECT 39.715 99.505 39.885 100.535 ;
        RECT 38.185 99.290 38.370 99.315 ;
        RECT 37.755 99.190 38.370 99.290 ;
        RECT 31.775 98.635 37.120 99.070 ;
        RECT 37.755 98.635 38.360 99.190 ;
        RECT 38.535 98.805 39.015 99.145 ;
        RECT 39.185 98.635 39.440 99.180 ;
        RECT 39.610 98.805 39.885 99.505 ;
        RECT 40.065 98.815 40.325 101.005 ;
        RECT 40.585 100.815 41.255 101.185 ;
        RECT 41.435 100.635 41.745 101.005 ;
        RECT 40.515 100.435 41.745 100.635 ;
        RECT 40.515 99.765 40.805 100.435 ;
        RECT 41.925 100.255 42.155 100.895 ;
        RECT 42.335 100.455 42.625 101.185 ;
        RECT 43.275 100.460 43.565 101.185 ;
        RECT 43.735 100.385 44.430 101.015 ;
        RECT 44.635 100.385 44.945 101.185 ;
        RECT 45.115 100.415 47.705 101.185 ;
        RECT 48.535 100.555 48.865 100.915 ;
        RECT 49.485 100.725 49.735 101.185 ;
        RECT 49.905 100.725 50.465 101.015 ;
        RECT 40.985 99.945 41.450 100.255 ;
        RECT 41.630 99.945 42.155 100.255 ;
        RECT 42.335 99.945 42.635 100.275 ;
        RECT 43.755 99.945 44.090 100.195 ;
        RECT 40.515 99.545 41.285 99.765 ;
        RECT 40.495 98.635 40.835 99.365 ;
        RECT 41.015 98.815 41.285 99.545 ;
        RECT 41.465 99.525 42.625 99.765 ;
        RECT 41.465 98.815 41.695 99.525 ;
        RECT 41.865 98.635 42.195 99.345 ;
        RECT 42.365 98.815 42.625 99.525 ;
        RECT 43.275 98.635 43.565 99.800 ;
        RECT 44.260 99.785 44.430 100.385 ;
        RECT 44.600 99.945 44.935 100.215 ;
        RECT 45.115 99.895 46.325 100.415 ;
        RECT 48.535 100.365 49.925 100.555 ;
        RECT 49.755 100.275 49.925 100.365 ;
        RECT 43.735 98.635 43.995 99.775 ;
        RECT 44.165 98.805 44.495 99.785 ;
        RECT 44.665 98.635 44.945 99.775 ;
        RECT 46.495 99.725 47.705 100.245 ;
        RECT 45.115 98.635 47.705 99.725 ;
        RECT 48.350 99.945 49.025 100.195 ;
        RECT 49.245 99.945 49.585 100.195 ;
        RECT 49.755 99.945 50.045 100.275 ;
        RECT 48.350 99.585 48.615 99.945 ;
        RECT 49.755 99.695 49.925 99.945 ;
        RECT 48.985 99.525 49.925 99.695 ;
        RECT 48.535 98.635 48.815 99.305 ;
        RECT 48.985 98.975 49.285 99.525 ;
        RECT 50.215 99.355 50.465 100.725 ;
        RECT 50.915 100.555 51.295 101.005 ;
        RECT 50.655 99.605 50.885 100.295 ;
        RECT 51.065 100.105 51.295 100.555 ;
        RECT 51.475 100.405 51.705 101.185 ;
        RECT 51.885 100.475 52.315 101.005 ;
        RECT 51.885 100.225 52.130 100.475 ;
        RECT 52.495 100.275 52.705 100.895 ;
        RECT 52.875 100.455 53.205 101.185 ;
        RECT 53.510 100.555 53.795 101.015 ;
        RECT 53.965 100.725 54.235 101.185 ;
        RECT 53.510 100.385 54.465 100.555 ;
        RECT 51.065 99.425 51.405 100.105 ;
        RECT 49.485 98.635 49.815 99.355 ;
        RECT 50.005 98.805 50.465 99.355 ;
        RECT 50.645 99.225 51.405 99.425 ;
        RECT 51.595 99.925 52.130 100.225 ;
        RECT 52.310 99.925 52.705 100.275 ;
        RECT 52.900 99.925 53.190 100.275 ;
        RECT 50.645 98.835 50.905 99.225 ;
        RECT 51.075 98.635 51.405 99.045 ;
        RECT 51.595 98.815 51.925 99.925 ;
        RECT 52.095 99.545 53.135 99.745 ;
        RECT 53.395 99.655 54.085 100.215 ;
        RECT 52.095 98.815 52.285 99.545 ;
        RECT 52.455 98.635 52.785 99.365 ;
        RECT 52.965 98.815 53.135 99.545 ;
        RECT 54.255 99.485 54.465 100.385 ;
        RECT 53.510 99.265 54.465 99.485 ;
        RECT 54.635 100.215 55.035 101.015 ;
        RECT 55.225 100.555 55.505 101.015 ;
        RECT 56.025 100.725 56.350 101.185 ;
        RECT 55.225 100.385 56.350 100.555 ;
        RECT 56.520 100.445 56.905 101.015 ;
        RECT 57.240 100.675 57.480 101.185 ;
        RECT 57.660 100.675 57.940 101.005 ;
        RECT 58.170 100.675 58.385 101.185 ;
        RECT 55.900 100.275 56.350 100.385 ;
        RECT 54.635 99.655 55.730 100.215 ;
        RECT 55.900 99.945 56.455 100.275 ;
        RECT 53.510 98.805 53.795 99.265 ;
        RECT 53.965 98.635 54.235 99.095 ;
        RECT 54.635 98.805 55.035 99.655 ;
        RECT 55.900 99.485 56.350 99.945 ;
        RECT 56.625 99.775 56.905 100.445 ;
        RECT 57.135 99.945 57.490 100.505 ;
        RECT 57.660 99.775 57.830 100.675 ;
        RECT 58.000 99.945 58.265 100.505 ;
        RECT 58.555 100.445 59.170 101.015 ;
        RECT 58.515 99.775 58.685 100.275 ;
        RECT 55.225 99.265 56.350 99.485 ;
        RECT 55.225 98.805 55.505 99.265 ;
        RECT 56.025 98.635 56.350 99.095 ;
        RECT 56.520 98.805 56.905 99.775 ;
        RECT 57.260 99.605 58.685 99.775 ;
        RECT 57.260 99.430 57.650 99.605 ;
        RECT 58.135 98.635 58.465 99.435 ;
        RECT 58.855 99.425 59.170 100.445 ;
        RECT 58.635 98.805 59.170 99.425 ;
        RECT 59.375 100.535 59.635 101.015 ;
        RECT 59.805 100.645 60.055 101.185 ;
        RECT 59.375 99.505 59.545 100.535 ;
        RECT 60.225 100.505 60.445 100.965 ;
        RECT 60.195 100.480 60.445 100.505 ;
        RECT 59.715 99.885 59.945 100.280 ;
        RECT 60.115 100.055 60.445 100.480 ;
        RECT 60.615 100.805 61.505 100.975 ;
        RECT 60.615 100.080 60.785 100.805 ;
        RECT 60.955 100.250 61.505 100.635 ;
        RECT 61.675 100.415 65.185 101.185 ;
        RECT 65.360 100.710 65.695 100.970 ;
        RECT 65.865 100.785 66.195 101.185 ;
        RECT 66.365 100.785 67.980 100.955 ;
        RECT 60.615 100.010 61.505 100.080 ;
        RECT 60.610 99.985 61.505 100.010 ;
        RECT 60.600 99.970 61.505 99.985 ;
        RECT 60.595 99.955 61.505 99.970 ;
        RECT 60.585 99.950 61.505 99.955 ;
        RECT 60.580 99.940 61.505 99.950 ;
        RECT 60.575 99.930 61.505 99.940 ;
        RECT 60.565 99.925 61.505 99.930 ;
        RECT 60.555 99.915 61.505 99.925 ;
        RECT 60.545 99.910 61.505 99.915 ;
        RECT 60.545 99.905 60.880 99.910 ;
        RECT 60.530 99.900 60.880 99.905 ;
        RECT 60.515 99.890 60.880 99.900 ;
        RECT 60.490 99.885 60.880 99.890 ;
        RECT 59.715 99.880 60.880 99.885 ;
        RECT 59.715 99.845 60.850 99.880 ;
        RECT 59.715 99.820 60.815 99.845 ;
        RECT 59.715 99.790 60.785 99.820 ;
        RECT 59.715 99.760 60.765 99.790 ;
        RECT 59.715 99.730 60.745 99.760 ;
        RECT 59.715 99.720 60.675 99.730 ;
        RECT 59.715 99.710 60.650 99.720 ;
        RECT 59.715 99.695 60.630 99.710 ;
        RECT 59.715 99.680 60.610 99.695 ;
        RECT 59.820 99.670 60.605 99.680 ;
        RECT 59.820 99.635 60.590 99.670 ;
        RECT 59.375 98.805 59.650 99.505 ;
        RECT 59.820 99.385 60.575 99.635 ;
        RECT 60.745 99.315 61.075 99.560 ;
        RECT 61.245 99.460 61.505 99.910 ;
        RECT 61.675 99.895 63.325 100.415 ;
        RECT 63.495 99.725 65.185 100.245 ;
        RECT 60.890 99.290 61.075 99.315 ;
        RECT 60.890 99.190 61.505 99.290 ;
        RECT 59.820 98.635 60.075 99.180 ;
        RECT 60.245 98.805 60.725 99.145 ;
        RECT 60.900 98.635 61.505 99.190 ;
        RECT 61.675 98.635 65.185 99.725 ;
        RECT 65.360 99.355 65.615 100.710 ;
        RECT 66.365 100.615 66.535 100.785 ;
        RECT 65.975 100.445 66.535 100.615 ;
        RECT 65.975 100.275 66.145 100.445 ;
        RECT 65.840 99.945 66.145 100.275 ;
        RECT 66.340 100.165 66.590 100.275 ;
        RECT 66.800 100.165 67.070 100.605 ;
        RECT 67.260 100.505 67.550 100.605 ;
        RECT 67.255 100.335 67.550 100.505 ;
        RECT 66.335 99.995 66.590 100.165 ;
        RECT 66.795 99.995 67.070 100.165 ;
        RECT 66.340 99.945 66.590 99.995 ;
        RECT 66.800 99.945 67.070 99.995 ;
        RECT 67.260 99.945 67.550 100.335 ;
        RECT 67.720 99.945 68.140 100.610 ;
        RECT 68.525 100.465 68.855 101.185 ;
        RECT 69.035 100.460 69.325 101.185 ;
        RECT 69.495 100.435 70.705 101.185 ;
        RECT 70.875 100.445 71.260 101.015 ;
        RECT 71.430 100.725 71.755 101.185 ;
        RECT 72.275 100.555 72.555 101.015 ;
        RECT 68.450 99.945 68.800 100.275 ;
        RECT 65.975 99.775 66.145 99.945 ;
        RECT 68.595 99.825 68.800 99.945 ;
        RECT 69.495 99.895 70.015 100.435 ;
        RECT 65.975 99.605 68.345 99.775 ;
        RECT 68.595 99.655 68.805 99.825 ;
        RECT 65.360 98.845 65.695 99.355 ;
        RECT 65.945 98.635 66.275 99.435 ;
        RECT 66.520 99.225 67.945 99.395 ;
        RECT 66.520 98.805 66.805 99.225 ;
        RECT 67.060 98.635 67.390 99.055 ;
        RECT 67.615 98.975 67.945 99.225 ;
        RECT 68.175 99.145 68.345 99.605 ;
        RECT 68.605 98.975 68.775 99.475 ;
        RECT 67.615 98.805 68.775 98.975 ;
        RECT 69.035 98.635 69.325 99.800 ;
        RECT 70.185 99.725 70.705 100.265 ;
        RECT 69.495 98.635 70.705 99.725 ;
        RECT 70.875 99.775 71.155 100.445 ;
        RECT 71.430 100.385 72.555 100.555 ;
        RECT 71.430 100.275 71.880 100.385 ;
        RECT 71.325 99.945 71.880 100.275 ;
        RECT 72.745 100.215 73.145 101.015 ;
        RECT 73.545 100.725 73.815 101.185 ;
        RECT 73.985 100.555 74.270 101.015 ;
        RECT 70.875 98.805 71.260 99.775 ;
        RECT 71.430 99.485 71.880 99.945 ;
        RECT 72.050 99.655 73.145 100.215 ;
        RECT 71.430 99.265 72.555 99.485 ;
        RECT 71.430 98.635 71.755 99.095 ;
        RECT 72.275 98.805 72.555 99.265 ;
        RECT 72.745 98.805 73.145 99.655 ;
        RECT 73.315 100.385 74.270 100.555 ;
        RECT 74.555 100.415 78.065 101.185 ;
        RECT 78.325 100.635 78.495 100.925 ;
        RECT 78.665 100.805 78.995 101.185 ;
        RECT 78.325 100.465 78.990 100.635 ;
        RECT 73.315 99.485 73.525 100.385 ;
        RECT 73.695 99.655 74.385 100.215 ;
        RECT 74.555 99.895 76.205 100.415 ;
        RECT 76.375 99.725 78.065 100.245 ;
        RECT 73.315 99.265 74.270 99.485 ;
        RECT 73.545 98.635 73.815 99.095 ;
        RECT 73.985 98.805 74.270 99.265 ;
        RECT 74.555 98.635 78.065 99.725 ;
        RECT 78.240 99.645 78.590 100.295 ;
        RECT 78.760 99.475 78.990 100.465 ;
        RECT 78.325 99.305 78.990 99.475 ;
        RECT 78.325 98.805 78.495 99.305 ;
        RECT 78.665 98.635 78.995 99.135 ;
        RECT 79.165 98.805 79.350 100.925 ;
        RECT 79.605 100.725 79.855 101.185 ;
        RECT 80.025 100.735 80.360 100.905 ;
        RECT 80.555 100.735 81.230 100.905 ;
        RECT 80.025 100.595 80.195 100.735 ;
        RECT 79.520 99.605 79.800 100.555 ;
        RECT 79.970 100.465 80.195 100.595 ;
        RECT 79.970 99.360 80.140 100.465 ;
        RECT 80.365 100.315 80.890 100.535 ;
        RECT 80.310 99.550 80.550 100.145 ;
        RECT 80.720 99.615 80.890 100.315 ;
        RECT 81.060 99.955 81.230 100.735 ;
        RECT 81.550 100.685 81.920 101.185 ;
        RECT 82.100 100.735 82.505 100.905 ;
        RECT 82.675 100.735 83.460 100.905 ;
        RECT 82.100 100.505 82.270 100.735 ;
        RECT 81.440 100.205 82.270 100.505 ;
        RECT 82.655 100.235 83.120 100.565 ;
        RECT 81.440 100.175 81.640 100.205 ;
        RECT 81.760 99.955 81.930 100.025 ;
        RECT 81.060 99.785 81.930 99.955 ;
        RECT 81.420 99.695 81.930 99.785 ;
        RECT 79.970 99.230 80.275 99.360 ;
        RECT 80.720 99.250 81.250 99.615 ;
        RECT 79.590 98.635 79.855 99.095 ;
        RECT 80.025 98.805 80.275 99.230 ;
        RECT 81.420 99.080 81.590 99.695 ;
        RECT 80.485 98.910 81.590 99.080 ;
        RECT 81.760 98.635 81.930 99.435 ;
        RECT 82.100 99.135 82.270 100.205 ;
        RECT 82.440 99.305 82.630 100.025 ;
        RECT 82.800 99.275 83.120 100.235 ;
        RECT 83.290 100.275 83.460 100.735 ;
        RECT 83.735 100.655 83.945 101.185 ;
        RECT 84.205 100.445 84.535 100.970 ;
        RECT 84.705 100.575 84.875 101.185 ;
        RECT 85.045 100.530 85.375 100.965 ;
        RECT 85.045 100.445 85.425 100.530 ;
        RECT 84.335 100.275 84.535 100.445 ;
        RECT 85.200 100.405 85.425 100.445 ;
        RECT 83.290 99.945 84.165 100.275 ;
        RECT 84.335 99.945 85.085 100.275 ;
        RECT 82.100 98.805 82.350 99.135 ;
        RECT 83.290 99.105 83.460 99.945 ;
        RECT 84.335 99.740 84.525 99.945 ;
        RECT 85.255 99.825 85.425 100.405 ;
        RECT 85.595 100.415 89.105 101.185 ;
        RECT 85.595 99.895 87.245 100.415 ;
        RECT 89.735 100.385 90.075 101.015 ;
        RECT 90.245 100.385 90.495 101.185 ;
        RECT 90.685 100.535 91.015 101.015 ;
        RECT 91.185 100.725 91.410 101.185 ;
        RECT 91.580 100.535 91.910 101.015 ;
        RECT 85.210 99.775 85.425 99.825 ;
        RECT 83.630 99.365 84.525 99.740 ;
        RECT 85.035 99.695 85.425 99.775 ;
        RECT 87.415 99.725 89.105 100.245 ;
        RECT 82.575 98.935 83.460 99.105 ;
        RECT 83.640 98.635 83.955 99.135 ;
        RECT 84.185 98.805 84.525 99.365 ;
        RECT 84.695 98.635 84.865 99.645 ;
        RECT 85.035 98.850 85.365 99.695 ;
        RECT 85.595 98.635 89.105 99.725 ;
        RECT 89.735 99.775 89.910 100.385 ;
        RECT 90.685 100.365 91.910 100.535 ;
        RECT 92.540 100.405 93.040 101.015 ;
        RECT 93.415 100.435 94.625 101.185 ;
        RECT 94.795 100.460 95.085 101.185 ;
        RECT 95.255 100.685 95.515 101.015 ;
        RECT 95.685 100.825 96.015 101.185 ;
        RECT 96.270 100.805 97.570 101.015 ;
        RECT 95.255 100.675 95.485 100.685 ;
        RECT 90.080 100.025 90.775 100.195 ;
        RECT 90.605 99.775 90.775 100.025 ;
        RECT 90.950 99.995 91.370 100.195 ;
        RECT 91.540 99.995 91.870 100.195 ;
        RECT 92.040 99.995 92.370 100.195 ;
        RECT 92.540 99.775 92.710 100.405 ;
        RECT 92.895 99.945 93.245 100.195 ;
        RECT 93.415 99.895 93.935 100.435 ;
        RECT 89.735 98.805 90.075 99.775 ;
        RECT 90.245 98.635 90.415 99.775 ;
        RECT 90.605 99.605 93.040 99.775 ;
        RECT 94.105 99.725 94.625 100.265 ;
        RECT 90.685 98.635 90.935 99.435 ;
        RECT 91.580 98.805 91.910 99.605 ;
        RECT 92.210 98.635 92.540 99.435 ;
        RECT 92.710 98.805 93.040 99.605 ;
        RECT 93.415 98.635 94.625 99.725 ;
        RECT 94.795 98.635 95.085 99.800 ;
        RECT 95.255 99.485 95.425 100.675 ;
        RECT 96.270 100.655 96.440 100.805 ;
        RECT 95.685 100.530 96.440 100.655 ;
        RECT 95.595 100.485 96.440 100.530 ;
        RECT 95.595 100.365 95.865 100.485 ;
        RECT 95.595 99.790 95.765 100.365 ;
        RECT 95.995 99.925 96.405 100.230 ;
        RECT 96.695 100.195 96.905 100.595 ;
        RECT 96.575 99.985 96.905 100.195 ;
        RECT 97.150 100.195 97.370 100.595 ;
        RECT 97.845 100.420 98.300 101.185 ;
        RECT 98.475 100.640 103.820 101.185 ;
        RECT 97.150 99.985 97.625 100.195 ;
        RECT 97.815 99.995 98.305 100.195 ;
        RECT 95.595 99.755 95.795 99.790 ;
        RECT 97.125 99.755 98.300 99.815 ;
        RECT 100.060 99.810 100.400 100.640 ;
        RECT 103.995 100.415 106.585 101.185 ;
        RECT 107.305 100.635 107.475 100.925 ;
        RECT 107.645 100.805 107.975 101.185 ;
        RECT 107.305 100.465 107.970 100.635 ;
        RECT 95.595 99.645 98.300 99.755 ;
        RECT 95.655 99.585 97.455 99.645 ;
        RECT 97.125 99.555 97.455 99.585 ;
        RECT 95.255 98.805 95.515 99.485 ;
        RECT 95.685 98.635 95.935 99.415 ;
        RECT 96.185 99.385 97.020 99.395 ;
        RECT 97.610 99.385 97.795 99.475 ;
        RECT 96.185 99.185 97.795 99.385 ;
        RECT 96.185 98.805 96.435 99.185 ;
        RECT 97.565 99.145 97.795 99.185 ;
        RECT 98.045 99.025 98.300 99.645 ;
        RECT 101.880 99.070 102.230 100.320 ;
        RECT 103.995 99.895 105.205 100.415 ;
        RECT 105.375 99.725 106.585 100.245 ;
        RECT 96.605 98.635 96.960 99.015 ;
        RECT 97.965 98.805 98.300 99.025 ;
        RECT 98.475 98.635 103.820 99.070 ;
        RECT 103.995 98.635 106.585 99.725 ;
        RECT 107.220 99.645 107.570 100.295 ;
        RECT 107.740 99.475 107.970 100.465 ;
        RECT 107.305 99.305 107.970 99.475 ;
        RECT 107.305 98.805 107.475 99.305 ;
        RECT 107.645 98.635 107.975 99.135 ;
        RECT 108.145 98.805 108.330 100.925 ;
        RECT 108.585 100.725 108.835 101.185 ;
        RECT 109.005 100.735 109.340 100.905 ;
        RECT 109.535 100.735 110.210 100.905 ;
        RECT 109.005 100.595 109.175 100.735 ;
        RECT 108.500 99.605 108.780 100.555 ;
        RECT 108.950 100.465 109.175 100.595 ;
        RECT 108.950 99.360 109.120 100.465 ;
        RECT 109.345 100.315 109.870 100.535 ;
        RECT 109.290 99.550 109.530 100.145 ;
        RECT 109.700 99.615 109.870 100.315 ;
        RECT 110.040 99.955 110.210 100.735 ;
        RECT 110.530 100.685 110.900 101.185 ;
        RECT 111.080 100.735 111.485 100.905 ;
        RECT 111.655 100.735 112.440 100.905 ;
        RECT 111.080 100.505 111.250 100.735 ;
        RECT 110.420 100.205 111.250 100.505 ;
        RECT 111.635 100.235 112.100 100.565 ;
        RECT 110.420 100.175 110.620 100.205 ;
        RECT 110.740 99.955 110.910 100.025 ;
        RECT 110.040 99.785 110.910 99.955 ;
        RECT 110.400 99.695 110.910 99.785 ;
        RECT 108.950 99.230 109.255 99.360 ;
        RECT 109.700 99.250 110.230 99.615 ;
        RECT 108.570 98.635 108.835 99.095 ;
        RECT 109.005 98.805 109.255 99.230 ;
        RECT 110.400 99.080 110.570 99.695 ;
        RECT 109.465 98.910 110.570 99.080 ;
        RECT 110.740 98.635 110.910 99.435 ;
        RECT 111.080 99.135 111.250 100.205 ;
        RECT 111.420 99.305 111.610 100.025 ;
        RECT 111.780 99.275 112.100 100.235 ;
        RECT 112.270 100.275 112.440 100.735 ;
        RECT 112.715 100.655 112.925 101.185 ;
        RECT 113.185 100.445 113.515 100.970 ;
        RECT 113.685 100.575 113.855 101.185 ;
        RECT 114.025 100.530 114.355 100.965 ;
        RECT 114.025 100.445 114.405 100.530 ;
        RECT 113.315 100.275 113.515 100.445 ;
        RECT 114.180 100.405 114.405 100.445 ;
        RECT 112.270 99.945 113.145 100.275 ;
        RECT 113.315 99.945 114.065 100.275 ;
        RECT 111.080 98.805 111.330 99.135 ;
        RECT 112.270 99.105 112.440 99.945 ;
        RECT 113.315 99.740 113.505 99.945 ;
        RECT 114.235 99.825 114.405 100.405 ;
        RECT 114.575 100.415 117.165 101.185 ;
        RECT 117.995 100.555 118.325 100.915 ;
        RECT 118.945 100.725 119.195 101.185 ;
        RECT 119.365 100.725 119.925 101.015 ;
        RECT 114.575 99.895 115.785 100.415 ;
        RECT 117.995 100.365 119.385 100.555 ;
        RECT 119.215 100.275 119.385 100.365 ;
        RECT 114.190 99.775 114.405 99.825 ;
        RECT 112.610 99.365 113.505 99.740 ;
        RECT 114.015 99.695 114.405 99.775 ;
        RECT 115.955 99.725 117.165 100.245 ;
        RECT 111.555 98.935 112.440 99.105 ;
        RECT 112.620 98.635 112.935 99.135 ;
        RECT 113.165 98.805 113.505 99.365 ;
        RECT 113.675 98.635 113.845 99.645 ;
        RECT 114.015 98.850 114.345 99.695 ;
        RECT 114.575 98.635 117.165 99.725 ;
        RECT 117.810 99.945 118.485 100.195 ;
        RECT 118.705 99.945 119.045 100.195 ;
        RECT 119.215 99.945 119.505 100.275 ;
        RECT 117.810 99.585 118.075 99.945 ;
        RECT 119.215 99.695 119.385 99.945 ;
        RECT 118.445 99.525 119.385 99.695 ;
        RECT 117.995 98.635 118.275 99.305 ;
        RECT 118.445 98.975 118.745 99.525 ;
        RECT 119.675 99.355 119.925 100.725 ;
        RECT 120.555 100.460 120.845 101.185 ;
        RECT 121.015 100.640 126.360 101.185 ;
        RECT 122.600 99.810 122.940 100.640 ;
        RECT 126.740 100.405 127.240 101.015 ;
        RECT 118.945 98.635 119.275 99.355 ;
        RECT 119.465 98.805 119.925 99.355 ;
        RECT 120.555 98.635 120.845 99.800 ;
        RECT 124.420 99.070 124.770 100.320 ;
        RECT 126.535 99.945 126.885 100.195 ;
        RECT 127.070 99.775 127.240 100.405 ;
        RECT 127.870 100.535 128.200 101.015 ;
        RECT 128.370 100.725 128.595 101.185 ;
        RECT 128.765 100.535 129.095 101.015 ;
        RECT 127.870 100.365 129.095 100.535 ;
        RECT 129.285 100.385 129.535 101.185 ;
        RECT 129.705 100.385 130.045 101.015 ;
        RECT 130.305 100.635 130.475 100.925 ;
        RECT 130.645 100.805 130.975 101.185 ;
        RECT 130.305 100.465 130.970 100.635 ;
        RECT 129.815 100.335 130.045 100.385 ;
        RECT 127.410 99.995 127.740 100.195 ;
        RECT 127.910 99.995 128.240 100.195 ;
        RECT 128.410 99.995 128.830 100.195 ;
        RECT 129.005 100.025 129.700 100.195 ;
        RECT 129.005 99.775 129.175 100.025 ;
        RECT 129.870 99.775 130.045 100.335 ;
        RECT 126.740 99.605 129.175 99.775 ;
        RECT 121.015 98.635 126.360 99.070 ;
        RECT 126.740 98.805 127.070 99.605 ;
        RECT 127.240 98.635 127.570 99.435 ;
        RECT 127.870 98.805 128.200 99.605 ;
        RECT 128.845 98.635 129.095 99.435 ;
        RECT 129.365 98.635 129.535 99.775 ;
        RECT 129.705 98.805 130.045 99.775 ;
        RECT 130.220 99.645 130.570 100.295 ;
        RECT 130.740 99.475 130.970 100.465 ;
        RECT 130.305 99.305 130.970 99.475 ;
        RECT 130.305 98.805 130.475 99.305 ;
        RECT 130.645 98.635 130.975 99.135 ;
        RECT 131.145 98.805 131.330 100.925 ;
        RECT 131.585 100.725 131.835 101.185 ;
        RECT 132.005 100.735 132.340 100.905 ;
        RECT 132.535 100.735 133.210 100.905 ;
        RECT 132.005 100.595 132.175 100.735 ;
        RECT 131.500 99.605 131.780 100.555 ;
        RECT 131.950 100.465 132.175 100.595 ;
        RECT 131.950 99.360 132.120 100.465 ;
        RECT 132.345 100.315 132.870 100.535 ;
        RECT 132.290 99.550 132.530 100.145 ;
        RECT 132.700 99.615 132.870 100.315 ;
        RECT 133.040 99.955 133.210 100.735 ;
        RECT 133.530 100.685 133.900 101.185 ;
        RECT 134.080 100.735 134.485 100.905 ;
        RECT 134.655 100.735 135.440 100.905 ;
        RECT 134.080 100.505 134.250 100.735 ;
        RECT 133.420 100.205 134.250 100.505 ;
        RECT 134.635 100.235 135.100 100.565 ;
        RECT 133.420 100.175 133.620 100.205 ;
        RECT 133.740 99.955 133.910 100.025 ;
        RECT 133.040 99.785 133.910 99.955 ;
        RECT 133.400 99.695 133.910 99.785 ;
        RECT 131.950 99.230 132.255 99.360 ;
        RECT 132.700 99.250 133.230 99.615 ;
        RECT 131.570 98.635 131.835 99.095 ;
        RECT 132.005 98.805 132.255 99.230 ;
        RECT 133.400 99.080 133.570 99.695 ;
        RECT 132.465 98.910 133.570 99.080 ;
        RECT 133.740 98.635 133.910 99.435 ;
        RECT 134.080 99.135 134.250 100.205 ;
        RECT 134.420 99.305 134.610 100.025 ;
        RECT 134.780 99.275 135.100 100.235 ;
        RECT 135.270 100.275 135.440 100.735 ;
        RECT 135.715 100.655 135.925 101.185 ;
        RECT 136.185 100.445 136.515 100.970 ;
        RECT 136.685 100.575 136.855 101.185 ;
        RECT 137.025 100.530 137.355 100.965 ;
        RECT 137.575 100.685 137.835 101.015 ;
        RECT 138.005 100.825 138.335 101.185 ;
        RECT 138.590 100.805 139.890 101.015 ;
        RECT 137.025 100.445 137.405 100.530 ;
        RECT 136.315 100.275 136.515 100.445 ;
        RECT 137.180 100.405 137.405 100.445 ;
        RECT 135.270 99.945 136.145 100.275 ;
        RECT 136.315 99.945 137.065 100.275 ;
        RECT 134.080 98.805 134.330 99.135 ;
        RECT 135.270 99.105 135.440 99.945 ;
        RECT 136.315 99.740 136.505 99.945 ;
        RECT 137.235 99.825 137.405 100.405 ;
        RECT 137.190 99.775 137.405 99.825 ;
        RECT 135.610 99.365 136.505 99.740 ;
        RECT 137.015 99.695 137.405 99.775 ;
        RECT 134.555 98.935 135.440 99.105 ;
        RECT 135.620 98.635 135.935 99.135 ;
        RECT 136.165 98.805 136.505 99.365 ;
        RECT 136.675 98.635 136.845 99.645 ;
        RECT 137.015 98.850 137.345 99.695 ;
        RECT 137.575 99.485 137.745 100.685 ;
        RECT 138.590 100.655 138.760 100.805 ;
        RECT 138.005 100.530 138.760 100.655 ;
        RECT 137.915 100.485 138.760 100.530 ;
        RECT 137.915 100.365 138.185 100.485 ;
        RECT 137.915 99.790 138.085 100.365 ;
        RECT 138.315 99.925 138.725 100.230 ;
        RECT 139.015 100.195 139.225 100.595 ;
        RECT 138.895 99.985 139.225 100.195 ;
        RECT 139.470 100.195 139.690 100.595 ;
        RECT 140.165 100.420 140.620 101.185 ;
        RECT 141.715 100.435 142.925 101.185 ;
        RECT 139.470 99.985 139.945 100.195 ;
        RECT 140.135 99.995 140.625 100.195 ;
        RECT 137.915 99.755 138.115 99.790 ;
        RECT 139.445 99.755 140.620 99.815 ;
        RECT 137.915 99.645 140.620 99.755 ;
        RECT 137.975 99.585 139.775 99.645 ;
        RECT 139.445 99.555 139.775 99.585 ;
        RECT 137.575 98.805 137.835 99.485 ;
        RECT 138.005 98.635 138.255 99.415 ;
        RECT 138.505 99.385 139.340 99.395 ;
        RECT 139.930 99.385 140.115 99.475 ;
        RECT 138.505 99.185 140.115 99.385 ;
        RECT 138.505 98.805 138.755 99.185 ;
        RECT 139.885 99.145 140.115 99.185 ;
        RECT 140.365 99.025 140.620 99.645 ;
        RECT 138.925 98.635 139.280 99.015 ;
        RECT 140.285 98.805 140.620 99.025 ;
        RECT 141.715 99.725 142.235 100.265 ;
        RECT 142.405 99.895 142.925 100.435 ;
        RECT 141.715 98.635 142.925 99.725 ;
        RECT 17.430 98.465 143.010 98.635 ;
        RECT 17.515 97.375 18.725 98.465 ;
        RECT 18.895 98.030 24.240 98.465 ;
        RECT 17.515 96.665 18.035 97.205 ;
        RECT 18.205 96.835 18.725 97.375 ;
        RECT 17.515 95.915 18.725 96.665 ;
        RECT 20.480 96.460 20.820 97.290 ;
        RECT 22.300 96.780 22.650 98.030 ;
        RECT 24.415 97.375 26.085 98.465 ;
        RECT 24.415 96.685 25.165 97.205 ;
        RECT 25.335 96.855 26.085 97.375 ;
        RECT 26.440 97.495 26.830 97.670 ;
        RECT 27.315 97.665 27.645 98.465 ;
        RECT 27.815 97.675 28.350 98.295 ;
        RECT 26.440 97.325 27.865 97.495 ;
        RECT 18.895 95.915 24.240 96.460 ;
        RECT 24.415 95.915 26.085 96.685 ;
        RECT 26.315 96.595 26.670 97.155 ;
        RECT 26.840 96.425 27.010 97.325 ;
        RECT 27.180 96.595 27.445 97.155 ;
        RECT 27.695 96.825 27.865 97.325 ;
        RECT 28.035 96.655 28.350 97.675 ;
        RECT 28.555 97.375 30.225 98.465 ;
        RECT 26.420 95.915 26.660 96.425 ;
        RECT 26.840 96.095 27.120 96.425 ;
        RECT 27.350 95.915 27.565 96.425 ;
        RECT 27.735 96.085 28.350 96.655 ;
        RECT 28.555 96.685 29.305 97.205 ;
        RECT 29.475 96.855 30.225 97.375 ;
        RECT 30.395 97.300 30.685 98.465 ;
        RECT 30.855 97.375 34.365 98.465 ;
        RECT 34.535 97.375 35.745 98.465 ;
        RECT 30.855 96.685 32.505 97.205 ;
        RECT 32.675 96.855 34.365 97.375 ;
        RECT 28.555 95.915 30.225 96.685 ;
        RECT 30.395 95.915 30.685 96.640 ;
        RECT 30.855 95.915 34.365 96.685 ;
        RECT 34.535 96.665 35.055 97.205 ;
        RECT 35.225 96.835 35.745 97.375 ;
        RECT 35.950 97.675 36.485 98.295 ;
        RECT 34.535 95.915 35.745 96.665 ;
        RECT 35.950 96.655 36.265 97.675 ;
        RECT 36.655 97.665 36.985 98.465 ;
        RECT 38.305 97.795 38.475 98.295 ;
        RECT 38.645 97.965 38.975 98.465 ;
        RECT 37.470 97.495 37.860 97.670 ;
        RECT 38.305 97.625 38.970 97.795 ;
        RECT 36.435 97.325 37.860 97.495 ;
        RECT 36.435 96.825 36.605 97.325 ;
        RECT 35.950 96.085 36.565 96.655 ;
        RECT 36.855 96.595 37.120 97.155 ;
        RECT 37.290 96.425 37.460 97.325 ;
        RECT 37.630 96.595 37.985 97.155 ;
        RECT 38.220 96.805 38.570 97.455 ;
        RECT 38.740 96.635 38.970 97.625 ;
        RECT 38.305 96.465 38.970 96.635 ;
        RECT 36.735 95.915 36.950 96.425 ;
        RECT 37.180 96.095 37.460 96.425 ;
        RECT 37.640 95.915 37.880 96.425 ;
        RECT 38.305 96.175 38.475 96.465 ;
        RECT 38.645 95.915 38.975 96.295 ;
        RECT 39.145 96.175 39.330 98.295 ;
        RECT 39.570 98.005 39.835 98.465 ;
        RECT 40.005 97.870 40.255 98.295 ;
        RECT 40.465 98.020 41.570 98.190 ;
        RECT 39.950 97.740 40.255 97.870 ;
        RECT 39.500 96.545 39.780 97.495 ;
        RECT 39.950 96.635 40.120 97.740 ;
        RECT 40.290 96.955 40.530 97.550 ;
        RECT 40.700 97.485 41.230 97.850 ;
        RECT 40.700 96.785 40.870 97.485 ;
        RECT 41.400 97.405 41.570 98.020 ;
        RECT 41.740 97.665 41.910 98.465 ;
        RECT 42.080 97.965 42.330 98.295 ;
        RECT 42.555 97.995 43.440 98.165 ;
        RECT 41.400 97.315 41.910 97.405 ;
        RECT 39.950 96.505 40.175 96.635 ;
        RECT 40.345 96.565 40.870 96.785 ;
        RECT 41.040 97.145 41.910 97.315 ;
        RECT 39.585 95.915 39.835 96.375 ;
        RECT 40.005 96.365 40.175 96.505 ;
        RECT 41.040 96.365 41.210 97.145 ;
        RECT 41.740 97.075 41.910 97.145 ;
        RECT 41.420 96.895 41.620 96.925 ;
        RECT 42.080 96.895 42.250 97.965 ;
        RECT 42.420 97.075 42.610 97.795 ;
        RECT 41.420 96.595 42.250 96.895 ;
        RECT 42.780 96.865 43.100 97.825 ;
        RECT 40.005 96.195 40.340 96.365 ;
        RECT 40.535 96.195 41.210 96.365 ;
        RECT 41.530 95.915 41.900 96.415 ;
        RECT 42.080 96.365 42.250 96.595 ;
        RECT 42.635 96.535 43.100 96.865 ;
        RECT 43.270 97.155 43.440 97.995 ;
        RECT 43.620 97.965 43.935 98.465 ;
        RECT 44.165 97.735 44.505 98.295 ;
        RECT 43.610 97.360 44.505 97.735 ;
        RECT 44.675 97.455 44.845 98.465 ;
        RECT 44.315 97.155 44.505 97.360 ;
        RECT 45.015 97.405 45.345 98.250 ;
        RECT 45.635 97.405 45.965 98.250 ;
        RECT 46.135 97.455 46.305 98.465 ;
        RECT 46.475 97.735 46.815 98.295 ;
        RECT 47.045 97.965 47.360 98.465 ;
        RECT 47.540 97.995 48.425 98.165 ;
        RECT 45.015 97.325 45.405 97.405 ;
        RECT 45.190 97.275 45.405 97.325 ;
        RECT 43.270 96.825 44.145 97.155 ;
        RECT 44.315 96.825 45.065 97.155 ;
        RECT 43.270 96.365 43.440 96.825 ;
        RECT 44.315 96.655 44.515 96.825 ;
        RECT 45.235 96.695 45.405 97.275 ;
        RECT 45.180 96.655 45.405 96.695 ;
        RECT 42.080 96.195 42.485 96.365 ;
        RECT 42.655 96.195 43.440 96.365 ;
        RECT 43.715 95.915 43.925 96.445 ;
        RECT 44.185 96.130 44.515 96.655 ;
        RECT 45.025 96.570 45.405 96.655 ;
        RECT 45.575 97.325 45.965 97.405 ;
        RECT 46.475 97.360 47.370 97.735 ;
        RECT 45.575 97.275 45.790 97.325 ;
        RECT 45.575 96.695 45.745 97.275 ;
        RECT 46.475 97.155 46.665 97.360 ;
        RECT 47.540 97.155 47.710 97.995 ;
        RECT 48.650 97.965 48.900 98.295 ;
        RECT 45.915 96.825 46.665 97.155 ;
        RECT 46.835 96.825 47.710 97.155 ;
        RECT 45.575 96.655 45.800 96.695 ;
        RECT 46.465 96.655 46.665 96.825 ;
        RECT 45.575 96.570 45.955 96.655 ;
        RECT 44.685 95.915 44.855 96.525 ;
        RECT 45.025 96.135 45.355 96.570 ;
        RECT 45.625 96.135 45.955 96.570 ;
        RECT 46.125 95.915 46.295 96.525 ;
        RECT 46.465 96.130 46.795 96.655 ;
        RECT 47.055 95.915 47.265 96.445 ;
        RECT 47.540 96.365 47.710 96.825 ;
        RECT 47.880 96.865 48.200 97.825 ;
        RECT 48.370 97.075 48.560 97.795 ;
        RECT 48.730 96.895 48.900 97.965 ;
        RECT 49.070 97.665 49.240 98.465 ;
        RECT 49.410 98.020 50.515 98.190 ;
        RECT 49.410 97.405 49.580 98.020 ;
        RECT 50.725 97.870 50.975 98.295 ;
        RECT 51.145 98.005 51.410 98.465 ;
        RECT 49.750 97.485 50.280 97.850 ;
        RECT 50.725 97.740 51.030 97.870 ;
        RECT 49.070 97.315 49.580 97.405 ;
        RECT 49.070 97.145 49.940 97.315 ;
        RECT 49.070 97.075 49.240 97.145 ;
        RECT 49.360 96.895 49.560 96.925 ;
        RECT 47.880 96.535 48.345 96.865 ;
        RECT 48.730 96.595 49.560 96.895 ;
        RECT 48.730 96.365 48.900 96.595 ;
        RECT 47.540 96.195 48.325 96.365 ;
        RECT 48.495 96.195 48.900 96.365 ;
        RECT 49.080 95.915 49.450 96.415 ;
        RECT 49.770 96.365 49.940 97.145 ;
        RECT 50.110 96.785 50.280 97.485 ;
        RECT 50.450 96.955 50.690 97.550 ;
        RECT 50.110 96.565 50.635 96.785 ;
        RECT 50.860 96.635 51.030 97.740 ;
        RECT 50.805 96.505 51.030 96.635 ;
        RECT 51.200 96.545 51.480 97.495 ;
        RECT 50.805 96.365 50.975 96.505 ;
        RECT 49.770 96.195 50.445 96.365 ;
        RECT 50.640 96.195 50.975 96.365 ;
        RECT 51.145 95.915 51.395 96.375 ;
        RECT 51.650 96.175 51.835 98.295 ;
        RECT 52.005 97.965 52.335 98.465 ;
        RECT 52.505 97.795 52.675 98.295 ;
        RECT 52.935 97.955 53.195 98.465 ;
        RECT 52.010 97.625 52.675 97.795 ;
        RECT 52.010 96.635 52.240 97.625 ;
        RECT 52.410 96.805 52.760 97.455 ;
        RECT 52.935 96.905 53.275 97.785 ;
        RECT 53.445 97.075 53.615 98.295 ;
        RECT 53.855 97.960 54.470 98.465 ;
        RECT 53.855 97.425 54.105 97.790 ;
        RECT 54.275 97.785 54.470 97.960 ;
        RECT 54.640 97.955 55.115 98.295 ;
        RECT 55.285 97.920 55.500 98.465 ;
        RECT 54.275 97.595 54.605 97.785 ;
        RECT 54.825 97.425 55.540 97.720 ;
        RECT 55.710 97.595 55.985 98.295 ;
        RECT 53.855 97.255 55.645 97.425 ;
        RECT 53.445 96.825 54.240 97.075 ;
        RECT 53.445 96.735 53.695 96.825 ;
        RECT 52.010 96.465 52.675 96.635 ;
        RECT 52.005 95.915 52.335 96.295 ;
        RECT 52.505 96.175 52.675 96.465 ;
        RECT 52.935 95.915 53.195 96.735 ;
        RECT 53.365 96.315 53.695 96.735 ;
        RECT 54.410 96.400 54.665 97.255 ;
        RECT 53.875 96.135 54.665 96.400 ;
        RECT 54.835 96.555 55.245 97.075 ;
        RECT 55.415 96.825 55.645 97.255 ;
        RECT 55.815 96.565 55.985 97.595 ;
        RECT 56.155 97.300 56.445 98.465 ;
        RECT 56.675 97.405 57.005 98.250 ;
        RECT 57.175 97.455 57.345 98.465 ;
        RECT 57.515 97.735 57.855 98.295 ;
        RECT 58.085 97.965 58.400 98.465 ;
        RECT 58.580 97.995 59.465 98.165 ;
        RECT 56.615 97.325 57.005 97.405 ;
        RECT 57.515 97.360 58.410 97.735 ;
        RECT 56.615 97.275 56.830 97.325 ;
        RECT 56.615 96.695 56.785 97.275 ;
        RECT 57.515 97.155 57.705 97.360 ;
        RECT 58.580 97.155 58.750 97.995 ;
        RECT 59.690 97.965 59.940 98.295 ;
        RECT 56.955 96.825 57.705 97.155 ;
        RECT 57.875 96.825 58.750 97.155 ;
        RECT 56.615 96.655 56.840 96.695 ;
        RECT 57.505 96.655 57.705 96.825 ;
        RECT 54.835 96.135 55.035 96.555 ;
        RECT 55.225 95.915 55.555 96.375 ;
        RECT 55.725 96.085 55.985 96.565 ;
        RECT 56.155 95.915 56.445 96.640 ;
        RECT 56.615 96.570 56.995 96.655 ;
        RECT 56.665 96.135 56.995 96.570 ;
        RECT 57.165 95.915 57.335 96.525 ;
        RECT 57.505 96.130 57.835 96.655 ;
        RECT 58.095 95.915 58.305 96.445 ;
        RECT 58.580 96.365 58.750 96.825 ;
        RECT 58.920 96.865 59.240 97.825 ;
        RECT 59.410 97.075 59.600 97.795 ;
        RECT 59.770 96.895 59.940 97.965 ;
        RECT 60.110 97.665 60.280 98.465 ;
        RECT 60.450 98.020 61.555 98.190 ;
        RECT 60.450 97.405 60.620 98.020 ;
        RECT 61.765 97.870 62.015 98.295 ;
        RECT 62.185 98.005 62.450 98.465 ;
        RECT 60.790 97.485 61.320 97.850 ;
        RECT 61.765 97.740 62.070 97.870 ;
        RECT 60.110 97.315 60.620 97.405 ;
        RECT 60.110 97.145 60.980 97.315 ;
        RECT 60.110 97.075 60.280 97.145 ;
        RECT 60.400 96.895 60.600 96.925 ;
        RECT 58.920 96.535 59.385 96.865 ;
        RECT 59.770 96.595 60.600 96.895 ;
        RECT 59.770 96.365 59.940 96.595 ;
        RECT 58.580 96.195 59.365 96.365 ;
        RECT 59.535 96.195 59.940 96.365 ;
        RECT 60.120 95.915 60.490 96.415 ;
        RECT 60.810 96.365 60.980 97.145 ;
        RECT 61.150 96.785 61.320 97.485 ;
        RECT 61.490 96.955 61.730 97.550 ;
        RECT 61.150 96.565 61.675 96.785 ;
        RECT 61.900 96.635 62.070 97.740 ;
        RECT 61.845 96.505 62.070 96.635 ;
        RECT 62.240 96.545 62.520 97.495 ;
        RECT 61.845 96.365 62.015 96.505 ;
        RECT 60.810 96.195 61.485 96.365 ;
        RECT 61.680 96.195 62.015 96.365 ;
        RECT 62.185 95.915 62.435 96.375 ;
        RECT 62.690 96.175 62.875 98.295 ;
        RECT 63.045 97.965 63.375 98.465 ;
        RECT 63.545 97.795 63.715 98.295 ;
        RECT 63.050 97.625 63.715 97.795 ;
        RECT 64.525 97.795 64.695 98.295 ;
        RECT 64.865 97.965 65.195 98.465 ;
        RECT 64.525 97.625 65.190 97.795 ;
        RECT 63.050 96.635 63.280 97.625 ;
        RECT 63.450 96.805 63.800 97.455 ;
        RECT 64.440 96.805 64.790 97.455 ;
        RECT 64.960 96.635 65.190 97.625 ;
        RECT 63.050 96.465 63.715 96.635 ;
        RECT 63.045 95.915 63.375 96.295 ;
        RECT 63.545 96.175 63.715 96.465 ;
        RECT 64.525 96.465 65.190 96.635 ;
        RECT 64.525 96.175 64.695 96.465 ;
        RECT 64.865 95.915 65.195 96.295 ;
        RECT 65.365 96.175 65.550 98.295 ;
        RECT 65.790 98.005 66.055 98.465 ;
        RECT 66.225 97.870 66.475 98.295 ;
        RECT 66.685 98.020 67.790 98.190 ;
        RECT 66.170 97.740 66.475 97.870 ;
        RECT 65.720 96.545 66.000 97.495 ;
        RECT 66.170 96.635 66.340 97.740 ;
        RECT 66.510 96.955 66.750 97.550 ;
        RECT 66.920 97.485 67.450 97.850 ;
        RECT 66.920 96.785 67.090 97.485 ;
        RECT 67.620 97.405 67.790 98.020 ;
        RECT 67.960 97.665 68.130 98.465 ;
        RECT 68.300 97.965 68.550 98.295 ;
        RECT 68.775 97.995 69.660 98.165 ;
        RECT 67.620 97.315 68.130 97.405 ;
        RECT 66.170 96.505 66.395 96.635 ;
        RECT 66.565 96.565 67.090 96.785 ;
        RECT 67.260 97.145 68.130 97.315 ;
        RECT 65.805 95.915 66.055 96.375 ;
        RECT 66.225 96.365 66.395 96.505 ;
        RECT 67.260 96.365 67.430 97.145 ;
        RECT 67.960 97.075 68.130 97.145 ;
        RECT 67.640 96.895 67.840 96.925 ;
        RECT 68.300 96.895 68.470 97.965 ;
        RECT 68.640 97.075 68.830 97.795 ;
        RECT 67.640 96.595 68.470 96.895 ;
        RECT 69.000 96.865 69.320 97.825 ;
        RECT 66.225 96.195 66.560 96.365 ;
        RECT 66.755 96.195 67.430 96.365 ;
        RECT 67.750 95.915 68.120 96.415 ;
        RECT 68.300 96.365 68.470 96.595 ;
        RECT 68.855 96.535 69.320 96.865 ;
        RECT 69.490 97.155 69.660 97.995 ;
        RECT 69.840 97.965 70.155 98.465 ;
        RECT 70.385 97.735 70.725 98.295 ;
        RECT 69.830 97.360 70.725 97.735 ;
        RECT 70.895 97.455 71.065 98.465 ;
        RECT 70.535 97.155 70.725 97.360 ;
        RECT 71.235 97.405 71.565 98.250 ;
        RECT 71.795 98.030 77.140 98.465 ;
        RECT 71.235 97.325 71.625 97.405 ;
        RECT 71.410 97.275 71.625 97.325 ;
        RECT 69.490 96.825 70.365 97.155 ;
        RECT 70.535 96.825 71.285 97.155 ;
        RECT 69.490 96.365 69.660 96.825 ;
        RECT 70.535 96.655 70.735 96.825 ;
        RECT 71.455 96.695 71.625 97.275 ;
        RECT 71.400 96.655 71.625 96.695 ;
        RECT 68.300 96.195 68.705 96.365 ;
        RECT 68.875 96.195 69.660 96.365 ;
        RECT 69.935 95.915 70.145 96.445 ;
        RECT 70.405 96.130 70.735 96.655 ;
        RECT 71.245 96.570 71.625 96.655 ;
        RECT 70.905 95.915 71.075 96.525 ;
        RECT 71.245 96.135 71.575 96.570 ;
        RECT 73.380 96.460 73.720 97.290 ;
        RECT 75.200 96.780 75.550 98.030 ;
        RECT 77.315 97.375 78.985 98.465 ;
        RECT 77.315 96.685 78.065 97.205 ;
        RECT 78.235 96.855 78.985 97.375 ;
        RECT 79.650 97.675 80.185 98.295 ;
        RECT 71.795 95.915 77.140 96.460 ;
        RECT 77.315 95.915 78.985 96.685 ;
        RECT 79.650 96.655 79.965 97.675 ;
        RECT 80.355 97.665 80.685 98.465 ;
        RECT 81.170 97.495 81.560 97.670 ;
        RECT 80.135 97.325 81.560 97.495 ;
        RECT 80.135 96.825 80.305 97.325 ;
        RECT 79.650 96.085 80.265 96.655 ;
        RECT 80.555 96.595 80.820 97.155 ;
        RECT 80.990 96.425 81.160 97.325 ;
        RECT 81.915 97.300 82.205 98.465 ;
        RECT 82.375 97.325 82.715 98.295 ;
        RECT 82.885 97.325 83.055 98.465 ;
        RECT 83.325 97.665 83.575 98.465 ;
        RECT 84.220 97.495 84.550 98.295 ;
        RECT 84.850 97.665 85.180 98.465 ;
        RECT 85.350 97.495 85.680 98.295 ;
        RECT 83.245 97.325 85.680 97.495 ;
        RECT 86.520 97.515 86.785 98.285 ;
        RECT 86.955 97.745 87.285 98.465 ;
        RECT 87.475 97.925 87.735 98.285 ;
        RECT 87.905 98.095 88.235 98.465 ;
        RECT 88.405 97.925 88.665 98.285 ;
        RECT 87.475 97.695 88.665 97.925 ;
        RECT 89.235 97.515 89.525 98.285 ;
        RECT 89.825 97.795 89.995 98.295 ;
        RECT 90.165 97.965 90.495 98.465 ;
        RECT 89.825 97.625 90.490 97.795 ;
        RECT 81.330 96.595 81.685 97.155 ;
        RECT 82.375 96.715 82.550 97.325 ;
        RECT 83.245 97.075 83.415 97.325 ;
        RECT 82.720 96.905 83.415 97.075 ;
        RECT 83.590 96.905 84.010 97.105 ;
        RECT 84.180 96.905 84.510 97.105 ;
        RECT 84.680 96.905 85.010 97.105 ;
        RECT 80.435 95.915 80.650 96.425 ;
        RECT 80.880 96.095 81.160 96.425 ;
        RECT 81.340 95.915 81.580 96.425 ;
        RECT 81.915 95.915 82.205 96.640 ;
        RECT 82.375 96.085 82.715 96.715 ;
        RECT 82.885 95.915 83.135 96.715 ;
        RECT 83.325 96.565 84.550 96.735 ;
        RECT 83.325 96.085 83.655 96.565 ;
        RECT 83.825 95.915 84.050 96.375 ;
        RECT 84.220 96.085 84.550 96.565 ;
        RECT 85.180 96.695 85.350 97.325 ;
        RECT 85.535 96.905 85.885 97.155 ;
        RECT 85.180 96.085 85.680 96.695 ;
        RECT 86.520 96.095 86.855 97.515 ;
        RECT 87.030 97.335 89.525 97.515 ;
        RECT 87.030 96.645 87.255 97.335 ;
        RECT 87.455 96.825 87.735 97.155 ;
        RECT 87.915 96.825 88.490 97.155 ;
        RECT 88.670 96.825 89.105 97.155 ;
        RECT 89.285 96.825 89.555 97.155 ;
        RECT 89.740 96.805 90.090 97.455 ;
        RECT 87.030 96.455 89.515 96.645 ;
        RECT 90.260 96.635 90.490 97.625 ;
        RECT 87.035 95.915 87.780 96.285 ;
        RECT 88.345 96.095 88.600 96.455 ;
        RECT 88.780 95.915 89.110 96.285 ;
        RECT 89.290 96.095 89.515 96.455 ;
        RECT 89.825 96.465 90.490 96.635 ;
        RECT 89.825 96.175 89.995 96.465 ;
        RECT 90.165 95.915 90.495 96.295 ;
        RECT 90.665 96.175 90.850 98.295 ;
        RECT 91.090 98.005 91.355 98.465 ;
        RECT 91.525 97.870 91.775 98.295 ;
        RECT 91.985 98.020 93.090 98.190 ;
        RECT 91.470 97.740 91.775 97.870 ;
        RECT 91.020 96.545 91.300 97.495 ;
        RECT 91.470 96.635 91.640 97.740 ;
        RECT 91.810 96.955 92.050 97.550 ;
        RECT 92.220 97.485 92.750 97.850 ;
        RECT 92.220 96.785 92.390 97.485 ;
        RECT 92.920 97.405 93.090 98.020 ;
        RECT 93.260 97.665 93.430 98.465 ;
        RECT 93.600 97.965 93.850 98.295 ;
        RECT 94.075 97.995 94.960 98.165 ;
        RECT 92.920 97.315 93.430 97.405 ;
        RECT 91.470 96.505 91.695 96.635 ;
        RECT 91.865 96.565 92.390 96.785 ;
        RECT 92.560 97.145 93.430 97.315 ;
        RECT 91.105 95.915 91.355 96.375 ;
        RECT 91.525 96.365 91.695 96.505 ;
        RECT 92.560 96.365 92.730 97.145 ;
        RECT 93.260 97.075 93.430 97.145 ;
        RECT 92.940 96.895 93.140 96.925 ;
        RECT 93.600 96.895 93.770 97.965 ;
        RECT 93.940 97.075 94.130 97.795 ;
        RECT 92.940 96.595 93.770 96.895 ;
        RECT 94.300 96.865 94.620 97.825 ;
        RECT 91.525 96.195 91.860 96.365 ;
        RECT 92.055 96.195 92.730 96.365 ;
        RECT 93.050 95.915 93.420 96.415 ;
        RECT 93.600 96.365 93.770 96.595 ;
        RECT 94.155 96.535 94.620 96.865 ;
        RECT 94.790 97.155 94.960 97.995 ;
        RECT 95.140 97.965 95.455 98.465 ;
        RECT 95.685 97.735 96.025 98.295 ;
        RECT 95.130 97.360 96.025 97.735 ;
        RECT 96.195 97.455 96.365 98.465 ;
        RECT 95.835 97.155 96.025 97.360 ;
        RECT 96.535 97.405 96.865 98.250 ;
        RECT 97.130 97.675 97.665 98.295 ;
        RECT 96.535 97.325 96.925 97.405 ;
        RECT 96.710 97.275 96.925 97.325 ;
        RECT 94.790 96.825 95.665 97.155 ;
        RECT 95.835 96.825 96.585 97.155 ;
        RECT 94.790 96.365 94.960 96.825 ;
        RECT 95.835 96.655 96.035 96.825 ;
        RECT 96.755 96.695 96.925 97.275 ;
        RECT 96.700 96.655 96.925 96.695 ;
        RECT 93.600 96.195 94.005 96.365 ;
        RECT 94.175 96.195 94.960 96.365 ;
        RECT 95.235 95.915 95.445 96.445 ;
        RECT 95.705 96.130 96.035 96.655 ;
        RECT 96.545 96.570 96.925 96.655 ;
        RECT 97.130 96.655 97.445 97.675 ;
        RECT 97.835 97.665 98.165 98.465 ;
        RECT 98.650 97.495 99.040 97.670 ;
        RECT 97.615 97.325 99.040 97.495 ;
        RECT 99.855 97.325 100.115 98.465 ;
        RECT 100.285 97.495 100.615 98.295 ;
        RECT 100.785 97.665 100.955 98.465 ;
        RECT 101.125 97.495 101.455 98.295 ;
        RECT 101.625 97.665 101.880 98.465 ;
        RECT 102.155 97.745 102.615 98.295 ;
        RECT 102.805 97.745 103.135 98.465 ;
        RECT 100.285 97.325 101.985 97.495 ;
        RECT 97.615 96.825 97.785 97.325 ;
        RECT 96.205 95.915 96.375 96.525 ;
        RECT 96.545 96.135 96.875 96.570 ;
        RECT 97.130 96.085 97.745 96.655 ;
        RECT 98.035 96.595 98.300 97.155 ;
        RECT 98.470 96.425 98.640 97.325 ;
        RECT 98.810 96.595 99.165 97.155 ;
        RECT 99.855 96.905 100.615 97.155 ;
        RECT 100.785 96.905 101.535 97.155 ;
        RECT 101.705 96.735 101.985 97.325 ;
        RECT 99.855 96.545 100.955 96.715 ;
        RECT 97.915 95.915 98.130 96.425 ;
        RECT 98.360 96.095 98.640 96.425 ;
        RECT 98.820 95.915 99.060 96.425 ;
        RECT 99.855 96.085 100.195 96.545 ;
        RECT 100.365 95.915 100.535 96.375 ;
        RECT 100.705 96.295 100.955 96.545 ;
        RECT 101.125 96.485 101.985 96.735 ;
        RECT 102.155 96.375 102.405 97.745 ;
        RECT 103.335 97.575 103.635 98.125 ;
        RECT 103.805 97.795 104.085 98.465 ;
        RECT 102.695 97.405 103.635 97.575 ;
        RECT 102.695 97.155 102.865 97.405 ;
        RECT 104.005 97.155 104.270 97.515 ;
        RECT 104.455 97.375 107.045 98.465 ;
        RECT 102.575 96.825 102.865 97.155 ;
        RECT 103.035 96.905 103.375 97.155 ;
        RECT 103.595 96.905 104.270 97.155 ;
        RECT 102.695 96.735 102.865 96.825 ;
        RECT 102.695 96.545 104.085 96.735 ;
        RECT 101.545 96.295 101.875 96.315 ;
        RECT 100.705 96.085 101.875 96.295 ;
        RECT 102.155 96.085 102.715 96.375 ;
        RECT 102.885 95.915 103.135 96.375 ;
        RECT 103.755 96.185 104.085 96.545 ;
        RECT 104.455 96.685 105.665 97.205 ;
        RECT 105.835 96.855 107.045 97.375 ;
        RECT 107.675 97.300 107.965 98.465 ;
        RECT 108.135 97.375 111.645 98.465 ;
        RECT 111.815 97.375 113.025 98.465 ;
        RECT 108.135 96.685 109.785 97.205 ;
        RECT 109.955 96.855 111.645 97.375 ;
        RECT 104.455 95.915 107.045 96.685 ;
        RECT 107.675 95.915 107.965 96.640 ;
        RECT 108.135 95.915 111.645 96.685 ;
        RECT 111.815 96.665 112.335 97.205 ;
        RECT 112.505 96.835 113.025 97.375 ;
        RECT 113.195 97.325 113.455 98.465 ;
        RECT 113.625 97.495 113.955 98.295 ;
        RECT 114.125 97.665 114.295 98.465 ;
        RECT 114.465 97.495 114.795 98.295 ;
        RECT 114.965 97.665 115.220 98.465 ;
        RECT 115.585 97.795 115.755 98.295 ;
        RECT 115.925 97.965 116.255 98.465 ;
        RECT 115.585 97.625 116.250 97.795 ;
        RECT 113.625 97.325 115.325 97.495 ;
        RECT 113.195 96.905 113.955 97.155 ;
        RECT 114.125 96.905 114.875 97.155 ;
        RECT 115.045 96.735 115.325 97.325 ;
        RECT 115.500 96.805 115.850 97.455 ;
        RECT 111.815 95.915 113.025 96.665 ;
        RECT 113.195 96.545 114.295 96.715 ;
        RECT 113.195 96.085 113.535 96.545 ;
        RECT 113.705 95.915 113.875 96.375 ;
        RECT 114.045 96.295 114.295 96.545 ;
        RECT 114.465 96.485 115.325 96.735 ;
        RECT 116.020 96.635 116.250 97.625 ;
        RECT 115.585 96.465 116.250 96.635 ;
        RECT 114.885 96.295 115.215 96.315 ;
        RECT 114.045 96.085 115.215 96.295 ;
        RECT 115.585 96.175 115.755 96.465 ;
        RECT 115.925 95.915 116.255 96.295 ;
        RECT 116.425 96.175 116.610 98.295 ;
        RECT 116.850 98.005 117.115 98.465 ;
        RECT 117.285 97.870 117.535 98.295 ;
        RECT 117.745 98.020 118.850 98.190 ;
        RECT 117.230 97.740 117.535 97.870 ;
        RECT 116.780 96.545 117.060 97.495 ;
        RECT 117.230 96.635 117.400 97.740 ;
        RECT 117.570 96.955 117.810 97.550 ;
        RECT 117.980 97.485 118.510 97.850 ;
        RECT 117.980 96.785 118.150 97.485 ;
        RECT 118.680 97.405 118.850 98.020 ;
        RECT 119.020 97.665 119.190 98.465 ;
        RECT 119.360 97.965 119.610 98.295 ;
        RECT 119.835 97.995 120.720 98.165 ;
        RECT 118.680 97.315 119.190 97.405 ;
        RECT 117.230 96.505 117.455 96.635 ;
        RECT 117.625 96.565 118.150 96.785 ;
        RECT 118.320 97.145 119.190 97.315 ;
        RECT 116.865 95.915 117.115 96.375 ;
        RECT 117.285 96.365 117.455 96.505 ;
        RECT 118.320 96.365 118.490 97.145 ;
        RECT 119.020 97.075 119.190 97.145 ;
        RECT 118.700 96.895 118.900 96.925 ;
        RECT 119.360 96.895 119.530 97.965 ;
        RECT 119.700 97.075 119.890 97.795 ;
        RECT 118.700 96.595 119.530 96.895 ;
        RECT 120.060 96.865 120.380 97.825 ;
        RECT 117.285 96.195 117.620 96.365 ;
        RECT 117.815 96.195 118.490 96.365 ;
        RECT 118.810 95.915 119.180 96.415 ;
        RECT 119.360 96.365 119.530 96.595 ;
        RECT 119.915 96.535 120.380 96.865 ;
        RECT 120.550 97.155 120.720 97.995 ;
        RECT 120.900 97.965 121.215 98.465 ;
        RECT 121.445 97.735 121.785 98.295 ;
        RECT 120.890 97.360 121.785 97.735 ;
        RECT 121.955 97.455 122.125 98.465 ;
        RECT 121.595 97.155 121.785 97.360 ;
        RECT 122.295 97.405 122.625 98.250 ;
        RECT 122.855 98.030 128.200 98.465 ;
        RECT 122.295 97.325 122.685 97.405 ;
        RECT 122.470 97.275 122.685 97.325 ;
        RECT 120.550 96.825 121.425 97.155 ;
        RECT 121.595 96.825 122.345 97.155 ;
        RECT 120.550 96.365 120.720 96.825 ;
        RECT 121.595 96.655 121.795 96.825 ;
        RECT 122.515 96.695 122.685 97.275 ;
        RECT 122.460 96.655 122.685 96.695 ;
        RECT 119.360 96.195 119.765 96.365 ;
        RECT 119.935 96.195 120.720 96.365 ;
        RECT 120.995 95.915 121.205 96.445 ;
        RECT 121.465 96.130 121.795 96.655 ;
        RECT 122.305 96.570 122.685 96.655 ;
        RECT 121.965 95.915 122.135 96.525 ;
        RECT 122.305 96.135 122.635 96.570 ;
        RECT 124.440 96.460 124.780 97.290 ;
        RECT 126.260 96.780 126.610 98.030 ;
        RECT 128.870 97.675 129.405 98.295 ;
        RECT 128.870 96.655 129.185 97.675 ;
        RECT 129.575 97.665 129.905 98.465 ;
        RECT 131.170 97.675 131.705 98.295 ;
        RECT 130.390 97.495 130.780 97.670 ;
        RECT 129.355 97.325 130.780 97.495 ;
        RECT 129.355 96.825 129.525 97.325 ;
        RECT 122.855 95.915 128.200 96.460 ;
        RECT 128.870 96.085 129.485 96.655 ;
        RECT 129.775 96.595 130.040 97.155 ;
        RECT 130.210 96.425 130.380 97.325 ;
        RECT 130.550 96.595 130.905 97.155 ;
        RECT 131.170 96.655 131.485 97.675 ;
        RECT 131.875 97.665 132.205 98.465 ;
        RECT 132.690 97.495 133.080 97.670 ;
        RECT 131.655 97.325 133.080 97.495 ;
        RECT 131.655 96.825 131.825 97.325 ;
        RECT 129.655 95.915 129.870 96.425 ;
        RECT 130.100 96.095 130.380 96.425 ;
        RECT 130.560 95.915 130.800 96.425 ;
        RECT 131.170 96.085 131.785 96.655 ;
        RECT 132.075 96.595 132.340 97.155 ;
        RECT 132.510 96.425 132.680 97.325 ;
        RECT 133.435 97.300 133.725 98.465 ;
        RECT 133.895 97.615 134.155 98.295 ;
        RECT 134.325 97.685 134.575 98.465 ;
        RECT 134.825 97.915 135.075 98.295 ;
        RECT 135.245 98.085 135.600 98.465 ;
        RECT 136.605 98.075 136.940 98.295 ;
        RECT 136.205 97.915 136.435 97.955 ;
        RECT 134.825 97.715 136.435 97.915 ;
        RECT 134.825 97.705 135.660 97.715 ;
        RECT 136.250 97.625 136.435 97.715 ;
        RECT 132.850 96.595 133.205 97.155 ;
        RECT 131.955 95.915 132.170 96.425 ;
        RECT 132.400 96.095 132.680 96.425 ;
        RECT 132.860 95.915 133.100 96.425 ;
        RECT 133.435 95.915 133.725 96.640 ;
        RECT 133.895 96.425 134.065 97.615 ;
        RECT 135.765 97.515 136.095 97.545 ;
        RECT 134.295 97.455 136.095 97.515 ;
        RECT 136.685 97.455 136.940 98.075 ;
        RECT 134.235 97.345 136.940 97.455 ;
        RECT 134.235 97.310 134.435 97.345 ;
        RECT 134.235 96.735 134.405 97.310 ;
        RECT 135.765 97.285 136.940 97.345 ;
        RECT 137.300 97.495 137.690 97.670 ;
        RECT 138.175 97.665 138.505 98.465 ;
        RECT 138.675 97.675 139.210 98.295 ;
        RECT 137.300 97.325 138.725 97.495 ;
        RECT 134.635 96.870 135.045 97.175 ;
        RECT 135.215 96.905 135.545 97.115 ;
        RECT 134.235 96.615 134.505 96.735 ;
        RECT 134.235 96.570 135.080 96.615 ;
        RECT 134.325 96.445 135.080 96.570 ;
        RECT 135.335 96.505 135.545 96.905 ;
        RECT 135.790 96.905 136.265 97.115 ;
        RECT 136.455 96.905 136.945 97.105 ;
        RECT 135.790 96.505 136.010 96.905 ;
        RECT 133.895 96.415 134.125 96.425 ;
        RECT 133.895 96.085 134.155 96.415 ;
        RECT 134.910 96.295 135.080 96.445 ;
        RECT 134.325 95.915 134.655 96.275 ;
        RECT 134.910 96.085 136.210 96.295 ;
        RECT 136.485 95.915 136.940 96.680 ;
        RECT 137.175 96.595 137.530 97.155 ;
        RECT 137.700 96.425 137.870 97.325 ;
        RECT 138.040 96.595 138.305 97.155 ;
        RECT 138.555 96.825 138.725 97.325 ;
        RECT 138.895 96.655 139.210 97.675 ;
        RECT 139.965 97.535 140.135 98.295 ;
        RECT 140.350 97.705 140.680 98.465 ;
        RECT 139.965 97.365 140.680 97.535 ;
        RECT 140.850 97.390 141.105 98.295 ;
        RECT 139.875 96.815 140.230 97.185 ;
        RECT 140.510 97.155 140.680 97.365 ;
        RECT 140.510 96.825 140.765 97.155 ;
        RECT 137.280 95.915 137.520 96.425 ;
        RECT 137.700 96.095 137.980 96.425 ;
        RECT 138.210 95.915 138.425 96.425 ;
        RECT 138.595 96.085 139.210 96.655 ;
        RECT 140.510 96.635 140.680 96.825 ;
        RECT 140.935 96.660 141.105 97.390 ;
        RECT 141.280 97.315 141.540 98.465 ;
        RECT 141.715 97.375 142.925 98.465 ;
        RECT 141.715 96.835 142.235 97.375 ;
        RECT 139.965 96.465 140.680 96.635 ;
        RECT 139.965 96.085 140.135 96.465 ;
        RECT 140.350 95.915 140.680 96.295 ;
        RECT 140.850 96.085 141.105 96.660 ;
        RECT 141.280 95.915 141.540 96.755 ;
        RECT 142.405 96.665 142.925 97.205 ;
        RECT 141.715 95.915 142.925 96.665 ;
        RECT 17.430 95.745 143.010 95.915 ;
        RECT 17.515 94.995 18.725 95.745 ;
        RECT 17.515 94.455 18.035 94.995 ;
        RECT 18.895 94.975 21.485 95.745 ;
        RECT 18.205 94.285 18.725 94.825 ;
        RECT 18.895 94.455 20.105 94.975 ;
        RECT 21.655 94.945 21.965 95.745 ;
        RECT 22.170 94.945 22.865 95.575 ;
        RECT 23.055 95.055 23.295 95.575 ;
        RECT 23.465 95.250 23.860 95.745 ;
        RECT 24.425 95.415 24.595 95.560 ;
        RECT 24.220 95.220 24.595 95.415 ;
        RECT 20.275 94.285 21.485 94.805 ;
        RECT 21.665 94.505 22.000 94.775 ;
        RECT 22.170 94.345 22.340 94.945 ;
        RECT 22.510 94.505 22.845 94.755 ;
        RECT 17.515 93.195 18.725 94.285 ;
        RECT 18.895 93.195 21.485 94.285 ;
        RECT 21.655 93.195 21.935 94.335 ;
        RECT 22.105 93.365 22.435 94.345 ;
        RECT 22.605 93.195 22.865 94.335 ;
        RECT 23.055 94.250 23.230 95.055 ;
        RECT 24.220 94.885 24.390 95.220 ;
        RECT 24.875 95.175 25.115 95.550 ;
        RECT 25.285 95.240 25.620 95.745 ;
        RECT 24.875 95.025 25.095 95.175 ;
        RECT 25.845 95.090 26.175 95.525 ;
        RECT 26.345 95.135 26.515 95.745 ;
        RECT 23.405 94.525 24.390 94.885 ;
        RECT 24.560 94.695 25.095 95.025 ;
        RECT 23.405 94.505 24.690 94.525 ;
        RECT 23.830 94.355 24.690 94.505 ;
        RECT 23.055 93.465 23.360 94.250 ;
        RECT 23.535 93.875 24.230 94.185 ;
        RECT 23.540 93.195 24.225 93.665 ;
        RECT 24.405 93.410 24.690 94.355 ;
        RECT 24.860 94.045 25.095 94.695 ;
        RECT 25.265 94.215 25.565 95.065 ;
        RECT 25.795 95.005 26.175 95.090 ;
        RECT 26.685 95.005 27.015 95.530 ;
        RECT 27.275 95.215 27.485 95.745 ;
        RECT 27.760 95.295 28.545 95.465 ;
        RECT 28.715 95.295 29.120 95.465 ;
        RECT 25.795 94.965 26.020 95.005 ;
        RECT 25.795 94.385 25.965 94.965 ;
        RECT 26.685 94.835 26.885 95.005 ;
        RECT 27.760 94.835 27.930 95.295 ;
        RECT 26.135 94.505 26.885 94.835 ;
        RECT 27.055 94.505 27.930 94.835 ;
        RECT 25.795 94.335 26.010 94.385 ;
        RECT 25.795 94.255 26.185 94.335 ;
        RECT 24.860 93.815 25.535 94.045 ;
        RECT 24.865 93.195 25.195 93.645 ;
        RECT 25.365 93.385 25.535 93.815 ;
        RECT 25.855 93.410 26.185 94.255 ;
        RECT 26.695 94.300 26.885 94.505 ;
        RECT 26.355 93.195 26.525 94.205 ;
        RECT 26.695 93.925 27.590 94.300 ;
        RECT 26.695 93.365 27.035 93.925 ;
        RECT 27.265 93.195 27.580 93.695 ;
        RECT 27.760 93.665 27.930 94.505 ;
        RECT 28.100 94.795 28.565 95.125 ;
        RECT 28.950 95.065 29.120 95.295 ;
        RECT 29.300 95.245 29.670 95.745 ;
        RECT 29.990 95.295 30.665 95.465 ;
        RECT 30.860 95.295 31.195 95.465 ;
        RECT 28.100 93.835 28.420 94.795 ;
        RECT 28.950 94.765 29.780 95.065 ;
        RECT 28.590 93.865 28.780 94.585 ;
        RECT 28.950 93.695 29.120 94.765 ;
        RECT 29.580 94.735 29.780 94.765 ;
        RECT 29.290 94.515 29.460 94.585 ;
        RECT 29.990 94.515 30.160 95.295 ;
        RECT 31.025 95.155 31.195 95.295 ;
        RECT 31.365 95.285 31.615 95.745 ;
        RECT 29.290 94.345 30.160 94.515 ;
        RECT 30.330 94.875 30.855 95.095 ;
        RECT 31.025 95.025 31.250 95.155 ;
        RECT 29.290 94.255 29.800 94.345 ;
        RECT 27.760 93.495 28.645 93.665 ;
        RECT 28.870 93.365 29.120 93.695 ;
        RECT 29.290 93.195 29.460 93.995 ;
        RECT 29.630 93.640 29.800 94.255 ;
        RECT 30.330 94.175 30.500 94.875 ;
        RECT 29.970 93.810 30.500 94.175 ;
        RECT 30.670 94.110 30.910 94.705 ;
        RECT 31.080 93.920 31.250 95.025 ;
        RECT 31.420 94.165 31.700 95.115 ;
        RECT 30.945 93.790 31.250 93.920 ;
        RECT 29.630 93.470 30.735 93.640 ;
        RECT 30.945 93.365 31.195 93.790 ;
        RECT 31.365 93.195 31.630 93.655 ;
        RECT 31.870 93.365 32.055 95.485 ;
        RECT 32.225 95.365 32.555 95.745 ;
        RECT 32.725 95.195 32.895 95.485 ;
        RECT 32.230 95.025 32.895 95.195 ;
        RECT 33.155 95.095 33.415 95.575 ;
        RECT 33.585 95.205 33.835 95.745 ;
        RECT 32.230 94.035 32.460 95.025 ;
        RECT 32.630 94.205 32.980 94.855 ;
        RECT 33.155 94.065 33.325 95.095 ;
        RECT 34.005 95.040 34.225 95.525 ;
        RECT 33.495 94.445 33.725 94.840 ;
        RECT 33.895 94.615 34.225 95.040 ;
        RECT 34.395 95.365 35.285 95.535 ;
        RECT 34.395 94.640 34.565 95.365 ;
        RECT 34.735 94.810 35.285 95.195 ;
        RECT 35.455 94.975 38.965 95.745 ;
        RECT 39.595 95.095 39.855 95.575 ;
        RECT 40.025 95.285 40.355 95.745 ;
        RECT 40.545 95.105 40.745 95.525 ;
        RECT 34.395 94.570 35.285 94.640 ;
        RECT 34.390 94.545 35.285 94.570 ;
        RECT 34.380 94.530 35.285 94.545 ;
        RECT 34.375 94.515 35.285 94.530 ;
        RECT 34.365 94.510 35.285 94.515 ;
        RECT 34.360 94.500 35.285 94.510 ;
        RECT 34.355 94.490 35.285 94.500 ;
        RECT 34.345 94.485 35.285 94.490 ;
        RECT 34.335 94.475 35.285 94.485 ;
        RECT 34.325 94.470 35.285 94.475 ;
        RECT 34.325 94.465 34.660 94.470 ;
        RECT 34.310 94.460 34.660 94.465 ;
        RECT 34.295 94.450 34.660 94.460 ;
        RECT 34.270 94.445 34.660 94.450 ;
        RECT 33.495 94.440 34.660 94.445 ;
        RECT 33.495 94.405 34.630 94.440 ;
        RECT 33.495 94.380 34.595 94.405 ;
        RECT 33.495 94.350 34.565 94.380 ;
        RECT 33.495 94.320 34.545 94.350 ;
        RECT 33.495 94.290 34.525 94.320 ;
        RECT 33.495 94.280 34.455 94.290 ;
        RECT 33.495 94.270 34.430 94.280 ;
        RECT 33.495 94.255 34.410 94.270 ;
        RECT 33.495 94.240 34.390 94.255 ;
        RECT 33.600 94.230 34.385 94.240 ;
        RECT 33.600 94.195 34.370 94.230 ;
        RECT 32.230 93.865 32.895 94.035 ;
        RECT 32.225 93.195 32.555 93.695 ;
        RECT 32.725 93.365 32.895 93.865 ;
        RECT 33.155 93.365 33.430 94.065 ;
        RECT 33.600 93.945 34.355 94.195 ;
        RECT 34.525 93.875 34.855 94.120 ;
        RECT 35.025 94.020 35.285 94.470 ;
        RECT 35.455 94.455 37.105 94.975 ;
        RECT 37.275 94.285 38.965 94.805 ;
        RECT 34.670 93.850 34.855 93.875 ;
        RECT 34.670 93.750 35.285 93.850 ;
        RECT 33.600 93.195 33.855 93.740 ;
        RECT 34.025 93.365 34.505 93.705 ;
        RECT 34.680 93.195 35.285 93.750 ;
        RECT 35.455 93.195 38.965 94.285 ;
        RECT 39.595 94.065 39.765 95.095 ;
        RECT 39.935 94.405 40.165 94.835 ;
        RECT 40.335 94.585 40.745 95.105 ;
        RECT 40.915 95.260 41.705 95.525 ;
        RECT 40.915 94.405 41.170 95.260 ;
        RECT 41.885 94.925 42.215 95.345 ;
        RECT 42.385 94.925 42.645 95.745 ;
        RECT 43.275 95.020 43.565 95.745 ;
        RECT 43.735 95.365 44.625 95.535 ;
        RECT 41.885 94.835 42.135 94.925 ;
        RECT 41.340 94.585 42.135 94.835 ;
        RECT 43.735 94.810 44.285 95.195 ;
        RECT 39.935 94.235 41.725 94.405 ;
        RECT 39.595 93.365 39.870 94.065 ;
        RECT 40.040 93.940 40.755 94.235 ;
        RECT 40.975 93.875 41.305 94.065 ;
        RECT 40.080 93.195 40.295 93.740 ;
        RECT 40.465 93.365 40.940 93.705 ;
        RECT 41.110 93.700 41.305 93.875 ;
        RECT 41.475 93.870 41.725 94.235 ;
        RECT 41.110 93.195 41.725 93.700 ;
        RECT 41.965 93.365 42.135 94.585 ;
        RECT 42.305 93.875 42.645 94.755 ;
        RECT 44.455 94.640 44.625 95.365 ;
        RECT 43.735 94.570 44.625 94.640 ;
        RECT 44.795 95.040 45.015 95.525 ;
        RECT 45.185 95.205 45.435 95.745 ;
        RECT 45.605 95.095 45.865 95.575 ;
        RECT 44.795 94.615 45.125 95.040 ;
        RECT 43.735 94.545 44.630 94.570 ;
        RECT 43.735 94.530 44.640 94.545 ;
        RECT 43.735 94.515 44.645 94.530 ;
        RECT 43.735 94.510 44.655 94.515 ;
        RECT 43.735 94.500 44.660 94.510 ;
        RECT 43.735 94.490 44.665 94.500 ;
        RECT 43.735 94.485 44.675 94.490 ;
        RECT 43.735 94.475 44.685 94.485 ;
        RECT 43.735 94.470 44.695 94.475 ;
        RECT 42.385 93.195 42.645 93.705 ;
        RECT 43.275 93.195 43.565 94.360 ;
        RECT 43.735 94.020 43.995 94.470 ;
        RECT 44.360 94.465 44.695 94.470 ;
        RECT 44.360 94.460 44.710 94.465 ;
        RECT 44.360 94.450 44.725 94.460 ;
        RECT 44.360 94.445 44.750 94.450 ;
        RECT 45.295 94.445 45.525 94.840 ;
        RECT 44.360 94.440 45.525 94.445 ;
        RECT 44.390 94.405 45.525 94.440 ;
        RECT 44.425 94.380 45.525 94.405 ;
        RECT 44.455 94.350 45.525 94.380 ;
        RECT 44.475 94.320 45.525 94.350 ;
        RECT 44.495 94.290 45.525 94.320 ;
        RECT 44.565 94.280 45.525 94.290 ;
        RECT 44.590 94.270 45.525 94.280 ;
        RECT 44.610 94.255 45.525 94.270 ;
        RECT 44.630 94.240 45.525 94.255 ;
        RECT 44.635 94.230 45.420 94.240 ;
        RECT 44.650 94.195 45.420 94.230 ;
        RECT 44.165 93.875 44.495 94.120 ;
        RECT 44.665 93.945 45.420 94.195 ;
        RECT 45.695 94.065 45.865 95.095 ;
        RECT 46.035 94.975 48.625 95.745 ;
        RECT 49.420 95.235 49.660 95.745 ;
        RECT 49.840 95.235 50.120 95.565 ;
        RECT 50.350 95.235 50.565 95.745 ;
        RECT 46.035 94.455 47.245 94.975 ;
        RECT 47.415 94.285 48.625 94.805 ;
        RECT 49.315 94.505 49.670 95.065 ;
        RECT 49.840 94.335 50.010 95.235 ;
        RECT 50.180 94.505 50.445 95.065 ;
        RECT 50.735 95.005 51.350 95.575 ;
        RECT 51.605 95.090 51.935 95.525 ;
        RECT 52.105 95.135 52.275 95.745 ;
        RECT 50.695 94.335 50.865 94.835 ;
        RECT 44.165 93.850 44.350 93.875 ;
        RECT 43.735 93.750 44.350 93.850 ;
        RECT 43.735 93.195 44.340 93.750 ;
        RECT 44.515 93.365 44.995 93.705 ;
        RECT 45.165 93.195 45.420 93.740 ;
        RECT 45.590 93.365 45.865 94.065 ;
        RECT 46.035 93.195 48.625 94.285 ;
        RECT 49.440 94.165 50.865 94.335 ;
        RECT 49.440 93.990 49.830 94.165 ;
        RECT 50.315 93.195 50.645 93.995 ;
        RECT 51.035 93.985 51.350 95.005 ;
        RECT 51.555 95.005 51.935 95.090 ;
        RECT 52.445 95.005 52.775 95.530 ;
        RECT 53.035 95.215 53.245 95.745 ;
        RECT 53.520 95.295 54.305 95.465 ;
        RECT 54.475 95.295 54.880 95.465 ;
        RECT 51.555 94.965 51.780 95.005 ;
        RECT 51.555 94.385 51.725 94.965 ;
        RECT 52.445 94.835 52.645 95.005 ;
        RECT 53.520 94.835 53.690 95.295 ;
        RECT 51.895 94.505 52.645 94.835 ;
        RECT 52.815 94.505 53.690 94.835 ;
        RECT 51.555 94.335 51.770 94.385 ;
        RECT 51.555 94.255 51.945 94.335 ;
        RECT 50.815 93.365 51.350 93.985 ;
        RECT 51.615 93.410 51.945 94.255 ;
        RECT 52.455 94.300 52.645 94.505 ;
        RECT 52.115 93.195 52.285 94.205 ;
        RECT 52.455 93.925 53.350 94.300 ;
        RECT 52.455 93.365 52.795 93.925 ;
        RECT 53.025 93.195 53.340 93.695 ;
        RECT 53.520 93.665 53.690 94.505 ;
        RECT 53.860 94.795 54.325 95.125 ;
        RECT 54.710 95.065 54.880 95.295 ;
        RECT 55.060 95.245 55.430 95.745 ;
        RECT 55.750 95.295 56.425 95.465 ;
        RECT 56.620 95.295 56.955 95.465 ;
        RECT 53.860 93.835 54.180 94.795 ;
        RECT 54.710 94.765 55.540 95.065 ;
        RECT 54.350 93.865 54.540 94.585 ;
        RECT 54.710 93.695 54.880 94.765 ;
        RECT 55.340 94.735 55.540 94.765 ;
        RECT 55.050 94.515 55.220 94.585 ;
        RECT 55.750 94.515 55.920 95.295 ;
        RECT 56.785 95.155 56.955 95.295 ;
        RECT 57.125 95.285 57.375 95.745 ;
        RECT 55.050 94.345 55.920 94.515 ;
        RECT 56.090 94.875 56.615 95.095 ;
        RECT 56.785 95.025 57.010 95.155 ;
        RECT 55.050 94.255 55.560 94.345 ;
        RECT 53.520 93.495 54.405 93.665 ;
        RECT 54.630 93.365 54.880 93.695 ;
        RECT 55.050 93.195 55.220 93.995 ;
        RECT 55.390 93.640 55.560 94.255 ;
        RECT 56.090 94.175 56.260 94.875 ;
        RECT 55.730 93.810 56.260 94.175 ;
        RECT 56.430 94.110 56.670 94.705 ;
        RECT 56.840 93.920 57.010 95.025 ;
        RECT 57.180 94.165 57.460 95.115 ;
        RECT 56.705 93.790 57.010 93.920 ;
        RECT 55.390 93.470 56.495 93.640 ;
        RECT 56.705 93.365 56.955 93.790 ;
        RECT 57.125 93.195 57.390 93.655 ;
        RECT 57.630 93.365 57.815 95.485 ;
        RECT 57.985 95.365 58.315 95.745 ;
        RECT 58.485 95.195 58.655 95.485 ;
        RECT 58.915 95.200 64.260 95.745 ;
        RECT 57.990 95.025 58.655 95.195 ;
        RECT 57.990 94.035 58.220 95.025 ;
        RECT 58.390 94.205 58.740 94.855 ;
        RECT 60.500 94.370 60.840 95.200 ;
        RECT 64.435 94.975 67.945 95.745 ;
        RECT 69.035 95.020 69.325 95.745 ;
        RECT 69.495 95.200 74.840 95.745 ;
        RECT 57.990 93.865 58.655 94.035 ;
        RECT 57.985 93.195 58.315 93.695 ;
        RECT 58.485 93.365 58.655 93.865 ;
        RECT 62.320 93.630 62.670 94.880 ;
        RECT 64.435 94.455 66.085 94.975 ;
        RECT 66.255 94.285 67.945 94.805 ;
        RECT 71.080 94.370 71.420 95.200 ;
        RECT 75.015 94.975 77.605 95.745 ;
        RECT 58.915 93.195 64.260 93.630 ;
        RECT 64.435 93.195 67.945 94.285 ;
        RECT 69.035 93.195 69.325 94.360 ;
        RECT 72.900 93.630 73.250 94.880 ;
        RECT 75.015 94.455 76.225 94.975 ;
        RECT 78.235 94.945 78.575 95.575 ;
        RECT 78.745 94.945 78.995 95.745 ;
        RECT 79.185 95.095 79.515 95.575 ;
        RECT 79.685 95.285 79.910 95.745 ;
        RECT 80.080 95.095 80.410 95.575 ;
        RECT 76.395 94.285 77.605 94.805 ;
        RECT 69.495 93.195 74.840 93.630 ;
        RECT 75.015 93.195 77.605 94.285 ;
        RECT 78.235 94.335 78.410 94.945 ;
        RECT 79.185 94.925 80.410 95.095 ;
        RECT 81.040 94.965 81.540 95.575 ;
        RECT 81.950 95.005 82.565 95.575 ;
        RECT 82.735 95.235 82.950 95.745 ;
        RECT 83.180 95.235 83.460 95.565 ;
        RECT 83.640 95.235 83.880 95.745 ;
        RECT 78.580 94.585 79.275 94.755 ;
        RECT 79.105 94.335 79.275 94.585 ;
        RECT 79.450 94.555 79.870 94.755 ;
        RECT 80.040 94.555 80.370 94.755 ;
        RECT 80.540 94.555 80.870 94.755 ;
        RECT 81.040 94.335 81.210 94.965 ;
        RECT 81.395 94.505 81.745 94.755 ;
        RECT 78.235 93.365 78.575 94.335 ;
        RECT 78.745 93.195 78.915 94.335 ;
        RECT 79.105 94.165 81.540 94.335 ;
        RECT 79.185 93.195 79.435 93.995 ;
        RECT 80.080 93.365 80.410 94.165 ;
        RECT 80.710 93.195 81.040 93.995 ;
        RECT 81.210 93.365 81.540 94.165 ;
        RECT 81.950 93.985 82.265 95.005 ;
        RECT 82.435 94.335 82.605 94.835 ;
        RECT 82.855 94.505 83.120 95.065 ;
        RECT 83.290 94.335 83.460 95.235 ;
        RECT 83.630 94.505 83.985 95.065 ;
        RECT 84.215 94.975 86.805 95.745 ;
        RECT 84.215 94.455 85.425 94.975 ;
        RECT 82.435 94.165 83.860 94.335 ;
        RECT 85.595 94.285 86.805 94.805 ;
        RECT 81.950 93.365 82.485 93.985 ;
        RECT 82.655 93.195 82.985 93.995 ;
        RECT 83.470 93.990 83.860 94.165 ;
        RECT 84.215 93.195 86.805 94.285 ;
        RECT 86.980 94.145 87.315 95.565 ;
        RECT 87.495 95.375 88.240 95.745 ;
        RECT 88.805 95.205 89.060 95.565 ;
        RECT 89.240 95.375 89.570 95.745 ;
        RECT 89.750 95.205 89.975 95.565 ;
        RECT 87.490 95.015 89.975 95.205 ;
        RECT 87.490 94.325 87.715 95.015 ;
        RECT 90.655 94.945 90.995 95.575 ;
        RECT 91.165 94.945 91.415 95.745 ;
        RECT 91.605 95.095 91.935 95.575 ;
        RECT 92.105 95.285 92.330 95.745 ;
        RECT 92.500 95.095 92.830 95.575 ;
        RECT 87.915 94.505 88.195 94.835 ;
        RECT 88.375 94.505 88.950 94.835 ;
        RECT 89.130 94.505 89.565 94.835 ;
        RECT 89.745 94.505 90.015 94.835 ;
        RECT 90.655 94.335 90.830 94.945 ;
        RECT 91.605 94.925 92.830 95.095 ;
        RECT 93.460 94.965 93.960 95.575 ;
        RECT 94.795 95.020 95.085 95.745 ;
        RECT 95.255 95.200 100.600 95.745 ;
        RECT 91.000 94.585 91.695 94.755 ;
        RECT 91.525 94.335 91.695 94.585 ;
        RECT 91.870 94.555 92.290 94.755 ;
        RECT 92.460 94.555 92.790 94.755 ;
        RECT 92.960 94.555 93.290 94.755 ;
        RECT 93.460 94.335 93.630 94.965 ;
        RECT 93.815 94.505 94.165 94.755 ;
        RECT 96.840 94.370 97.180 95.200 ;
        RECT 100.775 94.975 102.445 95.745 ;
        RECT 102.705 95.195 102.875 95.485 ;
        RECT 103.045 95.365 103.375 95.745 ;
        RECT 102.705 95.025 103.370 95.195 ;
        RECT 87.490 94.145 89.985 94.325 ;
        RECT 86.980 93.375 87.245 94.145 ;
        RECT 87.415 93.195 87.745 93.915 ;
        RECT 87.935 93.735 89.125 93.965 ;
        RECT 87.935 93.375 88.195 93.735 ;
        RECT 88.365 93.195 88.695 93.565 ;
        RECT 88.865 93.375 89.125 93.735 ;
        RECT 89.695 93.375 89.985 94.145 ;
        RECT 90.655 93.365 90.995 94.335 ;
        RECT 91.165 93.195 91.335 94.335 ;
        RECT 91.525 94.165 93.960 94.335 ;
        RECT 91.605 93.195 91.855 93.995 ;
        RECT 92.500 93.365 92.830 94.165 ;
        RECT 93.130 93.195 93.460 93.995 ;
        RECT 93.630 93.365 93.960 94.165 ;
        RECT 94.795 93.195 95.085 94.360 ;
        RECT 98.660 93.630 99.010 94.880 ;
        RECT 100.775 94.455 101.525 94.975 ;
        RECT 101.695 94.285 102.445 94.805 ;
        RECT 95.255 93.195 100.600 93.630 ;
        RECT 100.775 93.195 102.445 94.285 ;
        RECT 102.620 94.205 102.970 94.855 ;
        RECT 103.140 94.035 103.370 95.025 ;
        RECT 102.705 93.865 103.370 94.035 ;
        RECT 102.705 93.365 102.875 93.865 ;
        RECT 103.045 93.195 103.375 93.695 ;
        RECT 103.545 93.365 103.730 95.485 ;
        RECT 103.985 95.285 104.235 95.745 ;
        RECT 104.405 95.295 104.740 95.465 ;
        RECT 104.935 95.295 105.610 95.465 ;
        RECT 104.405 95.155 104.575 95.295 ;
        RECT 103.900 94.165 104.180 95.115 ;
        RECT 104.350 95.025 104.575 95.155 ;
        RECT 104.350 93.920 104.520 95.025 ;
        RECT 104.745 94.875 105.270 95.095 ;
        RECT 104.690 94.110 104.930 94.705 ;
        RECT 105.100 94.175 105.270 94.875 ;
        RECT 105.440 94.515 105.610 95.295 ;
        RECT 105.930 95.245 106.300 95.745 ;
        RECT 106.480 95.295 106.885 95.465 ;
        RECT 107.055 95.295 107.840 95.465 ;
        RECT 106.480 95.065 106.650 95.295 ;
        RECT 105.820 94.765 106.650 95.065 ;
        RECT 107.035 94.795 107.500 95.125 ;
        RECT 105.820 94.735 106.020 94.765 ;
        RECT 106.140 94.515 106.310 94.585 ;
        RECT 105.440 94.345 106.310 94.515 ;
        RECT 105.800 94.255 106.310 94.345 ;
        RECT 104.350 93.790 104.655 93.920 ;
        RECT 105.100 93.810 105.630 94.175 ;
        RECT 103.970 93.195 104.235 93.655 ;
        RECT 104.405 93.365 104.655 93.790 ;
        RECT 105.800 93.640 105.970 94.255 ;
        RECT 104.865 93.470 105.970 93.640 ;
        RECT 106.140 93.195 106.310 93.995 ;
        RECT 106.480 93.695 106.650 94.765 ;
        RECT 106.820 93.865 107.010 94.585 ;
        RECT 107.180 93.835 107.500 94.795 ;
        RECT 107.670 94.835 107.840 95.295 ;
        RECT 108.115 95.215 108.325 95.745 ;
        RECT 108.585 95.005 108.915 95.530 ;
        RECT 109.085 95.135 109.255 95.745 ;
        RECT 109.425 95.090 109.755 95.525 ;
        RECT 109.425 95.005 109.805 95.090 ;
        RECT 108.715 94.835 108.915 95.005 ;
        RECT 109.580 94.965 109.805 95.005 ;
        RECT 107.670 94.505 108.545 94.835 ;
        RECT 108.715 94.505 109.465 94.835 ;
        RECT 106.480 93.365 106.730 93.695 ;
        RECT 107.670 93.665 107.840 94.505 ;
        RECT 108.715 94.300 108.905 94.505 ;
        RECT 109.635 94.385 109.805 94.965 ;
        RECT 109.975 94.975 111.645 95.745 ;
        RECT 111.815 95.245 112.075 95.575 ;
        RECT 112.245 95.385 112.575 95.745 ;
        RECT 112.830 95.365 114.130 95.575 ;
        RECT 109.975 94.455 110.725 94.975 ;
        RECT 109.590 94.335 109.805 94.385 ;
        RECT 108.010 93.925 108.905 94.300 ;
        RECT 109.415 94.255 109.805 94.335 ;
        RECT 110.895 94.285 111.645 94.805 ;
        RECT 106.955 93.495 107.840 93.665 ;
        RECT 108.020 93.195 108.335 93.695 ;
        RECT 108.565 93.365 108.905 93.925 ;
        RECT 109.075 93.195 109.245 94.205 ;
        RECT 109.415 93.410 109.745 94.255 ;
        RECT 109.975 93.195 111.645 94.285 ;
        RECT 111.815 94.045 111.985 95.245 ;
        RECT 112.830 95.215 113.000 95.365 ;
        RECT 112.245 95.090 113.000 95.215 ;
        RECT 112.155 95.045 113.000 95.090 ;
        RECT 112.155 94.925 112.425 95.045 ;
        RECT 112.155 94.350 112.325 94.925 ;
        RECT 112.555 94.485 112.965 94.790 ;
        RECT 113.255 94.755 113.465 95.155 ;
        RECT 113.135 94.545 113.465 94.755 ;
        RECT 113.710 94.755 113.930 95.155 ;
        RECT 114.405 94.980 114.860 95.745 ;
        RECT 115.035 94.975 116.705 95.745 ;
        RECT 113.710 94.545 114.185 94.755 ;
        RECT 114.375 94.555 114.865 94.755 ;
        RECT 115.035 94.455 115.785 94.975 ;
        RECT 116.875 94.945 117.215 95.575 ;
        RECT 117.385 94.945 117.635 95.745 ;
        RECT 117.825 95.095 118.155 95.575 ;
        RECT 118.325 95.285 118.550 95.745 ;
        RECT 118.720 95.095 119.050 95.575 ;
        RECT 112.155 94.315 112.355 94.350 ;
        RECT 113.685 94.315 114.860 94.375 ;
        RECT 112.155 94.205 114.860 94.315 ;
        RECT 115.955 94.285 116.705 94.805 ;
        RECT 112.215 94.145 114.015 94.205 ;
        RECT 113.685 94.115 114.015 94.145 ;
        RECT 111.815 93.365 112.075 94.045 ;
        RECT 112.245 93.195 112.495 93.975 ;
        RECT 112.745 93.945 113.580 93.955 ;
        RECT 114.170 93.945 114.355 94.035 ;
        RECT 112.745 93.745 114.355 93.945 ;
        RECT 112.745 93.365 112.995 93.745 ;
        RECT 114.125 93.705 114.355 93.745 ;
        RECT 114.605 93.585 114.860 94.205 ;
        RECT 113.165 93.195 113.520 93.575 ;
        RECT 114.525 93.365 114.860 93.585 ;
        RECT 115.035 93.195 116.705 94.285 ;
        RECT 116.875 94.385 117.050 94.945 ;
        RECT 117.825 94.925 119.050 95.095 ;
        RECT 119.680 94.965 120.180 95.575 ;
        RECT 120.555 95.020 120.845 95.745 ;
        RECT 121.105 95.195 121.275 95.485 ;
        RECT 121.445 95.365 121.775 95.745 ;
        RECT 121.105 95.025 121.770 95.195 ;
        RECT 117.220 94.585 117.915 94.755 ;
        RECT 116.875 94.335 117.105 94.385 ;
        RECT 117.745 94.335 117.915 94.585 ;
        RECT 118.090 94.555 118.510 94.755 ;
        RECT 118.680 94.555 119.010 94.755 ;
        RECT 119.180 94.555 119.510 94.755 ;
        RECT 119.680 94.335 119.850 94.965 ;
        RECT 120.035 94.505 120.385 94.755 ;
        RECT 116.875 93.365 117.215 94.335 ;
        RECT 117.385 93.195 117.555 94.335 ;
        RECT 117.745 94.165 120.180 94.335 ;
        RECT 117.825 93.195 118.075 93.995 ;
        RECT 118.720 93.365 119.050 94.165 ;
        RECT 119.350 93.195 119.680 93.995 ;
        RECT 119.850 93.365 120.180 94.165 ;
        RECT 120.555 93.195 120.845 94.360 ;
        RECT 121.020 94.205 121.370 94.855 ;
        RECT 121.540 94.035 121.770 95.025 ;
        RECT 121.105 93.865 121.770 94.035 ;
        RECT 121.105 93.365 121.275 93.865 ;
        RECT 121.445 93.195 121.775 93.695 ;
        RECT 121.945 93.365 122.130 95.485 ;
        RECT 122.385 95.285 122.635 95.745 ;
        RECT 122.805 95.295 123.140 95.465 ;
        RECT 123.335 95.295 124.010 95.465 ;
        RECT 122.805 95.155 122.975 95.295 ;
        RECT 122.300 94.165 122.580 95.115 ;
        RECT 122.750 95.025 122.975 95.155 ;
        RECT 122.750 93.920 122.920 95.025 ;
        RECT 123.145 94.875 123.670 95.095 ;
        RECT 123.090 94.110 123.330 94.705 ;
        RECT 123.500 94.175 123.670 94.875 ;
        RECT 123.840 94.515 124.010 95.295 ;
        RECT 124.330 95.245 124.700 95.745 ;
        RECT 124.880 95.295 125.285 95.465 ;
        RECT 125.455 95.295 126.240 95.465 ;
        RECT 124.880 95.065 125.050 95.295 ;
        RECT 124.220 94.765 125.050 95.065 ;
        RECT 125.435 94.795 125.900 95.125 ;
        RECT 124.220 94.735 124.420 94.765 ;
        RECT 124.540 94.515 124.710 94.585 ;
        RECT 123.840 94.345 124.710 94.515 ;
        RECT 124.200 94.255 124.710 94.345 ;
        RECT 122.750 93.790 123.055 93.920 ;
        RECT 123.500 93.810 124.030 94.175 ;
        RECT 122.370 93.195 122.635 93.655 ;
        RECT 122.805 93.365 123.055 93.790 ;
        RECT 124.200 93.640 124.370 94.255 ;
        RECT 123.265 93.470 124.370 93.640 ;
        RECT 124.540 93.195 124.710 93.995 ;
        RECT 124.880 93.695 125.050 94.765 ;
        RECT 125.220 93.865 125.410 94.585 ;
        RECT 125.580 93.835 125.900 94.795 ;
        RECT 126.070 94.835 126.240 95.295 ;
        RECT 126.515 95.215 126.725 95.745 ;
        RECT 126.985 95.005 127.315 95.530 ;
        RECT 127.485 95.135 127.655 95.745 ;
        RECT 127.825 95.090 128.155 95.525 ;
        RECT 127.825 95.005 128.205 95.090 ;
        RECT 127.115 94.835 127.315 95.005 ;
        RECT 127.980 94.965 128.205 95.005 ;
        RECT 129.040 94.965 129.540 95.575 ;
        RECT 126.070 94.505 126.945 94.835 ;
        RECT 127.115 94.505 127.865 94.835 ;
        RECT 124.880 93.365 125.130 93.695 ;
        RECT 126.070 93.665 126.240 94.505 ;
        RECT 127.115 94.300 127.305 94.505 ;
        RECT 128.035 94.385 128.205 94.965 ;
        RECT 128.835 94.505 129.185 94.755 ;
        RECT 127.990 94.335 128.205 94.385 ;
        RECT 129.370 94.335 129.540 94.965 ;
        RECT 130.170 95.095 130.500 95.575 ;
        RECT 130.670 95.285 130.895 95.745 ;
        RECT 131.065 95.095 131.395 95.575 ;
        RECT 130.170 94.925 131.395 95.095 ;
        RECT 131.585 94.945 131.835 95.745 ;
        RECT 132.005 94.945 132.345 95.575 ;
        RECT 132.605 95.195 132.775 95.485 ;
        RECT 132.945 95.365 133.275 95.745 ;
        RECT 132.605 95.025 133.270 95.195 ;
        RECT 129.710 94.555 130.040 94.755 ;
        RECT 130.210 94.555 130.540 94.755 ;
        RECT 130.710 94.555 131.130 94.755 ;
        RECT 131.305 94.585 132.000 94.755 ;
        RECT 131.305 94.335 131.475 94.585 ;
        RECT 132.170 94.335 132.345 94.945 ;
        RECT 126.410 93.925 127.305 94.300 ;
        RECT 127.815 94.255 128.205 94.335 ;
        RECT 125.355 93.495 126.240 93.665 ;
        RECT 126.420 93.195 126.735 93.695 ;
        RECT 126.965 93.365 127.305 93.925 ;
        RECT 127.475 93.195 127.645 94.205 ;
        RECT 127.815 93.410 128.145 94.255 ;
        RECT 129.040 94.165 131.475 94.335 ;
        RECT 129.040 93.365 129.370 94.165 ;
        RECT 129.540 93.195 129.870 93.995 ;
        RECT 130.170 93.365 130.500 94.165 ;
        RECT 131.145 93.195 131.395 93.995 ;
        RECT 131.665 93.195 131.835 94.335 ;
        RECT 132.005 93.365 132.345 94.335 ;
        RECT 132.520 94.205 132.870 94.855 ;
        RECT 133.040 94.035 133.270 95.025 ;
        RECT 132.605 93.865 133.270 94.035 ;
        RECT 132.605 93.365 132.775 93.865 ;
        RECT 132.945 93.195 133.275 93.695 ;
        RECT 133.445 93.365 133.630 95.485 ;
        RECT 133.885 95.285 134.135 95.745 ;
        RECT 134.305 95.295 134.640 95.465 ;
        RECT 134.835 95.295 135.510 95.465 ;
        RECT 134.305 95.155 134.475 95.295 ;
        RECT 133.800 94.165 134.080 95.115 ;
        RECT 134.250 95.025 134.475 95.155 ;
        RECT 134.250 93.920 134.420 95.025 ;
        RECT 134.645 94.875 135.170 95.095 ;
        RECT 134.590 94.110 134.830 94.705 ;
        RECT 135.000 94.175 135.170 94.875 ;
        RECT 135.340 94.515 135.510 95.295 ;
        RECT 135.830 95.245 136.200 95.745 ;
        RECT 136.380 95.295 136.785 95.465 ;
        RECT 136.955 95.295 137.740 95.465 ;
        RECT 136.380 95.065 136.550 95.295 ;
        RECT 135.720 94.765 136.550 95.065 ;
        RECT 136.935 94.795 137.400 95.125 ;
        RECT 135.720 94.735 135.920 94.765 ;
        RECT 136.040 94.515 136.210 94.585 ;
        RECT 135.340 94.345 136.210 94.515 ;
        RECT 135.700 94.255 136.210 94.345 ;
        RECT 134.250 93.790 134.555 93.920 ;
        RECT 135.000 93.810 135.530 94.175 ;
        RECT 133.870 93.195 134.135 93.655 ;
        RECT 134.305 93.365 134.555 93.790 ;
        RECT 135.700 93.640 135.870 94.255 ;
        RECT 134.765 93.470 135.870 93.640 ;
        RECT 136.040 93.195 136.210 93.995 ;
        RECT 136.380 93.695 136.550 94.765 ;
        RECT 136.720 93.865 136.910 94.585 ;
        RECT 137.080 93.835 137.400 94.795 ;
        RECT 137.570 94.835 137.740 95.295 ;
        RECT 138.015 95.215 138.225 95.745 ;
        RECT 138.485 95.005 138.815 95.530 ;
        RECT 138.985 95.135 139.155 95.745 ;
        RECT 139.325 95.090 139.655 95.525 ;
        RECT 139.965 95.195 140.135 95.575 ;
        RECT 140.350 95.365 140.680 95.745 ;
        RECT 139.325 95.005 139.705 95.090 ;
        RECT 139.965 95.025 140.680 95.195 ;
        RECT 138.615 94.835 138.815 95.005 ;
        RECT 139.480 94.965 139.705 95.005 ;
        RECT 137.570 94.505 138.445 94.835 ;
        RECT 138.615 94.505 139.365 94.835 ;
        RECT 136.380 93.365 136.630 93.695 ;
        RECT 137.570 93.665 137.740 94.505 ;
        RECT 138.615 94.300 138.805 94.505 ;
        RECT 139.535 94.385 139.705 94.965 ;
        RECT 139.875 94.475 140.230 94.845 ;
        RECT 140.510 94.835 140.680 95.025 ;
        RECT 140.850 95.000 141.105 95.575 ;
        RECT 140.510 94.505 140.765 94.835 ;
        RECT 139.490 94.335 139.705 94.385 ;
        RECT 137.910 93.925 138.805 94.300 ;
        RECT 139.315 94.255 139.705 94.335 ;
        RECT 140.510 94.295 140.680 94.505 ;
        RECT 136.855 93.495 137.740 93.665 ;
        RECT 137.920 93.195 138.235 93.695 ;
        RECT 138.465 93.365 138.805 93.925 ;
        RECT 138.975 93.195 139.145 94.205 ;
        RECT 139.315 93.410 139.645 94.255 ;
        RECT 139.965 94.125 140.680 94.295 ;
        RECT 140.935 94.270 141.105 95.000 ;
        RECT 141.280 94.905 141.540 95.745 ;
        RECT 141.715 94.995 142.925 95.745 ;
        RECT 139.965 93.365 140.135 94.125 ;
        RECT 140.350 93.195 140.680 93.955 ;
        RECT 140.850 93.365 141.105 94.270 ;
        RECT 141.280 93.195 141.540 94.345 ;
        RECT 141.715 94.285 142.235 94.825 ;
        RECT 142.405 94.455 142.925 94.995 ;
        RECT 141.715 93.195 142.925 94.285 ;
        RECT 17.430 93.025 143.010 93.195 ;
        RECT 17.515 91.935 18.725 93.025 ;
        RECT 18.895 91.935 22.405 93.025 ;
        RECT 22.665 92.355 22.835 92.855 ;
        RECT 23.005 92.525 23.335 93.025 ;
        RECT 22.665 92.185 23.330 92.355 ;
        RECT 17.515 91.225 18.035 91.765 ;
        RECT 18.205 91.395 18.725 91.935 ;
        RECT 18.895 91.245 20.545 91.765 ;
        RECT 20.715 91.415 22.405 91.935 ;
        RECT 22.580 91.365 22.930 92.015 ;
        RECT 17.515 90.475 18.725 91.225 ;
        RECT 18.895 90.475 22.405 91.245 ;
        RECT 23.100 91.195 23.330 92.185 ;
        RECT 22.665 91.025 23.330 91.195 ;
        RECT 22.665 90.735 22.835 91.025 ;
        RECT 23.005 90.475 23.335 90.855 ;
        RECT 23.505 90.735 23.690 92.855 ;
        RECT 23.930 92.565 24.195 93.025 ;
        RECT 24.365 92.430 24.615 92.855 ;
        RECT 24.825 92.580 25.930 92.750 ;
        RECT 24.310 92.300 24.615 92.430 ;
        RECT 23.860 91.105 24.140 92.055 ;
        RECT 24.310 91.195 24.480 92.300 ;
        RECT 24.650 91.515 24.890 92.110 ;
        RECT 25.060 92.045 25.590 92.410 ;
        RECT 25.060 91.345 25.230 92.045 ;
        RECT 25.760 91.965 25.930 92.580 ;
        RECT 26.100 92.225 26.270 93.025 ;
        RECT 26.440 92.525 26.690 92.855 ;
        RECT 26.915 92.555 27.800 92.725 ;
        RECT 25.760 91.875 26.270 91.965 ;
        RECT 24.310 91.065 24.535 91.195 ;
        RECT 24.705 91.125 25.230 91.345 ;
        RECT 25.400 91.705 26.270 91.875 ;
        RECT 23.945 90.475 24.195 90.935 ;
        RECT 24.365 90.925 24.535 91.065 ;
        RECT 25.400 90.925 25.570 91.705 ;
        RECT 26.100 91.635 26.270 91.705 ;
        RECT 25.780 91.455 25.980 91.485 ;
        RECT 26.440 91.455 26.610 92.525 ;
        RECT 26.780 91.635 26.970 92.355 ;
        RECT 25.780 91.155 26.610 91.455 ;
        RECT 27.140 91.425 27.460 92.385 ;
        RECT 24.365 90.755 24.700 90.925 ;
        RECT 24.895 90.755 25.570 90.925 ;
        RECT 25.890 90.475 26.260 90.975 ;
        RECT 26.440 90.925 26.610 91.155 ;
        RECT 26.995 91.095 27.460 91.425 ;
        RECT 27.630 91.715 27.800 92.555 ;
        RECT 27.980 92.525 28.295 93.025 ;
        RECT 28.525 92.295 28.865 92.855 ;
        RECT 27.970 91.920 28.865 92.295 ;
        RECT 29.035 92.015 29.205 93.025 ;
        RECT 28.675 91.715 28.865 91.920 ;
        RECT 29.375 91.965 29.705 92.810 ;
        RECT 29.375 91.885 29.765 91.965 ;
        RECT 29.550 91.835 29.765 91.885 ;
        RECT 30.395 91.860 30.685 93.025 ;
        RECT 30.855 92.590 36.200 93.025 ;
        RECT 36.375 92.590 41.720 93.025 ;
        RECT 41.895 92.590 47.240 93.025 ;
        RECT 47.415 92.590 52.760 93.025 ;
        RECT 27.630 91.385 28.505 91.715 ;
        RECT 28.675 91.385 29.425 91.715 ;
        RECT 27.630 90.925 27.800 91.385 ;
        RECT 28.675 91.215 28.875 91.385 ;
        RECT 29.595 91.255 29.765 91.835 ;
        RECT 29.540 91.215 29.765 91.255 ;
        RECT 26.440 90.755 26.845 90.925 ;
        RECT 27.015 90.755 27.800 90.925 ;
        RECT 28.075 90.475 28.285 91.005 ;
        RECT 28.545 90.690 28.875 91.215 ;
        RECT 29.385 91.130 29.765 91.215 ;
        RECT 29.045 90.475 29.215 91.085 ;
        RECT 29.385 90.695 29.715 91.130 ;
        RECT 30.395 90.475 30.685 91.200 ;
        RECT 32.440 91.020 32.780 91.850 ;
        RECT 34.260 91.340 34.610 92.590 ;
        RECT 37.960 91.020 38.300 91.850 ;
        RECT 39.780 91.340 40.130 92.590 ;
        RECT 43.480 91.020 43.820 91.850 ;
        RECT 45.300 91.340 45.650 92.590 ;
        RECT 49.000 91.020 49.340 91.850 ;
        RECT 50.820 91.340 51.170 92.590 ;
        RECT 52.935 91.885 53.195 93.025 ;
        RECT 53.365 91.875 53.695 92.855 ;
        RECT 53.865 91.885 54.145 93.025 ;
        RECT 54.315 91.935 55.985 93.025 ;
        RECT 52.955 91.465 53.290 91.715 ;
        RECT 53.460 91.275 53.630 91.875 ;
        RECT 53.800 91.445 54.135 91.715 ;
        RECT 30.855 90.475 36.200 91.020 ;
        RECT 36.375 90.475 41.720 91.020 ;
        RECT 41.895 90.475 47.240 91.020 ;
        RECT 47.415 90.475 52.760 91.020 ;
        RECT 52.935 90.645 53.630 91.275 ;
        RECT 53.835 90.475 54.145 91.275 ;
        RECT 54.315 91.245 55.065 91.765 ;
        RECT 55.235 91.415 55.985 91.935 ;
        RECT 56.155 91.860 56.445 93.025 ;
        RECT 56.615 92.590 61.960 93.025 ;
        RECT 62.135 92.590 67.480 93.025 ;
        RECT 67.655 92.590 73.000 93.025 ;
        RECT 54.315 90.475 55.985 91.245 ;
        RECT 56.155 90.475 56.445 91.200 ;
        RECT 58.200 91.020 58.540 91.850 ;
        RECT 60.020 91.340 60.370 92.590 ;
        RECT 63.720 91.020 64.060 91.850 ;
        RECT 65.540 91.340 65.890 92.590 ;
        RECT 69.240 91.020 69.580 91.850 ;
        RECT 71.060 91.340 71.410 92.590 ;
        RECT 73.175 91.935 74.385 93.025 ;
        RECT 74.645 92.355 74.815 92.855 ;
        RECT 74.985 92.525 75.315 93.025 ;
        RECT 74.645 92.185 75.310 92.355 ;
        RECT 73.175 91.225 73.695 91.765 ;
        RECT 73.865 91.395 74.385 91.935 ;
        RECT 74.560 91.365 74.910 92.015 ;
        RECT 56.615 90.475 61.960 91.020 ;
        RECT 62.135 90.475 67.480 91.020 ;
        RECT 67.655 90.475 73.000 91.020 ;
        RECT 73.175 90.475 74.385 91.225 ;
        RECT 75.080 91.195 75.310 92.185 ;
        RECT 74.645 91.025 75.310 91.195 ;
        RECT 74.645 90.735 74.815 91.025 ;
        RECT 74.985 90.475 75.315 90.855 ;
        RECT 75.485 90.735 75.670 92.855 ;
        RECT 75.910 92.565 76.175 93.025 ;
        RECT 76.345 92.430 76.595 92.855 ;
        RECT 76.805 92.580 77.910 92.750 ;
        RECT 76.290 92.300 76.595 92.430 ;
        RECT 75.840 91.105 76.120 92.055 ;
        RECT 76.290 91.195 76.460 92.300 ;
        RECT 76.630 91.515 76.870 92.110 ;
        RECT 77.040 92.045 77.570 92.410 ;
        RECT 77.040 91.345 77.210 92.045 ;
        RECT 77.740 91.965 77.910 92.580 ;
        RECT 78.080 92.225 78.250 93.025 ;
        RECT 78.420 92.525 78.670 92.855 ;
        RECT 78.895 92.555 79.780 92.725 ;
        RECT 77.740 91.875 78.250 91.965 ;
        RECT 76.290 91.065 76.515 91.195 ;
        RECT 76.685 91.125 77.210 91.345 ;
        RECT 77.380 91.705 78.250 91.875 ;
        RECT 75.925 90.475 76.175 90.935 ;
        RECT 76.345 90.925 76.515 91.065 ;
        RECT 77.380 90.925 77.550 91.705 ;
        RECT 78.080 91.635 78.250 91.705 ;
        RECT 77.760 91.455 77.960 91.485 ;
        RECT 78.420 91.455 78.590 92.525 ;
        RECT 78.760 91.635 78.950 92.355 ;
        RECT 77.760 91.155 78.590 91.455 ;
        RECT 79.120 91.425 79.440 92.385 ;
        RECT 76.345 90.755 76.680 90.925 ;
        RECT 76.875 90.755 77.550 90.925 ;
        RECT 77.870 90.475 78.240 90.975 ;
        RECT 78.420 90.925 78.590 91.155 ;
        RECT 78.975 91.095 79.440 91.425 ;
        RECT 79.610 91.715 79.780 92.555 ;
        RECT 79.960 92.525 80.275 93.025 ;
        RECT 80.505 92.295 80.845 92.855 ;
        RECT 79.950 91.920 80.845 92.295 ;
        RECT 81.015 92.015 81.185 93.025 ;
        RECT 80.655 91.715 80.845 91.920 ;
        RECT 81.355 91.965 81.685 92.810 ;
        RECT 81.355 91.885 81.745 91.965 ;
        RECT 81.530 91.835 81.745 91.885 ;
        RECT 81.915 91.860 82.205 93.025 ;
        RECT 82.375 91.885 82.715 92.855 ;
        RECT 82.885 91.885 83.055 93.025 ;
        RECT 83.325 92.225 83.575 93.025 ;
        RECT 84.220 92.055 84.550 92.855 ;
        RECT 84.850 92.225 85.180 93.025 ;
        RECT 85.350 92.055 85.680 92.855 ;
        RECT 83.245 91.885 85.680 92.055 ;
        RECT 86.605 92.095 86.775 92.855 ;
        RECT 86.990 92.265 87.320 93.025 ;
        RECT 86.605 91.925 87.320 92.095 ;
        RECT 87.490 91.950 87.745 92.855 ;
        RECT 79.610 91.385 80.485 91.715 ;
        RECT 80.655 91.385 81.405 91.715 ;
        RECT 79.610 90.925 79.780 91.385 ;
        RECT 80.655 91.215 80.855 91.385 ;
        RECT 81.575 91.255 81.745 91.835 ;
        RECT 81.520 91.215 81.745 91.255 ;
        RECT 78.420 90.755 78.825 90.925 ;
        RECT 78.995 90.755 79.780 90.925 ;
        RECT 80.055 90.475 80.265 91.005 ;
        RECT 80.525 90.690 80.855 91.215 ;
        RECT 81.365 91.130 81.745 91.215 ;
        RECT 82.375 91.275 82.550 91.885 ;
        RECT 83.245 91.635 83.415 91.885 ;
        RECT 82.720 91.465 83.415 91.635 ;
        RECT 83.590 91.465 84.010 91.665 ;
        RECT 84.180 91.465 84.510 91.665 ;
        RECT 84.680 91.465 85.010 91.665 ;
        RECT 81.025 90.475 81.195 91.085 ;
        RECT 81.365 90.695 81.695 91.130 ;
        RECT 81.915 90.475 82.205 91.200 ;
        RECT 82.375 90.645 82.715 91.275 ;
        RECT 82.885 90.475 83.135 91.275 ;
        RECT 83.325 91.125 84.550 91.295 ;
        RECT 83.325 90.645 83.655 91.125 ;
        RECT 83.825 90.475 84.050 90.935 ;
        RECT 84.220 90.645 84.550 91.125 ;
        RECT 85.180 91.255 85.350 91.885 ;
        RECT 85.535 91.465 85.885 91.715 ;
        RECT 86.515 91.375 86.870 91.745 ;
        RECT 87.150 91.715 87.320 91.925 ;
        RECT 87.150 91.385 87.405 91.715 ;
        RECT 85.180 90.645 85.680 91.255 ;
        RECT 87.150 91.195 87.320 91.385 ;
        RECT 87.575 91.220 87.745 91.950 ;
        RECT 87.920 91.875 88.180 93.025 ;
        RECT 88.355 91.935 90.945 93.025 ;
        RECT 86.605 91.025 87.320 91.195 ;
        RECT 86.605 90.645 86.775 91.025 ;
        RECT 86.990 90.475 87.320 90.855 ;
        RECT 87.490 90.645 87.745 91.220 ;
        RECT 87.920 90.475 88.180 91.315 ;
        RECT 88.355 91.245 89.565 91.765 ;
        RECT 89.735 91.415 90.945 91.935 ;
        RECT 91.115 92.175 91.375 92.855 ;
        RECT 91.545 92.245 91.795 93.025 ;
        RECT 92.045 92.475 92.295 92.855 ;
        RECT 92.465 92.645 92.820 93.025 ;
        RECT 93.825 92.635 94.160 92.855 ;
        RECT 93.425 92.475 93.655 92.515 ;
        RECT 92.045 92.275 93.655 92.475 ;
        RECT 92.045 92.265 92.880 92.275 ;
        RECT 93.470 92.185 93.655 92.275 ;
        RECT 88.355 90.475 90.945 91.245 ;
        RECT 91.115 90.975 91.285 92.175 ;
        RECT 92.985 92.075 93.315 92.105 ;
        RECT 91.515 92.015 93.315 92.075 ;
        RECT 93.905 92.015 94.160 92.635 ;
        RECT 94.335 92.590 99.680 93.025 ;
        RECT 91.455 91.905 94.160 92.015 ;
        RECT 91.455 91.870 91.655 91.905 ;
        RECT 91.455 91.295 91.625 91.870 ;
        RECT 92.985 91.845 94.160 91.905 ;
        RECT 91.855 91.430 92.265 91.735 ;
        RECT 92.435 91.465 92.765 91.675 ;
        RECT 91.455 91.175 91.725 91.295 ;
        RECT 91.455 91.130 92.300 91.175 ;
        RECT 91.545 91.005 92.300 91.130 ;
        RECT 92.555 91.065 92.765 91.465 ;
        RECT 93.010 91.465 93.485 91.675 ;
        RECT 93.675 91.465 94.165 91.665 ;
        RECT 93.010 91.065 93.230 91.465 ;
        RECT 91.115 90.645 91.375 90.975 ;
        RECT 92.130 90.855 92.300 91.005 ;
        RECT 91.545 90.475 91.875 90.835 ;
        RECT 92.130 90.645 93.430 90.855 ;
        RECT 93.705 90.475 94.160 91.240 ;
        RECT 95.920 91.020 96.260 91.850 ;
        RECT 97.740 91.340 98.090 92.590 ;
        RECT 99.855 91.935 101.525 93.025 ;
        RECT 99.855 91.245 100.605 91.765 ;
        RECT 100.775 91.415 101.525 91.935 ;
        RECT 102.155 91.885 102.495 92.855 ;
        RECT 102.665 91.885 102.835 93.025 ;
        RECT 103.105 92.225 103.355 93.025 ;
        RECT 104.000 92.055 104.330 92.855 ;
        RECT 104.630 92.225 104.960 93.025 ;
        RECT 105.130 92.055 105.460 92.855 ;
        RECT 103.025 91.885 105.460 92.055 ;
        RECT 102.155 91.275 102.330 91.885 ;
        RECT 103.025 91.635 103.195 91.885 ;
        RECT 102.500 91.465 103.195 91.635 ;
        RECT 103.370 91.465 103.790 91.665 ;
        RECT 103.960 91.465 104.290 91.665 ;
        RECT 104.460 91.465 104.790 91.665 ;
        RECT 94.335 90.475 99.680 91.020 ;
        RECT 99.855 90.475 101.525 91.245 ;
        RECT 102.155 90.645 102.495 91.275 ;
        RECT 102.665 90.475 102.915 91.275 ;
        RECT 103.105 91.125 104.330 91.295 ;
        RECT 103.105 90.645 103.435 91.125 ;
        RECT 103.605 90.475 103.830 90.935 ;
        RECT 104.000 90.645 104.330 91.125 ;
        RECT 104.960 91.255 105.130 91.885 ;
        RECT 105.840 91.875 106.100 93.025 ;
        RECT 106.275 91.950 106.530 92.855 ;
        RECT 106.700 92.265 107.030 93.025 ;
        RECT 107.245 92.095 107.415 92.855 ;
        RECT 105.315 91.465 105.665 91.715 ;
        RECT 104.960 90.645 105.460 91.255 ;
        RECT 105.840 90.475 106.100 91.315 ;
        RECT 106.275 91.220 106.445 91.950 ;
        RECT 106.700 91.925 107.415 92.095 ;
        RECT 106.700 91.715 106.870 91.925 ;
        RECT 107.675 91.860 107.965 93.025 ;
        RECT 108.170 92.235 108.705 92.855 ;
        RECT 106.615 91.385 106.870 91.715 ;
        RECT 106.275 90.645 106.530 91.220 ;
        RECT 106.700 91.195 106.870 91.385 ;
        RECT 107.150 91.375 107.505 91.745 ;
        RECT 108.170 91.215 108.485 92.235 ;
        RECT 108.875 92.225 109.205 93.025 ;
        RECT 110.435 92.590 115.780 93.025 ;
        RECT 109.690 92.055 110.080 92.230 ;
        RECT 108.655 91.885 110.080 92.055 ;
        RECT 108.655 91.385 108.825 91.885 ;
        RECT 106.700 91.025 107.415 91.195 ;
        RECT 106.700 90.475 107.030 90.855 ;
        RECT 107.245 90.645 107.415 91.025 ;
        RECT 107.675 90.475 107.965 91.200 ;
        RECT 108.170 90.645 108.785 91.215 ;
        RECT 109.075 91.155 109.340 91.715 ;
        RECT 109.510 90.985 109.680 91.885 ;
        RECT 109.850 91.155 110.205 91.715 ;
        RECT 112.020 91.020 112.360 91.850 ;
        RECT 113.840 91.340 114.190 92.590 ;
        RECT 115.955 91.935 117.625 93.025 ;
        RECT 115.955 91.245 116.705 91.765 ;
        RECT 116.875 91.415 117.625 91.935 ;
        RECT 118.440 92.055 118.830 92.230 ;
        RECT 119.315 92.225 119.645 93.025 ;
        RECT 119.815 92.235 120.350 92.855 ;
        RECT 118.440 91.885 119.865 92.055 ;
        RECT 108.955 90.475 109.170 90.985 ;
        RECT 109.400 90.655 109.680 90.985 ;
        RECT 109.860 90.475 110.100 90.985 ;
        RECT 110.435 90.475 115.780 91.020 ;
        RECT 115.955 90.475 117.625 91.245 ;
        RECT 118.315 91.155 118.670 91.715 ;
        RECT 118.840 90.985 119.010 91.885 ;
        RECT 119.180 91.155 119.445 91.715 ;
        RECT 119.695 91.385 119.865 91.885 ;
        RECT 120.035 91.215 120.350 92.235 ;
        RECT 120.645 92.095 120.815 92.855 ;
        RECT 121.030 92.265 121.360 93.025 ;
        RECT 120.645 91.925 121.360 92.095 ;
        RECT 121.530 91.950 121.785 92.855 ;
        RECT 120.555 91.375 120.910 91.745 ;
        RECT 121.190 91.715 121.360 91.925 ;
        RECT 121.190 91.385 121.445 91.715 ;
        RECT 118.420 90.475 118.660 90.985 ;
        RECT 118.840 90.655 119.120 90.985 ;
        RECT 119.350 90.475 119.565 90.985 ;
        RECT 119.735 90.645 120.350 91.215 ;
        RECT 121.190 91.195 121.360 91.385 ;
        RECT 121.615 91.220 121.785 91.950 ;
        RECT 121.960 91.875 122.220 93.025 ;
        RECT 122.395 92.590 127.740 93.025 ;
        RECT 120.645 91.025 121.360 91.195 ;
        RECT 120.645 90.645 120.815 91.025 ;
        RECT 121.030 90.475 121.360 90.855 ;
        RECT 121.530 90.645 121.785 91.220 ;
        RECT 121.960 90.475 122.220 91.315 ;
        RECT 123.980 91.020 124.320 91.850 ;
        RECT 125.800 91.340 126.150 92.590 ;
        RECT 127.915 91.935 129.585 93.025 ;
        RECT 127.915 91.245 128.665 91.765 ;
        RECT 128.835 91.415 129.585 91.935 ;
        RECT 129.960 92.055 130.290 92.855 ;
        RECT 130.460 92.225 130.790 93.025 ;
        RECT 131.090 92.055 131.420 92.855 ;
        RECT 132.065 92.225 132.315 93.025 ;
        RECT 129.960 91.885 132.395 92.055 ;
        RECT 132.585 91.885 132.755 93.025 ;
        RECT 132.925 91.885 133.265 92.855 ;
        RECT 129.755 91.465 130.105 91.715 ;
        RECT 130.290 91.255 130.460 91.885 ;
        RECT 130.630 91.465 130.960 91.665 ;
        RECT 131.130 91.465 131.460 91.665 ;
        RECT 131.630 91.465 132.050 91.665 ;
        RECT 132.225 91.635 132.395 91.885 ;
        RECT 132.225 91.465 132.920 91.635 ;
        RECT 133.090 91.325 133.265 91.885 ;
        RECT 133.435 91.860 133.725 93.025 ;
        RECT 133.985 92.355 134.155 92.855 ;
        RECT 134.325 92.525 134.655 93.025 ;
        RECT 133.985 92.185 134.650 92.355 ;
        RECT 133.900 91.365 134.250 92.015 ;
        RECT 122.395 90.475 127.740 91.020 ;
        RECT 127.915 90.475 129.585 91.245 ;
        RECT 129.960 90.645 130.460 91.255 ;
        RECT 131.090 91.125 132.315 91.295 ;
        RECT 133.035 91.275 133.265 91.325 ;
        RECT 131.090 90.645 131.420 91.125 ;
        RECT 131.590 90.475 131.815 90.935 ;
        RECT 131.985 90.645 132.315 91.125 ;
        RECT 132.505 90.475 132.755 91.275 ;
        RECT 132.925 90.645 133.265 91.275 ;
        RECT 133.435 90.475 133.725 91.200 ;
        RECT 134.420 91.195 134.650 92.185 ;
        RECT 133.985 91.025 134.650 91.195 ;
        RECT 133.985 90.735 134.155 91.025 ;
        RECT 134.325 90.475 134.655 90.855 ;
        RECT 134.825 90.735 135.010 92.855 ;
        RECT 135.250 92.565 135.515 93.025 ;
        RECT 135.685 92.430 135.935 92.855 ;
        RECT 136.145 92.580 137.250 92.750 ;
        RECT 135.630 92.300 135.935 92.430 ;
        RECT 135.180 91.105 135.460 92.055 ;
        RECT 135.630 91.195 135.800 92.300 ;
        RECT 135.970 91.515 136.210 92.110 ;
        RECT 136.380 92.045 136.910 92.410 ;
        RECT 136.380 91.345 136.550 92.045 ;
        RECT 137.080 91.965 137.250 92.580 ;
        RECT 137.420 92.225 137.590 93.025 ;
        RECT 137.760 92.525 138.010 92.855 ;
        RECT 138.235 92.555 139.120 92.725 ;
        RECT 137.080 91.875 137.590 91.965 ;
        RECT 135.630 91.065 135.855 91.195 ;
        RECT 136.025 91.125 136.550 91.345 ;
        RECT 136.720 91.705 137.590 91.875 ;
        RECT 135.265 90.475 135.515 90.935 ;
        RECT 135.685 90.925 135.855 91.065 ;
        RECT 136.720 90.925 136.890 91.705 ;
        RECT 137.420 91.635 137.590 91.705 ;
        RECT 137.100 91.455 137.300 91.485 ;
        RECT 137.760 91.455 137.930 92.525 ;
        RECT 138.100 91.635 138.290 92.355 ;
        RECT 137.100 91.155 137.930 91.455 ;
        RECT 138.460 91.425 138.780 92.385 ;
        RECT 135.685 90.755 136.020 90.925 ;
        RECT 136.215 90.755 136.890 90.925 ;
        RECT 137.210 90.475 137.580 90.975 ;
        RECT 137.760 90.925 137.930 91.155 ;
        RECT 138.315 91.095 138.780 91.425 ;
        RECT 138.950 91.715 139.120 92.555 ;
        RECT 139.300 92.525 139.615 93.025 ;
        RECT 139.845 92.295 140.185 92.855 ;
        RECT 139.290 91.920 140.185 92.295 ;
        RECT 140.355 92.015 140.525 93.025 ;
        RECT 139.995 91.715 140.185 91.920 ;
        RECT 140.695 91.965 141.025 92.810 ;
        RECT 140.695 91.885 141.085 91.965 ;
        RECT 140.870 91.835 141.085 91.885 ;
        RECT 138.950 91.385 139.825 91.715 ;
        RECT 139.995 91.385 140.745 91.715 ;
        RECT 138.950 90.925 139.120 91.385 ;
        RECT 139.995 91.215 140.195 91.385 ;
        RECT 140.915 91.255 141.085 91.835 ;
        RECT 141.715 91.935 142.925 93.025 ;
        RECT 141.715 91.395 142.235 91.935 ;
        RECT 140.860 91.215 141.085 91.255 ;
        RECT 142.405 91.225 142.925 91.765 ;
        RECT 137.760 90.755 138.165 90.925 ;
        RECT 138.335 90.755 139.120 90.925 ;
        RECT 139.395 90.475 139.605 91.005 ;
        RECT 139.865 90.690 140.195 91.215 ;
        RECT 140.705 91.130 141.085 91.215 ;
        RECT 140.365 90.475 140.535 91.085 ;
        RECT 140.705 90.695 141.035 91.130 ;
        RECT 141.715 90.475 142.925 91.225 ;
        RECT 17.430 90.305 143.010 90.475 ;
        RECT 17.515 89.555 18.725 90.305 ;
        RECT 18.895 89.760 24.240 90.305 ;
        RECT 24.415 89.760 29.760 90.305 ;
        RECT 29.935 89.760 35.280 90.305 ;
        RECT 35.455 89.760 40.800 90.305 ;
        RECT 17.515 89.015 18.035 89.555 ;
        RECT 18.205 88.845 18.725 89.385 ;
        RECT 20.480 88.930 20.820 89.760 ;
        RECT 17.515 87.755 18.725 88.845 ;
        RECT 22.300 88.190 22.650 89.440 ;
        RECT 26.000 88.930 26.340 89.760 ;
        RECT 27.820 88.190 28.170 89.440 ;
        RECT 31.520 88.930 31.860 89.760 ;
        RECT 33.340 88.190 33.690 89.440 ;
        RECT 37.040 88.930 37.380 89.760 ;
        RECT 40.975 89.535 42.645 90.305 ;
        RECT 43.275 89.580 43.565 90.305 ;
        RECT 43.735 89.760 49.080 90.305 ;
        RECT 49.255 89.760 54.600 90.305 ;
        RECT 54.775 89.760 60.120 90.305 ;
        RECT 60.295 89.760 65.640 90.305 ;
        RECT 38.860 88.190 39.210 89.440 ;
        RECT 40.975 89.015 41.725 89.535 ;
        RECT 41.895 88.845 42.645 89.365 ;
        RECT 45.320 88.930 45.660 89.760 ;
        RECT 18.895 87.755 24.240 88.190 ;
        RECT 24.415 87.755 29.760 88.190 ;
        RECT 29.935 87.755 35.280 88.190 ;
        RECT 35.455 87.755 40.800 88.190 ;
        RECT 40.975 87.755 42.645 88.845 ;
        RECT 43.275 87.755 43.565 88.920 ;
        RECT 47.140 88.190 47.490 89.440 ;
        RECT 50.840 88.930 51.180 89.760 ;
        RECT 52.660 88.190 53.010 89.440 ;
        RECT 56.360 88.930 56.700 89.760 ;
        RECT 58.180 88.190 58.530 89.440 ;
        RECT 61.880 88.930 62.220 89.760 ;
        RECT 65.815 89.535 68.405 90.305 ;
        RECT 69.035 89.580 69.325 90.305 ;
        RECT 69.495 89.760 74.840 90.305 ;
        RECT 63.700 88.190 64.050 89.440 ;
        RECT 65.815 89.015 67.025 89.535 ;
        RECT 67.195 88.845 68.405 89.365 ;
        RECT 71.080 88.930 71.420 89.760 ;
        RECT 75.105 89.755 75.275 90.045 ;
        RECT 75.445 89.925 75.775 90.305 ;
        RECT 75.105 89.585 75.770 89.755 ;
        RECT 43.735 87.755 49.080 88.190 ;
        RECT 49.255 87.755 54.600 88.190 ;
        RECT 54.775 87.755 60.120 88.190 ;
        RECT 60.295 87.755 65.640 88.190 ;
        RECT 65.815 87.755 68.405 88.845 ;
        RECT 69.035 87.755 69.325 88.920 ;
        RECT 72.900 88.190 73.250 89.440 ;
        RECT 75.020 88.765 75.370 89.415 ;
        RECT 75.540 88.595 75.770 89.585 ;
        RECT 75.105 88.425 75.770 88.595 ;
        RECT 69.495 87.755 74.840 88.190 ;
        RECT 75.105 87.925 75.275 88.425 ;
        RECT 75.445 87.755 75.775 88.255 ;
        RECT 75.945 87.925 76.130 90.045 ;
        RECT 76.385 89.845 76.635 90.305 ;
        RECT 76.805 89.855 77.140 90.025 ;
        RECT 77.335 89.855 78.010 90.025 ;
        RECT 76.805 89.715 76.975 89.855 ;
        RECT 76.300 88.725 76.580 89.675 ;
        RECT 76.750 89.585 76.975 89.715 ;
        RECT 76.750 88.480 76.920 89.585 ;
        RECT 77.145 89.435 77.670 89.655 ;
        RECT 77.090 88.670 77.330 89.265 ;
        RECT 77.500 88.735 77.670 89.435 ;
        RECT 77.840 89.075 78.010 89.855 ;
        RECT 78.330 89.805 78.700 90.305 ;
        RECT 78.880 89.855 79.285 90.025 ;
        RECT 79.455 89.855 80.240 90.025 ;
        RECT 78.880 89.625 79.050 89.855 ;
        RECT 78.220 89.325 79.050 89.625 ;
        RECT 79.435 89.355 79.900 89.685 ;
        RECT 78.220 89.295 78.420 89.325 ;
        RECT 78.540 89.075 78.710 89.145 ;
        RECT 77.840 88.905 78.710 89.075 ;
        RECT 78.200 88.815 78.710 88.905 ;
        RECT 76.750 88.350 77.055 88.480 ;
        RECT 77.500 88.370 78.030 88.735 ;
        RECT 76.370 87.755 76.635 88.215 ;
        RECT 76.805 87.925 77.055 88.350 ;
        RECT 78.200 88.200 78.370 88.815 ;
        RECT 77.265 88.030 78.370 88.200 ;
        RECT 78.540 87.755 78.710 88.555 ;
        RECT 78.880 88.255 79.050 89.325 ;
        RECT 79.220 88.425 79.410 89.145 ;
        RECT 79.580 88.395 79.900 89.355 ;
        RECT 80.070 89.395 80.240 89.855 ;
        RECT 80.515 89.775 80.725 90.305 ;
        RECT 80.985 89.565 81.315 90.090 ;
        RECT 81.485 89.695 81.655 90.305 ;
        RECT 81.825 89.650 82.155 90.085 ;
        RECT 81.825 89.565 82.205 89.650 ;
        RECT 81.115 89.395 81.315 89.565 ;
        RECT 81.980 89.525 82.205 89.565 ;
        RECT 80.070 89.065 80.945 89.395 ;
        RECT 81.115 89.065 81.865 89.395 ;
        RECT 78.880 87.925 79.130 88.255 ;
        RECT 80.070 88.225 80.240 89.065 ;
        RECT 81.115 88.860 81.305 89.065 ;
        RECT 82.035 88.945 82.205 89.525 ;
        RECT 82.375 89.555 83.585 90.305 ;
        RECT 82.375 89.015 82.895 89.555 ;
        RECT 83.755 89.505 84.095 90.135 ;
        RECT 84.265 89.505 84.515 90.305 ;
        RECT 84.705 89.655 85.035 90.135 ;
        RECT 85.205 89.845 85.430 90.305 ;
        RECT 85.600 89.655 85.930 90.135 ;
        RECT 81.990 88.895 82.205 88.945 ;
        RECT 80.410 88.485 81.305 88.860 ;
        RECT 81.815 88.815 82.205 88.895 ;
        RECT 83.065 88.845 83.585 89.385 ;
        RECT 79.355 88.055 80.240 88.225 ;
        RECT 80.420 87.755 80.735 88.255 ;
        RECT 80.965 87.925 81.305 88.485 ;
        RECT 81.475 87.755 81.645 88.765 ;
        RECT 81.815 87.970 82.145 88.815 ;
        RECT 82.375 87.755 83.585 88.845 ;
        RECT 83.755 88.895 83.930 89.505 ;
        RECT 84.705 89.485 85.930 89.655 ;
        RECT 86.560 89.525 87.060 90.135 ;
        RECT 84.100 89.145 84.795 89.315 ;
        RECT 84.625 88.895 84.795 89.145 ;
        RECT 84.970 89.115 85.390 89.315 ;
        RECT 85.560 89.115 85.890 89.315 ;
        RECT 86.060 89.115 86.390 89.315 ;
        RECT 86.560 88.895 86.730 89.525 ;
        RECT 87.435 89.505 87.775 90.135 ;
        RECT 87.945 89.505 88.195 90.305 ;
        RECT 88.385 89.655 88.715 90.135 ;
        RECT 88.885 89.845 89.110 90.305 ;
        RECT 89.280 89.655 89.610 90.135 ;
        RECT 86.915 89.065 87.265 89.315 ;
        RECT 87.435 88.895 87.610 89.505 ;
        RECT 88.385 89.485 89.610 89.655 ;
        RECT 90.240 89.525 90.740 90.135 ;
        RECT 91.115 89.805 91.375 90.135 ;
        RECT 91.545 89.945 91.875 90.305 ;
        RECT 92.130 89.925 93.430 90.135 ;
        RECT 87.780 89.145 88.475 89.315 ;
        RECT 88.305 88.895 88.475 89.145 ;
        RECT 88.650 89.115 89.070 89.315 ;
        RECT 89.240 89.115 89.570 89.315 ;
        RECT 89.740 89.115 90.070 89.315 ;
        RECT 90.240 88.895 90.410 89.525 ;
        RECT 90.595 89.065 90.945 89.315 ;
        RECT 83.755 87.925 84.095 88.895 ;
        RECT 84.265 87.755 84.435 88.895 ;
        RECT 84.625 88.725 87.060 88.895 ;
        RECT 84.705 87.755 84.955 88.555 ;
        RECT 85.600 87.925 85.930 88.725 ;
        RECT 86.230 87.755 86.560 88.555 ;
        RECT 86.730 87.925 87.060 88.725 ;
        RECT 87.435 87.925 87.775 88.895 ;
        RECT 87.945 87.755 88.115 88.895 ;
        RECT 88.305 88.725 90.740 88.895 ;
        RECT 88.385 87.755 88.635 88.555 ;
        RECT 89.280 87.925 89.610 88.725 ;
        RECT 89.910 87.755 90.240 88.555 ;
        RECT 90.410 87.925 90.740 88.725 ;
        RECT 91.115 88.605 91.285 89.805 ;
        RECT 92.130 89.775 92.300 89.925 ;
        RECT 91.545 89.650 92.300 89.775 ;
        RECT 91.455 89.605 92.300 89.650 ;
        RECT 91.455 89.485 91.725 89.605 ;
        RECT 91.455 88.910 91.625 89.485 ;
        RECT 91.855 89.045 92.265 89.350 ;
        RECT 92.555 89.315 92.765 89.715 ;
        RECT 92.435 89.105 92.765 89.315 ;
        RECT 93.010 89.315 93.230 89.715 ;
        RECT 93.705 89.540 94.160 90.305 ;
        RECT 94.795 89.580 95.085 90.305 ;
        RECT 95.420 89.795 95.660 90.305 ;
        RECT 95.840 89.795 96.120 90.125 ;
        RECT 96.350 89.795 96.565 90.305 ;
        RECT 93.010 89.105 93.485 89.315 ;
        RECT 93.675 89.115 94.165 89.315 ;
        RECT 95.315 89.065 95.670 89.625 ;
        RECT 91.455 88.875 91.655 88.910 ;
        RECT 92.985 88.875 94.160 88.935 ;
        RECT 91.455 88.765 94.160 88.875 ;
        RECT 91.515 88.705 93.315 88.765 ;
        RECT 92.985 88.675 93.315 88.705 ;
        RECT 91.115 87.925 91.375 88.605 ;
        RECT 91.545 87.755 91.795 88.535 ;
        RECT 92.045 88.505 92.880 88.515 ;
        RECT 93.470 88.505 93.655 88.595 ;
        RECT 92.045 88.305 93.655 88.505 ;
        RECT 92.045 87.925 92.295 88.305 ;
        RECT 93.425 88.265 93.655 88.305 ;
        RECT 93.905 88.145 94.160 88.765 ;
        RECT 92.465 87.755 92.820 88.135 ;
        RECT 93.825 87.925 94.160 88.145 ;
        RECT 94.795 87.755 95.085 88.920 ;
        RECT 95.840 88.895 96.010 89.795 ;
        RECT 96.180 89.065 96.445 89.625 ;
        RECT 96.735 89.565 97.350 90.135 ;
        RECT 96.695 88.895 96.865 89.395 ;
        RECT 95.440 88.725 96.865 88.895 ;
        RECT 95.440 88.550 95.830 88.725 ;
        RECT 96.315 87.755 96.645 88.555 ;
        RECT 97.035 88.545 97.350 89.565 ;
        RECT 97.760 89.525 98.260 90.135 ;
        RECT 97.555 89.065 97.905 89.315 ;
        RECT 98.090 88.895 98.260 89.525 ;
        RECT 98.890 89.655 99.220 90.135 ;
        RECT 99.390 89.845 99.615 90.305 ;
        RECT 99.785 89.655 100.115 90.135 ;
        RECT 98.890 89.485 100.115 89.655 ;
        RECT 100.305 89.505 100.555 90.305 ;
        RECT 100.725 89.505 101.065 90.135 ;
        RECT 98.430 89.115 98.760 89.315 ;
        RECT 98.930 89.115 99.260 89.315 ;
        RECT 99.430 89.115 99.850 89.315 ;
        RECT 100.025 89.145 100.720 89.315 ;
        RECT 100.025 88.895 100.195 89.145 ;
        RECT 100.890 88.895 101.065 89.505 ;
        RECT 101.235 89.555 102.445 90.305 ;
        RECT 102.705 89.755 102.875 90.045 ;
        RECT 103.045 89.925 103.375 90.305 ;
        RECT 102.705 89.585 103.370 89.755 ;
        RECT 101.235 89.015 101.755 89.555 ;
        RECT 96.815 87.925 97.350 88.545 ;
        RECT 97.760 88.725 100.195 88.895 ;
        RECT 97.760 87.925 98.090 88.725 ;
        RECT 98.260 87.755 98.590 88.555 ;
        RECT 98.890 87.925 99.220 88.725 ;
        RECT 99.865 87.755 100.115 88.555 ;
        RECT 100.385 87.755 100.555 88.895 ;
        RECT 100.725 87.925 101.065 88.895 ;
        RECT 101.925 88.845 102.445 89.385 ;
        RECT 101.235 87.755 102.445 88.845 ;
        RECT 102.620 88.765 102.970 89.415 ;
        RECT 103.140 88.595 103.370 89.585 ;
        RECT 102.705 88.425 103.370 88.595 ;
        RECT 102.705 87.925 102.875 88.425 ;
        RECT 103.045 87.755 103.375 88.255 ;
        RECT 103.545 87.925 103.730 90.045 ;
        RECT 103.985 89.845 104.235 90.305 ;
        RECT 104.405 89.855 104.740 90.025 ;
        RECT 104.935 89.855 105.610 90.025 ;
        RECT 104.405 89.715 104.575 89.855 ;
        RECT 103.900 88.725 104.180 89.675 ;
        RECT 104.350 89.585 104.575 89.715 ;
        RECT 104.350 88.480 104.520 89.585 ;
        RECT 104.745 89.435 105.270 89.655 ;
        RECT 104.690 88.670 104.930 89.265 ;
        RECT 105.100 88.735 105.270 89.435 ;
        RECT 105.440 89.075 105.610 89.855 ;
        RECT 105.930 89.805 106.300 90.305 ;
        RECT 106.480 89.855 106.885 90.025 ;
        RECT 107.055 89.855 107.840 90.025 ;
        RECT 106.480 89.625 106.650 89.855 ;
        RECT 105.820 89.325 106.650 89.625 ;
        RECT 107.035 89.355 107.500 89.685 ;
        RECT 105.820 89.295 106.020 89.325 ;
        RECT 106.140 89.075 106.310 89.145 ;
        RECT 105.440 88.905 106.310 89.075 ;
        RECT 105.800 88.815 106.310 88.905 ;
        RECT 104.350 88.350 104.655 88.480 ;
        RECT 105.100 88.370 105.630 88.735 ;
        RECT 103.970 87.755 104.235 88.215 ;
        RECT 104.405 87.925 104.655 88.350 ;
        RECT 105.800 88.200 105.970 88.815 ;
        RECT 104.865 88.030 105.970 88.200 ;
        RECT 106.140 87.755 106.310 88.555 ;
        RECT 106.480 88.255 106.650 89.325 ;
        RECT 106.820 88.425 107.010 89.145 ;
        RECT 107.180 88.395 107.500 89.355 ;
        RECT 107.670 89.395 107.840 89.855 ;
        RECT 108.115 89.775 108.325 90.305 ;
        RECT 108.585 89.565 108.915 90.090 ;
        RECT 109.085 89.695 109.255 90.305 ;
        RECT 109.425 89.650 109.755 90.085 ;
        RECT 109.425 89.565 109.805 89.650 ;
        RECT 108.715 89.395 108.915 89.565 ;
        RECT 109.580 89.525 109.805 89.565 ;
        RECT 107.670 89.065 108.545 89.395 ;
        RECT 108.715 89.065 109.465 89.395 ;
        RECT 106.480 87.925 106.730 88.255 ;
        RECT 107.670 88.225 107.840 89.065 ;
        RECT 108.715 88.860 108.905 89.065 ;
        RECT 109.635 88.945 109.805 89.525 ;
        RECT 109.590 88.895 109.805 88.945 ;
        RECT 108.010 88.485 108.905 88.860 ;
        RECT 109.415 88.815 109.805 88.895 ;
        RECT 109.975 89.505 110.315 90.135 ;
        RECT 110.485 89.505 110.735 90.305 ;
        RECT 110.925 89.655 111.255 90.135 ;
        RECT 111.425 89.845 111.650 90.305 ;
        RECT 111.820 89.655 112.150 90.135 ;
        RECT 109.975 88.895 110.150 89.505 ;
        RECT 110.925 89.485 112.150 89.655 ;
        RECT 112.780 89.525 113.280 90.135 ;
        RECT 113.660 89.540 114.115 90.305 ;
        RECT 114.390 89.925 115.690 90.135 ;
        RECT 115.945 89.945 116.275 90.305 ;
        RECT 115.520 89.775 115.690 89.925 ;
        RECT 116.445 89.805 116.705 90.135 ;
        RECT 110.320 89.145 111.015 89.315 ;
        RECT 110.845 88.895 111.015 89.145 ;
        RECT 111.190 89.115 111.610 89.315 ;
        RECT 111.780 89.115 112.110 89.315 ;
        RECT 112.280 89.115 112.610 89.315 ;
        RECT 112.780 88.895 112.950 89.525 ;
        RECT 114.590 89.315 114.810 89.715 ;
        RECT 113.135 89.065 113.485 89.315 ;
        RECT 113.655 89.115 114.145 89.315 ;
        RECT 114.335 89.105 114.810 89.315 ;
        RECT 115.055 89.315 115.265 89.715 ;
        RECT 115.520 89.650 116.275 89.775 ;
        RECT 115.520 89.605 116.365 89.650 ;
        RECT 116.095 89.485 116.365 89.605 ;
        RECT 115.055 89.105 115.385 89.315 ;
        RECT 115.555 89.045 115.965 89.350 ;
        RECT 106.955 88.055 107.840 88.225 ;
        RECT 108.020 87.755 108.335 88.255 ;
        RECT 108.565 87.925 108.905 88.485 ;
        RECT 109.075 87.755 109.245 88.765 ;
        RECT 109.415 87.970 109.745 88.815 ;
        RECT 109.975 87.925 110.315 88.895 ;
        RECT 110.485 87.755 110.655 88.895 ;
        RECT 110.845 88.725 113.280 88.895 ;
        RECT 110.925 87.755 111.175 88.555 ;
        RECT 111.820 87.925 112.150 88.725 ;
        RECT 112.450 87.755 112.780 88.555 ;
        RECT 112.950 87.925 113.280 88.725 ;
        RECT 113.660 88.875 114.835 88.935 ;
        RECT 116.195 88.910 116.365 89.485 ;
        RECT 116.165 88.875 116.365 88.910 ;
        RECT 113.660 88.765 116.365 88.875 ;
        RECT 113.660 88.145 113.915 88.765 ;
        RECT 114.505 88.705 116.305 88.765 ;
        RECT 114.505 88.675 114.835 88.705 ;
        RECT 116.535 88.605 116.705 89.805 ;
        RECT 116.875 89.555 118.085 90.305 ;
        RECT 118.420 89.795 118.660 90.305 ;
        RECT 118.840 89.795 119.120 90.125 ;
        RECT 119.350 89.795 119.565 90.305 ;
        RECT 116.875 89.015 117.395 89.555 ;
        RECT 117.565 88.845 118.085 89.385 ;
        RECT 118.315 89.065 118.670 89.625 ;
        RECT 118.840 88.895 119.010 89.795 ;
        RECT 119.180 89.065 119.445 89.625 ;
        RECT 119.735 89.565 120.350 90.135 ;
        RECT 120.555 89.580 120.845 90.305 ;
        RECT 119.695 88.895 119.865 89.395 ;
        RECT 114.165 88.505 114.350 88.595 ;
        RECT 114.940 88.505 115.775 88.515 ;
        RECT 114.165 88.305 115.775 88.505 ;
        RECT 114.165 88.265 114.395 88.305 ;
        RECT 113.660 87.925 113.995 88.145 ;
        RECT 115.000 87.755 115.355 88.135 ;
        RECT 115.525 87.925 115.775 88.305 ;
        RECT 116.025 87.755 116.275 88.535 ;
        RECT 116.445 87.925 116.705 88.605 ;
        RECT 116.875 87.755 118.085 88.845 ;
        RECT 118.440 88.725 119.865 88.895 ;
        RECT 118.440 88.550 118.830 88.725 ;
        RECT 119.315 87.755 119.645 88.555 ;
        RECT 120.035 88.545 120.350 89.565 ;
        RECT 121.220 89.525 121.720 90.135 ;
        RECT 121.015 89.065 121.365 89.315 ;
        RECT 119.815 87.925 120.350 88.545 ;
        RECT 120.555 87.755 120.845 88.920 ;
        RECT 121.550 88.895 121.720 89.525 ;
        RECT 122.350 89.655 122.680 90.135 ;
        RECT 122.850 89.845 123.075 90.305 ;
        RECT 123.245 89.655 123.575 90.135 ;
        RECT 122.350 89.485 123.575 89.655 ;
        RECT 123.765 89.505 124.015 90.305 ;
        RECT 124.185 89.505 124.525 90.135 ;
        RECT 121.890 89.115 122.220 89.315 ;
        RECT 122.390 89.115 122.720 89.315 ;
        RECT 122.890 89.115 123.310 89.315 ;
        RECT 123.485 89.145 124.180 89.315 ;
        RECT 123.485 88.895 123.655 89.145 ;
        RECT 124.350 88.895 124.525 89.505 ;
        RECT 121.220 88.725 123.655 88.895 ;
        RECT 121.220 87.925 121.550 88.725 ;
        RECT 121.720 87.755 122.050 88.555 ;
        RECT 122.350 87.925 122.680 88.725 ;
        RECT 123.325 87.755 123.575 88.555 ;
        RECT 123.845 87.755 124.015 88.895 ;
        RECT 124.185 87.925 124.525 88.895 ;
        RECT 125.155 89.505 125.495 90.135 ;
        RECT 125.665 89.505 125.915 90.305 ;
        RECT 126.105 89.655 126.435 90.135 ;
        RECT 126.605 89.845 126.830 90.305 ;
        RECT 127.000 89.655 127.330 90.135 ;
        RECT 125.155 88.895 125.330 89.505 ;
        RECT 126.105 89.485 127.330 89.655 ;
        RECT 127.960 89.525 128.460 90.135 ;
        RECT 129.345 89.650 129.675 90.085 ;
        RECT 129.845 89.695 130.015 90.305 ;
        RECT 129.295 89.565 129.675 89.650 ;
        RECT 130.185 89.565 130.515 90.090 ;
        RECT 130.775 89.775 130.985 90.305 ;
        RECT 131.260 89.855 132.045 90.025 ;
        RECT 132.215 89.855 132.620 90.025 ;
        RECT 129.295 89.525 129.520 89.565 ;
        RECT 125.500 89.145 126.195 89.315 ;
        RECT 126.025 88.895 126.195 89.145 ;
        RECT 126.370 89.115 126.790 89.315 ;
        RECT 126.960 89.115 127.290 89.315 ;
        RECT 127.460 89.115 127.790 89.315 ;
        RECT 127.960 88.895 128.130 89.525 ;
        RECT 128.315 89.065 128.665 89.315 ;
        RECT 129.295 88.945 129.465 89.525 ;
        RECT 130.185 89.395 130.385 89.565 ;
        RECT 131.260 89.395 131.430 89.855 ;
        RECT 129.635 89.065 130.385 89.395 ;
        RECT 130.555 89.065 131.430 89.395 ;
        RECT 129.295 88.895 129.510 88.945 ;
        RECT 125.155 87.925 125.495 88.895 ;
        RECT 125.665 87.755 125.835 88.895 ;
        RECT 126.025 88.725 128.460 88.895 ;
        RECT 129.295 88.815 129.685 88.895 ;
        RECT 126.105 87.755 126.355 88.555 ;
        RECT 127.000 87.925 127.330 88.725 ;
        RECT 127.630 87.755 127.960 88.555 ;
        RECT 128.130 87.925 128.460 88.725 ;
        RECT 129.355 87.970 129.685 88.815 ;
        RECT 130.195 88.860 130.385 89.065 ;
        RECT 129.855 87.755 130.025 88.765 ;
        RECT 130.195 88.485 131.090 88.860 ;
        RECT 130.195 87.925 130.535 88.485 ;
        RECT 130.765 87.755 131.080 88.255 ;
        RECT 131.260 88.225 131.430 89.065 ;
        RECT 131.600 89.355 132.065 89.685 ;
        RECT 132.450 89.625 132.620 89.855 ;
        RECT 132.800 89.805 133.170 90.305 ;
        RECT 133.490 89.855 134.165 90.025 ;
        RECT 134.360 89.855 134.695 90.025 ;
        RECT 131.600 88.395 131.920 89.355 ;
        RECT 132.450 89.325 133.280 89.625 ;
        RECT 132.090 88.425 132.280 89.145 ;
        RECT 132.450 88.255 132.620 89.325 ;
        RECT 133.080 89.295 133.280 89.325 ;
        RECT 132.790 89.075 132.960 89.145 ;
        RECT 133.490 89.075 133.660 89.855 ;
        RECT 134.525 89.715 134.695 89.855 ;
        RECT 134.865 89.845 135.115 90.305 ;
        RECT 132.790 88.905 133.660 89.075 ;
        RECT 133.830 89.435 134.355 89.655 ;
        RECT 134.525 89.585 134.750 89.715 ;
        RECT 132.790 88.815 133.300 88.905 ;
        RECT 131.260 88.055 132.145 88.225 ;
        RECT 132.370 87.925 132.620 88.255 ;
        RECT 132.790 87.755 132.960 88.555 ;
        RECT 133.130 88.200 133.300 88.815 ;
        RECT 133.830 88.735 134.000 89.435 ;
        RECT 133.470 88.370 134.000 88.735 ;
        RECT 134.170 88.670 134.410 89.265 ;
        RECT 134.580 88.480 134.750 89.585 ;
        RECT 134.920 88.725 135.200 89.675 ;
        RECT 134.445 88.350 134.750 88.480 ;
        RECT 133.130 88.030 134.235 88.200 ;
        RECT 134.445 87.925 134.695 88.350 ;
        RECT 134.865 87.755 135.130 88.215 ;
        RECT 135.370 87.925 135.555 90.045 ;
        RECT 135.725 89.925 136.055 90.305 ;
        RECT 136.225 89.755 136.395 90.045 ;
        RECT 135.730 89.585 136.395 89.755 ;
        RECT 135.730 88.595 135.960 89.585 ;
        RECT 136.655 89.555 137.865 90.305 ;
        RECT 138.125 89.755 138.295 90.135 ;
        RECT 138.510 89.925 138.840 90.305 ;
        RECT 138.125 89.585 138.840 89.755 ;
        RECT 136.130 88.765 136.480 89.415 ;
        RECT 136.655 89.015 137.175 89.555 ;
        RECT 137.345 88.845 137.865 89.385 ;
        RECT 138.035 89.035 138.390 89.405 ;
        RECT 138.670 89.395 138.840 89.585 ;
        RECT 139.010 89.560 139.265 90.135 ;
        RECT 138.670 89.065 138.925 89.395 ;
        RECT 138.670 88.855 138.840 89.065 ;
        RECT 135.730 88.425 136.395 88.595 ;
        RECT 135.725 87.755 136.055 88.255 ;
        RECT 136.225 87.925 136.395 88.425 ;
        RECT 136.655 87.755 137.865 88.845 ;
        RECT 138.125 88.685 138.840 88.855 ;
        RECT 139.095 88.830 139.265 89.560 ;
        RECT 139.440 89.465 139.700 90.305 ;
        RECT 139.965 89.755 140.135 90.135 ;
        RECT 140.350 89.925 140.680 90.305 ;
        RECT 139.965 89.585 140.680 89.755 ;
        RECT 139.875 89.035 140.230 89.405 ;
        RECT 140.510 89.395 140.680 89.585 ;
        RECT 140.850 89.560 141.105 90.135 ;
        RECT 140.510 89.065 140.765 89.395 ;
        RECT 138.125 87.925 138.295 88.685 ;
        RECT 138.510 87.755 138.840 88.515 ;
        RECT 139.010 87.925 139.265 88.830 ;
        RECT 139.440 87.755 139.700 88.905 ;
        RECT 140.510 88.855 140.680 89.065 ;
        RECT 139.965 88.685 140.680 88.855 ;
        RECT 140.935 88.830 141.105 89.560 ;
        RECT 141.280 89.465 141.540 90.305 ;
        RECT 141.715 89.555 142.925 90.305 ;
        RECT 139.965 87.925 140.135 88.685 ;
        RECT 140.350 87.755 140.680 88.515 ;
        RECT 140.850 87.925 141.105 88.830 ;
        RECT 141.280 87.755 141.540 88.905 ;
        RECT 141.715 88.845 142.235 89.385 ;
        RECT 142.405 89.015 142.925 89.555 ;
        RECT 141.715 87.755 142.925 88.845 ;
        RECT 17.430 87.585 143.010 87.755 ;
        RECT 17.515 86.495 18.725 87.585 ;
        RECT 18.895 87.150 24.240 87.585 ;
        RECT 24.415 87.150 29.760 87.585 ;
        RECT 17.515 85.785 18.035 86.325 ;
        RECT 18.205 85.955 18.725 86.495 ;
        RECT 17.515 85.035 18.725 85.785 ;
        RECT 20.480 85.580 20.820 86.410 ;
        RECT 22.300 85.900 22.650 87.150 ;
        RECT 26.000 85.580 26.340 86.410 ;
        RECT 27.820 85.900 28.170 87.150 ;
        RECT 30.395 86.420 30.685 87.585 ;
        RECT 30.855 87.150 36.200 87.585 ;
        RECT 36.375 87.150 41.720 87.585 ;
        RECT 41.895 87.150 47.240 87.585 ;
        RECT 47.415 87.150 52.760 87.585 ;
        RECT 18.895 85.035 24.240 85.580 ;
        RECT 24.415 85.035 29.760 85.580 ;
        RECT 30.395 85.035 30.685 85.760 ;
        RECT 32.440 85.580 32.780 86.410 ;
        RECT 34.260 85.900 34.610 87.150 ;
        RECT 37.960 85.580 38.300 86.410 ;
        RECT 39.780 85.900 40.130 87.150 ;
        RECT 43.480 85.580 43.820 86.410 ;
        RECT 45.300 85.900 45.650 87.150 ;
        RECT 49.000 85.580 49.340 86.410 ;
        RECT 50.820 85.900 51.170 87.150 ;
        RECT 52.935 86.495 55.525 87.585 ;
        RECT 52.935 85.805 54.145 86.325 ;
        RECT 54.315 85.975 55.525 86.495 ;
        RECT 56.155 86.420 56.445 87.585 ;
        RECT 56.615 87.150 61.960 87.585 ;
        RECT 62.135 87.150 67.480 87.585 ;
        RECT 67.655 87.150 73.000 87.585 ;
        RECT 73.175 87.150 78.520 87.585 ;
        RECT 30.855 85.035 36.200 85.580 ;
        RECT 36.375 85.035 41.720 85.580 ;
        RECT 41.895 85.035 47.240 85.580 ;
        RECT 47.415 85.035 52.760 85.580 ;
        RECT 52.935 85.035 55.525 85.805 ;
        RECT 56.155 85.035 56.445 85.760 ;
        RECT 58.200 85.580 58.540 86.410 ;
        RECT 60.020 85.900 60.370 87.150 ;
        RECT 63.720 85.580 64.060 86.410 ;
        RECT 65.540 85.900 65.890 87.150 ;
        RECT 69.240 85.580 69.580 86.410 ;
        RECT 71.060 85.900 71.410 87.150 ;
        RECT 74.760 85.580 75.100 86.410 ;
        RECT 76.580 85.900 76.930 87.150 ;
        RECT 78.695 86.495 81.285 87.585 ;
        RECT 78.695 85.805 79.905 86.325 ;
        RECT 80.075 85.975 81.285 86.495 ;
        RECT 81.915 86.420 82.205 87.585 ;
        RECT 82.465 86.915 82.635 87.415 ;
        RECT 82.805 87.085 83.135 87.585 ;
        RECT 82.465 86.745 83.130 86.915 ;
        RECT 82.380 85.925 82.730 86.575 ;
        RECT 56.615 85.035 61.960 85.580 ;
        RECT 62.135 85.035 67.480 85.580 ;
        RECT 67.655 85.035 73.000 85.580 ;
        RECT 73.175 85.035 78.520 85.580 ;
        RECT 78.695 85.035 81.285 85.805 ;
        RECT 81.915 85.035 82.205 85.760 ;
        RECT 82.900 85.755 83.130 86.745 ;
        RECT 82.465 85.585 83.130 85.755 ;
        RECT 82.465 85.295 82.635 85.585 ;
        RECT 82.805 85.035 83.135 85.415 ;
        RECT 83.305 85.295 83.490 87.415 ;
        RECT 83.730 87.125 83.995 87.585 ;
        RECT 84.165 86.990 84.415 87.415 ;
        RECT 84.625 87.140 85.730 87.310 ;
        RECT 84.110 86.860 84.415 86.990 ;
        RECT 83.660 85.665 83.940 86.615 ;
        RECT 84.110 85.755 84.280 86.860 ;
        RECT 84.450 86.075 84.690 86.670 ;
        RECT 84.860 86.605 85.390 86.970 ;
        RECT 84.860 85.905 85.030 86.605 ;
        RECT 85.560 86.525 85.730 87.140 ;
        RECT 85.900 86.785 86.070 87.585 ;
        RECT 86.240 87.085 86.490 87.415 ;
        RECT 86.715 87.115 87.600 87.285 ;
        RECT 85.560 86.435 86.070 86.525 ;
        RECT 84.110 85.625 84.335 85.755 ;
        RECT 84.505 85.685 85.030 85.905 ;
        RECT 85.200 86.265 86.070 86.435 ;
        RECT 83.745 85.035 83.995 85.495 ;
        RECT 84.165 85.485 84.335 85.625 ;
        RECT 85.200 85.485 85.370 86.265 ;
        RECT 85.900 86.195 86.070 86.265 ;
        RECT 85.580 86.015 85.780 86.045 ;
        RECT 86.240 86.015 86.410 87.085 ;
        RECT 86.580 86.195 86.770 86.915 ;
        RECT 85.580 85.715 86.410 86.015 ;
        RECT 86.940 85.985 87.260 86.945 ;
        RECT 84.165 85.315 84.500 85.485 ;
        RECT 84.695 85.315 85.370 85.485 ;
        RECT 85.690 85.035 86.060 85.535 ;
        RECT 86.240 85.485 86.410 85.715 ;
        RECT 86.795 85.655 87.260 85.985 ;
        RECT 87.430 86.275 87.600 87.115 ;
        RECT 87.780 87.085 88.095 87.585 ;
        RECT 88.325 86.855 88.665 87.415 ;
        RECT 87.770 86.480 88.665 86.855 ;
        RECT 88.835 86.575 89.005 87.585 ;
        RECT 88.475 86.275 88.665 86.480 ;
        RECT 89.175 86.525 89.505 87.370 ;
        RECT 89.175 86.445 89.565 86.525 ;
        RECT 89.735 86.495 90.945 87.585 ;
        RECT 91.205 86.915 91.375 87.415 ;
        RECT 91.545 87.085 91.875 87.585 ;
        RECT 91.205 86.745 91.870 86.915 ;
        RECT 89.350 86.395 89.565 86.445 ;
        RECT 87.430 85.945 88.305 86.275 ;
        RECT 88.475 85.945 89.225 86.275 ;
        RECT 87.430 85.485 87.600 85.945 ;
        RECT 88.475 85.775 88.675 85.945 ;
        RECT 89.395 85.815 89.565 86.395 ;
        RECT 89.340 85.775 89.565 85.815 ;
        RECT 86.240 85.315 86.645 85.485 ;
        RECT 86.815 85.315 87.600 85.485 ;
        RECT 87.875 85.035 88.085 85.565 ;
        RECT 88.345 85.250 88.675 85.775 ;
        RECT 89.185 85.690 89.565 85.775 ;
        RECT 89.735 85.785 90.255 86.325 ;
        RECT 90.425 85.955 90.945 86.495 ;
        RECT 91.120 85.925 91.470 86.575 ;
        RECT 88.845 85.035 89.015 85.645 ;
        RECT 89.185 85.255 89.515 85.690 ;
        RECT 89.735 85.035 90.945 85.785 ;
        RECT 91.640 85.755 91.870 86.745 ;
        RECT 91.205 85.585 91.870 85.755 ;
        RECT 91.205 85.295 91.375 85.585 ;
        RECT 91.545 85.035 91.875 85.415 ;
        RECT 92.045 85.295 92.230 87.415 ;
        RECT 92.470 87.125 92.735 87.585 ;
        RECT 92.905 86.990 93.155 87.415 ;
        RECT 93.365 87.140 94.470 87.310 ;
        RECT 92.850 86.860 93.155 86.990 ;
        RECT 92.400 85.665 92.680 86.615 ;
        RECT 92.850 85.755 93.020 86.860 ;
        RECT 93.190 86.075 93.430 86.670 ;
        RECT 93.600 86.605 94.130 86.970 ;
        RECT 93.600 85.905 93.770 86.605 ;
        RECT 94.300 86.525 94.470 87.140 ;
        RECT 94.640 86.785 94.810 87.585 ;
        RECT 94.980 87.085 95.230 87.415 ;
        RECT 95.455 87.115 96.340 87.285 ;
        RECT 94.300 86.435 94.810 86.525 ;
        RECT 92.850 85.625 93.075 85.755 ;
        RECT 93.245 85.685 93.770 85.905 ;
        RECT 93.940 86.265 94.810 86.435 ;
        RECT 92.485 85.035 92.735 85.495 ;
        RECT 92.905 85.485 93.075 85.625 ;
        RECT 93.940 85.485 94.110 86.265 ;
        RECT 94.640 86.195 94.810 86.265 ;
        RECT 94.320 86.015 94.520 86.045 ;
        RECT 94.980 86.015 95.150 87.085 ;
        RECT 95.320 86.195 95.510 86.915 ;
        RECT 94.320 85.715 95.150 86.015 ;
        RECT 95.680 85.985 96.000 86.945 ;
        RECT 92.905 85.315 93.240 85.485 ;
        RECT 93.435 85.315 94.110 85.485 ;
        RECT 94.430 85.035 94.800 85.535 ;
        RECT 94.980 85.485 95.150 85.715 ;
        RECT 95.535 85.655 96.000 85.985 ;
        RECT 96.170 86.275 96.340 87.115 ;
        RECT 96.520 87.085 96.835 87.585 ;
        RECT 97.065 86.855 97.405 87.415 ;
        RECT 96.510 86.480 97.405 86.855 ;
        RECT 97.575 86.575 97.745 87.585 ;
        RECT 97.215 86.275 97.405 86.480 ;
        RECT 97.915 86.525 98.245 87.370 ;
        RECT 98.565 86.915 98.735 87.415 ;
        RECT 98.905 87.085 99.235 87.585 ;
        RECT 98.565 86.745 99.230 86.915 ;
        RECT 97.915 86.445 98.305 86.525 ;
        RECT 98.090 86.395 98.305 86.445 ;
        RECT 96.170 85.945 97.045 86.275 ;
        RECT 97.215 85.945 97.965 86.275 ;
        RECT 96.170 85.485 96.340 85.945 ;
        RECT 97.215 85.775 97.415 85.945 ;
        RECT 98.135 85.815 98.305 86.395 ;
        RECT 98.480 85.925 98.830 86.575 ;
        RECT 98.080 85.775 98.305 85.815 ;
        RECT 94.980 85.315 95.385 85.485 ;
        RECT 95.555 85.315 96.340 85.485 ;
        RECT 96.615 85.035 96.825 85.565 ;
        RECT 97.085 85.250 97.415 85.775 ;
        RECT 97.925 85.690 98.305 85.775 ;
        RECT 99.000 85.755 99.230 86.745 ;
        RECT 97.585 85.035 97.755 85.645 ;
        RECT 97.925 85.255 98.255 85.690 ;
        RECT 98.565 85.585 99.230 85.755 ;
        RECT 98.565 85.295 98.735 85.585 ;
        RECT 98.905 85.035 99.235 85.415 ;
        RECT 99.405 85.295 99.590 87.415 ;
        RECT 99.830 87.125 100.095 87.585 ;
        RECT 100.265 86.990 100.515 87.415 ;
        RECT 100.725 87.140 101.830 87.310 ;
        RECT 100.210 86.860 100.515 86.990 ;
        RECT 99.760 85.665 100.040 86.615 ;
        RECT 100.210 85.755 100.380 86.860 ;
        RECT 100.550 86.075 100.790 86.670 ;
        RECT 100.960 86.605 101.490 86.970 ;
        RECT 100.960 85.905 101.130 86.605 ;
        RECT 101.660 86.525 101.830 87.140 ;
        RECT 102.000 86.785 102.170 87.585 ;
        RECT 102.340 87.085 102.590 87.415 ;
        RECT 102.815 87.115 103.700 87.285 ;
        RECT 101.660 86.435 102.170 86.525 ;
        RECT 100.210 85.625 100.435 85.755 ;
        RECT 100.605 85.685 101.130 85.905 ;
        RECT 101.300 86.265 102.170 86.435 ;
        RECT 99.845 85.035 100.095 85.495 ;
        RECT 100.265 85.485 100.435 85.625 ;
        RECT 101.300 85.485 101.470 86.265 ;
        RECT 102.000 86.195 102.170 86.265 ;
        RECT 101.680 86.015 101.880 86.045 ;
        RECT 102.340 86.015 102.510 87.085 ;
        RECT 102.680 86.195 102.870 86.915 ;
        RECT 101.680 85.715 102.510 86.015 ;
        RECT 103.040 85.985 103.360 86.945 ;
        RECT 100.265 85.315 100.600 85.485 ;
        RECT 100.795 85.315 101.470 85.485 ;
        RECT 101.790 85.035 102.160 85.535 ;
        RECT 102.340 85.485 102.510 85.715 ;
        RECT 102.895 85.655 103.360 85.985 ;
        RECT 103.530 86.275 103.700 87.115 ;
        RECT 103.880 87.085 104.195 87.585 ;
        RECT 104.425 86.855 104.765 87.415 ;
        RECT 103.870 86.480 104.765 86.855 ;
        RECT 104.935 86.575 105.105 87.585 ;
        RECT 104.575 86.275 104.765 86.480 ;
        RECT 105.275 86.525 105.605 87.370 ;
        RECT 105.835 86.615 106.105 87.385 ;
        RECT 106.275 86.805 106.605 87.585 ;
        RECT 106.810 86.980 106.995 87.385 ;
        RECT 107.165 87.160 107.500 87.585 ;
        RECT 106.810 86.805 107.475 86.980 ;
        RECT 105.275 86.445 105.665 86.525 ;
        RECT 105.450 86.395 105.665 86.445 ;
        RECT 103.530 85.945 104.405 86.275 ;
        RECT 104.575 85.945 105.325 86.275 ;
        RECT 103.530 85.485 103.700 85.945 ;
        RECT 104.575 85.775 104.775 85.945 ;
        RECT 105.495 85.815 105.665 86.395 ;
        RECT 105.440 85.775 105.665 85.815 ;
        RECT 102.340 85.315 102.745 85.485 ;
        RECT 102.915 85.315 103.700 85.485 ;
        RECT 103.975 85.035 104.185 85.565 ;
        RECT 104.445 85.250 104.775 85.775 ;
        RECT 105.285 85.690 105.665 85.775 ;
        RECT 105.835 86.445 106.965 86.615 ;
        RECT 104.945 85.035 105.115 85.645 ;
        RECT 105.285 85.255 105.615 85.690 ;
        RECT 105.835 85.535 106.005 86.445 ;
        RECT 106.175 85.695 106.535 86.275 ;
        RECT 106.715 85.945 106.965 86.445 ;
        RECT 107.135 85.775 107.475 86.805 ;
        RECT 107.675 86.420 107.965 87.585 ;
        RECT 108.135 86.445 108.475 87.415 ;
        RECT 108.645 86.445 108.815 87.585 ;
        RECT 109.085 86.785 109.335 87.585 ;
        RECT 109.980 86.615 110.310 87.415 ;
        RECT 110.610 86.785 110.940 87.585 ;
        RECT 111.110 86.615 111.440 87.415 ;
        RECT 109.005 86.445 111.440 86.615 ;
        RECT 111.820 87.195 112.155 87.415 ;
        RECT 113.160 87.205 113.515 87.585 ;
        RECT 111.820 86.575 112.075 87.195 ;
        RECT 112.325 87.035 112.555 87.075 ;
        RECT 113.685 87.035 113.935 87.415 ;
        RECT 112.325 86.835 113.935 87.035 ;
        RECT 112.325 86.745 112.510 86.835 ;
        RECT 113.100 86.825 113.935 86.835 ;
        RECT 114.185 86.805 114.435 87.585 ;
        RECT 114.605 86.735 114.865 87.415 ;
        RECT 112.665 86.635 112.995 86.665 ;
        RECT 112.665 86.575 114.465 86.635 ;
        RECT 111.820 86.465 114.525 86.575 ;
        RECT 106.790 85.605 107.475 85.775 ;
        RECT 108.135 85.835 108.310 86.445 ;
        RECT 109.005 86.195 109.175 86.445 ;
        RECT 108.480 86.025 109.175 86.195 ;
        RECT 109.350 86.025 109.770 86.225 ;
        RECT 109.940 86.025 110.270 86.225 ;
        RECT 110.440 86.025 110.770 86.225 ;
        RECT 105.835 85.205 106.095 85.535 ;
        RECT 106.305 85.035 106.580 85.515 ;
        RECT 106.790 85.205 106.995 85.605 ;
        RECT 107.165 85.035 107.500 85.435 ;
        RECT 107.675 85.035 107.965 85.760 ;
        RECT 108.135 85.205 108.475 85.835 ;
        RECT 108.645 85.035 108.895 85.835 ;
        RECT 109.085 85.685 110.310 85.855 ;
        RECT 109.085 85.205 109.415 85.685 ;
        RECT 109.585 85.035 109.810 85.495 ;
        RECT 109.980 85.205 110.310 85.685 ;
        RECT 110.940 85.815 111.110 86.445 ;
        RECT 111.820 86.405 112.995 86.465 ;
        RECT 114.325 86.430 114.525 86.465 ;
        RECT 111.295 86.025 111.645 86.275 ;
        RECT 111.815 86.025 112.305 86.225 ;
        RECT 112.495 86.025 112.970 86.235 ;
        RECT 110.940 85.205 111.440 85.815 ;
        RECT 111.820 85.035 112.275 85.800 ;
        RECT 112.750 85.625 112.970 86.025 ;
        RECT 113.215 86.025 113.545 86.235 ;
        RECT 113.215 85.625 113.425 86.025 ;
        RECT 113.715 85.990 114.125 86.295 ;
        RECT 114.355 85.855 114.525 86.430 ;
        RECT 114.255 85.735 114.525 85.855 ;
        RECT 113.680 85.690 114.525 85.735 ;
        RECT 113.680 85.565 114.435 85.690 ;
        RECT 113.680 85.415 113.850 85.565 ;
        RECT 114.695 85.545 114.865 86.735 ;
        RECT 115.555 86.525 115.885 87.370 ;
        RECT 116.055 86.575 116.225 87.585 ;
        RECT 116.395 86.855 116.735 87.415 ;
        RECT 116.965 87.085 117.280 87.585 ;
        RECT 117.460 87.115 118.345 87.285 ;
        RECT 115.495 86.445 115.885 86.525 ;
        RECT 116.395 86.480 117.290 86.855 ;
        RECT 115.495 86.395 115.710 86.445 ;
        RECT 115.495 85.815 115.665 86.395 ;
        RECT 116.395 86.275 116.585 86.480 ;
        RECT 117.460 86.275 117.630 87.115 ;
        RECT 118.570 87.085 118.820 87.415 ;
        RECT 115.835 85.945 116.585 86.275 ;
        RECT 116.755 85.945 117.630 86.275 ;
        RECT 115.495 85.775 115.720 85.815 ;
        RECT 116.385 85.775 116.585 85.945 ;
        RECT 115.495 85.690 115.875 85.775 ;
        RECT 114.635 85.535 114.865 85.545 ;
        RECT 112.550 85.205 113.850 85.415 ;
        RECT 114.105 85.035 114.435 85.395 ;
        RECT 114.605 85.205 114.865 85.535 ;
        RECT 115.545 85.255 115.875 85.690 ;
        RECT 116.045 85.035 116.215 85.645 ;
        RECT 116.385 85.250 116.715 85.775 ;
        RECT 116.975 85.035 117.185 85.565 ;
        RECT 117.460 85.485 117.630 85.945 ;
        RECT 117.800 85.985 118.120 86.945 ;
        RECT 118.290 86.195 118.480 86.915 ;
        RECT 118.650 86.015 118.820 87.085 ;
        RECT 118.990 86.785 119.160 87.585 ;
        RECT 119.330 87.140 120.435 87.310 ;
        RECT 119.330 86.525 119.500 87.140 ;
        RECT 120.645 86.990 120.895 87.415 ;
        RECT 121.065 87.125 121.330 87.585 ;
        RECT 119.670 86.605 120.200 86.970 ;
        RECT 120.645 86.860 120.950 86.990 ;
        RECT 118.990 86.435 119.500 86.525 ;
        RECT 118.990 86.265 119.860 86.435 ;
        RECT 118.990 86.195 119.160 86.265 ;
        RECT 119.280 86.015 119.480 86.045 ;
        RECT 117.800 85.655 118.265 85.985 ;
        RECT 118.650 85.715 119.480 86.015 ;
        RECT 118.650 85.485 118.820 85.715 ;
        RECT 117.460 85.315 118.245 85.485 ;
        RECT 118.415 85.315 118.820 85.485 ;
        RECT 119.000 85.035 119.370 85.535 ;
        RECT 119.690 85.485 119.860 86.265 ;
        RECT 120.030 85.905 120.200 86.605 ;
        RECT 120.370 86.075 120.610 86.670 ;
        RECT 120.030 85.685 120.555 85.905 ;
        RECT 120.780 85.755 120.950 86.860 ;
        RECT 120.725 85.625 120.950 85.755 ;
        RECT 121.120 85.665 121.400 86.615 ;
        RECT 120.725 85.485 120.895 85.625 ;
        RECT 119.690 85.315 120.365 85.485 ;
        RECT 120.560 85.315 120.895 85.485 ;
        RECT 121.065 85.035 121.315 85.495 ;
        RECT 121.570 85.295 121.755 87.415 ;
        RECT 121.925 87.085 122.255 87.585 ;
        RECT 122.425 86.915 122.595 87.415 ;
        RECT 121.930 86.745 122.595 86.915 ;
        RECT 122.945 86.915 123.115 87.415 ;
        RECT 123.285 87.085 123.615 87.585 ;
        RECT 122.945 86.745 123.610 86.915 ;
        RECT 121.930 85.755 122.160 86.745 ;
        RECT 122.330 85.925 122.680 86.575 ;
        RECT 122.860 85.925 123.210 86.575 ;
        RECT 123.380 85.755 123.610 86.745 ;
        RECT 121.930 85.585 122.595 85.755 ;
        RECT 121.925 85.035 122.255 85.415 ;
        RECT 122.425 85.295 122.595 85.585 ;
        RECT 122.945 85.585 123.610 85.755 ;
        RECT 122.945 85.295 123.115 85.585 ;
        RECT 123.285 85.035 123.615 85.415 ;
        RECT 123.785 85.295 123.970 87.415 ;
        RECT 124.210 87.125 124.475 87.585 ;
        RECT 124.645 86.990 124.895 87.415 ;
        RECT 125.105 87.140 126.210 87.310 ;
        RECT 124.590 86.860 124.895 86.990 ;
        RECT 124.140 85.665 124.420 86.615 ;
        RECT 124.590 85.755 124.760 86.860 ;
        RECT 124.930 86.075 125.170 86.670 ;
        RECT 125.340 86.605 125.870 86.970 ;
        RECT 125.340 85.905 125.510 86.605 ;
        RECT 126.040 86.525 126.210 87.140 ;
        RECT 126.380 86.785 126.550 87.585 ;
        RECT 126.720 87.085 126.970 87.415 ;
        RECT 127.195 87.115 128.080 87.285 ;
        RECT 126.040 86.435 126.550 86.525 ;
        RECT 124.590 85.625 124.815 85.755 ;
        RECT 124.985 85.685 125.510 85.905 ;
        RECT 125.680 86.265 126.550 86.435 ;
        RECT 124.225 85.035 124.475 85.495 ;
        RECT 124.645 85.485 124.815 85.625 ;
        RECT 125.680 85.485 125.850 86.265 ;
        RECT 126.380 86.195 126.550 86.265 ;
        RECT 126.060 86.015 126.260 86.045 ;
        RECT 126.720 86.015 126.890 87.085 ;
        RECT 127.060 86.195 127.250 86.915 ;
        RECT 126.060 85.715 126.890 86.015 ;
        RECT 127.420 85.985 127.740 86.945 ;
        RECT 124.645 85.315 124.980 85.485 ;
        RECT 125.175 85.315 125.850 85.485 ;
        RECT 126.170 85.035 126.540 85.535 ;
        RECT 126.720 85.485 126.890 85.715 ;
        RECT 127.275 85.655 127.740 85.985 ;
        RECT 127.910 86.275 128.080 87.115 ;
        RECT 128.260 87.085 128.575 87.585 ;
        RECT 128.805 86.855 129.145 87.415 ;
        RECT 128.250 86.480 129.145 86.855 ;
        RECT 129.315 86.575 129.485 87.585 ;
        RECT 128.955 86.275 129.145 86.480 ;
        RECT 129.655 86.525 129.985 87.370 ;
        RECT 130.250 86.795 130.785 87.415 ;
        RECT 129.655 86.445 130.045 86.525 ;
        RECT 129.830 86.395 130.045 86.445 ;
        RECT 127.910 85.945 128.785 86.275 ;
        RECT 128.955 85.945 129.705 86.275 ;
        RECT 127.910 85.485 128.080 85.945 ;
        RECT 128.955 85.775 129.155 85.945 ;
        RECT 129.875 85.815 130.045 86.395 ;
        RECT 129.820 85.775 130.045 85.815 ;
        RECT 126.720 85.315 127.125 85.485 ;
        RECT 127.295 85.315 128.080 85.485 ;
        RECT 128.355 85.035 128.565 85.565 ;
        RECT 128.825 85.250 129.155 85.775 ;
        RECT 129.665 85.690 130.045 85.775 ;
        RECT 130.250 85.775 130.565 86.795 ;
        RECT 130.955 86.785 131.285 87.585 ;
        RECT 131.770 86.615 132.160 86.790 ;
        RECT 130.735 86.445 132.160 86.615 ;
        RECT 130.735 85.945 130.905 86.445 ;
        RECT 129.325 85.035 129.495 85.645 ;
        RECT 129.665 85.255 129.995 85.690 ;
        RECT 130.250 85.205 130.865 85.775 ;
        RECT 131.155 85.715 131.420 86.275 ;
        RECT 131.590 85.545 131.760 86.445 ;
        RECT 133.435 86.420 133.725 87.585 ;
        RECT 134.100 86.615 134.430 87.415 ;
        RECT 134.600 86.785 134.930 87.585 ;
        RECT 135.230 86.615 135.560 87.415 ;
        RECT 136.205 86.785 136.455 87.585 ;
        RECT 134.100 86.445 136.535 86.615 ;
        RECT 136.725 86.445 136.895 87.585 ;
        RECT 137.065 86.445 137.405 87.415 ;
        RECT 137.575 86.495 139.245 87.585 ;
        RECT 131.930 85.715 132.285 86.275 ;
        RECT 133.895 86.025 134.245 86.275 ;
        RECT 134.430 85.815 134.600 86.445 ;
        RECT 134.770 86.025 135.100 86.225 ;
        RECT 135.270 86.025 135.600 86.225 ;
        RECT 135.770 86.025 136.190 86.225 ;
        RECT 136.365 86.195 136.535 86.445 ;
        RECT 136.365 86.025 137.060 86.195 ;
        RECT 131.035 85.035 131.250 85.545 ;
        RECT 131.480 85.215 131.760 85.545 ;
        RECT 131.940 85.035 132.180 85.545 ;
        RECT 133.435 85.035 133.725 85.760 ;
        RECT 134.100 85.205 134.600 85.815 ;
        RECT 135.230 85.685 136.455 85.855 ;
        RECT 137.230 85.835 137.405 86.445 ;
        RECT 135.230 85.205 135.560 85.685 ;
        RECT 135.730 85.035 135.955 85.495 ;
        RECT 136.125 85.205 136.455 85.685 ;
        RECT 136.645 85.035 136.895 85.835 ;
        RECT 137.065 85.205 137.405 85.835 ;
        RECT 137.575 85.805 138.325 86.325 ;
        RECT 138.495 85.975 139.245 86.495 ;
        RECT 139.965 86.655 140.135 87.415 ;
        RECT 140.350 86.825 140.680 87.585 ;
        RECT 139.965 86.485 140.680 86.655 ;
        RECT 140.850 86.510 141.105 87.415 ;
        RECT 139.875 85.935 140.230 86.305 ;
        RECT 140.510 86.275 140.680 86.485 ;
        RECT 140.510 85.945 140.765 86.275 ;
        RECT 137.575 85.035 139.245 85.805 ;
        RECT 140.510 85.755 140.680 85.945 ;
        RECT 140.935 85.780 141.105 86.510 ;
        RECT 141.280 86.435 141.540 87.585 ;
        RECT 141.715 86.495 142.925 87.585 ;
        RECT 141.715 85.955 142.235 86.495 ;
        RECT 139.965 85.585 140.680 85.755 ;
        RECT 139.965 85.205 140.135 85.585 ;
        RECT 140.350 85.035 140.680 85.415 ;
        RECT 140.850 85.205 141.105 85.780 ;
        RECT 141.280 85.035 141.540 85.875 ;
        RECT 142.405 85.785 142.925 86.325 ;
        RECT 141.715 85.035 142.925 85.785 ;
        RECT 17.430 84.865 143.010 85.035 ;
        RECT 17.515 84.115 18.725 84.865 ;
        RECT 18.895 84.320 24.240 84.865 ;
        RECT 24.415 84.320 29.760 84.865 ;
        RECT 29.935 84.320 35.280 84.865 ;
        RECT 35.455 84.320 40.800 84.865 ;
        RECT 17.515 83.575 18.035 84.115 ;
        RECT 18.205 83.405 18.725 83.945 ;
        RECT 20.480 83.490 20.820 84.320 ;
        RECT 17.515 82.315 18.725 83.405 ;
        RECT 22.300 82.750 22.650 84.000 ;
        RECT 26.000 83.490 26.340 84.320 ;
        RECT 27.820 82.750 28.170 84.000 ;
        RECT 31.520 83.490 31.860 84.320 ;
        RECT 33.340 82.750 33.690 84.000 ;
        RECT 37.040 83.490 37.380 84.320 ;
        RECT 40.975 84.095 42.645 84.865 ;
        RECT 43.275 84.140 43.565 84.865 ;
        RECT 43.735 84.320 49.080 84.865 ;
        RECT 49.255 84.320 54.600 84.865 ;
        RECT 54.775 84.320 60.120 84.865 ;
        RECT 60.295 84.320 65.640 84.865 ;
        RECT 38.860 82.750 39.210 84.000 ;
        RECT 40.975 83.575 41.725 84.095 ;
        RECT 41.895 83.405 42.645 83.925 ;
        RECT 45.320 83.490 45.660 84.320 ;
        RECT 18.895 82.315 24.240 82.750 ;
        RECT 24.415 82.315 29.760 82.750 ;
        RECT 29.935 82.315 35.280 82.750 ;
        RECT 35.455 82.315 40.800 82.750 ;
        RECT 40.975 82.315 42.645 83.405 ;
        RECT 43.275 82.315 43.565 83.480 ;
        RECT 47.140 82.750 47.490 84.000 ;
        RECT 50.840 83.490 51.180 84.320 ;
        RECT 52.660 82.750 53.010 84.000 ;
        RECT 56.360 83.490 56.700 84.320 ;
        RECT 58.180 82.750 58.530 84.000 ;
        RECT 61.880 83.490 62.220 84.320 ;
        RECT 65.815 84.095 68.405 84.865 ;
        RECT 69.035 84.140 69.325 84.865 ;
        RECT 69.495 84.320 74.840 84.865 ;
        RECT 75.015 84.320 80.360 84.865 ;
        RECT 63.700 82.750 64.050 84.000 ;
        RECT 65.815 83.575 67.025 84.095 ;
        RECT 67.195 83.405 68.405 83.925 ;
        RECT 71.080 83.490 71.420 84.320 ;
        RECT 43.735 82.315 49.080 82.750 ;
        RECT 49.255 82.315 54.600 82.750 ;
        RECT 54.775 82.315 60.120 82.750 ;
        RECT 60.295 82.315 65.640 82.750 ;
        RECT 65.815 82.315 68.405 83.405 ;
        RECT 69.035 82.315 69.325 83.480 ;
        RECT 72.900 82.750 73.250 84.000 ;
        RECT 76.600 83.490 76.940 84.320 ;
        RECT 80.625 84.315 80.795 84.605 ;
        RECT 80.965 84.485 81.295 84.865 ;
        RECT 80.625 84.145 81.290 84.315 ;
        RECT 78.420 82.750 78.770 84.000 ;
        RECT 80.540 83.325 80.890 83.975 ;
        RECT 81.060 83.155 81.290 84.145 ;
        RECT 80.625 82.985 81.290 83.155 ;
        RECT 69.495 82.315 74.840 82.750 ;
        RECT 75.015 82.315 80.360 82.750 ;
        RECT 80.625 82.485 80.795 82.985 ;
        RECT 80.965 82.315 81.295 82.815 ;
        RECT 81.465 82.485 81.650 84.605 ;
        RECT 81.905 84.405 82.155 84.865 ;
        RECT 82.325 84.415 82.660 84.585 ;
        RECT 82.855 84.415 83.530 84.585 ;
        RECT 82.325 84.275 82.495 84.415 ;
        RECT 81.820 83.285 82.100 84.235 ;
        RECT 82.270 84.145 82.495 84.275 ;
        RECT 82.270 83.040 82.440 84.145 ;
        RECT 82.665 83.995 83.190 84.215 ;
        RECT 82.610 83.230 82.850 83.825 ;
        RECT 83.020 83.295 83.190 83.995 ;
        RECT 83.360 83.635 83.530 84.415 ;
        RECT 83.850 84.365 84.220 84.865 ;
        RECT 84.400 84.415 84.805 84.585 ;
        RECT 84.975 84.415 85.760 84.585 ;
        RECT 84.400 84.185 84.570 84.415 ;
        RECT 83.740 83.885 84.570 84.185 ;
        RECT 84.955 83.915 85.420 84.245 ;
        RECT 83.740 83.855 83.940 83.885 ;
        RECT 84.060 83.635 84.230 83.705 ;
        RECT 83.360 83.465 84.230 83.635 ;
        RECT 83.720 83.375 84.230 83.465 ;
        RECT 82.270 82.910 82.575 83.040 ;
        RECT 83.020 82.930 83.550 83.295 ;
        RECT 81.890 82.315 82.155 82.775 ;
        RECT 82.325 82.485 82.575 82.910 ;
        RECT 83.720 82.760 83.890 83.375 ;
        RECT 82.785 82.590 83.890 82.760 ;
        RECT 84.060 82.315 84.230 83.115 ;
        RECT 84.400 82.815 84.570 83.885 ;
        RECT 84.740 82.985 84.930 83.705 ;
        RECT 85.100 82.955 85.420 83.915 ;
        RECT 85.590 83.955 85.760 84.415 ;
        RECT 86.035 84.335 86.245 84.865 ;
        RECT 86.505 84.125 86.835 84.650 ;
        RECT 87.005 84.255 87.175 84.865 ;
        RECT 87.345 84.210 87.675 84.645 ;
        RECT 87.345 84.125 87.725 84.210 ;
        RECT 86.635 83.955 86.835 84.125 ;
        RECT 87.500 84.085 87.725 84.125 ;
        RECT 85.590 83.625 86.465 83.955 ;
        RECT 86.635 83.625 87.385 83.955 ;
        RECT 84.400 82.485 84.650 82.815 ;
        RECT 85.590 82.785 85.760 83.625 ;
        RECT 86.635 83.420 86.825 83.625 ;
        RECT 87.555 83.505 87.725 84.085 ;
        RECT 87.510 83.455 87.725 83.505 ;
        RECT 85.930 83.045 86.825 83.420 ;
        RECT 87.335 83.375 87.725 83.455 ;
        RECT 87.930 84.125 88.545 84.695 ;
        RECT 88.715 84.355 88.930 84.865 ;
        RECT 89.160 84.355 89.440 84.685 ;
        RECT 89.620 84.355 89.860 84.865 ;
        RECT 84.875 82.615 85.760 82.785 ;
        RECT 85.940 82.315 86.255 82.815 ;
        RECT 86.485 82.485 86.825 83.045 ;
        RECT 86.995 82.315 87.165 83.325 ;
        RECT 87.335 82.530 87.665 83.375 ;
        RECT 87.930 83.105 88.245 84.125 ;
        RECT 88.415 83.455 88.585 83.955 ;
        RECT 88.835 83.625 89.100 84.185 ;
        RECT 89.270 83.455 89.440 84.355 ;
        RECT 89.610 83.625 89.965 84.185 ;
        RECT 90.230 84.125 90.845 84.695 ;
        RECT 91.015 84.355 91.230 84.865 ;
        RECT 91.460 84.355 91.740 84.685 ;
        RECT 91.920 84.355 92.160 84.865 ;
        RECT 88.415 83.285 89.840 83.455 ;
        RECT 87.930 82.485 88.465 83.105 ;
        RECT 88.635 82.315 88.965 83.115 ;
        RECT 89.450 83.110 89.840 83.285 ;
        RECT 90.230 83.105 90.545 84.125 ;
        RECT 90.715 83.455 90.885 83.955 ;
        RECT 91.135 83.625 91.400 84.185 ;
        RECT 91.570 83.455 91.740 84.355 ;
        RECT 91.910 83.625 92.265 84.185 ;
        RECT 92.495 84.095 94.165 84.865 ;
        RECT 94.795 84.140 95.085 84.865 ;
        RECT 92.495 83.575 93.245 84.095 ;
        RECT 95.255 84.065 95.595 84.695 ;
        RECT 95.765 84.065 96.015 84.865 ;
        RECT 96.205 84.215 96.535 84.695 ;
        RECT 96.705 84.405 96.930 84.865 ;
        RECT 97.100 84.215 97.430 84.695 ;
        RECT 90.715 83.285 92.140 83.455 ;
        RECT 93.415 83.405 94.165 83.925 ;
        RECT 90.230 82.485 90.765 83.105 ;
        RECT 90.935 82.315 91.265 83.115 ;
        RECT 91.750 83.110 92.140 83.285 ;
        RECT 92.495 82.315 94.165 83.405 ;
        RECT 94.795 82.315 95.085 83.480 ;
        RECT 95.255 83.455 95.430 84.065 ;
        RECT 96.205 84.045 97.430 84.215 ;
        RECT 98.060 84.085 98.560 84.695 ;
        RECT 99.430 84.125 100.045 84.695 ;
        RECT 100.215 84.355 100.430 84.865 ;
        RECT 100.660 84.355 100.940 84.685 ;
        RECT 101.120 84.355 101.360 84.865 ;
        RECT 95.600 83.705 96.295 83.875 ;
        RECT 96.125 83.455 96.295 83.705 ;
        RECT 96.470 83.675 96.890 83.875 ;
        RECT 97.060 83.675 97.390 83.875 ;
        RECT 97.560 83.675 97.890 83.875 ;
        RECT 98.060 83.455 98.230 84.085 ;
        RECT 98.415 83.625 98.765 83.875 ;
        RECT 95.255 82.485 95.595 83.455 ;
        RECT 95.765 82.315 95.935 83.455 ;
        RECT 96.125 83.285 98.560 83.455 ;
        RECT 96.205 82.315 96.455 83.115 ;
        RECT 97.100 82.485 97.430 83.285 ;
        RECT 97.730 82.315 98.060 83.115 ;
        RECT 98.230 82.485 98.560 83.285 ;
        RECT 99.430 83.105 99.745 84.125 ;
        RECT 99.915 83.455 100.085 83.955 ;
        RECT 100.335 83.625 100.600 84.185 ;
        RECT 100.770 83.455 100.940 84.355 ;
        RECT 101.745 84.210 102.075 84.645 ;
        RECT 102.245 84.255 102.415 84.865 ;
        RECT 101.110 83.625 101.465 84.185 ;
        RECT 101.695 84.125 102.075 84.210 ;
        RECT 102.585 84.125 102.915 84.650 ;
        RECT 103.175 84.335 103.385 84.865 ;
        RECT 103.660 84.415 104.445 84.585 ;
        RECT 104.615 84.415 105.020 84.585 ;
        RECT 101.695 84.085 101.920 84.125 ;
        RECT 101.695 83.505 101.865 84.085 ;
        RECT 102.585 83.955 102.785 84.125 ;
        RECT 103.660 83.955 103.830 84.415 ;
        RECT 102.035 83.625 102.785 83.955 ;
        RECT 102.955 83.625 103.830 83.955 ;
        RECT 101.695 83.455 101.910 83.505 ;
        RECT 99.915 83.285 101.340 83.455 ;
        RECT 101.695 83.375 102.085 83.455 ;
        RECT 99.430 82.485 99.965 83.105 ;
        RECT 100.135 82.315 100.465 83.115 ;
        RECT 100.950 83.110 101.340 83.285 ;
        RECT 101.755 82.530 102.085 83.375 ;
        RECT 102.595 83.420 102.785 83.625 ;
        RECT 102.255 82.315 102.425 83.325 ;
        RECT 102.595 83.045 103.490 83.420 ;
        RECT 102.595 82.485 102.935 83.045 ;
        RECT 103.165 82.315 103.480 82.815 ;
        RECT 103.660 82.785 103.830 83.625 ;
        RECT 104.000 83.915 104.465 84.245 ;
        RECT 104.850 84.185 105.020 84.415 ;
        RECT 105.200 84.365 105.570 84.865 ;
        RECT 105.890 84.415 106.565 84.585 ;
        RECT 106.760 84.415 107.095 84.585 ;
        RECT 104.000 82.955 104.320 83.915 ;
        RECT 104.850 83.885 105.680 84.185 ;
        RECT 104.490 82.985 104.680 83.705 ;
        RECT 104.850 82.815 105.020 83.885 ;
        RECT 105.480 83.855 105.680 83.885 ;
        RECT 105.190 83.635 105.360 83.705 ;
        RECT 105.890 83.635 106.060 84.415 ;
        RECT 106.925 84.275 107.095 84.415 ;
        RECT 107.265 84.405 107.515 84.865 ;
        RECT 105.190 83.465 106.060 83.635 ;
        RECT 106.230 83.995 106.755 84.215 ;
        RECT 106.925 84.145 107.150 84.275 ;
        RECT 105.190 83.375 105.700 83.465 ;
        RECT 103.660 82.615 104.545 82.785 ;
        RECT 104.770 82.485 105.020 82.815 ;
        RECT 105.190 82.315 105.360 83.115 ;
        RECT 105.530 82.760 105.700 83.375 ;
        RECT 106.230 83.295 106.400 83.995 ;
        RECT 105.870 82.930 106.400 83.295 ;
        RECT 106.570 83.230 106.810 83.825 ;
        RECT 106.980 83.040 107.150 84.145 ;
        RECT 107.320 83.285 107.600 84.235 ;
        RECT 106.845 82.910 107.150 83.040 ;
        RECT 105.530 82.590 106.635 82.760 ;
        RECT 106.845 82.485 107.095 82.910 ;
        RECT 107.265 82.315 107.530 82.775 ;
        RECT 107.770 82.485 107.955 84.605 ;
        RECT 108.125 84.485 108.455 84.865 ;
        RECT 108.625 84.315 108.795 84.605 ;
        RECT 109.220 84.355 109.460 84.865 ;
        RECT 109.640 84.355 109.920 84.685 ;
        RECT 110.150 84.355 110.365 84.865 ;
        RECT 108.130 84.145 108.795 84.315 ;
        RECT 108.130 83.155 108.360 84.145 ;
        RECT 108.530 83.325 108.880 83.975 ;
        RECT 109.115 83.625 109.470 84.185 ;
        RECT 109.640 83.455 109.810 84.355 ;
        RECT 109.980 83.625 110.245 84.185 ;
        RECT 110.535 84.125 111.150 84.695 ;
        RECT 110.495 83.455 110.665 83.955 ;
        RECT 109.240 83.285 110.665 83.455 ;
        RECT 108.130 82.985 108.795 83.155 ;
        RECT 109.240 83.110 109.630 83.285 ;
        RECT 108.125 82.315 108.455 82.815 ;
        RECT 108.625 82.485 108.795 82.985 ;
        RECT 110.115 82.315 110.445 83.115 ;
        RECT 110.835 83.105 111.150 84.125 ;
        RECT 111.355 84.095 113.025 84.865 ;
        RECT 113.195 84.365 113.455 84.695 ;
        RECT 113.625 84.505 113.955 84.865 ;
        RECT 114.210 84.485 115.510 84.695 ;
        RECT 113.195 84.355 113.425 84.365 ;
        RECT 111.355 83.575 112.105 84.095 ;
        RECT 112.275 83.405 113.025 83.925 ;
        RECT 110.615 82.485 111.150 83.105 ;
        RECT 111.355 82.315 113.025 83.405 ;
        RECT 113.195 83.165 113.365 84.355 ;
        RECT 114.210 84.335 114.380 84.485 ;
        RECT 113.625 84.210 114.380 84.335 ;
        RECT 113.535 84.165 114.380 84.210 ;
        RECT 113.535 84.045 113.805 84.165 ;
        RECT 113.535 83.470 113.705 84.045 ;
        RECT 113.935 83.605 114.345 83.910 ;
        RECT 114.635 83.875 114.845 84.275 ;
        RECT 114.515 83.665 114.845 83.875 ;
        RECT 115.090 83.875 115.310 84.275 ;
        RECT 115.785 84.100 116.240 84.865 ;
        RECT 116.420 84.100 116.875 84.865 ;
        RECT 117.150 84.485 118.450 84.695 ;
        RECT 118.705 84.505 119.035 84.865 ;
        RECT 118.280 84.335 118.450 84.485 ;
        RECT 119.205 84.365 119.465 84.695 ;
        RECT 119.235 84.355 119.465 84.365 ;
        RECT 117.350 83.875 117.570 84.275 ;
        RECT 115.090 83.665 115.565 83.875 ;
        RECT 115.755 83.675 116.245 83.875 ;
        RECT 116.415 83.675 116.905 83.875 ;
        RECT 117.095 83.665 117.570 83.875 ;
        RECT 117.815 83.875 118.025 84.275 ;
        RECT 118.280 84.210 119.035 84.335 ;
        RECT 118.280 84.165 119.125 84.210 ;
        RECT 118.855 84.045 119.125 84.165 ;
        RECT 117.815 83.665 118.145 83.875 ;
        RECT 118.315 83.605 118.725 83.910 ;
        RECT 113.535 83.435 113.735 83.470 ;
        RECT 115.065 83.435 116.240 83.495 ;
        RECT 113.535 83.325 116.240 83.435 ;
        RECT 113.595 83.265 115.395 83.325 ;
        RECT 115.065 83.235 115.395 83.265 ;
        RECT 113.195 82.485 113.455 83.165 ;
        RECT 113.625 82.315 113.875 83.095 ;
        RECT 114.125 83.065 114.960 83.075 ;
        RECT 115.550 83.065 115.735 83.155 ;
        RECT 114.125 82.865 115.735 83.065 ;
        RECT 114.125 82.485 114.375 82.865 ;
        RECT 115.505 82.825 115.735 82.865 ;
        RECT 115.985 82.705 116.240 83.325 ;
        RECT 114.545 82.315 114.900 82.695 ;
        RECT 115.905 82.485 116.240 82.705 ;
        RECT 116.420 83.435 117.595 83.495 ;
        RECT 118.955 83.470 119.125 84.045 ;
        RECT 118.925 83.435 119.125 83.470 ;
        RECT 116.420 83.325 119.125 83.435 ;
        RECT 116.420 82.705 116.675 83.325 ;
        RECT 117.265 83.265 119.065 83.325 ;
        RECT 117.265 83.235 117.595 83.265 ;
        RECT 119.295 83.165 119.465 84.355 ;
        RECT 120.555 84.140 120.845 84.865 ;
        RECT 121.015 84.065 121.355 84.695 ;
        RECT 121.525 84.065 121.775 84.865 ;
        RECT 121.965 84.215 122.295 84.695 ;
        RECT 122.465 84.405 122.690 84.865 ;
        RECT 122.860 84.215 123.190 84.695 ;
        RECT 116.925 83.065 117.110 83.155 ;
        RECT 117.700 83.065 118.535 83.075 ;
        RECT 116.925 82.865 118.535 83.065 ;
        RECT 116.925 82.825 117.155 82.865 ;
        RECT 116.420 82.485 116.755 82.705 ;
        RECT 117.760 82.315 118.115 82.695 ;
        RECT 118.285 82.485 118.535 82.865 ;
        RECT 118.785 82.315 119.035 83.095 ;
        RECT 119.205 82.485 119.465 83.165 ;
        RECT 120.555 82.315 120.845 83.480 ;
        RECT 121.015 83.455 121.190 84.065 ;
        RECT 121.965 84.045 123.190 84.215 ;
        RECT 123.820 84.085 124.320 84.695 ;
        RECT 125.245 84.315 125.415 84.605 ;
        RECT 125.585 84.485 125.915 84.865 ;
        RECT 125.245 84.145 125.910 84.315 ;
        RECT 121.360 83.705 122.055 83.875 ;
        RECT 121.885 83.455 122.055 83.705 ;
        RECT 122.230 83.675 122.650 83.875 ;
        RECT 122.820 83.675 123.150 83.875 ;
        RECT 123.320 83.675 123.650 83.875 ;
        RECT 123.820 83.455 123.990 84.085 ;
        RECT 124.175 83.625 124.525 83.875 ;
        RECT 121.015 82.485 121.355 83.455 ;
        RECT 121.525 82.315 121.695 83.455 ;
        RECT 121.885 83.285 124.320 83.455 ;
        RECT 125.160 83.325 125.510 83.975 ;
        RECT 121.965 82.315 122.215 83.115 ;
        RECT 122.860 82.485 123.190 83.285 ;
        RECT 123.490 82.315 123.820 83.115 ;
        RECT 123.990 82.485 124.320 83.285 ;
        RECT 125.680 83.155 125.910 84.145 ;
        RECT 125.245 82.985 125.910 83.155 ;
        RECT 125.245 82.485 125.415 82.985 ;
        RECT 125.585 82.315 125.915 82.815 ;
        RECT 126.085 82.485 126.270 84.605 ;
        RECT 126.525 84.405 126.775 84.865 ;
        RECT 126.945 84.415 127.280 84.585 ;
        RECT 127.475 84.415 128.150 84.585 ;
        RECT 126.945 84.275 127.115 84.415 ;
        RECT 126.440 83.285 126.720 84.235 ;
        RECT 126.890 84.145 127.115 84.275 ;
        RECT 126.890 83.040 127.060 84.145 ;
        RECT 127.285 83.995 127.810 84.215 ;
        RECT 127.230 83.230 127.470 83.825 ;
        RECT 127.640 83.295 127.810 83.995 ;
        RECT 127.980 83.635 128.150 84.415 ;
        RECT 128.470 84.365 128.840 84.865 ;
        RECT 129.020 84.415 129.425 84.585 ;
        RECT 129.595 84.415 130.380 84.585 ;
        RECT 129.020 84.185 129.190 84.415 ;
        RECT 128.360 83.885 129.190 84.185 ;
        RECT 129.575 83.915 130.040 84.245 ;
        RECT 128.360 83.855 128.560 83.885 ;
        RECT 128.680 83.635 128.850 83.705 ;
        RECT 127.980 83.465 128.850 83.635 ;
        RECT 128.340 83.375 128.850 83.465 ;
        RECT 126.890 82.910 127.195 83.040 ;
        RECT 127.640 82.930 128.170 83.295 ;
        RECT 126.510 82.315 126.775 82.775 ;
        RECT 126.945 82.485 127.195 82.910 ;
        RECT 128.340 82.760 128.510 83.375 ;
        RECT 127.405 82.590 128.510 82.760 ;
        RECT 128.680 82.315 128.850 83.115 ;
        RECT 129.020 82.815 129.190 83.885 ;
        RECT 129.360 82.985 129.550 83.705 ;
        RECT 129.720 82.955 130.040 83.915 ;
        RECT 130.210 83.955 130.380 84.415 ;
        RECT 130.655 84.335 130.865 84.865 ;
        RECT 131.125 84.125 131.455 84.650 ;
        RECT 131.625 84.255 131.795 84.865 ;
        RECT 131.965 84.210 132.295 84.645 ;
        RECT 132.680 84.355 132.920 84.865 ;
        RECT 133.100 84.355 133.380 84.685 ;
        RECT 133.610 84.355 133.825 84.865 ;
        RECT 131.965 84.125 132.345 84.210 ;
        RECT 131.255 83.955 131.455 84.125 ;
        RECT 132.120 84.085 132.345 84.125 ;
        RECT 130.210 83.625 131.085 83.955 ;
        RECT 131.255 83.625 132.005 83.955 ;
        RECT 129.020 82.485 129.270 82.815 ;
        RECT 130.210 82.785 130.380 83.625 ;
        RECT 131.255 83.420 131.445 83.625 ;
        RECT 132.175 83.505 132.345 84.085 ;
        RECT 132.575 83.625 132.930 84.185 ;
        RECT 132.130 83.455 132.345 83.505 ;
        RECT 133.100 83.455 133.270 84.355 ;
        RECT 133.440 83.625 133.705 84.185 ;
        RECT 133.995 84.125 134.610 84.695 ;
        RECT 133.955 83.455 134.125 83.955 ;
        RECT 130.550 83.045 131.445 83.420 ;
        RECT 131.955 83.375 132.345 83.455 ;
        RECT 129.495 82.615 130.380 82.785 ;
        RECT 130.560 82.315 130.875 82.815 ;
        RECT 131.105 82.485 131.445 83.045 ;
        RECT 131.615 82.315 131.785 83.325 ;
        RECT 131.955 82.530 132.285 83.375 ;
        RECT 132.700 83.285 134.125 83.455 ;
        RECT 132.700 83.110 133.090 83.285 ;
        RECT 133.575 82.315 133.905 83.115 ;
        RECT 134.295 83.105 134.610 84.125 ;
        RECT 134.815 84.095 138.325 84.865 ;
        RECT 138.495 84.115 139.705 84.865 ;
        RECT 139.965 84.315 140.135 84.695 ;
        RECT 140.350 84.485 140.680 84.865 ;
        RECT 139.965 84.145 140.680 84.315 ;
        RECT 134.815 83.575 136.465 84.095 ;
        RECT 136.635 83.405 138.325 83.925 ;
        RECT 138.495 83.575 139.015 84.115 ;
        RECT 139.185 83.405 139.705 83.945 ;
        RECT 139.875 83.595 140.230 83.965 ;
        RECT 140.510 83.955 140.680 84.145 ;
        RECT 140.850 84.120 141.105 84.695 ;
        RECT 140.510 83.625 140.765 83.955 ;
        RECT 140.510 83.415 140.680 83.625 ;
        RECT 134.075 82.485 134.610 83.105 ;
        RECT 134.815 82.315 138.325 83.405 ;
        RECT 138.495 82.315 139.705 83.405 ;
        RECT 139.965 83.245 140.680 83.415 ;
        RECT 140.935 83.390 141.105 84.120 ;
        RECT 141.280 84.025 141.540 84.865 ;
        RECT 141.715 84.115 142.925 84.865 ;
        RECT 139.965 82.485 140.135 83.245 ;
        RECT 140.350 82.315 140.680 83.075 ;
        RECT 140.850 82.485 141.105 83.390 ;
        RECT 141.280 82.315 141.540 83.465 ;
        RECT 141.715 83.405 142.235 83.945 ;
        RECT 142.405 83.575 142.925 84.115 ;
        RECT 141.715 82.315 142.925 83.405 ;
        RECT 17.430 82.145 143.010 82.315 ;
        RECT 17.515 81.055 18.725 82.145 ;
        RECT 18.895 81.710 24.240 82.145 ;
        RECT 24.415 81.710 29.760 82.145 ;
        RECT 17.515 80.345 18.035 80.885 ;
        RECT 18.205 80.515 18.725 81.055 ;
        RECT 17.515 79.595 18.725 80.345 ;
        RECT 20.480 80.140 20.820 80.970 ;
        RECT 22.300 80.460 22.650 81.710 ;
        RECT 26.000 80.140 26.340 80.970 ;
        RECT 27.820 80.460 28.170 81.710 ;
        RECT 30.395 80.980 30.685 82.145 ;
        RECT 30.855 81.710 36.200 82.145 ;
        RECT 36.375 81.710 41.720 82.145 ;
        RECT 18.895 79.595 24.240 80.140 ;
        RECT 24.415 79.595 29.760 80.140 ;
        RECT 30.395 79.595 30.685 80.320 ;
        RECT 32.440 80.140 32.780 80.970 ;
        RECT 34.260 80.460 34.610 81.710 ;
        RECT 37.960 80.140 38.300 80.970 ;
        RECT 39.780 80.460 40.130 81.710 ;
        RECT 41.895 81.055 43.105 82.145 ;
        RECT 41.895 80.345 42.415 80.885 ;
        RECT 42.585 80.515 43.105 81.055 ;
        RECT 43.275 80.980 43.565 82.145 ;
        RECT 43.735 81.710 49.080 82.145 ;
        RECT 49.255 81.710 54.600 82.145 ;
        RECT 30.855 79.595 36.200 80.140 ;
        RECT 36.375 79.595 41.720 80.140 ;
        RECT 41.895 79.595 43.105 80.345 ;
        RECT 43.275 79.595 43.565 80.320 ;
        RECT 45.320 80.140 45.660 80.970 ;
        RECT 47.140 80.460 47.490 81.710 ;
        RECT 50.840 80.140 51.180 80.970 ;
        RECT 52.660 80.460 53.010 81.710 ;
        RECT 54.775 81.055 55.985 82.145 ;
        RECT 54.775 80.345 55.295 80.885 ;
        RECT 55.465 80.515 55.985 81.055 ;
        RECT 56.155 80.980 56.445 82.145 ;
        RECT 56.615 81.710 61.960 82.145 ;
        RECT 43.735 79.595 49.080 80.140 ;
        RECT 49.255 79.595 54.600 80.140 ;
        RECT 54.775 79.595 55.985 80.345 ;
        RECT 56.155 79.595 56.445 80.320 ;
        RECT 58.200 80.140 58.540 80.970 ;
        RECT 60.020 80.460 60.370 81.710 ;
        RECT 62.135 81.055 63.805 82.145 ;
        RECT 62.135 80.365 62.885 80.885 ;
        RECT 63.055 80.535 63.805 81.055 ;
        RECT 64.065 81.215 64.235 81.975 ;
        RECT 64.450 81.385 64.780 82.145 ;
        RECT 64.065 81.045 64.780 81.215 ;
        RECT 64.950 81.070 65.205 81.975 ;
        RECT 63.975 80.495 64.330 80.865 ;
        RECT 64.610 80.835 64.780 81.045 ;
        RECT 64.610 80.505 64.865 80.835 ;
        RECT 56.615 79.595 61.960 80.140 ;
        RECT 62.135 79.595 63.805 80.365 ;
        RECT 64.610 80.315 64.780 80.505 ;
        RECT 65.035 80.340 65.205 81.070 ;
        RECT 65.380 80.995 65.640 82.145 ;
        RECT 65.815 81.055 68.405 82.145 ;
        RECT 64.065 80.145 64.780 80.315 ;
        RECT 64.065 79.765 64.235 80.145 ;
        RECT 64.450 79.595 64.780 79.975 ;
        RECT 64.950 79.765 65.205 80.340 ;
        RECT 65.380 79.595 65.640 80.435 ;
        RECT 65.815 80.365 67.025 80.885 ;
        RECT 67.195 80.535 68.405 81.055 ;
        RECT 69.035 80.980 69.325 82.145 ;
        RECT 70.420 80.995 70.680 82.145 ;
        RECT 70.855 81.070 71.110 81.975 ;
        RECT 71.280 81.385 71.610 82.145 ;
        RECT 71.825 81.215 71.995 81.975 ;
        RECT 65.815 79.595 68.405 80.365 ;
        RECT 69.035 79.595 69.325 80.320 ;
        RECT 70.420 79.595 70.680 80.435 ;
        RECT 70.855 80.340 71.025 81.070 ;
        RECT 71.280 81.045 71.995 81.215 ;
        RECT 72.255 81.055 73.465 82.145 ;
        RECT 73.635 81.550 74.070 81.975 ;
        RECT 74.240 81.720 74.625 82.145 ;
        RECT 73.635 81.380 74.625 81.550 ;
        RECT 71.280 80.835 71.450 81.045 ;
        RECT 71.195 80.505 71.450 80.835 ;
        RECT 70.855 79.765 71.110 80.340 ;
        RECT 71.280 80.315 71.450 80.505 ;
        RECT 71.730 80.495 72.085 80.865 ;
        RECT 72.255 80.345 72.775 80.885 ;
        RECT 72.945 80.515 73.465 81.055 ;
        RECT 73.635 80.505 74.120 81.210 ;
        RECT 74.290 80.835 74.625 81.380 ;
        RECT 74.795 81.185 75.220 81.975 ;
        RECT 75.390 81.550 75.665 81.975 ;
        RECT 75.835 81.720 76.220 82.145 ;
        RECT 75.390 81.355 76.220 81.550 ;
        RECT 74.795 81.005 75.700 81.185 ;
        RECT 74.290 80.505 74.700 80.835 ;
        RECT 74.870 80.505 75.700 81.005 ;
        RECT 75.870 80.835 76.220 81.355 ;
        RECT 76.390 81.185 76.635 81.975 ;
        RECT 76.825 81.550 77.080 81.975 ;
        RECT 77.250 81.720 77.635 82.145 ;
        RECT 76.825 81.355 77.635 81.550 ;
        RECT 76.390 81.005 77.115 81.185 ;
        RECT 75.870 80.505 76.295 80.835 ;
        RECT 76.465 80.505 77.115 81.005 ;
        RECT 77.285 80.835 77.635 81.355 ;
        RECT 77.805 81.005 78.065 81.975 ;
        RECT 77.285 80.505 77.710 80.835 ;
        RECT 71.280 80.145 71.995 80.315 ;
        RECT 71.280 79.595 71.610 79.975 ;
        RECT 71.825 79.765 71.995 80.145 ;
        RECT 72.255 79.595 73.465 80.345 ;
        RECT 74.290 80.335 74.625 80.505 ;
        RECT 74.870 80.335 75.220 80.505 ;
        RECT 75.870 80.335 76.220 80.505 ;
        RECT 76.465 80.335 76.635 80.505 ;
        RECT 77.285 80.335 77.635 80.505 ;
        RECT 77.880 80.335 78.065 81.005 ;
        RECT 78.240 80.995 78.500 82.145 ;
        RECT 78.675 81.070 78.930 81.975 ;
        RECT 79.100 81.385 79.430 82.145 ;
        RECT 79.645 81.215 79.815 81.975 ;
        RECT 73.635 80.165 74.625 80.335 ;
        RECT 73.635 79.765 74.070 80.165 ;
        RECT 74.240 79.595 74.625 79.995 ;
        RECT 74.795 79.765 75.220 80.335 ;
        RECT 75.410 80.165 76.220 80.335 ;
        RECT 75.410 79.765 75.665 80.165 ;
        RECT 75.835 79.595 76.220 79.995 ;
        RECT 76.390 79.765 76.635 80.335 ;
        RECT 76.825 80.165 77.635 80.335 ;
        RECT 76.825 79.765 77.080 80.165 ;
        RECT 77.250 79.595 77.635 79.995 ;
        RECT 77.805 79.765 78.065 80.335 ;
        RECT 78.240 79.595 78.500 80.435 ;
        RECT 78.675 80.340 78.845 81.070 ;
        RECT 79.100 81.045 79.815 81.215 ;
        RECT 79.100 80.835 79.270 81.045 ;
        RECT 80.080 80.995 80.340 82.145 ;
        RECT 80.515 81.070 80.770 81.975 ;
        RECT 80.940 81.385 81.270 82.145 ;
        RECT 81.485 81.215 81.655 81.975 ;
        RECT 79.015 80.505 79.270 80.835 ;
        RECT 78.675 79.765 78.930 80.340 ;
        RECT 79.100 80.315 79.270 80.505 ;
        RECT 79.550 80.495 79.905 80.865 ;
        RECT 79.100 80.145 79.815 80.315 ;
        RECT 79.100 79.595 79.430 79.975 ;
        RECT 79.645 79.765 79.815 80.145 ;
        RECT 80.080 79.595 80.340 80.435 ;
        RECT 80.515 80.340 80.685 81.070 ;
        RECT 80.940 81.045 81.655 81.215 ;
        RECT 80.940 80.835 81.110 81.045 ;
        RECT 81.915 80.980 82.205 82.145 ;
        RECT 83.300 80.995 83.560 82.145 ;
        RECT 83.735 81.070 83.990 81.975 ;
        RECT 84.160 81.385 84.490 82.145 ;
        RECT 84.705 81.215 84.875 81.975 ;
        RECT 80.855 80.505 81.110 80.835 ;
        RECT 80.515 79.765 80.770 80.340 ;
        RECT 80.940 80.315 81.110 80.505 ;
        RECT 81.390 80.495 81.745 80.865 ;
        RECT 80.940 80.145 81.655 80.315 ;
        RECT 80.940 79.595 81.270 79.975 ;
        RECT 81.485 79.765 81.655 80.145 ;
        RECT 81.915 79.595 82.205 80.320 ;
        RECT 83.300 79.595 83.560 80.435 ;
        RECT 83.735 80.340 83.905 81.070 ;
        RECT 84.160 81.045 84.875 81.215 ;
        RECT 85.135 81.055 86.345 82.145 ;
        RECT 84.160 80.835 84.330 81.045 ;
        RECT 84.075 80.505 84.330 80.835 ;
        RECT 83.735 79.765 83.990 80.340 ;
        RECT 84.160 80.315 84.330 80.505 ;
        RECT 84.610 80.495 84.965 80.865 ;
        RECT 85.135 80.345 85.655 80.885 ;
        RECT 85.825 80.515 86.345 81.055 ;
        RECT 86.520 80.995 86.780 82.145 ;
        RECT 86.955 81.070 87.210 81.975 ;
        RECT 87.380 81.385 87.710 82.145 ;
        RECT 87.925 81.215 88.095 81.975 ;
        RECT 84.160 80.145 84.875 80.315 ;
        RECT 84.160 79.595 84.490 79.975 ;
        RECT 84.705 79.765 84.875 80.145 ;
        RECT 85.135 79.595 86.345 80.345 ;
        RECT 86.520 79.595 86.780 80.435 ;
        RECT 86.955 80.340 87.125 81.070 ;
        RECT 87.380 81.045 88.095 81.215 ;
        RECT 88.355 81.055 89.565 82.145 ;
        RECT 87.380 80.835 87.550 81.045 ;
        RECT 87.295 80.505 87.550 80.835 ;
        RECT 86.955 79.765 87.210 80.340 ;
        RECT 87.380 80.315 87.550 80.505 ;
        RECT 87.830 80.495 88.185 80.865 ;
        RECT 88.355 80.345 88.875 80.885 ;
        RECT 89.045 80.515 89.565 81.055 ;
        RECT 89.740 80.995 90.000 82.145 ;
        RECT 90.175 81.070 90.430 81.975 ;
        RECT 90.600 81.385 90.930 82.145 ;
        RECT 91.145 81.215 91.315 81.975 ;
        RECT 87.380 80.145 88.095 80.315 ;
        RECT 87.380 79.595 87.710 79.975 ;
        RECT 87.925 79.765 88.095 80.145 ;
        RECT 88.355 79.595 89.565 80.345 ;
        RECT 89.740 79.595 90.000 80.435 ;
        RECT 90.175 80.340 90.345 81.070 ;
        RECT 90.600 81.045 91.315 81.215 ;
        RECT 91.575 81.055 92.785 82.145 ;
        RECT 90.600 80.835 90.770 81.045 ;
        RECT 90.515 80.505 90.770 80.835 ;
        RECT 90.175 79.765 90.430 80.340 ;
        RECT 90.600 80.315 90.770 80.505 ;
        RECT 91.050 80.495 91.405 80.865 ;
        RECT 91.575 80.345 92.095 80.885 ;
        RECT 92.265 80.515 92.785 81.055 ;
        RECT 92.960 80.995 93.220 82.145 ;
        RECT 93.395 81.070 93.650 81.975 ;
        RECT 93.820 81.385 94.150 82.145 ;
        RECT 94.365 81.215 94.535 81.975 ;
        RECT 90.600 80.145 91.315 80.315 ;
        RECT 90.600 79.595 90.930 79.975 ;
        RECT 91.145 79.765 91.315 80.145 ;
        RECT 91.575 79.595 92.785 80.345 ;
        RECT 92.960 79.595 93.220 80.435 ;
        RECT 93.395 80.340 93.565 81.070 ;
        RECT 93.820 81.045 94.535 81.215 ;
        RECT 93.820 80.835 93.990 81.045 ;
        RECT 94.795 80.980 95.085 82.145 ;
        RECT 96.180 80.995 96.440 82.145 ;
        RECT 96.615 81.070 96.870 81.975 ;
        RECT 97.040 81.385 97.370 82.145 ;
        RECT 97.585 81.215 97.755 81.975 ;
        RECT 93.735 80.505 93.990 80.835 ;
        RECT 93.395 79.765 93.650 80.340 ;
        RECT 93.820 80.315 93.990 80.505 ;
        RECT 94.270 80.495 94.625 80.865 ;
        RECT 93.820 80.145 94.535 80.315 ;
        RECT 93.820 79.595 94.150 79.975 ;
        RECT 94.365 79.765 94.535 80.145 ;
        RECT 94.795 79.595 95.085 80.320 ;
        RECT 96.180 79.595 96.440 80.435 ;
        RECT 96.615 80.340 96.785 81.070 ;
        RECT 97.040 81.045 97.755 81.215 ;
        RECT 98.015 81.055 99.225 82.145 ;
        RECT 97.040 80.835 97.210 81.045 ;
        RECT 96.955 80.505 97.210 80.835 ;
        RECT 96.615 79.765 96.870 80.340 ;
        RECT 97.040 80.315 97.210 80.505 ;
        RECT 97.490 80.495 97.845 80.865 ;
        RECT 98.015 80.345 98.535 80.885 ;
        RECT 98.705 80.515 99.225 81.055 ;
        RECT 99.400 80.995 99.660 82.145 ;
        RECT 99.835 81.070 100.090 81.975 ;
        RECT 100.260 81.385 100.590 82.145 ;
        RECT 100.805 81.215 100.975 81.975 ;
        RECT 97.040 80.145 97.755 80.315 ;
        RECT 97.040 79.595 97.370 79.975 ;
        RECT 97.585 79.765 97.755 80.145 ;
        RECT 98.015 79.595 99.225 80.345 ;
        RECT 99.400 79.595 99.660 80.435 ;
        RECT 99.835 80.340 100.005 81.070 ;
        RECT 100.260 81.045 100.975 81.215 ;
        RECT 100.260 80.835 100.430 81.045 ;
        RECT 102.160 80.995 102.420 82.145 ;
        RECT 102.595 81.070 102.850 81.975 ;
        RECT 103.020 81.385 103.350 82.145 ;
        RECT 103.565 81.215 103.735 81.975 ;
        RECT 100.175 80.505 100.430 80.835 ;
        RECT 99.835 79.765 100.090 80.340 ;
        RECT 100.260 80.315 100.430 80.505 ;
        RECT 100.710 80.495 101.065 80.865 ;
        RECT 100.260 80.145 100.975 80.315 ;
        RECT 100.260 79.595 100.590 79.975 ;
        RECT 100.805 79.765 100.975 80.145 ;
        RECT 102.160 79.595 102.420 80.435 ;
        RECT 102.595 80.340 102.765 81.070 ;
        RECT 103.020 81.045 103.735 81.215 ;
        RECT 104.180 81.175 104.570 81.350 ;
        RECT 105.055 81.345 105.385 82.145 ;
        RECT 105.555 81.355 106.090 81.975 ;
        RECT 103.020 80.835 103.190 81.045 ;
        RECT 104.180 81.005 105.605 81.175 ;
        RECT 102.935 80.505 103.190 80.835 ;
        RECT 102.595 79.765 102.850 80.340 ;
        RECT 103.020 80.315 103.190 80.505 ;
        RECT 103.470 80.495 103.825 80.865 ;
        RECT 103.020 80.145 103.735 80.315 ;
        RECT 104.055 80.275 104.410 80.835 ;
        RECT 103.020 79.595 103.350 79.975 ;
        RECT 103.565 79.765 103.735 80.145 ;
        RECT 104.580 80.105 104.750 81.005 ;
        RECT 104.920 80.275 105.185 80.835 ;
        RECT 105.435 80.505 105.605 81.005 ;
        RECT 105.775 80.335 106.090 81.355 ;
        RECT 106.295 81.055 107.505 82.145 ;
        RECT 104.160 79.595 104.400 80.105 ;
        RECT 104.580 79.775 104.860 80.105 ;
        RECT 105.090 79.595 105.305 80.105 ;
        RECT 105.475 79.765 106.090 80.335 ;
        RECT 106.295 80.345 106.815 80.885 ;
        RECT 106.985 80.515 107.505 81.055 ;
        RECT 107.675 80.980 107.965 82.145 ;
        RECT 108.140 80.995 108.400 82.145 ;
        RECT 108.575 81.070 108.830 81.975 ;
        RECT 109.000 81.385 109.330 82.145 ;
        RECT 109.545 81.215 109.715 81.975 ;
        RECT 106.295 79.595 107.505 80.345 ;
        RECT 107.675 79.595 107.965 80.320 ;
        RECT 108.140 79.595 108.400 80.435 ;
        RECT 108.575 80.340 108.745 81.070 ;
        RECT 109.000 81.045 109.715 81.215 ;
        RECT 109.000 80.835 109.170 81.045 ;
        RECT 109.980 80.995 110.240 82.145 ;
        RECT 110.415 81.070 110.670 81.975 ;
        RECT 110.840 81.385 111.170 82.145 ;
        RECT 111.385 81.215 111.555 81.975 ;
        RECT 108.915 80.505 109.170 80.835 ;
        RECT 108.575 79.765 108.830 80.340 ;
        RECT 109.000 80.315 109.170 80.505 ;
        RECT 109.450 80.495 109.805 80.865 ;
        RECT 109.000 80.145 109.715 80.315 ;
        RECT 109.000 79.595 109.330 79.975 ;
        RECT 109.545 79.765 109.715 80.145 ;
        RECT 109.980 79.595 110.240 80.435 ;
        RECT 110.415 80.340 110.585 81.070 ;
        RECT 110.840 81.045 111.555 81.215 ;
        RECT 110.840 80.835 111.010 81.045 ;
        RECT 112.280 80.995 112.540 82.145 ;
        RECT 112.715 81.070 112.970 81.975 ;
        RECT 113.140 81.385 113.470 82.145 ;
        RECT 113.685 81.215 113.855 81.975 ;
        RECT 110.755 80.505 111.010 80.835 ;
        RECT 110.415 79.765 110.670 80.340 ;
        RECT 110.840 80.315 111.010 80.505 ;
        RECT 111.290 80.495 111.645 80.865 ;
        RECT 110.840 80.145 111.555 80.315 ;
        RECT 110.840 79.595 111.170 79.975 ;
        RECT 111.385 79.765 111.555 80.145 ;
        RECT 112.280 79.595 112.540 80.435 ;
        RECT 112.715 80.340 112.885 81.070 ;
        RECT 113.140 81.045 113.855 81.215 ;
        RECT 114.115 81.055 115.325 82.145 ;
        RECT 113.140 80.835 113.310 81.045 ;
        RECT 113.055 80.505 113.310 80.835 ;
        RECT 112.715 79.765 112.970 80.340 ;
        RECT 113.140 80.315 113.310 80.505 ;
        RECT 113.590 80.495 113.945 80.865 ;
        RECT 114.115 80.345 114.635 80.885 ;
        RECT 114.805 80.515 115.325 81.055 ;
        RECT 115.585 81.215 115.755 81.975 ;
        RECT 115.970 81.385 116.300 82.145 ;
        RECT 115.585 81.045 116.300 81.215 ;
        RECT 116.470 81.070 116.725 81.975 ;
        RECT 115.495 80.495 115.850 80.865 ;
        RECT 116.130 80.835 116.300 81.045 ;
        RECT 116.130 80.505 116.385 80.835 ;
        RECT 113.140 80.145 113.855 80.315 ;
        RECT 113.140 79.595 113.470 79.975 ;
        RECT 113.685 79.765 113.855 80.145 ;
        RECT 114.115 79.595 115.325 80.345 ;
        RECT 116.130 80.315 116.300 80.505 ;
        RECT 116.555 80.340 116.725 81.070 ;
        RECT 116.900 80.995 117.160 82.145 ;
        RECT 117.980 81.175 118.370 81.350 ;
        RECT 118.855 81.345 119.185 82.145 ;
        RECT 119.355 81.355 119.890 81.975 ;
        RECT 117.980 81.005 119.405 81.175 ;
        RECT 115.585 80.145 116.300 80.315 ;
        RECT 115.585 79.765 115.755 80.145 ;
        RECT 115.970 79.595 116.300 79.975 ;
        RECT 116.470 79.765 116.725 80.340 ;
        RECT 116.900 79.595 117.160 80.435 ;
        RECT 117.855 80.275 118.210 80.835 ;
        RECT 118.380 80.105 118.550 81.005 ;
        RECT 118.720 80.275 118.985 80.835 ;
        RECT 119.235 80.505 119.405 81.005 ;
        RECT 119.575 80.335 119.890 81.355 ;
        RECT 120.555 80.980 120.845 82.145 ;
        RECT 121.105 81.215 121.275 81.975 ;
        RECT 121.490 81.385 121.820 82.145 ;
        RECT 121.105 81.045 121.820 81.215 ;
        RECT 121.990 81.070 122.245 81.975 ;
        RECT 121.015 80.495 121.370 80.865 ;
        RECT 121.650 80.835 121.820 81.045 ;
        RECT 121.650 80.505 121.905 80.835 ;
        RECT 117.960 79.595 118.200 80.105 ;
        RECT 118.380 79.775 118.660 80.105 ;
        RECT 118.890 79.595 119.105 80.105 ;
        RECT 119.275 79.765 119.890 80.335 ;
        RECT 120.555 79.595 120.845 80.320 ;
        RECT 121.650 80.315 121.820 80.505 ;
        RECT 122.075 80.340 122.245 81.070 ;
        RECT 122.420 80.995 122.680 82.145 ;
        RECT 122.945 81.215 123.115 81.975 ;
        RECT 123.330 81.385 123.660 82.145 ;
        RECT 122.945 81.045 123.660 81.215 ;
        RECT 123.830 81.070 124.085 81.975 ;
        RECT 122.855 80.495 123.210 80.865 ;
        RECT 123.490 80.835 123.660 81.045 ;
        RECT 123.490 80.505 123.745 80.835 ;
        RECT 121.105 80.145 121.820 80.315 ;
        RECT 121.105 79.765 121.275 80.145 ;
        RECT 121.490 79.595 121.820 79.975 ;
        RECT 121.990 79.765 122.245 80.340 ;
        RECT 122.420 79.595 122.680 80.435 ;
        RECT 123.490 80.315 123.660 80.505 ;
        RECT 123.915 80.340 124.085 81.070 ;
        RECT 124.260 80.995 124.520 82.145 ;
        RECT 125.160 80.995 125.420 82.145 ;
        RECT 125.595 81.070 125.850 81.975 ;
        RECT 126.020 81.385 126.350 82.145 ;
        RECT 126.565 81.215 126.735 81.975 ;
        RECT 122.945 80.145 123.660 80.315 ;
        RECT 122.945 79.765 123.115 80.145 ;
        RECT 123.330 79.595 123.660 79.975 ;
        RECT 123.830 79.765 124.085 80.340 ;
        RECT 124.260 79.595 124.520 80.435 ;
        RECT 125.160 79.595 125.420 80.435 ;
        RECT 125.595 80.340 125.765 81.070 ;
        RECT 126.020 81.045 126.735 81.215 ;
        RECT 126.995 81.055 128.205 82.145 ;
        RECT 126.020 80.835 126.190 81.045 ;
        RECT 125.935 80.505 126.190 80.835 ;
        RECT 125.595 79.765 125.850 80.340 ;
        RECT 126.020 80.315 126.190 80.505 ;
        RECT 126.470 80.495 126.825 80.865 ;
        RECT 126.995 80.345 127.515 80.885 ;
        RECT 127.685 80.515 128.205 81.055 ;
        RECT 128.465 81.215 128.635 81.975 ;
        RECT 128.850 81.385 129.180 82.145 ;
        RECT 128.465 81.045 129.180 81.215 ;
        RECT 129.350 81.070 129.605 81.975 ;
        RECT 128.375 80.495 128.730 80.865 ;
        RECT 129.010 80.835 129.180 81.045 ;
        RECT 129.010 80.505 129.265 80.835 ;
        RECT 126.020 80.145 126.735 80.315 ;
        RECT 126.020 79.595 126.350 79.975 ;
        RECT 126.565 79.765 126.735 80.145 ;
        RECT 126.995 79.595 128.205 80.345 ;
        RECT 129.010 80.315 129.180 80.505 ;
        RECT 129.435 80.340 129.605 81.070 ;
        RECT 129.780 80.995 130.040 82.145 ;
        RECT 130.215 81.055 131.425 82.145 ;
        RECT 128.465 80.145 129.180 80.315 ;
        RECT 128.465 79.765 128.635 80.145 ;
        RECT 128.850 79.595 129.180 79.975 ;
        RECT 129.350 79.765 129.605 80.340 ;
        RECT 129.780 79.595 130.040 80.435 ;
        RECT 130.215 80.345 130.735 80.885 ;
        RECT 130.905 80.515 131.425 81.055 ;
        RECT 131.685 81.215 131.855 81.975 ;
        RECT 132.070 81.385 132.400 82.145 ;
        RECT 131.685 81.045 132.400 81.215 ;
        RECT 132.570 81.070 132.825 81.975 ;
        RECT 131.595 80.495 131.950 80.865 ;
        RECT 132.230 80.835 132.400 81.045 ;
        RECT 132.230 80.505 132.485 80.835 ;
        RECT 130.215 79.595 131.425 80.345 ;
        RECT 132.230 80.315 132.400 80.505 ;
        RECT 132.655 80.340 132.825 81.070 ;
        RECT 133.000 80.995 133.260 82.145 ;
        RECT 133.435 80.980 133.725 82.145 ;
        RECT 134.820 80.995 135.080 82.145 ;
        RECT 135.255 81.070 135.510 81.975 ;
        RECT 135.680 81.385 136.010 82.145 ;
        RECT 136.225 81.215 136.395 81.975 ;
        RECT 131.685 80.145 132.400 80.315 ;
        RECT 131.685 79.765 131.855 80.145 ;
        RECT 132.070 79.595 132.400 79.975 ;
        RECT 132.570 79.765 132.825 80.340 ;
        RECT 133.000 79.595 133.260 80.435 ;
        RECT 133.435 79.595 133.725 80.320 ;
        RECT 134.820 79.595 135.080 80.435 ;
        RECT 135.255 80.340 135.425 81.070 ;
        RECT 135.680 81.045 136.395 81.215 ;
        RECT 136.655 81.055 140.165 82.145 ;
        RECT 140.335 81.055 141.545 82.145 ;
        RECT 135.680 80.835 135.850 81.045 ;
        RECT 135.595 80.505 135.850 80.835 ;
        RECT 135.255 79.765 135.510 80.340 ;
        RECT 135.680 80.315 135.850 80.505 ;
        RECT 136.130 80.495 136.485 80.865 ;
        RECT 136.655 80.365 138.305 80.885 ;
        RECT 138.475 80.535 140.165 81.055 ;
        RECT 135.680 80.145 136.395 80.315 ;
        RECT 135.680 79.595 136.010 79.975 ;
        RECT 136.225 79.765 136.395 80.145 ;
        RECT 136.655 79.595 140.165 80.365 ;
        RECT 140.335 80.345 140.855 80.885 ;
        RECT 141.025 80.515 141.545 81.055 ;
        RECT 141.715 81.055 142.925 82.145 ;
        RECT 141.715 80.515 142.235 81.055 ;
        RECT 142.405 80.345 142.925 80.885 ;
        RECT 140.335 79.595 141.545 80.345 ;
        RECT 141.715 79.595 142.925 80.345 ;
        RECT 17.430 79.425 143.010 79.595 ;
        RECT 12.750 48.645 48.630 48.815 ;
        RECT 12.835 47.555 14.045 48.645 ;
        RECT 14.215 48.210 19.560 48.645 ;
        RECT 12.835 46.845 13.355 47.385 ;
        RECT 13.525 47.015 14.045 47.555 ;
        RECT 12.835 46.095 14.045 46.845 ;
        RECT 15.800 46.640 16.140 47.470 ;
        RECT 17.620 46.960 17.970 48.210 ;
        RECT 20.745 47.715 20.915 48.475 ;
        RECT 21.130 47.885 21.460 48.645 ;
        RECT 20.745 47.545 21.460 47.715 ;
        RECT 21.630 47.570 21.885 48.475 ;
        RECT 20.655 46.995 21.010 47.365 ;
        RECT 21.290 47.335 21.460 47.545 ;
        RECT 21.290 47.005 21.545 47.335 ;
        RECT 21.290 46.815 21.460 47.005 ;
        RECT 21.715 46.840 21.885 47.570 ;
        RECT 22.060 47.495 22.320 48.645 ;
        RECT 22.505 47.845 22.835 48.645 ;
        RECT 23.015 48.305 24.445 48.475 ;
        RECT 23.015 47.675 23.265 48.305 ;
        RECT 22.495 47.505 23.265 47.675 ;
        RECT 20.745 46.645 21.460 46.815 ;
        RECT 14.215 46.095 19.560 46.640 ;
        RECT 20.745 46.265 20.915 46.645 ;
        RECT 21.130 46.095 21.460 46.475 ;
        RECT 21.630 46.265 21.885 46.840 ;
        RECT 22.060 46.095 22.320 46.935 ;
        RECT 22.495 46.835 22.665 47.505 ;
        RECT 22.835 47.005 23.240 47.335 ;
        RECT 23.455 47.005 23.705 48.135 ;
        RECT 23.905 47.335 24.105 48.135 ;
        RECT 24.275 47.625 24.445 48.305 ;
        RECT 24.615 47.795 24.930 48.645 ;
        RECT 25.105 47.845 25.545 48.475 ;
        RECT 24.275 47.455 25.065 47.625 ;
        RECT 23.905 47.005 24.150 47.335 ;
        RECT 24.335 47.005 24.725 47.285 ;
        RECT 24.895 47.005 25.065 47.455 ;
        RECT 25.235 46.835 25.545 47.845 ;
        RECT 25.715 47.480 26.005 48.645 ;
        RECT 27.210 48.015 27.495 48.475 ;
        RECT 27.665 48.185 27.935 48.645 ;
        RECT 27.210 47.795 28.165 48.015 ;
        RECT 27.095 47.065 27.785 47.625 ;
        RECT 27.955 46.895 28.165 47.795 ;
        RECT 22.495 46.265 22.985 46.835 ;
        RECT 23.155 46.665 24.315 46.835 ;
        RECT 23.155 46.265 23.385 46.665 ;
        RECT 23.555 46.095 23.975 46.495 ;
        RECT 24.145 46.265 24.315 46.665 ;
        RECT 24.485 46.095 24.935 46.835 ;
        RECT 25.105 46.275 25.545 46.835 ;
        RECT 25.715 46.095 26.005 46.820 ;
        RECT 27.210 46.725 28.165 46.895 ;
        RECT 28.335 47.625 28.735 48.475 ;
        RECT 28.925 48.015 29.205 48.475 ;
        RECT 29.725 48.185 30.050 48.645 ;
        RECT 28.925 47.795 30.050 48.015 ;
        RECT 28.335 47.065 29.430 47.625 ;
        RECT 29.600 47.335 30.050 47.795 ;
        RECT 30.220 47.505 30.605 48.475 ;
        RECT 27.210 46.265 27.495 46.725 ;
        RECT 27.665 46.095 27.935 46.555 ;
        RECT 28.335 46.265 28.735 47.065 ;
        RECT 29.600 47.005 30.155 47.335 ;
        RECT 29.600 46.895 30.050 47.005 ;
        RECT 28.925 46.725 30.050 46.895 ;
        RECT 30.325 46.835 30.605 47.505 ;
        RECT 31.700 47.495 31.960 48.645 ;
        RECT 32.135 47.570 32.390 48.475 ;
        RECT 32.560 47.885 32.890 48.645 ;
        RECT 33.105 47.715 33.275 48.475 ;
        RECT 33.650 48.015 33.935 48.475 ;
        RECT 34.105 48.185 34.375 48.645 ;
        RECT 33.650 47.795 34.605 48.015 ;
        RECT 28.925 46.265 29.205 46.725 ;
        RECT 29.725 46.095 30.050 46.555 ;
        RECT 30.220 46.265 30.605 46.835 ;
        RECT 31.700 46.095 31.960 46.935 ;
        RECT 32.135 46.840 32.305 47.570 ;
        RECT 32.560 47.545 33.275 47.715 ;
        RECT 32.560 47.335 32.730 47.545 ;
        RECT 32.475 47.005 32.730 47.335 ;
        RECT 32.135 46.265 32.390 46.840 ;
        RECT 32.560 46.815 32.730 47.005 ;
        RECT 33.010 46.995 33.365 47.365 ;
        RECT 33.535 47.065 34.225 47.625 ;
        RECT 34.395 46.895 34.605 47.795 ;
        RECT 32.560 46.645 33.275 46.815 ;
        RECT 32.560 46.095 32.890 46.475 ;
        RECT 33.105 46.265 33.275 46.645 ;
        RECT 33.650 46.725 34.605 46.895 ;
        RECT 34.775 47.625 35.175 48.475 ;
        RECT 35.365 48.015 35.645 48.475 ;
        RECT 36.165 48.185 36.490 48.645 ;
        RECT 35.365 47.795 36.490 48.015 ;
        RECT 34.775 47.065 35.870 47.625 ;
        RECT 36.040 47.335 36.490 47.795 ;
        RECT 36.660 47.505 37.045 48.475 ;
        RECT 37.295 47.715 37.475 48.475 ;
        RECT 37.655 47.885 37.985 48.645 ;
        RECT 37.295 47.545 37.970 47.715 ;
        RECT 38.155 47.570 38.425 48.475 ;
        RECT 33.650 46.265 33.935 46.725 ;
        RECT 34.105 46.095 34.375 46.555 ;
        RECT 34.775 46.265 35.175 47.065 ;
        RECT 36.040 47.005 36.595 47.335 ;
        RECT 36.040 46.895 36.490 47.005 ;
        RECT 35.365 46.725 36.490 46.895 ;
        RECT 36.765 46.835 37.045 47.505 ;
        RECT 37.800 47.400 37.970 47.545 ;
        RECT 37.235 46.995 37.575 47.365 ;
        RECT 37.800 47.070 38.075 47.400 ;
        RECT 35.365 46.265 35.645 46.725 ;
        RECT 36.165 46.095 36.490 46.555 ;
        RECT 36.660 46.265 37.045 46.835 ;
        RECT 37.800 46.815 37.970 47.070 ;
        RECT 37.305 46.645 37.970 46.815 ;
        RECT 38.245 46.770 38.425 47.570 ;
        RECT 38.595 47.480 38.885 48.645 ;
        RECT 39.980 47.495 40.240 48.645 ;
        RECT 40.415 47.570 40.670 48.475 ;
        RECT 40.840 47.885 41.170 48.645 ;
        RECT 41.385 47.715 41.555 48.475 ;
        RECT 37.305 46.265 37.475 46.645 ;
        RECT 37.655 46.095 37.985 46.475 ;
        RECT 38.165 46.265 38.425 46.770 ;
        RECT 38.595 46.095 38.885 46.820 ;
        RECT 39.980 46.095 40.240 46.935 ;
        RECT 40.415 46.840 40.585 47.570 ;
        RECT 40.840 47.545 41.555 47.715 ;
        RECT 41.815 47.555 43.025 48.645 ;
        RECT 40.840 47.335 41.010 47.545 ;
        RECT 40.755 47.005 41.010 47.335 ;
        RECT 40.415 46.265 40.670 46.840 ;
        RECT 40.840 46.815 41.010 47.005 ;
        RECT 41.290 46.995 41.645 47.365 ;
        RECT 41.815 46.845 42.335 47.385 ;
        RECT 42.505 47.015 43.025 47.555 ;
        RECT 43.195 47.570 43.465 48.475 ;
        RECT 43.635 47.885 43.965 48.645 ;
        RECT 44.145 47.715 44.315 48.475 ;
        RECT 40.840 46.645 41.555 46.815 ;
        RECT 40.840 46.095 41.170 46.475 ;
        RECT 41.385 46.265 41.555 46.645 ;
        RECT 41.815 46.095 43.025 46.845 ;
        RECT 43.195 46.770 43.365 47.570 ;
        RECT 43.650 47.545 44.315 47.715 ;
        RECT 44.575 47.570 44.845 48.475 ;
        RECT 45.015 47.885 45.345 48.645 ;
        RECT 45.525 47.715 45.695 48.475 ;
        RECT 43.650 47.400 43.820 47.545 ;
        RECT 43.535 47.070 43.820 47.400 ;
        RECT 43.650 46.815 43.820 47.070 ;
        RECT 44.055 46.995 44.385 47.365 ;
        RECT 43.195 46.265 43.455 46.770 ;
        RECT 43.650 46.645 44.315 46.815 ;
        RECT 43.635 46.095 43.965 46.475 ;
        RECT 44.145 46.265 44.315 46.645 ;
        RECT 44.575 46.770 44.745 47.570 ;
        RECT 45.030 47.545 45.695 47.715 ;
        RECT 45.955 47.570 46.225 48.475 ;
        RECT 46.395 47.885 46.725 48.645 ;
        RECT 46.905 47.715 47.085 48.475 ;
        RECT 45.030 47.400 45.200 47.545 ;
        RECT 44.915 47.070 45.200 47.400 ;
        RECT 45.030 46.815 45.200 47.070 ;
        RECT 45.435 46.995 45.765 47.365 ;
        RECT 44.575 46.265 44.835 46.770 ;
        RECT 45.030 46.645 45.695 46.815 ;
        RECT 45.015 46.095 45.345 46.475 ;
        RECT 45.525 46.265 45.695 46.645 ;
        RECT 45.955 46.770 46.135 47.570 ;
        RECT 46.410 47.545 47.085 47.715 ;
        RECT 47.335 47.555 48.545 48.645 ;
        RECT 46.410 47.400 46.580 47.545 ;
        RECT 46.305 47.070 46.580 47.400 ;
        RECT 46.410 46.815 46.580 47.070 ;
        RECT 46.805 46.995 47.145 47.365 ;
        RECT 47.335 47.015 47.855 47.555 ;
        RECT 48.025 46.845 48.545 47.385 ;
        RECT 45.955 46.265 46.215 46.770 ;
        RECT 46.410 46.645 47.075 46.815 ;
        RECT 46.395 46.095 46.725 46.475 ;
        RECT 46.905 46.265 47.075 46.645 ;
        RECT 47.335 46.095 48.545 46.845 ;
        RECT 12.750 45.925 48.630 46.095 ;
        RECT 12.835 45.175 14.045 45.925 ;
        RECT 12.835 44.635 13.355 45.175 ;
        RECT 14.215 45.155 17.725 45.925 ;
        RECT 18.405 45.270 18.735 45.705 ;
        RECT 18.905 45.315 19.075 45.925 ;
        RECT 18.355 45.185 18.735 45.270 ;
        RECT 19.245 45.185 19.575 45.710 ;
        RECT 19.835 45.395 20.045 45.925 ;
        RECT 20.320 45.475 21.105 45.645 ;
        RECT 21.275 45.475 21.680 45.645 ;
        RECT 13.525 44.465 14.045 45.005 ;
        RECT 14.215 44.635 15.865 45.155 ;
        RECT 18.355 45.145 18.580 45.185 ;
        RECT 16.035 44.465 17.725 44.985 ;
        RECT 12.835 43.375 14.045 44.465 ;
        RECT 14.215 43.375 17.725 44.465 ;
        RECT 18.355 44.565 18.525 45.145 ;
        RECT 19.245 45.015 19.445 45.185 ;
        RECT 20.320 45.015 20.490 45.475 ;
        RECT 18.695 44.685 19.445 45.015 ;
        RECT 19.615 44.685 20.490 45.015 ;
        RECT 18.355 44.515 18.570 44.565 ;
        RECT 18.355 44.435 18.745 44.515 ;
        RECT 18.415 43.590 18.745 44.435 ;
        RECT 19.255 44.480 19.445 44.685 ;
        RECT 18.915 43.375 19.085 44.385 ;
        RECT 19.255 44.105 20.150 44.480 ;
        RECT 19.255 43.545 19.595 44.105 ;
        RECT 19.825 43.375 20.140 43.875 ;
        RECT 20.320 43.845 20.490 44.685 ;
        RECT 20.660 44.975 21.125 45.305 ;
        RECT 21.510 45.245 21.680 45.475 ;
        RECT 21.860 45.425 22.230 45.925 ;
        RECT 22.550 45.475 23.225 45.645 ;
        RECT 23.420 45.475 23.755 45.645 ;
        RECT 20.660 44.015 20.980 44.975 ;
        RECT 21.510 44.945 22.340 45.245 ;
        RECT 21.150 44.045 21.340 44.765 ;
        RECT 21.510 43.875 21.680 44.945 ;
        RECT 22.140 44.915 22.340 44.945 ;
        RECT 21.850 44.695 22.020 44.765 ;
        RECT 22.550 44.695 22.720 45.475 ;
        RECT 23.585 45.335 23.755 45.475 ;
        RECT 23.925 45.465 24.175 45.925 ;
        RECT 21.850 44.525 22.720 44.695 ;
        RECT 22.890 45.055 23.415 45.275 ;
        RECT 23.585 45.205 23.810 45.335 ;
        RECT 21.850 44.435 22.360 44.525 ;
        RECT 20.320 43.675 21.205 43.845 ;
        RECT 21.430 43.545 21.680 43.875 ;
        RECT 21.850 43.375 22.020 44.175 ;
        RECT 22.190 43.820 22.360 44.435 ;
        RECT 22.890 44.355 23.060 45.055 ;
        RECT 22.530 43.990 23.060 44.355 ;
        RECT 23.230 44.290 23.470 44.885 ;
        RECT 23.640 44.100 23.810 45.205 ;
        RECT 23.980 44.345 24.260 45.295 ;
        RECT 23.505 43.970 23.810 44.100 ;
        RECT 22.190 43.650 23.295 43.820 ;
        RECT 23.505 43.545 23.755 43.970 ;
        RECT 23.925 43.375 24.190 43.835 ;
        RECT 24.430 43.545 24.615 45.665 ;
        RECT 24.785 45.545 25.115 45.925 ;
        RECT 25.285 45.375 25.455 45.665 ;
        RECT 24.790 45.205 25.455 45.375 ;
        RECT 25.805 45.375 25.975 45.665 ;
        RECT 26.145 45.545 26.475 45.925 ;
        RECT 25.805 45.205 26.470 45.375 ;
        RECT 24.790 44.215 25.020 45.205 ;
        RECT 25.190 44.385 25.540 45.035 ;
        RECT 25.720 44.385 26.070 45.035 ;
        RECT 26.240 44.215 26.470 45.205 ;
        RECT 24.790 44.045 25.455 44.215 ;
        RECT 24.785 43.375 25.115 43.875 ;
        RECT 25.285 43.545 25.455 44.045 ;
        RECT 25.805 44.045 26.470 44.215 ;
        RECT 25.805 43.545 25.975 44.045 ;
        RECT 26.145 43.375 26.475 43.875 ;
        RECT 26.645 43.545 26.830 45.665 ;
        RECT 27.085 45.465 27.335 45.925 ;
        RECT 27.505 45.475 27.840 45.645 ;
        RECT 28.035 45.475 28.710 45.645 ;
        RECT 27.505 45.335 27.675 45.475 ;
        RECT 27.000 44.345 27.280 45.295 ;
        RECT 27.450 45.205 27.675 45.335 ;
        RECT 27.450 44.100 27.620 45.205 ;
        RECT 27.845 45.055 28.370 45.275 ;
        RECT 27.790 44.290 28.030 44.885 ;
        RECT 28.200 44.355 28.370 45.055 ;
        RECT 28.540 44.695 28.710 45.475 ;
        RECT 29.030 45.425 29.400 45.925 ;
        RECT 29.580 45.475 29.985 45.645 ;
        RECT 30.155 45.475 30.940 45.645 ;
        RECT 29.580 45.245 29.750 45.475 ;
        RECT 28.920 44.945 29.750 45.245 ;
        RECT 30.135 44.975 30.600 45.305 ;
        RECT 28.920 44.915 29.120 44.945 ;
        RECT 29.240 44.695 29.410 44.765 ;
        RECT 28.540 44.525 29.410 44.695 ;
        RECT 28.900 44.435 29.410 44.525 ;
        RECT 27.450 43.970 27.755 44.100 ;
        RECT 28.200 43.990 28.730 44.355 ;
        RECT 27.070 43.375 27.335 43.835 ;
        RECT 27.505 43.545 27.755 43.970 ;
        RECT 28.900 43.820 29.070 44.435 ;
        RECT 27.965 43.650 29.070 43.820 ;
        RECT 29.240 43.375 29.410 44.175 ;
        RECT 29.580 43.875 29.750 44.945 ;
        RECT 29.920 44.045 30.110 44.765 ;
        RECT 30.280 44.015 30.600 44.975 ;
        RECT 30.770 45.015 30.940 45.475 ;
        RECT 31.215 45.395 31.425 45.925 ;
        RECT 31.685 45.185 32.015 45.710 ;
        RECT 32.185 45.315 32.355 45.925 ;
        RECT 32.525 45.270 32.855 45.705 ;
        RECT 32.525 45.185 32.905 45.270 ;
        RECT 31.815 45.015 32.015 45.185 ;
        RECT 32.680 45.145 32.905 45.185 ;
        RECT 30.770 44.685 31.645 45.015 ;
        RECT 31.815 44.685 32.565 45.015 ;
        RECT 29.580 43.545 29.830 43.875 ;
        RECT 30.770 43.845 30.940 44.685 ;
        RECT 31.815 44.480 32.005 44.685 ;
        RECT 32.735 44.565 32.905 45.145 ;
        RECT 32.690 44.515 32.905 44.565 ;
        RECT 31.110 44.105 32.005 44.480 ;
        RECT 32.515 44.435 32.905 44.515 ;
        RECT 33.110 45.185 33.725 45.755 ;
        RECT 33.895 45.415 34.110 45.925 ;
        RECT 34.340 45.415 34.620 45.745 ;
        RECT 34.800 45.415 35.040 45.925 ;
        RECT 30.055 43.675 30.940 43.845 ;
        RECT 31.120 43.375 31.435 43.875 ;
        RECT 31.665 43.545 32.005 44.105 ;
        RECT 32.175 43.375 32.345 44.385 ;
        RECT 32.515 43.590 32.845 44.435 ;
        RECT 33.110 44.165 33.425 45.185 ;
        RECT 33.595 44.515 33.765 45.015 ;
        RECT 34.015 44.685 34.280 45.245 ;
        RECT 34.450 44.515 34.620 45.415 ;
        RECT 35.465 45.375 35.635 45.755 ;
        RECT 35.850 45.545 36.180 45.925 ;
        RECT 34.790 44.685 35.145 45.245 ;
        RECT 35.465 45.205 36.180 45.375 ;
        RECT 35.375 44.655 35.730 45.025 ;
        RECT 36.010 45.015 36.180 45.205 ;
        RECT 36.350 45.180 36.605 45.755 ;
        RECT 36.010 44.685 36.265 45.015 ;
        RECT 33.595 44.345 35.020 44.515 ;
        RECT 36.010 44.475 36.180 44.685 ;
        RECT 33.110 43.545 33.645 44.165 ;
        RECT 33.815 43.375 34.145 44.175 ;
        RECT 34.630 44.170 35.020 44.345 ;
        RECT 35.465 44.305 36.180 44.475 ;
        RECT 36.435 44.450 36.605 45.180 ;
        RECT 36.780 45.085 37.040 45.925 ;
        RECT 37.255 45.105 37.485 45.925 ;
        RECT 37.655 45.125 37.985 45.755 ;
        RECT 37.235 44.685 37.565 44.935 ;
        RECT 37.735 44.525 37.985 45.125 ;
        RECT 38.155 45.105 38.365 45.925 ;
        RECT 38.595 45.200 38.885 45.925 ;
        RECT 39.055 45.185 39.495 45.745 ;
        RECT 39.665 45.185 40.115 45.925 ;
        RECT 40.285 45.355 40.455 45.755 ;
        RECT 40.625 45.525 41.045 45.925 ;
        RECT 41.215 45.355 41.445 45.755 ;
        RECT 40.285 45.185 41.445 45.355 ;
        RECT 41.615 45.185 42.105 45.755 ;
        RECT 35.465 43.545 35.635 44.305 ;
        RECT 35.850 43.375 36.180 44.135 ;
        RECT 36.350 43.545 36.605 44.450 ;
        RECT 36.780 43.375 37.040 44.525 ;
        RECT 37.255 43.375 37.485 44.515 ;
        RECT 37.655 43.545 37.985 44.525 ;
        RECT 38.155 43.375 38.365 44.515 ;
        RECT 38.595 43.375 38.885 44.540 ;
        RECT 39.055 44.175 39.365 45.185 ;
        RECT 39.535 44.565 39.705 45.015 ;
        RECT 39.875 44.735 40.265 45.015 ;
        RECT 40.450 44.685 40.695 45.015 ;
        RECT 39.535 44.395 40.325 44.565 ;
        RECT 39.055 43.545 39.495 44.175 ;
        RECT 39.670 43.375 39.985 44.225 ;
        RECT 40.155 43.715 40.325 44.395 ;
        RECT 40.495 43.885 40.695 44.685 ;
        RECT 40.895 43.885 41.145 45.015 ;
        RECT 41.360 44.685 41.765 45.015 ;
        RECT 41.935 44.515 42.105 45.185 ;
        RECT 42.390 45.295 42.675 45.755 ;
        RECT 42.845 45.465 43.115 45.925 ;
        RECT 42.390 45.125 43.345 45.295 ;
        RECT 41.335 44.345 42.105 44.515 ;
        RECT 42.275 44.395 42.965 44.955 ;
        RECT 41.335 43.715 41.585 44.345 ;
        RECT 43.135 44.225 43.345 45.125 ;
        RECT 40.155 43.545 41.585 43.715 ;
        RECT 41.765 43.375 42.095 44.175 ;
        RECT 42.390 44.005 43.345 44.225 ;
        RECT 43.515 44.955 43.915 45.755 ;
        RECT 44.105 45.295 44.385 45.755 ;
        RECT 44.905 45.465 45.230 45.925 ;
        RECT 44.105 45.125 45.230 45.295 ;
        RECT 45.400 45.185 45.785 45.755 ;
        RECT 44.780 45.015 45.230 45.125 ;
        RECT 43.515 44.395 44.610 44.955 ;
        RECT 44.780 44.685 45.335 45.015 ;
        RECT 42.390 43.545 42.675 44.005 ;
        RECT 42.845 43.375 43.115 43.835 ;
        RECT 43.515 43.545 43.915 44.395 ;
        RECT 44.780 44.225 45.230 44.685 ;
        RECT 45.505 44.515 45.785 45.185 ;
        RECT 44.105 44.005 45.230 44.225 ;
        RECT 44.105 43.545 44.385 44.005 ;
        RECT 44.905 43.375 45.230 43.835 ;
        RECT 45.400 43.545 45.785 44.515 ;
        RECT 45.955 45.250 46.215 45.755 ;
        RECT 46.395 45.545 46.725 45.925 ;
        RECT 46.905 45.375 47.075 45.755 ;
        RECT 45.955 44.450 46.135 45.250 ;
        RECT 46.410 45.205 47.075 45.375 ;
        RECT 46.410 44.950 46.580 45.205 ;
        RECT 47.335 45.175 48.545 45.925 ;
        RECT 46.305 44.620 46.580 44.950 ;
        RECT 46.805 44.655 47.145 45.025 ;
        RECT 46.410 44.475 46.580 44.620 ;
        RECT 45.955 43.545 46.225 44.450 ;
        RECT 46.410 44.305 47.085 44.475 ;
        RECT 46.395 43.375 46.725 44.135 ;
        RECT 46.905 43.545 47.085 44.305 ;
        RECT 47.335 44.465 47.855 45.005 ;
        RECT 48.025 44.635 48.545 45.175 ;
        RECT 47.335 43.375 48.545 44.465 ;
        RECT 12.750 43.205 48.630 43.375 ;
        RECT 12.835 42.115 14.045 43.205 ;
        RECT 14.305 42.535 14.475 43.035 ;
        RECT 14.645 42.705 14.975 43.205 ;
        RECT 14.305 42.365 14.970 42.535 ;
        RECT 12.835 41.405 13.355 41.945 ;
        RECT 13.525 41.575 14.045 42.115 ;
        RECT 14.220 41.545 14.570 42.195 ;
        RECT 12.835 40.655 14.045 41.405 ;
        RECT 14.740 41.375 14.970 42.365 ;
        RECT 14.305 41.205 14.970 41.375 ;
        RECT 14.305 40.915 14.475 41.205 ;
        RECT 14.645 40.655 14.975 41.035 ;
        RECT 15.145 40.915 15.330 43.035 ;
        RECT 15.570 42.745 15.835 43.205 ;
        RECT 16.005 42.610 16.255 43.035 ;
        RECT 16.465 42.760 17.570 42.930 ;
        RECT 15.950 42.480 16.255 42.610 ;
        RECT 15.500 41.285 15.780 42.235 ;
        RECT 15.950 41.375 16.120 42.480 ;
        RECT 16.290 41.695 16.530 42.290 ;
        RECT 16.700 42.225 17.230 42.590 ;
        RECT 16.700 41.525 16.870 42.225 ;
        RECT 17.400 42.145 17.570 42.760 ;
        RECT 17.740 42.405 17.910 43.205 ;
        RECT 18.080 42.705 18.330 43.035 ;
        RECT 18.555 42.735 19.440 42.905 ;
        RECT 17.400 42.055 17.910 42.145 ;
        RECT 15.950 41.245 16.175 41.375 ;
        RECT 16.345 41.305 16.870 41.525 ;
        RECT 17.040 41.885 17.910 42.055 ;
        RECT 15.585 40.655 15.835 41.115 ;
        RECT 16.005 41.105 16.175 41.245 ;
        RECT 17.040 41.105 17.210 41.885 ;
        RECT 17.740 41.815 17.910 41.885 ;
        RECT 17.420 41.635 17.620 41.665 ;
        RECT 18.080 41.635 18.250 42.705 ;
        RECT 18.420 41.815 18.610 42.535 ;
        RECT 17.420 41.335 18.250 41.635 ;
        RECT 18.780 41.605 19.100 42.565 ;
        RECT 16.005 40.935 16.340 41.105 ;
        RECT 16.535 40.935 17.210 41.105 ;
        RECT 17.530 40.655 17.900 41.155 ;
        RECT 18.080 41.105 18.250 41.335 ;
        RECT 18.635 41.275 19.100 41.605 ;
        RECT 19.270 41.895 19.440 42.735 ;
        RECT 19.620 42.705 19.935 43.205 ;
        RECT 20.165 42.475 20.505 43.035 ;
        RECT 19.610 42.100 20.505 42.475 ;
        RECT 20.675 42.195 20.845 43.205 ;
        RECT 20.315 41.895 20.505 42.100 ;
        RECT 21.015 42.145 21.345 42.990 ;
        RECT 21.015 42.065 21.405 42.145 ;
        RECT 21.190 42.015 21.405 42.065 ;
        RECT 19.270 41.565 20.145 41.895 ;
        RECT 20.315 41.565 21.065 41.895 ;
        RECT 19.270 41.105 19.440 41.565 ;
        RECT 20.315 41.395 20.515 41.565 ;
        RECT 21.235 41.435 21.405 42.015 ;
        RECT 21.180 41.395 21.405 41.435 ;
        RECT 18.080 40.935 18.485 41.105 ;
        RECT 18.655 40.935 19.440 41.105 ;
        RECT 19.715 40.655 19.925 41.185 ;
        RECT 20.185 40.870 20.515 41.395 ;
        RECT 21.025 41.310 21.405 41.395 ;
        RECT 21.575 42.065 21.960 43.035 ;
        RECT 22.130 42.745 22.455 43.205 ;
        RECT 22.975 42.575 23.255 43.035 ;
        RECT 22.130 42.355 23.255 42.575 ;
        RECT 21.575 41.395 21.855 42.065 ;
        RECT 22.130 41.895 22.580 42.355 ;
        RECT 23.445 42.185 23.845 43.035 ;
        RECT 24.245 42.745 24.515 43.205 ;
        RECT 24.685 42.575 24.970 43.035 ;
        RECT 22.025 41.565 22.580 41.895 ;
        RECT 22.750 41.625 23.845 42.185 ;
        RECT 22.130 41.455 22.580 41.565 ;
        RECT 20.685 40.655 20.855 41.265 ;
        RECT 21.025 40.875 21.355 41.310 ;
        RECT 21.575 40.825 21.960 41.395 ;
        RECT 22.130 41.285 23.255 41.455 ;
        RECT 22.130 40.655 22.455 41.115 ;
        RECT 22.975 40.825 23.255 41.285 ;
        RECT 23.445 40.825 23.845 41.625 ;
        RECT 24.015 42.355 24.970 42.575 ;
        RECT 24.015 41.455 24.225 42.355 ;
        RECT 24.395 41.625 25.085 42.185 ;
        RECT 25.715 42.040 26.005 43.205 ;
        RECT 26.180 42.065 26.515 43.035 ;
        RECT 26.685 42.065 26.855 43.205 ;
        RECT 27.025 42.865 29.055 43.035 ;
        RECT 24.015 41.285 24.970 41.455 ;
        RECT 26.180 41.395 26.350 42.065 ;
        RECT 27.025 41.895 27.195 42.865 ;
        RECT 26.520 41.565 26.775 41.895 ;
        RECT 27.000 41.565 27.195 41.895 ;
        RECT 27.365 42.525 28.490 42.695 ;
        RECT 26.605 41.395 26.775 41.565 ;
        RECT 27.365 41.395 27.535 42.525 ;
        RECT 24.245 40.655 24.515 41.115 ;
        RECT 24.685 40.825 24.970 41.285 ;
        RECT 25.715 40.655 26.005 41.380 ;
        RECT 26.180 40.825 26.435 41.395 ;
        RECT 26.605 41.225 27.535 41.395 ;
        RECT 27.705 42.185 28.715 42.355 ;
        RECT 27.705 41.385 27.875 42.185 ;
        RECT 28.080 41.845 28.355 41.985 ;
        RECT 28.075 41.675 28.355 41.845 ;
        RECT 27.360 41.190 27.535 41.225 ;
        RECT 26.605 40.655 26.935 41.055 ;
        RECT 27.360 40.825 27.890 41.190 ;
        RECT 28.080 40.825 28.355 41.675 ;
        RECT 28.525 40.825 28.715 42.185 ;
        RECT 28.885 42.200 29.055 42.865 ;
        RECT 29.225 42.445 29.395 43.205 ;
        RECT 29.630 42.445 30.145 42.855 ;
        RECT 28.885 42.010 29.635 42.200 ;
        RECT 29.805 41.635 30.145 42.445 ;
        RECT 30.960 42.235 31.350 42.410 ;
        RECT 31.835 42.405 32.165 43.205 ;
        RECT 32.335 42.415 32.870 43.035 ;
        RECT 30.960 42.065 32.385 42.235 ;
        RECT 28.915 41.465 30.145 41.635 ;
        RECT 28.895 40.655 29.405 41.190 ;
        RECT 29.625 40.860 29.870 41.465 ;
        RECT 30.835 41.335 31.190 41.895 ;
        RECT 31.360 41.165 31.530 42.065 ;
        RECT 31.700 41.335 31.965 41.895 ;
        RECT 32.215 41.565 32.385 42.065 ;
        RECT 32.555 41.395 32.870 42.415 ;
        RECT 33.135 42.065 33.345 43.205 ;
        RECT 33.515 42.055 33.845 43.035 ;
        RECT 34.015 42.065 34.245 43.205 ;
        RECT 34.545 42.535 34.715 43.035 ;
        RECT 34.885 42.705 35.215 43.205 ;
        RECT 34.545 42.365 35.210 42.535 ;
        RECT 30.940 40.655 31.180 41.165 ;
        RECT 31.360 40.835 31.640 41.165 ;
        RECT 31.870 40.655 32.085 41.165 ;
        RECT 32.255 40.825 32.870 41.395 ;
        RECT 33.135 40.655 33.345 41.475 ;
        RECT 33.515 41.455 33.765 42.055 ;
        RECT 33.935 41.645 34.265 41.895 ;
        RECT 34.460 41.545 34.810 42.195 ;
        RECT 33.515 40.825 33.845 41.455 ;
        RECT 34.015 40.655 34.245 41.475 ;
        RECT 34.980 41.375 35.210 42.365 ;
        RECT 34.545 41.205 35.210 41.375 ;
        RECT 34.545 40.915 34.715 41.205 ;
        RECT 34.885 40.655 35.215 41.035 ;
        RECT 35.385 40.915 35.570 43.035 ;
        RECT 35.810 42.745 36.075 43.205 ;
        RECT 36.245 42.610 36.495 43.035 ;
        RECT 36.705 42.760 37.810 42.930 ;
        RECT 36.190 42.480 36.495 42.610 ;
        RECT 35.740 41.285 36.020 42.235 ;
        RECT 36.190 41.375 36.360 42.480 ;
        RECT 36.530 41.695 36.770 42.290 ;
        RECT 36.940 42.225 37.470 42.590 ;
        RECT 36.940 41.525 37.110 42.225 ;
        RECT 37.640 42.145 37.810 42.760 ;
        RECT 37.980 42.405 38.150 43.205 ;
        RECT 38.320 42.705 38.570 43.035 ;
        RECT 38.795 42.735 39.680 42.905 ;
        RECT 37.640 42.055 38.150 42.145 ;
        RECT 36.190 41.245 36.415 41.375 ;
        RECT 36.585 41.305 37.110 41.525 ;
        RECT 37.280 41.885 38.150 42.055 ;
        RECT 35.825 40.655 36.075 41.115 ;
        RECT 36.245 41.105 36.415 41.245 ;
        RECT 37.280 41.105 37.450 41.885 ;
        RECT 37.980 41.815 38.150 41.885 ;
        RECT 37.660 41.635 37.860 41.665 ;
        RECT 38.320 41.635 38.490 42.705 ;
        RECT 38.660 41.815 38.850 42.535 ;
        RECT 37.660 41.335 38.490 41.635 ;
        RECT 39.020 41.605 39.340 42.565 ;
        RECT 36.245 40.935 36.580 41.105 ;
        RECT 36.775 40.935 37.450 41.105 ;
        RECT 37.770 40.655 38.140 41.155 ;
        RECT 38.320 41.105 38.490 41.335 ;
        RECT 38.875 41.275 39.340 41.605 ;
        RECT 39.510 41.895 39.680 42.735 ;
        RECT 39.860 42.705 40.175 43.205 ;
        RECT 40.405 42.475 40.745 43.035 ;
        RECT 39.850 42.100 40.745 42.475 ;
        RECT 40.915 42.195 41.085 43.205 ;
        RECT 40.555 41.895 40.745 42.100 ;
        RECT 41.255 42.145 41.585 42.990 ;
        RECT 42.460 42.235 42.850 42.410 ;
        RECT 43.335 42.405 43.665 43.205 ;
        RECT 43.835 42.415 44.370 43.035 ;
        RECT 41.255 42.065 41.645 42.145 ;
        RECT 42.460 42.065 43.885 42.235 ;
        RECT 41.430 42.015 41.645 42.065 ;
        RECT 39.510 41.565 40.385 41.895 ;
        RECT 40.555 41.565 41.305 41.895 ;
        RECT 39.510 41.105 39.680 41.565 ;
        RECT 40.555 41.395 40.755 41.565 ;
        RECT 41.475 41.435 41.645 42.015 ;
        RECT 41.420 41.395 41.645 41.435 ;
        RECT 38.320 40.935 38.725 41.105 ;
        RECT 38.895 40.935 39.680 41.105 ;
        RECT 39.955 40.655 40.165 41.185 ;
        RECT 40.425 40.870 40.755 41.395 ;
        RECT 41.265 41.310 41.645 41.395 ;
        RECT 42.335 41.335 42.690 41.895 ;
        RECT 40.925 40.655 41.095 41.265 ;
        RECT 41.265 40.875 41.595 41.310 ;
        RECT 42.860 41.165 43.030 42.065 ;
        RECT 43.200 41.335 43.465 41.895 ;
        RECT 43.715 41.565 43.885 42.065 ;
        RECT 44.055 41.395 44.370 42.415 ;
        RECT 44.665 42.275 44.835 43.035 ;
        RECT 45.015 42.445 45.345 43.205 ;
        RECT 44.665 42.105 45.330 42.275 ;
        RECT 45.515 42.130 45.785 43.035 ;
        RECT 45.160 41.960 45.330 42.105 ;
        RECT 44.595 41.555 44.925 41.925 ;
        RECT 45.160 41.630 45.445 41.960 ;
        RECT 42.440 40.655 42.680 41.165 ;
        RECT 42.860 40.835 43.140 41.165 ;
        RECT 43.370 40.655 43.585 41.165 ;
        RECT 43.755 40.825 44.370 41.395 ;
        RECT 45.160 41.375 45.330 41.630 ;
        RECT 44.665 41.205 45.330 41.375 ;
        RECT 45.615 41.330 45.785 42.130 ;
        RECT 44.665 40.825 44.835 41.205 ;
        RECT 45.015 40.655 45.345 41.035 ;
        RECT 45.525 40.825 45.785 41.330 ;
        RECT 45.955 42.130 46.225 43.035 ;
        RECT 46.395 42.445 46.725 43.205 ;
        RECT 46.905 42.275 47.085 43.035 ;
        RECT 45.955 41.330 46.135 42.130 ;
        RECT 46.410 42.105 47.085 42.275 ;
        RECT 47.335 42.115 48.545 43.205 ;
        RECT 46.410 41.960 46.580 42.105 ;
        RECT 46.305 41.630 46.580 41.960 ;
        RECT 46.410 41.375 46.580 41.630 ;
        RECT 46.805 41.555 47.145 41.925 ;
        RECT 47.335 41.575 47.855 42.115 ;
        RECT 48.025 41.405 48.545 41.945 ;
        RECT 45.955 40.825 46.215 41.330 ;
        RECT 46.410 41.205 47.075 41.375 ;
        RECT 46.395 40.655 46.725 41.035 ;
        RECT 46.905 40.825 47.075 41.205 ;
        RECT 47.335 40.655 48.545 41.405 ;
        RECT 12.750 40.485 48.630 40.655 ;
        RECT 12.835 39.735 14.045 40.485 ;
        RECT 12.835 39.195 13.355 39.735 ;
        RECT 14.220 39.645 14.480 40.485 ;
        RECT 14.655 39.740 14.910 40.315 ;
        RECT 15.080 40.105 15.410 40.485 ;
        RECT 15.625 39.935 15.795 40.315 ;
        RECT 15.080 39.765 15.795 39.935 ;
        RECT 13.525 39.025 14.045 39.565 ;
        RECT 12.835 37.935 14.045 39.025 ;
        RECT 14.220 37.935 14.480 39.085 ;
        RECT 14.655 39.010 14.825 39.740 ;
        RECT 15.080 39.575 15.250 39.765 ;
        RECT 16.060 39.745 16.315 40.315 ;
        RECT 16.485 40.085 16.815 40.485 ;
        RECT 17.240 39.950 17.770 40.315 ;
        RECT 17.960 40.145 18.235 40.315 ;
        RECT 17.955 39.975 18.235 40.145 ;
        RECT 17.240 39.915 17.415 39.950 ;
        RECT 16.485 39.745 17.415 39.915 ;
        RECT 14.995 39.245 15.250 39.575 ;
        RECT 15.080 39.035 15.250 39.245 ;
        RECT 15.530 39.215 15.885 39.585 ;
        RECT 16.060 39.075 16.230 39.745 ;
        RECT 16.485 39.575 16.655 39.745 ;
        RECT 16.400 39.245 16.655 39.575 ;
        RECT 16.880 39.245 17.075 39.575 ;
        RECT 14.655 38.105 14.910 39.010 ;
        RECT 15.080 38.865 15.795 39.035 ;
        RECT 15.080 37.935 15.410 38.695 ;
        RECT 15.625 38.105 15.795 38.865 ;
        RECT 16.060 38.105 16.395 39.075 ;
        RECT 16.565 37.935 16.735 39.075 ;
        RECT 16.905 38.275 17.075 39.245 ;
        RECT 17.245 38.615 17.415 39.745 ;
        RECT 17.585 38.955 17.755 39.755 ;
        RECT 17.960 39.155 18.235 39.975 ;
        RECT 18.405 38.955 18.595 40.315 ;
        RECT 18.775 39.950 19.285 40.485 ;
        RECT 19.505 39.675 19.750 40.280 ;
        RECT 20.195 39.735 21.405 40.485 ;
        RECT 21.665 40.005 21.965 40.485 ;
        RECT 22.135 39.835 22.395 40.290 ;
        RECT 22.565 40.005 22.825 40.485 ;
        RECT 23.005 39.835 23.265 40.290 ;
        RECT 23.435 40.005 23.685 40.485 ;
        RECT 23.865 39.835 24.125 40.290 ;
        RECT 24.295 40.005 24.545 40.485 ;
        RECT 24.725 39.835 24.985 40.290 ;
        RECT 25.155 40.005 25.400 40.485 ;
        RECT 25.570 39.835 25.845 40.290 ;
        RECT 26.015 40.005 26.260 40.485 ;
        RECT 26.430 39.835 26.690 40.290 ;
        RECT 26.860 40.005 27.120 40.485 ;
        RECT 27.290 39.835 27.550 40.290 ;
        RECT 27.720 40.005 27.980 40.485 ;
        RECT 28.150 39.835 28.410 40.290 ;
        RECT 28.580 39.925 28.840 40.485 ;
        RECT 18.795 39.505 20.025 39.675 ;
        RECT 17.585 38.785 18.595 38.955 ;
        RECT 18.765 38.940 19.515 39.130 ;
        RECT 17.245 38.445 18.370 38.615 ;
        RECT 18.765 38.275 18.935 38.940 ;
        RECT 19.685 38.695 20.025 39.505 ;
        RECT 20.195 39.195 20.715 39.735 ;
        RECT 21.665 39.665 28.410 39.835 ;
        RECT 20.885 39.025 21.405 39.565 ;
        RECT 16.905 38.105 18.935 38.275 ;
        RECT 19.105 37.935 19.275 38.695 ;
        RECT 19.510 38.285 20.025 38.695 ;
        RECT 20.195 37.935 21.405 39.025 ;
        RECT 21.665 39.075 22.830 39.665 ;
        RECT 29.010 39.495 29.260 40.305 ;
        RECT 29.440 39.960 29.700 40.485 ;
        RECT 29.870 39.495 30.120 40.305 ;
        RECT 30.300 39.975 30.605 40.485 ;
        RECT 23.000 39.245 30.120 39.495 ;
        RECT 30.290 39.245 30.605 39.805 ;
        RECT 30.775 39.745 31.160 40.315 ;
        RECT 31.330 40.025 31.655 40.485 ;
        RECT 32.175 39.855 32.455 40.315 ;
        RECT 21.665 38.850 28.410 39.075 ;
        RECT 21.665 37.935 21.935 38.680 ;
        RECT 22.105 38.110 22.395 38.850 ;
        RECT 23.005 38.835 28.410 38.850 ;
        RECT 22.565 37.940 22.820 38.665 ;
        RECT 23.005 38.110 23.265 38.835 ;
        RECT 23.435 37.940 23.680 38.665 ;
        RECT 23.865 38.110 24.125 38.835 ;
        RECT 24.295 37.940 24.540 38.665 ;
        RECT 24.725 38.110 24.985 38.835 ;
        RECT 25.155 37.940 25.400 38.665 ;
        RECT 25.570 38.110 25.830 38.835 ;
        RECT 26.000 37.940 26.260 38.665 ;
        RECT 26.430 38.110 26.690 38.835 ;
        RECT 26.860 37.940 27.120 38.665 ;
        RECT 27.290 38.110 27.550 38.835 ;
        RECT 27.720 37.940 27.980 38.665 ;
        RECT 28.150 38.110 28.410 38.835 ;
        RECT 28.580 37.940 28.840 38.735 ;
        RECT 29.010 38.110 29.260 39.245 ;
        RECT 22.565 37.935 28.840 37.940 ;
        RECT 29.440 37.935 29.700 38.745 ;
        RECT 29.875 38.105 30.120 39.245 ;
        RECT 30.775 39.075 31.055 39.745 ;
        RECT 31.330 39.685 32.455 39.855 ;
        RECT 31.330 39.575 31.780 39.685 ;
        RECT 31.225 39.245 31.780 39.575 ;
        RECT 32.645 39.515 33.045 40.315 ;
        RECT 33.445 40.025 33.715 40.485 ;
        RECT 33.885 39.855 34.170 40.315 ;
        RECT 30.300 37.935 30.595 38.745 ;
        RECT 30.775 38.105 31.160 39.075 ;
        RECT 31.330 38.785 31.780 39.245 ;
        RECT 31.950 38.955 33.045 39.515 ;
        RECT 31.330 38.565 32.455 38.785 ;
        RECT 31.330 37.935 31.655 38.395 ;
        RECT 32.175 38.105 32.455 38.565 ;
        RECT 32.645 38.105 33.045 38.955 ;
        RECT 33.215 39.685 34.170 39.855 ;
        RECT 34.455 39.735 35.665 40.485 ;
        RECT 35.845 39.985 36.175 40.485 ;
        RECT 36.375 39.915 36.545 40.265 ;
        RECT 36.745 40.085 37.075 40.485 ;
        RECT 37.245 39.915 37.415 40.265 ;
        RECT 37.585 40.085 37.965 40.485 ;
        RECT 33.215 38.785 33.425 39.685 ;
        RECT 33.595 38.955 34.285 39.515 ;
        RECT 34.455 39.195 34.975 39.735 ;
        RECT 35.145 39.025 35.665 39.565 ;
        RECT 35.840 39.245 36.190 39.815 ;
        RECT 36.375 39.745 37.985 39.915 ;
        RECT 38.155 39.810 38.425 40.155 ;
        RECT 37.815 39.575 37.985 39.745 ;
        RECT 33.215 38.565 34.170 38.785 ;
        RECT 33.445 37.935 33.715 38.395 ;
        RECT 33.885 38.105 34.170 38.565 ;
        RECT 34.455 37.935 35.665 39.025 ;
        RECT 35.840 38.785 36.160 39.075 ;
        RECT 36.360 38.955 37.070 39.575 ;
        RECT 37.240 39.245 37.645 39.575 ;
        RECT 37.815 39.245 38.085 39.575 ;
        RECT 37.815 39.075 37.985 39.245 ;
        RECT 38.255 39.075 38.425 39.810 ;
        RECT 38.595 39.760 38.885 40.485 ;
        RECT 39.055 39.745 39.415 40.120 ;
        RECT 39.680 39.745 39.850 40.485 ;
        RECT 40.130 39.915 40.300 40.120 ;
        RECT 40.130 39.745 40.670 39.915 ;
        RECT 37.260 38.905 37.985 39.075 ;
        RECT 37.260 38.785 37.430 38.905 ;
        RECT 35.840 38.615 37.430 38.785 ;
        RECT 35.840 38.155 37.495 38.445 ;
        RECT 37.665 37.935 37.945 38.735 ;
        RECT 38.155 38.105 38.425 39.075 ;
        RECT 38.595 37.935 38.885 39.100 ;
        RECT 39.055 39.090 39.310 39.745 ;
        RECT 39.480 39.245 39.830 39.575 ;
        RECT 40.000 39.245 40.330 39.575 ;
        RECT 39.055 38.105 39.395 39.090 ;
        RECT 39.565 38.705 39.830 39.245 ;
        RECT 40.500 39.045 40.670 39.745 ;
        RECT 40.045 38.875 40.670 39.045 ;
        RECT 40.840 39.115 41.010 40.315 ;
        RECT 41.240 39.835 41.570 40.315 ;
        RECT 41.740 40.015 41.910 40.485 ;
        RECT 42.080 39.835 42.410 40.300 ;
        RECT 41.240 39.665 42.410 39.835 ;
        RECT 42.735 39.745 43.095 40.120 ;
        RECT 43.360 39.745 43.530 40.485 ;
        RECT 43.810 39.915 43.980 40.120 ;
        RECT 43.810 39.745 44.350 39.915 ;
        RECT 41.180 39.285 41.750 39.495 ;
        RECT 41.920 39.285 42.565 39.495 ;
        RECT 40.840 38.705 41.545 39.115 ;
        RECT 42.735 39.090 42.990 39.745 ;
        RECT 43.160 39.245 43.510 39.575 ;
        RECT 43.680 39.245 44.010 39.575 ;
        RECT 39.565 38.535 41.545 38.705 ;
        RECT 39.565 37.935 39.975 38.365 ;
        RECT 40.720 37.935 41.050 38.355 ;
        RECT 41.220 38.105 41.545 38.535 ;
        RECT 42.020 37.935 42.350 39.035 ;
        RECT 42.735 38.105 43.075 39.090 ;
        RECT 43.245 38.705 43.510 39.245 ;
        RECT 44.180 39.045 44.350 39.745 ;
        RECT 43.725 38.875 44.350 39.045 ;
        RECT 44.520 39.115 44.690 40.315 ;
        RECT 44.920 39.835 45.250 40.315 ;
        RECT 45.420 40.015 45.590 40.485 ;
        RECT 45.760 39.835 46.090 40.300 ;
        RECT 44.920 39.665 46.090 39.835 ;
        RECT 47.335 39.735 48.545 40.485 ;
        RECT 44.860 39.285 45.430 39.495 ;
        RECT 45.600 39.285 46.245 39.495 ;
        RECT 44.520 38.705 45.225 39.115 ;
        RECT 43.245 38.535 45.225 38.705 ;
        RECT 43.245 37.935 43.655 38.365 ;
        RECT 44.400 37.935 44.730 38.355 ;
        RECT 44.900 38.105 45.225 38.535 ;
        RECT 45.700 37.935 46.030 39.035 ;
        RECT 47.335 39.025 47.855 39.565 ;
        RECT 48.025 39.195 48.545 39.735 ;
        RECT 47.335 37.935 48.545 39.025 ;
        RECT 12.750 37.765 48.630 37.935 ;
        RECT 12.835 36.675 14.045 37.765 ;
        RECT 12.835 35.965 13.355 36.505 ;
        RECT 13.525 36.135 14.045 36.675 ;
        RECT 14.220 36.625 14.555 37.595 ;
        RECT 14.725 36.625 14.895 37.765 ;
        RECT 15.065 37.425 17.095 37.595 ;
        RECT 12.835 35.215 14.045 35.965 ;
        RECT 14.220 35.955 14.390 36.625 ;
        RECT 15.065 36.455 15.235 37.425 ;
        RECT 14.560 36.125 14.815 36.455 ;
        RECT 15.040 36.125 15.235 36.455 ;
        RECT 15.405 37.085 16.530 37.255 ;
        RECT 14.645 35.955 14.815 36.125 ;
        RECT 15.405 35.955 15.575 37.085 ;
        RECT 14.220 35.385 14.475 35.955 ;
        RECT 14.645 35.785 15.575 35.955 ;
        RECT 15.745 36.745 16.755 36.915 ;
        RECT 15.745 35.945 15.915 36.745 ;
        RECT 15.400 35.750 15.575 35.785 ;
        RECT 14.645 35.215 14.975 35.615 ;
        RECT 15.400 35.385 15.930 35.750 ;
        RECT 16.120 35.725 16.395 36.545 ;
        RECT 16.115 35.555 16.395 35.725 ;
        RECT 16.120 35.385 16.395 35.555 ;
        RECT 16.565 35.385 16.755 36.745 ;
        RECT 16.925 36.760 17.095 37.425 ;
        RECT 17.265 37.005 17.435 37.765 ;
        RECT 17.670 37.005 18.185 37.415 ;
        RECT 16.925 36.570 17.675 36.760 ;
        RECT 17.845 36.195 18.185 37.005 ;
        RECT 18.445 37.095 18.615 37.595 ;
        RECT 18.785 37.265 19.115 37.765 ;
        RECT 18.445 36.925 19.110 37.095 ;
        RECT 16.955 36.025 18.185 36.195 ;
        RECT 18.360 36.105 18.710 36.755 ;
        RECT 16.935 35.215 17.445 35.750 ;
        RECT 17.665 35.420 17.910 36.025 ;
        RECT 18.880 35.935 19.110 36.925 ;
        RECT 18.445 35.765 19.110 35.935 ;
        RECT 18.445 35.475 18.615 35.765 ;
        RECT 18.785 35.215 19.115 35.595 ;
        RECT 19.285 35.475 19.470 37.595 ;
        RECT 19.710 37.305 19.975 37.765 ;
        RECT 20.145 37.170 20.395 37.595 ;
        RECT 20.605 37.320 21.710 37.490 ;
        RECT 20.090 37.040 20.395 37.170 ;
        RECT 19.640 35.845 19.920 36.795 ;
        RECT 20.090 35.935 20.260 37.040 ;
        RECT 20.430 36.255 20.670 36.850 ;
        RECT 20.840 36.785 21.370 37.150 ;
        RECT 20.840 36.085 21.010 36.785 ;
        RECT 21.540 36.705 21.710 37.320 ;
        RECT 21.880 36.965 22.050 37.765 ;
        RECT 22.220 37.265 22.470 37.595 ;
        RECT 22.695 37.295 23.580 37.465 ;
        RECT 21.540 36.615 22.050 36.705 ;
        RECT 20.090 35.805 20.315 35.935 ;
        RECT 20.485 35.865 21.010 36.085 ;
        RECT 21.180 36.445 22.050 36.615 ;
        RECT 19.725 35.215 19.975 35.675 ;
        RECT 20.145 35.665 20.315 35.805 ;
        RECT 21.180 35.665 21.350 36.445 ;
        RECT 21.880 36.375 22.050 36.445 ;
        RECT 21.560 36.195 21.760 36.225 ;
        RECT 22.220 36.195 22.390 37.265 ;
        RECT 22.560 36.375 22.750 37.095 ;
        RECT 21.560 35.895 22.390 36.195 ;
        RECT 22.920 36.165 23.240 37.125 ;
        RECT 20.145 35.495 20.480 35.665 ;
        RECT 20.675 35.495 21.350 35.665 ;
        RECT 21.670 35.215 22.040 35.715 ;
        RECT 22.220 35.665 22.390 35.895 ;
        RECT 22.775 35.835 23.240 36.165 ;
        RECT 23.410 36.455 23.580 37.295 ;
        RECT 23.760 37.265 24.075 37.765 ;
        RECT 24.305 37.035 24.645 37.595 ;
        RECT 23.750 36.660 24.645 37.035 ;
        RECT 24.815 36.755 24.985 37.765 ;
        RECT 24.455 36.455 24.645 36.660 ;
        RECT 25.155 36.705 25.485 37.550 ;
        RECT 25.155 36.625 25.545 36.705 ;
        RECT 25.330 36.575 25.545 36.625 ;
        RECT 25.715 36.600 26.005 37.765 ;
        RECT 26.265 37.095 26.435 37.595 ;
        RECT 26.605 37.265 26.935 37.765 ;
        RECT 26.265 36.925 26.930 37.095 ;
        RECT 23.410 36.125 24.285 36.455 ;
        RECT 24.455 36.125 25.205 36.455 ;
        RECT 23.410 35.665 23.580 36.125 ;
        RECT 24.455 35.955 24.655 36.125 ;
        RECT 25.375 35.995 25.545 36.575 ;
        RECT 26.180 36.105 26.530 36.755 ;
        RECT 25.320 35.955 25.545 35.995 ;
        RECT 22.220 35.495 22.625 35.665 ;
        RECT 22.795 35.495 23.580 35.665 ;
        RECT 23.855 35.215 24.065 35.745 ;
        RECT 24.325 35.430 24.655 35.955 ;
        RECT 25.165 35.870 25.545 35.955 ;
        RECT 24.825 35.215 24.995 35.825 ;
        RECT 25.165 35.435 25.495 35.870 ;
        RECT 25.715 35.215 26.005 35.940 ;
        RECT 26.700 35.935 26.930 36.925 ;
        RECT 26.265 35.765 26.930 35.935 ;
        RECT 26.265 35.475 26.435 35.765 ;
        RECT 26.605 35.215 26.935 35.595 ;
        RECT 27.105 35.475 27.290 37.595 ;
        RECT 27.530 37.305 27.795 37.765 ;
        RECT 27.965 37.170 28.215 37.595 ;
        RECT 28.425 37.320 29.530 37.490 ;
        RECT 27.910 37.040 28.215 37.170 ;
        RECT 27.460 35.845 27.740 36.795 ;
        RECT 27.910 35.935 28.080 37.040 ;
        RECT 28.250 36.255 28.490 36.850 ;
        RECT 28.660 36.785 29.190 37.150 ;
        RECT 28.660 36.085 28.830 36.785 ;
        RECT 29.360 36.705 29.530 37.320 ;
        RECT 29.700 36.965 29.870 37.765 ;
        RECT 30.040 37.265 30.290 37.595 ;
        RECT 30.515 37.295 31.400 37.465 ;
        RECT 29.360 36.615 29.870 36.705 ;
        RECT 27.910 35.805 28.135 35.935 ;
        RECT 28.305 35.865 28.830 36.085 ;
        RECT 29.000 36.445 29.870 36.615 ;
        RECT 27.545 35.215 27.795 35.675 ;
        RECT 27.965 35.665 28.135 35.805 ;
        RECT 29.000 35.665 29.170 36.445 ;
        RECT 29.700 36.375 29.870 36.445 ;
        RECT 29.380 36.195 29.580 36.225 ;
        RECT 30.040 36.195 30.210 37.265 ;
        RECT 30.380 36.375 30.570 37.095 ;
        RECT 29.380 35.895 30.210 36.195 ;
        RECT 30.740 36.165 31.060 37.125 ;
        RECT 27.965 35.495 28.300 35.665 ;
        RECT 28.495 35.495 29.170 35.665 ;
        RECT 29.490 35.215 29.860 35.715 ;
        RECT 30.040 35.665 30.210 35.895 ;
        RECT 30.595 35.835 31.060 36.165 ;
        RECT 31.230 36.455 31.400 37.295 ;
        RECT 31.580 37.265 31.895 37.765 ;
        RECT 32.125 37.035 32.465 37.595 ;
        RECT 31.570 36.660 32.465 37.035 ;
        RECT 32.635 36.755 32.805 37.765 ;
        RECT 32.275 36.455 32.465 36.660 ;
        RECT 32.975 36.705 33.305 37.550 ;
        RECT 33.995 36.810 34.265 37.765 ;
        RECT 34.450 36.710 34.755 37.495 ;
        RECT 34.935 37.295 35.620 37.765 ;
        RECT 34.930 36.775 35.625 37.085 ;
        RECT 32.975 36.625 33.365 36.705 ;
        RECT 33.150 36.575 33.365 36.625 ;
        RECT 31.230 36.125 32.105 36.455 ;
        RECT 32.275 36.125 33.025 36.455 ;
        RECT 31.230 35.665 31.400 36.125 ;
        RECT 32.275 35.955 32.475 36.125 ;
        RECT 33.195 35.995 33.365 36.575 ;
        RECT 33.140 35.955 33.365 35.995 ;
        RECT 30.040 35.495 30.445 35.665 ;
        RECT 30.615 35.495 31.400 35.665 ;
        RECT 31.675 35.215 31.885 35.745 ;
        RECT 32.145 35.430 32.475 35.955 ;
        RECT 32.985 35.870 33.365 35.955 ;
        RECT 34.450 35.905 34.625 36.710 ;
        RECT 35.800 36.605 36.085 37.550 ;
        RECT 36.285 37.315 36.615 37.765 ;
        RECT 36.785 37.145 36.955 37.575 ;
        RECT 35.225 36.455 36.085 36.605 ;
        RECT 34.795 36.435 36.085 36.455 ;
        RECT 36.275 36.915 36.955 37.145 ;
        RECT 38.135 36.965 38.575 37.595 ;
        RECT 34.795 36.075 35.785 36.435 ;
        RECT 36.275 36.265 36.510 36.915 ;
        RECT 32.645 35.215 32.815 35.825 ;
        RECT 32.985 35.435 33.315 35.870 ;
        RECT 33.995 35.215 34.265 35.850 ;
        RECT 34.450 35.385 34.685 35.905 ;
        RECT 35.615 35.740 35.785 36.075 ;
        RECT 35.955 35.935 36.510 36.265 ;
        RECT 36.295 35.785 36.510 35.935 ;
        RECT 36.680 36.065 36.980 36.745 ;
        RECT 36.680 35.895 36.985 36.065 ;
        RECT 38.135 35.955 38.445 36.965 ;
        RECT 38.750 36.915 39.065 37.765 ;
        RECT 39.235 37.425 40.665 37.595 ;
        RECT 39.235 36.745 39.405 37.425 ;
        RECT 38.615 36.575 39.405 36.745 ;
        RECT 38.615 36.125 38.785 36.575 ;
        RECT 39.575 36.455 39.775 37.255 ;
        RECT 38.955 36.125 39.345 36.405 ;
        RECT 39.530 36.125 39.775 36.455 ;
        RECT 39.975 36.125 40.225 37.255 ;
        RECT 40.415 36.795 40.665 37.425 ;
        RECT 40.845 36.965 41.175 37.765 ;
        RECT 41.365 36.795 41.695 37.580 ;
        RECT 40.415 36.625 41.185 36.795 ;
        RECT 41.365 36.625 42.045 36.795 ;
        RECT 42.225 36.625 42.555 37.765 ;
        RECT 40.440 36.125 40.845 36.455 ;
        RECT 41.015 35.955 41.185 36.625 ;
        RECT 41.355 36.205 41.705 36.455 ;
        RECT 41.875 36.025 42.045 36.625 ;
        RECT 43.195 36.610 43.535 37.595 ;
        RECT 43.705 37.335 44.115 37.765 ;
        RECT 44.860 37.345 45.190 37.765 ;
        RECT 45.360 37.165 45.685 37.595 ;
        RECT 43.705 36.995 45.685 37.165 ;
        RECT 42.215 36.205 42.565 36.455 ;
        RECT 34.855 35.215 35.255 35.710 ;
        RECT 35.615 35.545 36.015 35.740 ;
        RECT 35.845 35.400 36.015 35.545 ;
        RECT 36.295 35.410 36.535 35.785 ;
        RECT 36.705 35.215 37.035 35.720 ;
        RECT 38.135 35.395 38.575 35.955 ;
        RECT 38.745 35.215 39.195 35.955 ;
        RECT 39.365 35.785 40.525 35.955 ;
        RECT 39.365 35.385 39.535 35.785 ;
        RECT 39.705 35.215 40.125 35.615 ;
        RECT 40.295 35.385 40.525 35.785 ;
        RECT 40.695 35.385 41.185 35.955 ;
        RECT 41.375 35.215 41.615 36.025 ;
        RECT 41.785 35.385 42.115 36.025 ;
        RECT 42.285 35.215 42.555 36.025 ;
        RECT 43.195 35.955 43.450 36.610 ;
        RECT 43.705 36.455 43.970 36.995 ;
        RECT 44.185 36.655 44.810 36.825 ;
        RECT 43.620 36.125 43.970 36.455 ;
        RECT 44.140 36.125 44.470 36.455 ;
        RECT 44.640 35.955 44.810 36.655 ;
        RECT 43.195 35.580 43.555 35.955 ;
        RECT 43.820 35.215 43.990 35.955 ;
        RECT 44.270 35.785 44.810 35.955 ;
        RECT 44.980 36.585 45.685 36.995 ;
        RECT 46.160 36.665 46.490 37.765 ;
        RECT 47.335 36.675 48.545 37.765 ;
        RECT 44.270 35.580 44.440 35.785 ;
        RECT 44.980 35.385 45.150 36.585 ;
        RECT 45.320 36.205 45.890 36.415 ;
        RECT 46.060 36.205 46.705 36.415 ;
        RECT 47.335 36.135 47.855 36.675 ;
        RECT 45.380 35.865 46.550 36.035 ;
        RECT 48.025 35.965 48.545 36.505 ;
        RECT 45.380 35.385 45.710 35.865 ;
        RECT 45.880 35.215 46.050 35.685 ;
        RECT 46.220 35.400 46.550 35.865 ;
        RECT 47.335 35.215 48.545 35.965 ;
        RECT 12.750 35.045 48.630 35.215 ;
        RECT 12.835 34.295 14.045 35.045 ;
        RECT 14.265 34.390 14.595 34.825 ;
        RECT 14.765 34.435 14.935 35.045 ;
        RECT 14.215 34.305 14.595 34.390 ;
        RECT 15.105 34.305 15.435 34.830 ;
        RECT 15.695 34.515 15.905 35.045 ;
        RECT 16.180 34.595 16.965 34.765 ;
        RECT 17.135 34.595 17.540 34.765 ;
        RECT 12.835 33.755 13.355 34.295 ;
        RECT 14.215 34.265 14.440 34.305 ;
        RECT 13.525 33.585 14.045 34.125 ;
        RECT 12.835 32.495 14.045 33.585 ;
        RECT 14.215 33.685 14.385 34.265 ;
        RECT 15.105 34.135 15.305 34.305 ;
        RECT 16.180 34.135 16.350 34.595 ;
        RECT 14.555 33.805 15.305 34.135 ;
        RECT 15.475 33.805 16.350 34.135 ;
        RECT 14.215 33.635 14.430 33.685 ;
        RECT 14.215 33.555 14.605 33.635 ;
        RECT 14.275 32.710 14.605 33.555 ;
        RECT 15.115 33.600 15.305 33.805 ;
        RECT 14.775 32.495 14.945 33.505 ;
        RECT 15.115 33.225 16.010 33.600 ;
        RECT 15.115 32.665 15.455 33.225 ;
        RECT 15.685 32.495 16.000 32.995 ;
        RECT 16.180 32.965 16.350 33.805 ;
        RECT 16.520 34.095 16.985 34.425 ;
        RECT 17.370 34.365 17.540 34.595 ;
        RECT 17.720 34.545 18.090 35.045 ;
        RECT 18.410 34.595 19.085 34.765 ;
        RECT 19.280 34.595 19.615 34.765 ;
        RECT 16.520 33.135 16.840 34.095 ;
        RECT 17.370 34.065 18.200 34.365 ;
        RECT 17.010 33.165 17.200 33.885 ;
        RECT 17.370 32.995 17.540 34.065 ;
        RECT 18.000 34.035 18.200 34.065 ;
        RECT 17.710 33.815 17.880 33.885 ;
        RECT 18.410 33.815 18.580 34.595 ;
        RECT 19.445 34.455 19.615 34.595 ;
        RECT 19.785 34.585 20.035 35.045 ;
        RECT 17.710 33.645 18.580 33.815 ;
        RECT 18.750 34.175 19.275 34.395 ;
        RECT 19.445 34.325 19.670 34.455 ;
        RECT 17.710 33.555 18.220 33.645 ;
        RECT 16.180 32.795 17.065 32.965 ;
        RECT 17.290 32.665 17.540 32.995 ;
        RECT 17.710 32.495 17.880 33.295 ;
        RECT 18.050 32.940 18.220 33.555 ;
        RECT 18.750 33.475 18.920 34.175 ;
        RECT 18.390 33.110 18.920 33.475 ;
        RECT 19.090 33.410 19.330 34.005 ;
        RECT 19.500 33.220 19.670 34.325 ;
        RECT 19.840 33.465 20.120 34.415 ;
        RECT 19.365 33.090 19.670 33.220 ;
        RECT 18.050 32.770 19.155 32.940 ;
        RECT 19.365 32.665 19.615 33.090 ;
        RECT 19.785 32.495 20.050 32.955 ;
        RECT 20.290 32.665 20.475 34.785 ;
        RECT 20.645 34.665 20.975 35.045 ;
        RECT 21.145 34.495 21.315 34.785 ;
        RECT 20.650 34.325 21.315 34.495 ;
        RECT 20.650 33.335 20.880 34.325 ;
        RECT 21.575 34.275 24.165 35.045 ;
        RECT 24.795 34.535 25.100 35.045 ;
        RECT 21.050 33.505 21.400 34.155 ;
        RECT 21.575 33.755 22.785 34.275 ;
        RECT 22.955 33.585 24.165 34.105 ;
        RECT 24.795 33.805 25.110 34.365 ;
        RECT 25.280 34.055 25.530 34.865 ;
        RECT 25.700 34.520 25.960 35.045 ;
        RECT 26.140 34.055 26.390 34.865 ;
        RECT 26.560 34.485 26.820 35.045 ;
        RECT 26.990 34.395 27.250 34.850 ;
        RECT 27.420 34.565 27.680 35.045 ;
        RECT 27.850 34.395 28.110 34.850 ;
        RECT 28.280 34.565 28.540 35.045 ;
        RECT 28.710 34.395 28.970 34.850 ;
        RECT 29.140 34.565 29.385 35.045 ;
        RECT 29.555 34.395 29.830 34.850 ;
        RECT 30.000 34.565 30.245 35.045 ;
        RECT 30.415 34.395 30.675 34.850 ;
        RECT 30.855 34.565 31.105 35.045 ;
        RECT 31.275 34.395 31.535 34.850 ;
        RECT 31.715 34.565 31.965 35.045 ;
        RECT 32.135 34.395 32.395 34.850 ;
        RECT 32.575 34.565 32.835 35.045 ;
        RECT 33.005 34.395 33.265 34.850 ;
        RECT 33.435 34.565 33.735 35.045 ;
        RECT 26.990 34.225 33.735 34.395 ;
        RECT 25.280 33.805 32.400 34.055 ;
        RECT 20.650 33.165 21.315 33.335 ;
        RECT 20.645 32.495 20.975 32.995 ;
        RECT 21.145 32.665 21.315 33.165 ;
        RECT 21.575 32.495 24.165 33.585 ;
        RECT 24.805 32.495 25.100 33.305 ;
        RECT 25.280 32.665 25.525 33.805 ;
        RECT 25.700 32.495 25.960 33.305 ;
        RECT 26.140 32.670 26.390 33.805 ;
        RECT 32.570 33.635 33.735 34.225 ;
        RECT 26.990 33.410 33.735 33.635 ;
        RECT 33.995 34.305 34.380 34.875 ;
        RECT 34.550 34.585 34.875 35.045 ;
        RECT 35.395 34.415 35.675 34.875 ;
        RECT 33.995 33.635 34.275 34.305 ;
        RECT 34.550 34.245 35.675 34.415 ;
        RECT 34.550 34.135 35.000 34.245 ;
        RECT 34.445 33.805 35.000 34.135 ;
        RECT 35.865 34.075 36.265 34.875 ;
        RECT 36.665 34.585 36.935 35.045 ;
        RECT 37.105 34.415 37.390 34.875 ;
        RECT 26.990 33.395 32.395 33.410 ;
        RECT 26.560 32.500 26.820 33.295 ;
        RECT 26.990 32.670 27.250 33.395 ;
        RECT 27.420 32.500 27.680 33.225 ;
        RECT 27.850 32.670 28.110 33.395 ;
        RECT 28.280 32.500 28.540 33.225 ;
        RECT 28.710 32.670 28.970 33.395 ;
        RECT 29.140 32.500 29.400 33.225 ;
        RECT 29.570 32.670 29.830 33.395 ;
        RECT 30.000 32.500 30.245 33.225 ;
        RECT 30.415 32.670 30.675 33.395 ;
        RECT 30.860 32.500 31.105 33.225 ;
        RECT 31.275 32.670 31.535 33.395 ;
        RECT 31.720 32.500 31.965 33.225 ;
        RECT 32.135 32.670 32.395 33.395 ;
        RECT 32.580 32.500 32.835 33.225 ;
        RECT 33.005 32.670 33.295 33.410 ;
        RECT 26.560 32.495 32.835 32.500 ;
        RECT 33.465 32.495 33.735 33.240 ;
        RECT 33.995 32.665 34.380 33.635 ;
        RECT 34.550 33.345 35.000 33.805 ;
        RECT 35.170 33.515 36.265 34.075 ;
        RECT 34.550 33.125 35.675 33.345 ;
        RECT 34.550 32.495 34.875 32.955 ;
        RECT 35.395 32.665 35.675 33.125 ;
        RECT 35.865 32.665 36.265 33.515 ;
        RECT 36.435 34.245 37.390 34.415 ;
        RECT 38.595 34.320 38.885 35.045 ;
        RECT 39.070 34.475 39.325 34.825 ;
        RECT 39.495 34.645 39.825 35.045 ;
        RECT 39.995 34.475 40.165 34.825 ;
        RECT 40.335 34.645 40.715 35.045 ;
        RECT 39.070 34.305 40.735 34.475 ;
        RECT 40.905 34.370 41.180 34.715 ;
        RECT 36.435 33.345 36.645 34.245 ;
        RECT 40.565 34.135 40.735 34.305 ;
        RECT 36.815 33.515 37.505 34.075 ;
        RECT 39.055 33.805 39.400 34.135 ;
        RECT 39.570 33.805 40.395 34.135 ;
        RECT 40.565 33.805 40.840 34.135 ;
        RECT 36.435 33.125 37.390 33.345 ;
        RECT 36.665 32.495 36.935 32.955 ;
        RECT 37.105 32.665 37.390 33.125 ;
        RECT 38.595 32.495 38.885 33.660 ;
        RECT 39.075 33.345 39.400 33.635 ;
        RECT 39.570 33.515 39.765 33.805 ;
        RECT 40.565 33.635 40.735 33.805 ;
        RECT 41.010 33.635 41.180 34.370 ;
        RECT 41.355 34.275 43.945 35.045 ;
        RECT 41.355 33.755 42.565 34.275 ;
        RECT 44.585 34.235 44.855 35.045 ;
        RECT 45.025 34.235 45.355 34.875 ;
        RECT 45.525 34.235 45.765 35.045 ;
        RECT 45.955 34.370 46.215 34.875 ;
        RECT 46.395 34.665 46.725 35.045 ;
        RECT 46.905 34.495 47.075 34.875 ;
        RECT 40.075 33.465 40.735 33.635 ;
        RECT 40.075 33.345 40.245 33.465 ;
        RECT 39.075 33.175 40.245 33.345 ;
        RECT 39.055 32.715 40.245 33.005 ;
        RECT 40.415 32.495 40.695 33.295 ;
        RECT 40.905 32.665 41.180 33.635 ;
        RECT 42.735 33.585 43.945 34.105 ;
        RECT 44.575 33.805 44.925 34.055 ;
        RECT 45.095 33.635 45.265 34.235 ;
        RECT 45.435 33.805 45.785 34.055 ;
        RECT 41.355 32.495 43.945 33.585 ;
        RECT 44.585 32.495 44.915 33.635 ;
        RECT 45.095 33.465 45.775 33.635 ;
        RECT 45.445 32.680 45.775 33.465 ;
        RECT 45.955 33.570 46.125 34.370 ;
        RECT 46.410 34.325 47.075 34.495 ;
        RECT 46.410 34.070 46.580 34.325 ;
        RECT 47.335 34.295 48.545 35.045 ;
        RECT 46.295 33.740 46.580 34.070 ;
        RECT 46.815 33.775 47.145 34.145 ;
        RECT 46.410 33.595 46.580 33.740 ;
        RECT 45.955 32.665 46.225 33.570 ;
        RECT 46.410 33.425 47.075 33.595 ;
        RECT 46.395 32.495 46.725 33.255 ;
        RECT 46.905 32.665 47.075 33.425 ;
        RECT 47.335 33.585 47.855 34.125 ;
        RECT 48.025 33.755 48.545 34.295 ;
        RECT 47.335 32.495 48.545 33.585 ;
        RECT 12.750 32.325 48.630 32.495 ;
        RECT 12.835 31.235 14.045 32.325 ;
        RECT 14.215 31.235 15.425 32.325 ;
        RECT 15.710 31.695 15.995 32.155 ;
        RECT 16.165 31.865 16.435 32.325 ;
        RECT 15.710 31.475 16.665 31.695 ;
        RECT 12.835 30.525 13.355 31.065 ;
        RECT 13.525 30.695 14.045 31.235 ;
        RECT 14.215 30.525 14.735 31.065 ;
        RECT 14.905 30.695 15.425 31.235 ;
        RECT 15.595 30.745 16.285 31.305 ;
        RECT 16.455 30.575 16.665 31.475 ;
        RECT 12.835 29.775 14.045 30.525 ;
        RECT 14.215 29.775 15.425 30.525 ;
        RECT 15.710 30.405 16.665 30.575 ;
        RECT 16.835 31.305 17.235 32.155 ;
        RECT 17.425 31.695 17.705 32.155 ;
        RECT 18.225 31.865 18.550 32.325 ;
        RECT 17.425 31.475 18.550 31.695 ;
        RECT 16.835 30.745 17.930 31.305 ;
        RECT 18.100 31.015 18.550 31.475 ;
        RECT 18.720 31.185 19.105 32.155 ;
        RECT 15.710 29.945 15.995 30.405 ;
        RECT 16.165 29.775 16.435 30.235 ;
        RECT 16.835 29.945 17.235 30.745 ;
        RECT 18.100 30.685 18.655 31.015 ;
        RECT 18.100 30.575 18.550 30.685 ;
        RECT 17.425 30.405 18.550 30.575 ;
        RECT 18.825 30.515 19.105 31.185 ;
        RECT 17.425 29.945 17.705 30.405 ;
        RECT 18.225 29.775 18.550 30.235 ;
        RECT 18.720 29.945 19.105 30.515 ;
        RECT 19.275 31.185 19.660 32.155 ;
        RECT 19.830 31.865 20.155 32.325 ;
        RECT 20.675 31.695 20.955 32.155 ;
        RECT 19.830 31.475 20.955 31.695 ;
        RECT 19.275 30.515 19.555 31.185 ;
        RECT 19.830 31.015 20.280 31.475 ;
        RECT 21.145 31.305 21.545 32.155 ;
        RECT 21.945 31.865 22.215 32.325 ;
        RECT 22.385 31.695 22.670 32.155 ;
        RECT 19.725 30.685 20.280 31.015 ;
        RECT 20.450 30.745 21.545 31.305 ;
        RECT 19.830 30.575 20.280 30.685 ;
        RECT 19.275 29.945 19.660 30.515 ;
        RECT 19.830 30.405 20.955 30.575 ;
        RECT 19.830 29.775 20.155 30.235 ;
        RECT 20.675 29.945 20.955 30.405 ;
        RECT 21.145 29.945 21.545 30.745 ;
        RECT 21.715 31.475 22.670 31.695 ;
        RECT 21.715 30.575 21.925 31.475 ;
        RECT 22.095 30.745 22.785 31.305 ;
        RECT 22.955 31.235 25.545 32.325 ;
        RECT 21.715 30.405 22.670 30.575 ;
        RECT 21.945 29.775 22.215 30.235 ;
        RECT 22.385 29.945 22.670 30.405 ;
        RECT 22.955 30.545 24.165 31.065 ;
        RECT 24.335 30.715 25.545 31.235 ;
        RECT 25.715 31.160 26.005 32.325 ;
        RECT 26.185 31.185 26.515 32.325 ;
        RECT 27.045 31.355 27.375 32.140 ;
        RECT 26.695 31.185 27.375 31.355 ;
        RECT 27.675 31.205 28.005 32.325 ;
        RECT 26.175 30.765 26.525 31.015 ;
        RECT 26.695 30.585 26.865 31.185 ;
        RECT 27.035 30.765 27.385 31.015 ;
        RECT 27.615 30.765 28.125 31.015 ;
        RECT 28.335 30.765 28.705 32.080 ;
        RECT 28.875 30.765 29.205 32.080 ;
        RECT 29.415 30.765 29.745 32.080 ;
        RECT 30.015 31.435 30.265 32.155 ;
        RECT 30.435 31.605 30.765 32.325 ;
        RECT 30.015 31.145 30.765 31.435 ;
        RECT 31.000 31.145 31.525 32.155 ;
        RECT 30.505 30.975 30.765 31.145 ;
        RECT 29.915 30.765 30.335 30.975 ;
        RECT 30.505 30.765 31.085 30.975 ;
        RECT 30.505 30.595 30.875 30.765 ;
        RECT 22.955 29.775 25.545 30.545 ;
        RECT 25.715 29.775 26.005 30.500 ;
        RECT 26.185 29.775 26.455 30.585 ;
        RECT 26.625 29.945 26.955 30.585 ;
        RECT 27.125 29.775 27.365 30.585 ;
        RECT 27.655 30.425 29.955 30.595 ;
        RECT 27.655 29.945 27.985 30.425 ;
        RECT 28.155 29.775 28.485 30.235 ;
        RECT 28.700 29.945 29.030 30.425 ;
        RECT 29.230 29.775 29.560 30.235 ;
        RECT 29.785 30.105 29.955 30.425 ;
        RECT 30.125 30.405 30.875 30.595 ;
        RECT 31.255 30.575 31.525 31.145 ;
        RECT 30.125 29.960 30.455 30.405 ;
        RECT 30.725 29.775 30.895 30.235 ;
        RECT 31.185 29.945 31.525 30.575 ;
        RECT 31.695 31.185 32.080 32.155 ;
        RECT 32.250 31.865 32.575 32.325 ;
        RECT 33.095 31.695 33.375 32.155 ;
        RECT 32.250 31.475 33.375 31.695 ;
        RECT 31.695 30.515 31.975 31.185 ;
        RECT 32.250 31.015 32.700 31.475 ;
        RECT 33.565 31.305 33.965 32.155 ;
        RECT 34.365 31.865 34.635 32.325 ;
        RECT 34.805 31.695 35.090 32.155 ;
        RECT 32.145 30.685 32.700 31.015 ;
        RECT 32.870 30.745 33.965 31.305 ;
        RECT 32.250 30.575 32.700 30.685 ;
        RECT 31.695 29.945 32.080 30.515 ;
        RECT 32.250 30.405 33.375 30.575 ;
        RECT 32.250 29.775 32.575 30.235 ;
        RECT 33.095 29.945 33.375 30.405 ;
        RECT 33.565 29.945 33.965 30.745 ;
        RECT 34.135 31.475 35.090 31.695 ;
        RECT 34.135 30.575 34.345 31.475 ;
        RECT 34.515 30.745 35.205 31.305 ;
        RECT 35.375 31.235 36.585 32.325 ;
        RECT 34.135 30.405 35.090 30.575 ;
        RECT 34.365 29.775 34.635 30.235 ;
        RECT 34.805 29.945 35.090 30.405 ;
        RECT 35.375 30.525 35.895 31.065 ;
        RECT 36.065 30.695 36.585 31.235 ;
        RECT 36.755 31.185 37.030 32.155 ;
        RECT 37.240 31.525 37.520 32.325 ;
        RECT 37.690 31.815 39.740 32.105 ;
        RECT 37.690 31.475 39.320 31.645 ;
        RECT 37.690 31.355 37.860 31.475 ;
        RECT 37.200 31.185 37.860 31.355 ;
        RECT 35.375 29.775 36.585 30.525 ;
        RECT 36.755 30.450 36.925 31.185 ;
        RECT 37.200 31.015 37.370 31.185 ;
        RECT 37.095 30.685 37.370 31.015 ;
        RECT 37.540 30.685 37.920 31.015 ;
        RECT 38.090 30.685 38.830 31.305 ;
        RECT 39.000 31.185 39.320 31.475 ;
        RECT 39.515 31.015 39.755 31.610 ;
        RECT 39.925 31.250 40.265 32.325 ;
        RECT 40.445 31.355 40.775 32.140 ;
        RECT 40.445 31.185 41.125 31.355 ;
        RECT 41.305 31.185 41.635 32.325 ;
        RECT 41.895 31.395 42.075 32.155 ;
        RECT 42.255 31.565 42.585 32.325 ;
        RECT 41.895 31.225 42.570 31.395 ;
        RECT 42.755 31.250 43.025 32.155 ;
        RECT 39.100 30.685 39.755 31.015 ;
        RECT 37.200 30.515 37.370 30.685 ;
        RECT 36.755 30.105 37.030 30.450 ;
        RECT 37.200 30.345 38.785 30.515 ;
        RECT 37.220 29.775 37.600 30.175 ;
        RECT 37.770 29.995 37.940 30.345 ;
        RECT 38.110 29.775 38.440 30.175 ;
        RECT 38.615 29.995 38.785 30.345 ;
        RECT 38.985 29.775 39.315 30.275 ;
        RECT 39.510 29.995 39.755 30.685 ;
        RECT 39.925 30.445 40.265 31.015 ;
        RECT 40.435 30.765 40.785 31.015 ;
        RECT 40.955 30.585 41.125 31.185 ;
        RECT 42.400 31.080 42.570 31.225 ;
        RECT 41.295 30.765 41.645 31.015 ;
        RECT 41.835 30.675 42.175 31.045 ;
        RECT 42.400 30.750 42.675 31.080 ;
        RECT 39.925 29.775 40.265 30.275 ;
        RECT 40.455 29.775 40.695 30.585 ;
        RECT 40.865 29.945 41.195 30.585 ;
        RECT 41.365 29.775 41.635 30.585 ;
        RECT 42.400 30.495 42.570 30.750 ;
        RECT 41.905 30.325 42.570 30.495 ;
        RECT 42.845 30.450 43.025 31.250 ;
        RECT 43.410 31.225 43.740 32.325 ;
        RECT 44.215 31.725 44.540 32.155 ;
        RECT 44.710 31.905 45.040 32.325 ;
        RECT 45.785 31.895 46.195 32.325 ;
        RECT 44.215 31.555 46.195 31.725 ;
        RECT 44.215 31.145 44.920 31.555 ;
        RECT 43.195 30.765 43.840 30.975 ;
        RECT 44.010 30.765 44.580 30.975 ;
        RECT 41.905 29.945 42.075 30.325 ;
        RECT 42.255 29.775 42.585 30.155 ;
        RECT 42.765 29.945 43.025 30.450 ;
        RECT 43.350 30.425 44.520 30.595 ;
        RECT 43.350 29.960 43.680 30.425 ;
        RECT 43.850 29.775 44.020 30.245 ;
        RECT 44.190 29.945 44.520 30.425 ;
        RECT 44.750 29.945 44.920 31.145 ;
        RECT 45.090 31.215 45.715 31.385 ;
        RECT 45.090 30.515 45.260 31.215 ;
        RECT 45.930 31.015 46.195 31.555 ;
        RECT 46.365 31.170 46.705 32.155 ;
        RECT 45.430 30.685 45.760 31.015 ;
        RECT 45.930 30.685 46.280 31.015 ;
        RECT 46.450 30.515 46.705 31.170 ;
        RECT 47.335 31.235 48.545 32.325 ;
        RECT 47.335 30.695 47.855 31.235 ;
        RECT 48.025 30.525 48.545 31.065 ;
        RECT 45.090 30.345 45.630 30.515 ;
        RECT 45.460 30.140 45.630 30.345 ;
        RECT 45.910 29.775 46.080 30.515 ;
        RECT 46.345 30.140 46.705 30.515 ;
        RECT 47.335 29.775 48.545 30.525 ;
        RECT 12.750 29.605 48.630 29.775 ;
        RECT 12.835 28.855 14.045 29.605 ;
        RECT 12.835 28.315 13.355 28.855 ;
        RECT 14.220 28.765 14.480 29.605 ;
        RECT 14.655 28.860 14.910 29.435 ;
        RECT 15.080 29.225 15.410 29.605 ;
        RECT 15.625 29.055 15.795 29.435 ;
        RECT 15.080 28.885 15.795 29.055 ;
        RECT 13.525 28.145 14.045 28.685 ;
        RECT 12.835 27.055 14.045 28.145 ;
        RECT 14.220 27.055 14.480 28.205 ;
        RECT 14.655 28.130 14.825 28.860 ;
        RECT 15.080 28.695 15.250 28.885 ;
        RECT 16.520 28.865 16.775 29.435 ;
        RECT 16.945 29.205 17.275 29.605 ;
        RECT 17.700 29.070 18.230 29.435 ;
        RECT 18.420 29.265 18.695 29.435 ;
        RECT 18.415 29.095 18.695 29.265 ;
        RECT 17.700 29.035 17.875 29.070 ;
        RECT 16.945 28.865 17.875 29.035 ;
        RECT 14.995 28.365 15.250 28.695 ;
        RECT 15.080 28.155 15.250 28.365 ;
        RECT 15.530 28.335 15.885 28.705 ;
        RECT 16.520 28.195 16.690 28.865 ;
        RECT 16.945 28.695 17.115 28.865 ;
        RECT 16.860 28.365 17.115 28.695 ;
        RECT 17.340 28.365 17.535 28.695 ;
        RECT 14.655 27.225 14.910 28.130 ;
        RECT 15.080 27.985 15.795 28.155 ;
        RECT 15.080 27.055 15.410 27.815 ;
        RECT 15.625 27.225 15.795 27.985 ;
        RECT 16.520 27.225 16.855 28.195 ;
        RECT 17.025 27.055 17.195 28.195 ;
        RECT 17.365 27.395 17.535 28.365 ;
        RECT 17.705 27.735 17.875 28.865 ;
        RECT 18.045 28.075 18.215 28.875 ;
        RECT 18.420 28.275 18.695 29.095 ;
        RECT 18.865 28.075 19.055 29.435 ;
        RECT 19.235 29.070 19.745 29.605 ;
        RECT 19.965 28.795 20.210 29.400 ;
        RECT 20.745 29.055 20.915 29.345 ;
        RECT 21.085 29.225 21.415 29.605 ;
        RECT 20.745 28.885 21.410 29.055 ;
        RECT 19.255 28.625 20.485 28.795 ;
        RECT 18.045 27.905 19.055 28.075 ;
        RECT 19.225 28.060 19.975 28.250 ;
        RECT 17.705 27.565 18.830 27.735 ;
        RECT 19.225 27.395 19.395 28.060 ;
        RECT 20.145 27.815 20.485 28.625 ;
        RECT 20.660 28.065 21.010 28.715 ;
        RECT 21.180 27.895 21.410 28.885 ;
        RECT 17.365 27.225 19.395 27.395 ;
        RECT 19.565 27.055 19.735 27.815 ;
        RECT 19.970 27.405 20.485 27.815 ;
        RECT 20.745 27.725 21.410 27.895 ;
        RECT 20.745 27.225 20.915 27.725 ;
        RECT 21.085 27.055 21.415 27.555 ;
        RECT 21.585 27.225 21.770 29.345 ;
        RECT 22.025 29.145 22.275 29.605 ;
        RECT 22.445 29.155 22.780 29.325 ;
        RECT 22.975 29.155 23.650 29.325 ;
        RECT 22.445 29.015 22.615 29.155 ;
        RECT 21.940 28.025 22.220 28.975 ;
        RECT 22.390 28.885 22.615 29.015 ;
        RECT 22.390 27.780 22.560 28.885 ;
        RECT 22.785 28.735 23.310 28.955 ;
        RECT 22.730 27.970 22.970 28.565 ;
        RECT 23.140 28.035 23.310 28.735 ;
        RECT 23.480 28.375 23.650 29.155 ;
        RECT 23.970 29.105 24.340 29.605 ;
        RECT 24.520 29.155 24.925 29.325 ;
        RECT 25.095 29.155 25.880 29.325 ;
        RECT 24.520 28.925 24.690 29.155 ;
        RECT 23.860 28.625 24.690 28.925 ;
        RECT 25.075 28.655 25.540 28.985 ;
        RECT 23.860 28.595 24.060 28.625 ;
        RECT 24.180 28.375 24.350 28.445 ;
        RECT 23.480 28.205 24.350 28.375 ;
        RECT 23.840 28.115 24.350 28.205 ;
        RECT 22.390 27.650 22.695 27.780 ;
        RECT 23.140 27.670 23.670 28.035 ;
        RECT 22.010 27.055 22.275 27.515 ;
        RECT 22.445 27.225 22.695 27.650 ;
        RECT 23.840 27.500 24.010 28.115 ;
        RECT 22.905 27.330 24.010 27.500 ;
        RECT 24.180 27.055 24.350 27.855 ;
        RECT 24.520 27.555 24.690 28.625 ;
        RECT 24.860 27.725 25.050 28.445 ;
        RECT 25.220 27.695 25.540 28.655 ;
        RECT 25.710 28.695 25.880 29.155 ;
        RECT 26.155 29.075 26.365 29.605 ;
        RECT 26.625 28.865 26.955 29.390 ;
        RECT 27.125 28.995 27.295 29.605 ;
        RECT 27.465 28.950 27.795 29.385 ;
        RECT 27.465 28.865 27.845 28.950 ;
        RECT 26.755 28.695 26.955 28.865 ;
        RECT 27.620 28.825 27.845 28.865 ;
        RECT 25.710 28.365 26.585 28.695 ;
        RECT 26.755 28.365 27.505 28.695 ;
        RECT 24.520 27.225 24.770 27.555 ;
        RECT 25.710 27.525 25.880 28.365 ;
        RECT 26.755 28.160 26.945 28.365 ;
        RECT 27.675 28.245 27.845 28.825 ;
        RECT 27.630 28.195 27.845 28.245 ;
        RECT 26.050 27.785 26.945 28.160 ;
        RECT 27.455 28.115 27.845 28.195 ;
        RECT 28.020 28.865 28.275 29.435 ;
        RECT 28.445 29.205 28.775 29.605 ;
        RECT 29.200 29.070 29.730 29.435 ;
        RECT 29.200 29.035 29.375 29.070 ;
        RECT 28.445 28.865 29.375 29.035 ;
        RECT 28.020 28.195 28.190 28.865 ;
        RECT 28.445 28.695 28.615 28.865 ;
        RECT 28.360 28.365 28.615 28.695 ;
        RECT 28.840 28.365 29.035 28.695 ;
        RECT 24.995 27.355 25.880 27.525 ;
        RECT 26.060 27.055 26.375 27.555 ;
        RECT 26.605 27.225 26.945 27.785 ;
        RECT 27.115 27.055 27.285 28.065 ;
        RECT 27.455 27.270 27.785 28.115 ;
        RECT 28.020 27.225 28.355 28.195 ;
        RECT 28.525 27.055 28.695 28.195 ;
        RECT 28.865 27.395 29.035 28.365 ;
        RECT 29.205 27.735 29.375 28.865 ;
        RECT 29.545 28.075 29.715 28.875 ;
        RECT 29.920 28.585 30.195 29.435 ;
        RECT 29.915 28.415 30.195 28.585 ;
        RECT 29.920 28.275 30.195 28.415 ;
        RECT 30.365 28.075 30.555 29.435 ;
        RECT 30.735 29.070 31.245 29.605 ;
        RECT 31.465 28.795 31.710 29.400 ;
        RECT 32.155 28.865 32.540 29.435 ;
        RECT 32.710 29.145 33.035 29.605 ;
        RECT 33.555 28.975 33.835 29.435 ;
        RECT 30.755 28.625 31.985 28.795 ;
        RECT 29.545 27.905 30.555 28.075 ;
        RECT 30.725 28.060 31.475 28.250 ;
        RECT 29.205 27.565 30.330 27.735 ;
        RECT 30.725 27.395 30.895 28.060 ;
        RECT 31.645 27.815 31.985 28.625 ;
        RECT 28.865 27.225 30.895 27.395 ;
        RECT 31.065 27.055 31.235 27.815 ;
        RECT 31.470 27.405 31.985 27.815 ;
        RECT 32.155 28.195 32.435 28.865 ;
        RECT 32.710 28.805 33.835 28.975 ;
        RECT 32.710 28.695 33.160 28.805 ;
        RECT 32.605 28.365 33.160 28.695 ;
        RECT 34.025 28.635 34.425 29.435 ;
        RECT 34.825 29.145 35.095 29.605 ;
        RECT 35.265 28.975 35.550 29.435 ;
        RECT 32.155 27.225 32.540 28.195 ;
        RECT 32.710 27.905 33.160 28.365 ;
        RECT 33.330 28.075 34.425 28.635 ;
        RECT 32.710 27.685 33.835 27.905 ;
        RECT 32.710 27.055 33.035 27.515 ;
        RECT 33.555 27.225 33.835 27.685 ;
        RECT 34.025 27.225 34.425 28.075 ;
        RECT 34.595 28.805 35.550 28.975 ;
        RECT 35.835 28.835 38.425 29.605 ;
        RECT 38.595 28.880 38.885 29.605 ;
        RECT 39.385 29.205 39.715 29.605 ;
        RECT 39.885 29.035 40.215 29.375 ;
        RECT 41.265 29.205 41.595 29.605 ;
        RECT 39.230 28.865 41.595 29.035 ;
        RECT 41.765 28.880 42.095 29.390 ;
        RECT 34.595 27.905 34.805 28.805 ;
        RECT 34.975 28.075 35.665 28.635 ;
        RECT 35.835 28.315 37.045 28.835 ;
        RECT 37.215 28.145 38.425 28.665 ;
        RECT 34.595 27.685 35.550 27.905 ;
        RECT 34.825 27.055 35.095 27.515 ;
        RECT 35.265 27.225 35.550 27.685 ;
        RECT 35.835 27.055 38.425 28.145 ;
        RECT 38.595 27.055 38.885 28.220 ;
        RECT 39.230 27.865 39.400 28.865 ;
        RECT 41.425 28.695 41.595 28.865 ;
        RECT 39.570 28.035 39.815 28.695 ;
        RECT 40.030 28.035 40.295 28.695 ;
        RECT 40.490 28.035 40.775 28.695 ;
        RECT 40.950 28.365 41.255 28.695 ;
        RECT 41.425 28.365 41.735 28.695 ;
        RECT 40.950 28.035 41.165 28.365 ;
        RECT 39.230 27.695 39.685 27.865 ;
        RECT 39.355 27.265 39.685 27.695 ;
        RECT 39.865 27.695 41.155 27.865 ;
        RECT 39.865 27.275 40.115 27.695 ;
        RECT 40.345 27.055 40.675 27.525 ;
        RECT 40.905 27.275 41.155 27.695 ;
        RECT 41.345 27.055 41.595 28.195 ;
        RECT 41.905 28.115 42.095 28.880 ;
        RECT 43.350 28.955 43.680 29.420 ;
        RECT 43.850 29.135 44.020 29.605 ;
        RECT 44.190 28.955 44.520 29.435 ;
        RECT 43.350 28.785 44.520 28.955 ;
        RECT 43.195 28.405 43.840 28.615 ;
        RECT 44.010 28.405 44.580 28.615 ;
        RECT 44.750 28.235 44.920 29.435 ;
        RECT 45.460 29.035 45.630 29.240 ;
        RECT 41.765 27.265 42.095 28.115 ;
        RECT 43.410 27.055 43.740 28.155 ;
        RECT 44.215 27.825 44.920 28.235 ;
        RECT 45.090 28.865 45.630 29.035 ;
        RECT 45.910 28.865 46.080 29.605 ;
        RECT 46.475 29.240 46.645 29.265 ;
        RECT 46.345 28.865 46.705 29.240 ;
        RECT 45.090 28.165 45.260 28.865 ;
        RECT 45.430 28.365 45.760 28.695 ;
        RECT 45.930 28.365 46.280 28.695 ;
        RECT 45.090 27.995 45.715 28.165 ;
        RECT 45.930 27.825 46.195 28.365 ;
        RECT 46.450 28.210 46.705 28.865 ;
        RECT 47.335 28.855 48.545 29.605 ;
        RECT 44.215 27.655 46.195 27.825 ;
        RECT 44.215 27.225 44.540 27.655 ;
        RECT 44.710 27.055 45.040 27.475 ;
        RECT 45.785 27.055 46.195 27.485 ;
        RECT 46.365 27.225 46.705 28.210 ;
        RECT 47.335 28.145 47.855 28.685 ;
        RECT 48.025 28.315 48.545 28.855 ;
        RECT 47.335 27.055 48.545 28.145 ;
        RECT 12.750 26.885 48.630 27.055 ;
        RECT 12.835 25.795 14.045 26.885 ;
        RECT 14.305 26.215 14.475 26.715 ;
        RECT 14.645 26.385 14.975 26.885 ;
        RECT 14.305 26.045 14.970 26.215 ;
        RECT 12.835 25.085 13.355 25.625 ;
        RECT 13.525 25.255 14.045 25.795 ;
        RECT 14.220 25.225 14.570 25.875 ;
        RECT 12.835 24.335 14.045 25.085 ;
        RECT 14.740 25.055 14.970 26.045 ;
        RECT 14.305 24.885 14.970 25.055 ;
        RECT 14.305 24.595 14.475 24.885 ;
        RECT 14.645 24.335 14.975 24.715 ;
        RECT 15.145 24.595 15.330 26.715 ;
        RECT 15.570 26.425 15.835 26.885 ;
        RECT 16.005 26.290 16.255 26.715 ;
        RECT 16.465 26.440 17.570 26.610 ;
        RECT 15.950 26.160 16.255 26.290 ;
        RECT 15.500 24.965 15.780 25.915 ;
        RECT 15.950 25.055 16.120 26.160 ;
        RECT 16.290 25.375 16.530 25.970 ;
        RECT 16.700 25.905 17.230 26.270 ;
        RECT 16.700 25.205 16.870 25.905 ;
        RECT 17.400 25.825 17.570 26.440 ;
        RECT 17.740 26.085 17.910 26.885 ;
        RECT 18.080 26.385 18.330 26.715 ;
        RECT 18.555 26.415 19.440 26.585 ;
        RECT 17.400 25.735 17.910 25.825 ;
        RECT 15.950 24.925 16.175 25.055 ;
        RECT 16.345 24.985 16.870 25.205 ;
        RECT 17.040 25.565 17.910 25.735 ;
        RECT 15.585 24.335 15.835 24.795 ;
        RECT 16.005 24.785 16.175 24.925 ;
        RECT 17.040 24.785 17.210 25.565 ;
        RECT 17.740 25.495 17.910 25.565 ;
        RECT 17.420 25.315 17.620 25.345 ;
        RECT 18.080 25.315 18.250 26.385 ;
        RECT 18.420 25.495 18.610 26.215 ;
        RECT 17.420 25.015 18.250 25.315 ;
        RECT 18.780 25.285 19.100 26.245 ;
        RECT 16.005 24.615 16.340 24.785 ;
        RECT 16.535 24.615 17.210 24.785 ;
        RECT 17.530 24.335 17.900 24.835 ;
        RECT 18.080 24.785 18.250 25.015 ;
        RECT 18.635 24.955 19.100 25.285 ;
        RECT 19.270 25.575 19.440 26.415 ;
        RECT 19.620 26.385 19.935 26.885 ;
        RECT 20.165 26.155 20.505 26.715 ;
        RECT 19.610 25.780 20.505 26.155 ;
        RECT 20.675 25.875 20.845 26.885 ;
        RECT 20.315 25.575 20.505 25.780 ;
        RECT 21.015 25.825 21.345 26.670 ;
        RECT 21.015 25.745 21.405 25.825 ;
        RECT 21.575 25.795 25.085 26.885 ;
        RECT 21.190 25.695 21.405 25.745 ;
        RECT 19.270 25.245 20.145 25.575 ;
        RECT 20.315 25.245 21.065 25.575 ;
        RECT 19.270 24.785 19.440 25.245 ;
        RECT 20.315 25.075 20.515 25.245 ;
        RECT 21.235 25.115 21.405 25.695 ;
        RECT 21.180 25.075 21.405 25.115 ;
        RECT 18.080 24.615 18.485 24.785 ;
        RECT 18.655 24.615 19.440 24.785 ;
        RECT 19.715 24.335 19.925 24.865 ;
        RECT 20.185 24.550 20.515 25.075 ;
        RECT 21.025 24.990 21.405 25.075 ;
        RECT 21.575 25.105 23.225 25.625 ;
        RECT 23.395 25.275 25.085 25.795 ;
        RECT 25.715 25.720 26.005 26.885 ;
        RECT 26.265 26.215 26.435 26.715 ;
        RECT 26.605 26.385 26.935 26.885 ;
        RECT 26.265 26.045 26.930 26.215 ;
        RECT 26.180 25.225 26.530 25.875 ;
        RECT 20.685 24.335 20.855 24.945 ;
        RECT 21.025 24.555 21.355 24.990 ;
        RECT 21.575 24.335 25.085 25.105 ;
        RECT 25.715 24.335 26.005 25.060 ;
        RECT 26.700 25.055 26.930 26.045 ;
        RECT 26.265 24.885 26.930 25.055 ;
        RECT 26.265 24.595 26.435 24.885 ;
        RECT 26.605 24.335 26.935 24.715 ;
        RECT 27.105 24.595 27.290 26.715 ;
        RECT 27.530 26.425 27.795 26.885 ;
        RECT 27.965 26.290 28.215 26.715 ;
        RECT 28.425 26.440 29.530 26.610 ;
        RECT 27.910 26.160 28.215 26.290 ;
        RECT 27.460 24.965 27.740 25.915 ;
        RECT 27.910 25.055 28.080 26.160 ;
        RECT 28.250 25.375 28.490 25.970 ;
        RECT 28.660 25.905 29.190 26.270 ;
        RECT 28.660 25.205 28.830 25.905 ;
        RECT 29.360 25.825 29.530 26.440 ;
        RECT 29.700 26.085 29.870 26.885 ;
        RECT 30.040 26.385 30.290 26.715 ;
        RECT 30.515 26.415 31.400 26.585 ;
        RECT 29.360 25.735 29.870 25.825 ;
        RECT 27.910 24.925 28.135 25.055 ;
        RECT 28.305 24.985 28.830 25.205 ;
        RECT 29.000 25.565 29.870 25.735 ;
        RECT 27.545 24.335 27.795 24.795 ;
        RECT 27.965 24.785 28.135 24.925 ;
        RECT 29.000 24.785 29.170 25.565 ;
        RECT 29.700 25.495 29.870 25.565 ;
        RECT 29.380 25.315 29.580 25.345 ;
        RECT 30.040 25.315 30.210 26.385 ;
        RECT 30.380 25.495 30.570 26.215 ;
        RECT 29.380 25.015 30.210 25.315 ;
        RECT 30.740 25.285 31.060 26.245 ;
        RECT 27.965 24.615 28.300 24.785 ;
        RECT 28.495 24.615 29.170 24.785 ;
        RECT 29.490 24.335 29.860 24.835 ;
        RECT 30.040 24.785 30.210 25.015 ;
        RECT 30.595 24.955 31.060 25.285 ;
        RECT 31.230 25.575 31.400 26.415 ;
        RECT 31.580 26.385 31.895 26.885 ;
        RECT 32.125 26.155 32.465 26.715 ;
        RECT 31.570 25.780 32.465 26.155 ;
        RECT 32.635 25.875 32.805 26.885 ;
        RECT 32.275 25.575 32.465 25.780 ;
        RECT 32.975 25.825 33.305 26.670 ;
        RECT 33.625 26.265 33.795 26.695 ;
        RECT 33.965 26.435 34.295 26.885 ;
        RECT 33.625 26.035 34.305 26.265 ;
        RECT 32.975 25.745 33.365 25.825 ;
        RECT 33.150 25.695 33.365 25.745 ;
        RECT 33.595 25.695 33.900 25.865 ;
        RECT 31.230 25.245 32.105 25.575 ;
        RECT 32.275 25.245 33.025 25.575 ;
        RECT 31.230 24.785 31.400 25.245 ;
        RECT 32.275 25.075 32.475 25.245 ;
        RECT 33.195 25.115 33.365 25.695 ;
        RECT 33.140 25.075 33.365 25.115 ;
        RECT 30.040 24.615 30.445 24.785 ;
        RECT 30.615 24.615 31.400 24.785 ;
        RECT 31.675 24.335 31.885 24.865 ;
        RECT 32.145 24.550 32.475 25.075 ;
        RECT 32.985 24.990 33.365 25.075 ;
        RECT 33.600 25.015 33.900 25.695 ;
        RECT 34.070 25.385 34.305 26.035 ;
        RECT 34.495 25.725 34.780 26.670 ;
        RECT 34.960 26.415 35.645 26.885 ;
        RECT 34.955 25.895 35.650 26.205 ;
        RECT 35.825 25.830 36.130 26.615 ;
        RECT 36.315 25.930 36.585 26.885 ;
        RECT 34.495 25.575 35.355 25.725 ;
        RECT 34.495 25.555 35.785 25.575 ;
        RECT 34.070 25.055 34.625 25.385 ;
        RECT 34.795 25.195 35.785 25.555 ;
        RECT 32.645 24.335 32.815 24.945 ;
        RECT 32.985 24.555 33.315 24.990 ;
        RECT 34.070 24.905 34.285 25.055 ;
        RECT 33.545 24.335 33.875 24.840 ;
        RECT 34.045 24.530 34.285 24.905 ;
        RECT 34.795 24.860 34.965 25.195 ;
        RECT 35.955 25.025 36.130 25.830 ;
        RECT 36.755 25.795 39.345 26.885 ;
        RECT 40.090 26.255 40.375 26.715 ;
        RECT 40.545 26.425 40.815 26.885 ;
        RECT 40.090 26.035 41.045 26.255 ;
        RECT 34.565 24.665 34.965 24.860 ;
        RECT 34.565 24.520 34.735 24.665 ;
        RECT 35.325 24.335 35.725 24.830 ;
        RECT 35.895 24.505 36.130 25.025 ;
        RECT 36.755 25.105 37.965 25.625 ;
        RECT 38.135 25.275 39.345 25.795 ;
        RECT 39.975 25.305 40.665 25.865 ;
        RECT 40.835 25.135 41.045 26.035 ;
        RECT 36.315 24.335 36.585 24.970 ;
        RECT 36.755 24.335 39.345 25.105 ;
        RECT 40.090 24.965 41.045 25.135 ;
        RECT 41.215 25.865 41.615 26.715 ;
        RECT 41.805 26.255 42.085 26.715 ;
        RECT 42.605 26.425 42.930 26.885 ;
        RECT 41.805 26.035 42.930 26.255 ;
        RECT 41.215 25.305 42.310 25.865 ;
        RECT 42.480 25.575 42.930 26.035 ;
        RECT 43.100 25.745 43.485 26.715 ;
        RECT 40.090 24.505 40.375 24.965 ;
        RECT 40.545 24.335 40.815 24.795 ;
        RECT 41.215 24.505 41.615 25.305 ;
        RECT 42.480 25.245 43.035 25.575 ;
        RECT 42.480 25.135 42.930 25.245 ;
        RECT 41.805 24.965 42.930 25.135 ;
        RECT 43.205 25.075 43.485 25.745 ;
        RECT 41.805 24.505 42.085 24.965 ;
        RECT 42.605 24.335 42.930 24.795 ;
        RECT 43.100 24.505 43.485 25.075 ;
        RECT 43.655 26.085 44.095 26.715 ;
        RECT 43.655 25.075 43.965 26.085 ;
        RECT 44.270 26.035 44.585 26.885 ;
        RECT 44.755 26.545 46.185 26.715 ;
        RECT 44.755 25.865 44.925 26.545 ;
        RECT 44.135 25.695 44.925 25.865 ;
        RECT 44.135 25.245 44.305 25.695 ;
        RECT 45.095 25.575 45.295 26.375 ;
        RECT 44.475 25.245 44.865 25.525 ;
        RECT 45.050 25.245 45.295 25.575 ;
        RECT 45.495 25.245 45.745 26.375 ;
        RECT 45.935 25.915 46.185 26.545 ;
        RECT 46.365 26.085 46.695 26.885 ;
        RECT 45.935 25.745 46.705 25.915 ;
        RECT 45.960 25.245 46.365 25.575 ;
        RECT 46.535 25.075 46.705 25.745 ;
        RECT 47.335 25.795 48.545 26.885 ;
        RECT 47.335 25.255 47.855 25.795 ;
        RECT 48.025 25.085 48.545 25.625 ;
        RECT 43.655 24.515 44.095 25.075 ;
        RECT 44.265 24.335 44.715 25.075 ;
        RECT 44.885 24.905 46.045 25.075 ;
        RECT 44.885 24.505 45.055 24.905 ;
        RECT 45.225 24.335 45.645 24.735 ;
        RECT 45.815 24.505 46.045 24.905 ;
        RECT 46.215 24.505 46.705 25.075 ;
        RECT 47.335 24.335 48.545 25.085 ;
        RECT 12.750 24.165 48.630 24.335 ;
        RECT 12.835 23.415 14.045 24.165 ;
        RECT 12.835 22.875 13.355 23.415 ;
        RECT 14.220 23.325 14.480 24.165 ;
        RECT 14.655 23.420 14.910 23.995 ;
        RECT 15.080 23.785 15.410 24.165 ;
        RECT 15.625 23.615 15.795 23.995 ;
        RECT 15.080 23.445 15.795 23.615 ;
        RECT 17.090 23.535 17.375 23.995 ;
        RECT 17.545 23.705 17.815 24.165 ;
        RECT 13.525 22.705 14.045 23.245 ;
        RECT 12.835 21.615 14.045 22.705 ;
        RECT 14.220 21.615 14.480 22.765 ;
        RECT 14.655 22.690 14.825 23.420 ;
        RECT 15.080 23.255 15.250 23.445 ;
        RECT 17.090 23.365 18.045 23.535 ;
        RECT 14.995 22.925 15.250 23.255 ;
        RECT 15.080 22.715 15.250 22.925 ;
        RECT 15.530 22.895 15.885 23.265 ;
        RECT 14.655 21.785 14.910 22.690 ;
        RECT 15.080 22.545 15.795 22.715 ;
        RECT 16.975 22.635 17.665 23.195 ;
        RECT 15.080 21.615 15.410 22.375 ;
        RECT 15.625 21.785 15.795 22.545 ;
        RECT 17.835 22.465 18.045 23.365 ;
        RECT 17.090 22.245 18.045 22.465 ;
        RECT 18.215 23.195 18.615 23.995 ;
        RECT 18.805 23.535 19.085 23.995 ;
        RECT 19.605 23.705 19.930 24.165 ;
        RECT 18.805 23.365 19.930 23.535 ;
        RECT 20.100 23.425 20.485 23.995 ;
        RECT 19.480 23.255 19.930 23.365 ;
        RECT 18.215 22.635 19.310 23.195 ;
        RECT 19.480 22.925 20.035 23.255 ;
        RECT 17.090 21.785 17.375 22.245 ;
        RECT 17.545 21.615 17.815 22.075 ;
        RECT 18.215 21.785 18.615 22.635 ;
        RECT 19.480 22.465 19.930 22.925 ;
        RECT 20.205 22.755 20.485 23.425 ;
        RECT 21.690 23.535 21.975 23.995 ;
        RECT 22.145 23.705 22.415 24.165 ;
        RECT 21.690 23.365 22.645 23.535 ;
        RECT 18.805 22.245 19.930 22.465 ;
        RECT 18.805 21.785 19.085 22.245 ;
        RECT 19.605 21.615 19.930 22.075 ;
        RECT 20.100 21.785 20.485 22.755 ;
        RECT 21.575 22.635 22.265 23.195 ;
        RECT 22.435 22.465 22.645 23.365 ;
        RECT 21.690 22.245 22.645 22.465 ;
        RECT 22.815 23.195 23.215 23.995 ;
        RECT 23.405 23.535 23.685 23.995 ;
        RECT 24.205 23.705 24.530 24.165 ;
        RECT 23.405 23.365 24.530 23.535 ;
        RECT 24.700 23.425 25.085 23.995 ;
        RECT 24.080 23.255 24.530 23.365 ;
        RECT 22.815 22.635 23.910 23.195 ;
        RECT 24.080 22.925 24.635 23.255 ;
        RECT 21.690 21.785 21.975 22.245 ;
        RECT 22.145 21.615 22.415 22.075 ;
        RECT 22.815 21.785 23.215 22.635 ;
        RECT 24.080 22.465 24.530 22.925 ;
        RECT 24.805 22.755 25.085 23.425 ;
        RECT 25.530 23.355 25.775 23.960 ;
        RECT 25.995 23.630 26.505 24.165 ;
        RECT 23.405 22.245 24.530 22.465 ;
        RECT 23.405 21.785 23.685 22.245 ;
        RECT 24.205 21.615 24.530 22.075 ;
        RECT 24.700 21.785 25.085 22.755 ;
        RECT 25.255 23.185 26.485 23.355 ;
        RECT 25.255 22.375 25.595 23.185 ;
        RECT 25.765 22.620 26.515 22.810 ;
        RECT 25.255 21.965 25.770 22.375 ;
        RECT 26.005 21.615 26.175 22.375 ;
        RECT 26.345 21.955 26.515 22.620 ;
        RECT 26.685 22.635 26.875 23.995 ;
        RECT 27.045 23.145 27.320 23.995 ;
        RECT 27.510 23.630 28.040 23.995 ;
        RECT 28.465 23.765 28.795 24.165 ;
        RECT 27.865 23.595 28.040 23.630 ;
        RECT 27.045 22.975 27.325 23.145 ;
        RECT 27.045 22.835 27.320 22.975 ;
        RECT 27.525 22.635 27.695 23.435 ;
        RECT 26.685 22.465 27.695 22.635 ;
        RECT 27.865 23.425 28.795 23.595 ;
        RECT 28.965 23.425 29.220 23.995 ;
        RECT 27.865 22.295 28.035 23.425 ;
        RECT 28.625 23.255 28.795 23.425 ;
        RECT 26.910 22.125 28.035 22.295 ;
        RECT 28.205 22.925 28.400 23.255 ;
        RECT 28.625 22.925 28.880 23.255 ;
        RECT 28.205 21.955 28.375 22.925 ;
        RECT 29.050 22.755 29.220 23.425 ;
        RECT 29.395 23.395 31.065 24.165 ;
        RECT 31.325 23.615 31.495 23.905 ;
        RECT 31.665 23.785 31.995 24.165 ;
        RECT 31.325 23.445 31.990 23.615 ;
        RECT 29.395 22.875 30.145 23.395 ;
        RECT 26.345 21.785 28.375 21.955 ;
        RECT 28.545 21.615 28.715 22.755 ;
        RECT 28.885 21.785 29.220 22.755 ;
        RECT 30.315 22.705 31.065 23.225 ;
        RECT 29.395 21.615 31.065 22.705 ;
        RECT 31.240 22.625 31.590 23.275 ;
        RECT 31.760 22.455 31.990 23.445 ;
        RECT 31.325 22.285 31.990 22.455 ;
        RECT 31.325 21.785 31.495 22.285 ;
        RECT 31.665 21.615 31.995 22.115 ;
        RECT 32.165 21.785 32.350 23.905 ;
        RECT 32.605 23.705 32.855 24.165 ;
        RECT 33.025 23.715 33.360 23.885 ;
        RECT 33.555 23.715 34.230 23.885 ;
        RECT 33.025 23.575 33.195 23.715 ;
        RECT 32.520 22.585 32.800 23.535 ;
        RECT 32.970 23.445 33.195 23.575 ;
        RECT 32.970 22.340 33.140 23.445 ;
        RECT 33.365 23.295 33.890 23.515 ;
        RECT 33.310 22.530 33.550 23.125 ;
        RECT 33.720 22.595 33.890 23.295 ;
        RECT 34.060 22.935 34.230 23.715 ;
        RECT 34.550 23.665 34.920 24.165 ;
        RECT 35.100 23.715 35.505 23.885 ;
        RECT 35.675 23.715 36.460 23.885 ;
        RECT 35.100 23.485 35.270 23.715 ;
        RECT 34.440 23.185 35.270 23.485 ;
        RECT 35.655 23.215 36.120 23.545 ;
        RECT 34.440 23.155 34.640 23.185 ;
        RECT 34.760 22.935 34.930 23.005 ;
        RECT 34.060 22.765 34.930 22.935 ;
        RECT 34.420 22.675 34.930 22.765 ;
        RECT 32.970 22.210 33.275 22.340 ;
        RECT 33.720 22.230 34.250 22.595 ;
        RECT 32.590 21.615 32.855 22.075 ;
        RECT 33.025 21.785 33.275 22.210 ;
        RECT 34.420 22.060 34.590 22.675 ;
        RECT 33.485 21.890 34.590 22.060 ;
        RECT 34.760 21.615 34.930 22.415 ;
        RECT 35.100 22.115 35.270 23.185 ;
        RECT 35.440 22.285 35.630 23.005 ;
        RECT 35.800 22.255 36.120 23.215 ;
        RECT 36.290 23.255 36.460 23.715 ;
        RECT 36.735 23.635 36.945 24.165 ;
        RECT 37.205 23.425 37.535 23.950 ;
        RECT 37.705 23.555 37.875 24.165 ;
        RECT 38.045 23.510 38.375 23.945 ;
        RECT 38.045 23.425 38.425 23.510 ;
        RECT 38.595 23.440 38.885 24.165 ;
        RECT 37.335 23.255 37.535 23.425 ;
        RECT 38.200 23.385 38.425 23.425 ;
        RECT 36.290 22.925 37.165 23.255 ;
        RECT 37.335 22.925 38.085 23.255 ;
        RECT 35.100 21.785 35.350 22.115 ;
        RECT 36.290 22.085 36.460 22.925 ;
        RECT 37.335 22.720 37.525 22.925 ;
        RECT 38.255 22.805 38.425 23.385 ;
        RECT 38.210 22.755 38.425 22.805 ;
        RECT 39.060 23.425 39.315 23.995 ;
        RECT 39.485 23.765 39.815 24.165 ;
        RECT 40.240 23.630 40.770 23.995 ;
        RECT 40.960 23.825 41.235 23.995 ;
        RECT 40.955 23.655 41.235 23.825 ;
        RECT 40.240 23.595 40.415 23.630 ;
        RECT 39.485 23.425 40.415 23.595 ;
        RECT 36.630 22.345 37.525 22.720 ;
        RECT 38.035 22.675 38.425 22.755 ;
        RECT 35.575 21.915 36.460 22.085 ;
        RECT 36.640 21.615 36.955 22.115 ;
        RECT 37.185 21.785 37.525 22.345 ;
        RECT 37.695 21.615 37.865 22.625 ;
        RECT 38.035 21.830 38.365 22.675 ;
        RECT 38.595 21.615 38.885 22.780 ;
        RECT 39.060 22.755 39.230 23.425 ;
        RECT 39.485 23.255 39.655 23.425 ;
        RECT 39.400 22.925 39.655 23.255 ;
        RECT 39.880 22.925 40.075 23.255 ;
        RECT 39.060 21.785 39.395 22.755 ;
        RECT 39.565 21.615 39.735 22.755 ;
        RECT 39.905 21.955 40.075 22.925 ;
        RECT 40.245 22.295 40.415 23.425 ;
        RECT 40.585 22.635 40.755 23.435 ;
        RECT 40.960 22.835 41.235 23.655 ;
        RECT 41.405 22.635 41.595 23.995 ;
        RECT 41.775 23.630 42.285 24.165 ;
        RECT 42.505 23.355 42.750 23.960 ;
        RECT 43.285 23.615 43.455 23.995 ;
        RECT 43.635 23.785 43.965 24.165 ;
        RECT 43.285 23.445 43.950 23.615 ;
        RECT 44.145 23.490 44.405 23.995 ;
        RECT 41.795 23.185 43.025 23.355 ;
        RECT 40.585 22.465 41.595 22.635 ;
        RECT 41.765 22.620 42.515 22.810 ;
        RECT 40.245 22.125 41.370 22.295 ;
        RECT 41.765 21.955 41.935 22.620 ;
        RECT 42.685 22.375 43.025 23.185 ;
        RECT 43.215 22.895 43.545 23.265 ;
        RECT 43.780 23.190 43.950 23.445 ;
        RECT 43.780 22.860 44.065 23.190 ;
        RECT 43.780 22.715 43.950 22.860 ;
        RECT 39.905 21.785 41.935 21.955 ;
        RECT 42.105 21.615 42.275 22.375 ;
        RECT 42.510 21.965 43.025 22.375 ;
        RECT 43.285 22.545 43.950 22.715 ;
        RECT 44.235 22.690 44.405 23.490 ;
        RECT 43.285 21.785 43.455 22.545 ;
        RECT 43.635 21.615 43.965 22.375 ;
        RECT 44.135 21.785 44.405 22.690 ;
        RECT 44.575 23.490 44.845 23.835 ;
        RECT 45.035 23.765 45.415 24.165 ;
        RECT 45.585 23.595 45.755 23.945 ;
        RECT 45.925 23.765 46.255 24.165 ;
        RECT 46.455 23.595 46.625 23.945 ;
        RECT 46.825 23.665 47.155 24.165 ;
        RECT 44.575 22.755 44.745 23.490 ;
        RECT 45.015 23.425 46.625 23.595 ;
        RECT 45.015 23.255 45.185 23.425 ;
        RECT 44.915 22.925 45.185 23.255 ;
        RECT 45.355 22.925 45.760 23.255 ;
        RECT 45.015 22.755 45.185 22.925 ;
        RECT 44.575 21.785 44.845 22.755 ;
        RECT 45.015 22.585 45.740 22.755 ;
        RECT 45.930 22.635 46.640 23.255 ;
        RECT 46.810 22.925 47.160 23.495 ;
        RECT 47.335 23.415 48.545 24.165 ;
        RECT 45.570 22.465 45.740 22.585 ;
        RECT 46.840 22.465 47.160 22.755 ;
        RECT 45.055 21.615 45.335 22.415 ;
        RECT 45.570 22.295 47.160 22.465 ;
        RECT 47.335 22.705 47.855 23.245 ;
        RECT 48.025 22.875 48.545 23.415 ;
        RECT 45.505 21.835 47.160 22.125 ;
        RECT 47.335 21.615 48.545 22.705 ;
        RECT 12.750 21.445 48.630 21.615 ;
        RECT 12.835 20.355 14.045 21.445 ;
        RECT 14.275 20.385 14.605 21.230 ;
        RECT 14.775 20.435 14.945 21.445 ;
        RECT 15.115 20.715 15.455 21.275 ;
        RECT 15.685 20.945 16.000 21.445 ;
        RECT 16.180 20.975 17.065 21.145 ;
        RECT 12.835 19.645 13.355 20.185 ;
        RECT 13.525 19.815 14.045 20.355 ;
        RECT 14.215 20.305 14.605 20.385 ;
        RECT 15.115 20.340 16.010 20.715 ;
        RECT 14.215 20.255 14.430 20.305 ;
        RECT 14.215 19.675 14.385 20.255 ;
        RECT 15.115 20.135 15.305 20.340 ;
        RECT 16.180 20.135 16.350 20.975 ;
        RECT 17.290 20.945 17.540 21.275 ;
        RECT 14.555 19.805 15.305 20.135 ;
        RECT 15.475 19.805 16.350 20.135 ;
        RECT 12.835 18.895 14.045 19.645 ;
        RECT 14.215 19.635 14.440 19.675 ;
        RECT 15.105 19.635 15.305 19.805 ;
        RECT 14.215 19.550 14.595 19.635 ;
        RECT 14.265 19.115 14.595 19.550 ;
        RECT 14.765 18.895 14.935 19.505 ;
        RECT 15.105 19.110 15.435 19.635 ;
        RECT 15.695 18.895 15.905 19.425 ;
        RECT 16.180 19.345 16.350 19.805 ;
        RECT 16.520 19.845 16.840 20.805 ;
        RECT 17.010 20.055 17.200 20.775 ;
        RECT 17.370 19.875 17.540 20.945 ;
        RECT 17.710 20.645 17.880 21.445 ;
        RECT 18.050 21.000 19.155 21.170 ;
        RECT 18.050 20.385 18.220 21.000 ;
        RECT 19.365 20.850 19.615 21.275 ;
        RECT 19.785 20.985 20.050 21.445 ;
        RECT 18.390 20.465 18.920 20.830 ;
        RECT 19.365 20.720 19.670 20.850 ;
        RECT 17.710 20.295 18.220 20.385 ;
        RECT 17.710 20.125 18.580 20.295 ;
        RECT 17.710 20.055 17.880 20.125 ;
        RECT 18.000 19.875 18.200 19.905 ;
        RECT 16.520 19.515 16.985 19.845 ;
        RECT 17.370 19.575 18.200 19.875 ;
        RECT 17.370 19.345 17.540 19.575 ;
        RECT 16.180 19.175 16.965 19.345 ;
        RECT 17.135 19.175 17.540 19.345 ;
        RECT 17.720 18.895 18.090 19.395 ;
        RECT 18.410 19.345 18.580 20.125 ;
        RECT 18.750 19.765 18.920 20.465 ;
        RECT 19.090 19.935 19.330 20.530 ;
        RECT 18.750 19.545 19.275 19.765 ;
        RECT 19.500 19.615 19.670 20.720 ;
        RECT 19.445 19.485 19.670 19.615 ;
        RECT 19.840 19.525 20.120 20.475 ;
        RECT 19.445 19.345 19.615 19.485 ;
        RECT 18.410 19.175 19.085 19.345 ;
        RECT 19.280 19.175 19.615 19.345 ;
        RECT 19.785 18.895 20.035 19.355 ;
        RECT 20.290 19.155 20.475 21.275 ;
        RECT 20.645 20.945 20.975 21.445 ;
        RECT 21.145 20.775 21.315 21.275 ;
        RECT 20.650 20.605 21.315 20.775 ;
        RECT 20.650 19.615 20.880 20.605 ;
        RECT 21.050 19.785 21.400 20.435 ;
        RECT 21.575 20.355 25.085 21.445 ;
        RECT 21.575 19.665 23.225 20.185 ;
        RECT 23.395 19.835 25.085 20.355 ;
        RECT 25.715 20.280 26.005 21.445 ;
        RECT 26.185 20.635 26.480 21.445 ;
        RECT 26.660 20.135 26.905 21.275 ;
        RECT 27.080 20.635 27.340 21.445 ;
        RECT 27.940 21.440 34.215 21.445 ;
        RECT 27.520 20.135 27.770 21.270 ;
        RECT 27.940 20.645 28.200 21.440 ;
        RECT 28.370 20.545 28.630 21.270 ;
        RECT 28.800 20.715 29.060 21.440 ;
        RECT 29.230 20.545 29.490 21.270 ;
        RECT 29.660 20.715 29.920 21.440 ;
        RECT 30.090 20.545 30.350 21.270 ;
        RECT 30.520 20.715 30.780 21.440 ;
        RECT 30.950 20.545 31.210 21.270 ;
        RECT 31.380 20.715 31.625 21.440 ;
        RECT 31.795 20.545 32.055 21.270 ;
        RECT 32.240 20.715 32.485 21.440 ;
        RECT 32.655 20.545 32.915 21.270 ;
        RECT 33.100 20.715 33.345 21.440 ;
        RECT 33.515 20.545 33.775 21.270 ;
        RECT 33.960 20.715 34.215 21.440 ;
        RECT 28.370 20.530 33.775 20.545 ;
        RECT 34.385 20.530 34.675 21.270 ;
        RECT 34.845 20.700 35.115 21.445 ;
        RECT 28.370 20.305 35.115 20.530 ;
        RECT 35.375 20.355 36.585 21.445 ;
        RECT 20.650 19.445 21.315 19.615 ;
        RECT 20.645 18.895 20.975 19.275 ;
        RECT 21.145 19.155 21.315 19.445 ;
        RECT 21.575 18.895 25.085 19.665 ;
        RECT 25.715 18.895 26.005 19.620 ;
        RECT 26.175 19.575 26.490 20.135 ;
        RECT 26.660 19.885 33.780 20.135 ;
        RECT 26.175 18.895 26.480 19.405 ;
        RECT 26.660 19.075 26.910 19.885 ;
        RECT 27.080 18.895 27.340 19.420 ;
        RECT 27.520 19.075 27.770 19.885 ;
        RECT 33.950 19.715 35.115 20.305 ;
        RECT 28.370 19.545 35.115 19.715 ;
        RECT 35.375 19.645 35.895 20.185 ;
        RECT 36.065 19.815 36.585 20.355 ;
        RECT 36.845 20.515 37.015 21.275 ;
        RECT 37.195 20.685 37.525 21.445 ;
        RECT 36.845 20.345 37.510 20.515 ;
        RECT 37.695 20.370 37.965 21.275 ;
        RECT 37.340 20.200 37.510 20.345 ;
        RECT 36.775 19.795 37.105 20.165 ;
        RECT 37.340 19.870 37.625 20.200 ;
        RECT 27.940 18.895 28.200 19.455 ;
        RECT 28.370 19.090 28.630 19.545 ;
        RECT 28.800 18.895 29.060 19.375 ;
        RECT 29.230 19.090 29.490 19.545 ;
        RECT 29.660 18.895 29.920 19.375 ;
        RECT 30.090 19.090 30.350 19.545 ;
        RECT 30.520 18.895 30.765 19.375 ;
        RECT 30.935 19.090 31.210 19.545 ;
        RECT 31.380 18.895 31.625 19.375 ;
        RECT 31.795 19.090 32.055 19.545 ;
        RECT 32.235 18.895 32.485 19.375 ;
        RECT 32.655 19.090 32.915 19.545 ;
        RECT 33.095 18.895 33.345 19.375 ;
        RECT 33.515 19.090 33.775 19.545 ;
        RECT 33.955 18.895 34.215 19.375 ;
        RECT 34.385 19.090 34.645 19.545 ;
        RECT 34.815 18.895 35.115 19.375 ;
        RECT 35.375 18.895 36.585 19.645 ;
        RECT 37.340 19.615 37.510 19.870 ;
        RECT 36.845 19.445 37.510 19.615 ;
        RECT 37.795 19.570 37.965 20.370 ;
        RECT 38.225 20.515 38.395 21.275 ;
        RECT 38.575 20.685 38.905 21.445 ;
        RECT 38.225 20.345 38.890 20.515 ;
        RECT 39.075 20.370 39.345 21.275 ;
        RECT 38.720 20.200 38.890 20.345 ;
        RECT 38.155 19.795 38.485 20.165 ;
        RECT 38.720 19.870 39.005 20.200 ;
        RECT 38.720 19.615 38.890 19.870 ;
        RECT 36.845 19.065 37.015 19.445 ;
        RECT 37.195 18.895 37.525 19.275 ;
        RECT 37.705 19.065 37.965 19.570 ;
        RECT 38.225 19.445 38.890 19.615 ;
        RECT 39.175 19.570 39.345 20.370 ;
        RECT 39.605 20.515 39.775 21.275 ;
        RECT 39.955 20.685 40.285 21.445 ;
        RECT 39.605 20.345 40.270 20.515 ;
        RECT 40.455 20.370 40.725 21.275 ;
        RECT 40.100 20.200 40.270 20.345 ;
        RECT 39.535 19.795 39.865 20.165 ;
        RECT 40.100 19.870 40.385 20.200 ;
        RECT 40.100 19.615 40.270 19.870 ;
        RECT 38.225 19.065 38.395 19.445 ;
        RECT 38.575 18.895 38.905 19.275 ;
        RECT 39.085 19.065 39.345 19.570 ;
        RECT 39.605 19.445 40.270 19.615 ;
        RECT 40.555 19.570 40.725 20.370 ;
        RECT 40.985 20.515 41.155 21.275 ;
        RECT 41.335 20.685 41.665 21.445 ;
        RECT 40.985 20.345 41.650 20.515 ;
        RECT 41.835 20.370 42.105 21.275 ;
        RECT 41.480 20.200 41.650 20.345 ;
        RECT 40.915 19.795 41.245 20.165 ;
        RECT 41.480 19.870 41.765 20.200 ;
        RECT 41.480 19.615 41.650 19.870 ;
        RECT 39.605 19.065 39.775 19.445 ;
        RECT 39.955 18.895 40.285 19.275 ;
        RECT 40.465 19.065 40.725 19.570 ;
        RECT 40.985 19.445 41.650 19.615 ;
        RECT 41.935 19.570 42.105 20.370 ;
        RECT 42.285 20.305 42.615 21.445 ;
        RECT 43.145 20.475 43.475 21.260 ;
        RECT 42.795 20.305 43.475 20.475 ;
        RECT 42.275 19.885 42.625 20.135 ;
        RECT 42.795 19.705 42.965 20.305 ;
        RECT 43.655 20.290 43.995 21.275 ;
        RECT 44.165 21.015 44.575 21.445 ;
        RECT 45.320 21.025 45.650 21.445 ;
        RECT 45.820 20.845 46.145 21.275 ;
        RECT 44.165 20.675 46.145 20.845 ;
        RECT 43.135 19.885 43.485 20.135 ;
        RECT 40.985 19.065 41.155 19.445 ;
        RECT 41.335 18.895 41.665 19.275 ;
        RECT 41.845 19.065 42.105 19.570 ;
        RECT 42.285 18.895 42.555 19.705 ;
        RECT 42.725 19.065 43.055 19.705 ;
        RECT 43.225 18.895 43.465 19.705 ;
        RECT 43.655 19.635 43.910 20.290 ;
        RECT 44.165 20.135 44.430 20.675 ;
        RECT 44.645 20.335 45.270 20.505 ;
        RECT 44.080 19.805 44.430 20.135 ;
        RECT 44.600 19.805 44.930 20.135 ;
        RECT 45.100 19.635 45.270 20.335 ;
        RECT 43.655 19.260 44.015 19.635 ;
        RECT 44.280 18.895 44.450 19.635 ;
        RECT 44.730 19.465 45.270 19.635 ;
        RECT 45.440 20.265 46.145 20.675 ;
        RECT 46.620 20.345 46.950 21.445 ;
        RECT 47.335 20.355 48.545 21.445 ;
        RECT 44.730 19.260 44.900 19.465 ;
        RECT 45.440 19.065 45.610 20.265 ;
        RECT 45.780 19.885 46.350 20.095 ;
        RECT 46.520 19.885 47.165 20.095 ;
        RECT 47.335 19.815 47.855 20.355 ;
        RECT 45.840 19.545 47.010 19.715 ;
        RECT 48.025 19.645 48.545 20.185 ;
        RECT 45.840 19.065 46.170 19.545 ;
        RECT 46.340 18.895 46.510 19.365 ;
        RECT 46.680 19.080 47.010 19.545 ;
        RECT 47.335 18.895 48.545 19.645 ;
        RECT 12.750 18.725 48.630 18.895 ;
        RECT 12.835 17.975 14.045 18.725 ;
        RECT 12.835 17.435 13.355 17.975 ;
        RECT 14.220 17.885 14.480 18.725 ;
        RECT 14.655 17.980 14.910 18.555 ;
        RECT 15.080 18.345 15.410 18.725 ;
        RECT 15.625 18.175 15.795 18.555 ;
        RECT 15.080 18.005 15.795 18.175 ;
        RECT 13.525 17.265 14.045 17.805 ;
        RECT 12.835 16.175 14.045 17.265 ;
        RECT 14.220 16.175 14.480 17.325 ;
        RECT 14.655 17.250 14.825 17.980 ;
        RECT 15.080 17.815 15.250 18.005 ;
        RECT 16.980 17.985 17.235 18.555 ;
        RECT 17.405 18.325 17.735 18.725 ;
        RECT 18.160 18.190 18.690 18.555 ;
        RECT 18.880 18.385 19.155 18.555 ;
        RECT 18.875 18.215 19.155 18.385 ;
        RECT 18.160 18.155 18.335 18.190 ;
        RECT 17.405 17.985 18.335 18.155 ;
        RECT 14.995 17.485 15.250 17.815 ;
        RECT 15.080 17.275 15.250 17.485 ;
        RECT 15.530 17.455 15.885 17.825 ;
        RECT 16.980 17.315 17.150 17.985 ;
        RECT 17.405 17.815 17.575 17.985 ;
        RECT 17.320 17.485 17.575 17.815 ;
        RECT 17.800 17.485 17.995 17.815 ;
        RECT 14.655 16.345 14.910 17.250 ;
        RECT 15.080 17.105 15.795 17.275 ;
        RECT 15.080 16.175 15.410 16.935 ;
        RECT 15.625 16.345 15.795 17.105 ;
        RECT 16.980 16.345 17.315 17.315 ;
        RECT 17.485 16.175 17.655 17.315 ;
        RECT 17.825 16.515 17.995 17.485 ;
        RECT 18.165 16.855 18.335 17.985 ;
        RECT 18.505 17.195 18.675 17.995 ;
        RECT 18.880 17.395 19.155 18.215 ;
        RECT 19.325 17.195 19.515 18.555 ;
        RECT 19.695 18.190 20.205 18.725 ;
        RECT 20.425 17.915 20.670 18.520 ;
        RECT 21.115 17.955 24.625 18.725 ;
        RECT 24.795 17.975 26.005 18.725 ;
        RECT 26.225 18.070 26.555 18.505 ;
        RECT 26.725 18.115 26.895 18.725 ;
        RECT 26.175 17.985 26.555 18.070 ;
        RECT 27.065 17.985 27.395 18.510 ;
        RECT 27.655 18.195 27.865 18.725 ;
        RECT 28.140 18.275 28.925 18.445 ;
        RECT 29.095 18.275 29.500 18.445 ;
        RECT 19.715 17.745 20.945 17.915 ;
        RECT 18.505 17.025 19.515 17.195 ;
        RECT 19.685 17.180 20.435 17.370 ;
        RECT 18.165 16.685 19.290 16.855 ;
        RECT 19.685 16.515 19.855 17.180 ;
        RECT 20.605 16.935 20.945 17.745 ;
        RECT 21.115 17.435 22.765 17.955 ;
        RECT 22.935 17.265 24.625 17.785 ;
        RECT 24.795 17.435 25.315 17.975 ;
        RECT 26.175 17.945 26.400 17.985 ;
        RECT 25.485 17.265 26.005 17.805 ;
        RECT 17.825 16.345 19.855 16.515 ;
        RECT 20.025 16.175 20.195 16.935 ;
        RECT 20.430 16.525 20.945 16.935 ;
        RECT 21.115 16.175 24.625 17.265 ;
        RECT 24.795 16.175 26.005 17.265 ;
        RECT 26.175 17.365 26.345 17.945 ;
        RECT 27.065 17.815 27.265 17.985 ;
        RECT 28.140 17.815 28.310 18.275 ;
        RECT 26.515 17.485 27.265 17.815 ;
        RECT 27.435 17.485 28.310 17.815 ;
        RECT 26.175 17.315 26.390 17.365 ;
        RECT 26.175 17.235 26.565 17.315 ;
        RECT 26.235 16.390 26.565 17.235 ;
        RECT 27.075 17.280 27.265 17.485 ;
        RECT 26.735 16.175 26.905 17.185 ;
        RECT 27.075 16.905 27.970 17.280 ;
        RECT 27.075 16.345 27.415 16.905 ;
        RECT 27.645 16.175 27.960 16.675 ;
        RECT 28.140 16.645 28.310 17.485 ;
        RECT 28.480 17.775 28.945 18.105 ;
        RECT 29.330 18.045 29.500 18.275 ;
        RECT 29.680 18.225 30.050 18.725 ;
        RECT 30.370 18.275 31.045 18.445 ;
        RECT 31.240 18.275 31.575 18.445 ;
        RECT 28.480 16.815 28.800 17.775 ;
        RECT 29.330 17.745 30.160 18.045 ;
        RECT 28.970 16.845 29.160 17.565 ;
        RECT 29.330 16.675 29.500 17.745 ;
        RECT 29.960 17.715 30.160 17.745 ;
        RECT 29.670 17.495 29.840 17.565 ;
        RECT 30.370 17.495 30.540 18.275 ;
        RECT 31.405 18.135 31.575 18.275 ;
        RECT 31.745 18.265 31.995 18.725 ;
        RECT 29.670 17.325 30.540 17.495 ;
        RECT 30.710 17.855 31.235 18.075 ;
        RECT 31.405 18.005 31.630 18.135 ;
        RECT 29.670 17.235 30.180 17.325 ;
        RECT 28.140 16.475 29.025 16.645 ;
        RECT 29.250 16.345 29.500 16.675 ;
        RECT 29.670 16.175 29.840 16.975 ;
        RECT 30.010 16.620 30.180 17.235 ;
        RECT 30.710 17.155 30.880 17.855 ;
        RECT 30.350 16.790 30.880 17.155 ;
        RECT 31.050 17.090 31.290 17.685 ;
        RECT 31.460 16.900 31.630 18.005 ;
        RECT 31.800 17.145 32.080 18.095 ;
        RECT 31.325 16.770 31.630 16.900 ;
        RECT 30.010 16.450 31.115 16.620 ;
        RECT 31.325 16.345 31.575 16.770 ;
        RECT 31.745 16.175 32.010 16.635 ;
        RECT 32.250 16.345 32.435 18.465 ;
        RECT 32.605 18.345 32.935 18.725 ;
        RECT 33.105 18.175 33.275 18.465 ;
        RECT 32.610 18.005 33.275 18.175 ;
        RECT 32.610 17.015 32.840 18.005 ;
        RECT 33.540 17.985 33.795 18.555 ;
        RECT 33.965 18.325 34.295 18.725 ;
        RECT 34.720 18.190 35.250 18.555 ;
        RECT 34.720 18.155 34.895 18.190 ;
        RECT 33.965 17.985 34.895 18.155 ;
        RECT 33.010 17.185 33.360 17.835 ;
        RECT 33.540 17.315 33.710 17.985 ;
        RECT 33.965 17.815 34.135 17.985 ;
        RECT 33.880 17.485 34.135 17.815 ;
        RECT 34.360 17.485 34.555 17.815 ;
        RECT 32.610 16.845 33.275 17.015 ;
        RECT 32.605 16.175 32.935 16.675 ;
        RECT 33.105 16.345 33.275 16.845 ;
        RECT 33.540 16.345 33.875 17.315 ;
        RECT 34.045 16.175 34.215 17.315 ;
        RECT 34.385 16.515 34.555 17.485 ;
        RECT 34.725 16.855 34.895 17.985 ;
        RECT 35.065 17.195 35.235 17.995 ;
        RECT 35.440 17.705 35.715 18.555 ;
        RECT 35.435 17.535 35.715 17.705 ;
        RECT 35.440 17.395 35.715 17.535 ;
        RECT 35.885 17.195 36.075 18.555 ;
        RECT 36.255 18.190 36.765 18.725 ;
        RECT 36.985 17.915 37.230 18.520 ;
        RECT 38.595 18.000 38.885 18.725 ;
        RECT 39.055 17.985 39.440 18.555 ;
        RECT 39.610 18.265 39.935 18.725 ;
        RECT 40.455 18.095 40.735 18.555 ;
        RECT 36.275 17.745 37.505 17.915 ;
        RECT 35.065 17.025 36.075 17.195 ;
        RECT 36.245 17.180 36.995 17.370 ;
        RECT 34.725 16.685 35.850 16.855 ;
        RECT 36.245 16.515 36.415 17.180 ;
        RECT 37.165 16.935 37.505 17.745 ;
        RECT 34.385 16.345 36.415 16.515 ;
        RECT 36.585 16.175 36.755 16.935 ;
        RECT 36.990 16.525 37.505 16.935 ;
        RECT 38.595 16.175 38.885 17.340 ;
        RECT 39.055 17.315 39.335 17.985 ;
        RECT 39.610 17.925 40.735 18.095 ;
        RECT 39.610 17.815 40.060 17.925 ;
        RECT 39.505 17.485 40.060 17.815 ;
        RECT 40.925 17.755 41.325 18.555 ;
        RECT 41.725 18.265 41.995 18.725 ;
        RECT 42.165 18.095 42.450 18.555 ;
        RECT 39.055 16.345 39.440 17.315 ;
        RECT 39.610 17.025 40.060 17.485 ;
        RECT 40.230 17.195 41.325 17.755 ;
        RECT 39.610 16.805 40.735 17.025 ;
        RECT 39.610 16.175 39.935 16.635 ;
        RECT 40.455 16.345 40.735 16.805 ;
        RECT 40.925 16.345 41.325 17.195 ;
        RECT 41.495 17.925 42.450 18.095 ;
        RECT 43.655 18.095 43.995 18.555 ;
        RECT 44.165 18.265 44.335 18.725 ;
        RECT 44.965 18.290 45.325 18.555 ;
        RECT 44.970 18.285 45.325 18.290 ;
        RECT 44.975 18.275 45.325 18.285 ;
        RECT 44.980 18.270 45.325 18.275 ;
        RECT 44.985 18.260 45.325 18.270 ;
        RECT 45.565 18.265 45.735 18.725 ;
        RECT 44.990 18.255 45.325 18.260 ;
        RECT 45.000 18.245 45.325 18.255 ;
        RECT 45.010 18.235 45.325 18.245 ;
        RECT 44.505 18.095 44.835 18.175 ;
        RECT 41.495 17.025 41.705 17.925 ;
        RECT 43.655 17.905 44.835 18.095 ;
        RECT 45.025 18.095 45.325 18.235 ;
        RECT 45.025 17.905 45.735 18.095 ;
        RECT 41.875 17.195 42.565 17.755 ;
        RECT 43.655 17.535 43.985 17.735 ;
        RECT 44.295 17.715 44.625 17.735 ;
        RECT 44.175 17.535 44.625 17.715 ;
        RECT 43.655 17.195 43.885 17.535 ;
        RECT 41.495 16.805 42.450 17.025 ;
        RECT 41.725 16.175 41.995 16.635 ;
        RECT 42.165 16.345 42.450 16.805 ;
        RECT 43.665 16.175 43.995 16.895 ;
        RECT 44.175 16.420 44.390 17.535 ;
        RECT 44.795 17.505 45.265 17.735 ;
        RECT 45.450 17.335 45.735 17.905 ;
        RECT 45.905 17.780 46.245 18.555 ;
        RECT 47.335 17.975 48.545 18.725 ;
        RECT 44.585 17.120 45.735 17.335 ;
        RECT 44.585 16.345 44.915 17.120 ;
        RECT 45.085 16.175 45.795 16.950 ;
        RECT 45.965 16.345 46.245 17.780 ;
        RECT 47.335 17.265 47.855 17.805 ;
        RECT 48.025 17.435 48.545 17.975 ;
        RECT 47.335 16.175 48.545 17.265 ;
        RECT 12.750 16.005 48.630 16.175 ;
        RECT 12.835 14.915 14.045 16.005 ;
        RECT 14.215 15.570 19.560 16.005 ;
        RECT 12.835 14.205 13.355 14.745 ;
        RECT 13.525 14.375 14.045 14.915 ;
        RECT 12.835 13.455 14.045 14.205 ;
        RECT 15.800 14.000 16.140 14.830 ;
        RECT 17.620 14.320 17.970 15.570 ;
        RECT 19.735 14.915 23.245 16.005 ;
        RECT 19.735 14.225 21.385 14.745 ;
        RECT 21.555 14.395 23.245 14.915 ;
        RECT 23.965 15.075 24.135 15.835 ;
        RECT 24.350 15.245 24.680 16.005 ;
        RECT 23.965 14.905 24.680 15.075 ;
        RECT 24.850 14.930 25.105 15.835 ;
        RECT 23.875 14.355 24.230 14.725 ;
        RECT 24.510 14.695 24.680 14.905 ;
        RECT 24.510 14.365 24.765 14.695 ;
        RECT 14.215 13.455 19.560 14.000 ;
        RECT 19.735 13.455 23.245 14.225 ;
        RECT 24.510 14.175 24.680 14.365 ;
        RECT 24.935 14.200 25.105 14.930 ;
        RECT 25.280 14.855 25.540 16.005 ;
        RECT 25.715 14.840 26.005 16.005 ;
        RECT 26.640 14.855 26.900 16.005 ;
        RECT 27.075 14.930 27.330 15.835 ;
        RECT 27.500 15.245 27.830 16.005 ;
        RECT 28.045 15.075 28.215 15.835 ;
        RECT 28.565 15.335 28.735 15.835 ;
        RECT 28.905 15.505 29.235 16.005 ;
        RECT 28.565 15.165 29.230 15.335 ;
        RECT 23.965 14.005 24.680 14.175 ;
        RECT 23.965 13.625 24.135 14.005 ;
        RECT 24.350 13.455 24.680 13.835 ;
        RECT 24.850 13.625 25.105 14.200 ;
        RECT 25.280 13.455 25.540 14.295 ;
        RECT 25.715 13.455 26.005 14.180 ;
        RECT 26.640 13.455 26.900 14.295 ;
        RECT 27.075 14.200 27.245 14.930 ;
        RECT 27.500 14.905 28.215 15.075 ;
        RECT 27.500 14.695 27.670 14.905 ;
        RECT 27.415 14.365 27.670 14.695 ;
        RECT 27.075 13.625 27.330 14.200 ;
        RECT 27.500 14.175 27.670 14.365 ;
        RECT 27.950 14.355 28.305 14.725 ;
        RECT 28.480 14.345 28.830 14.995 ;
        RECT 29.000 14.175 29.230 15.165 ;
        RECT 27.500 14.005 28.215 14.175 ;
        RECT 27.500 13.455 27.830 13.835 ;
        RECT 28.045 13.625 28.215 14.005 ;
        RECT 28.565 14.005 29.230 14.175 ;
        RECT 28.565 13.715 28.735 14.005 ;
        RECT 28.905 13.455 29.235 13.835 ;
        RECT 29.405 13.715 29.590 15.835 ;
        RECT 29.830 15.545 30.095 16.005 ;
        RECT 30.265 15.410 30.515 15.835 ;
        RECT 30.725 15.560 31.830 15.730 ;
        RECT 30.210 15.280 30.515 15.410 ;
        RECT 29.760 14.085 30.040 15.035 ;
        RECT 30.210 14.175 30.380 15.280 ;
        RECT 30.550 14.495 30.790 15.090 ;
        RECT 30.960 15.025 31.490 15.390 ;
        RECT 30.960 14.325 31.130 15.025 ;
        RECT 31.660 14.945 31.830 15.560 ;
        RECT 32.000 15.205 32.170 16.005 ;
        RECT 32.340 15.505 32.590 15.835 ;
        RECT 32.815 15.535 33.700 15.705 ;
        RECT 31.660 14.855 32.170 14.945 ;
        RECT 30.210 14.045 30.435 14.175 ;
        RECT 30.605 14.105 31.130 14.325 ;
        RECT 31.300 14.685 32.170 14.855 ;
        RECT 29.845 13.455 30.095 13.915 ;
        RECT 30.265 13.905 30.435 14.045 ;
        RECT 31.300 13.905 31.470 14.685 ;
        RECT 32.000 14.615 32.170 14.685 ;
        RECT 31.680 14.435 31.880 14.465 ;
        RECT 32.340 14.435 32.510 15.505 ;
        RECT 32.680 14.615 32.870 15.335 ;
        RECT 31.680 14.135 32.510 14.435 ;
        RECT 33.040 14.405 33.360 15.365 ;
        RECT 30.265 13.735 30.600 13.905 ;
        RECT 30.795 13.735 31.470 13.905 ;
        RECT 31.790 13.455 32.160 13.955 ;
        RECT 32.340 13.905 32.510 14.135 ;
        RECT 32.895 14.075 33.360 14.405 ;
        RECT 33.530 14.695 33.700 15.535 ;
        RECT 33.880 15.505 34.195 16.005 ;
        RECT 34.425 15.275 34.765 15.835 ;
        RECT 33.870 14.900 34.765 15.275 ;
        RECT 34.935 14.995 35.105 16.005 ;
        RECT 34.575 14.695 34.765 14.900 ;
        RECT 35.275 14.945 35.605 15.790 ;
        RECT 35.275 14.865 35.665 14.945 ;
        RECT 35.450 14.815 35.665 14.865 ;
        RECT 35.840 14.855 36.100 16.005 ;
        RECT 36.275 14.930 36.530 15.835 ;
        RECT 36.700 15.245 37.030 16.005 ;
        RECT 37.245 15.075 37.415 15.835 ;
        RECT 33.530 14.365 34.405 14.695 ;
        RECT 34.575 14.365 35.325 14.695 ;
        RECT 33.530 13.905 33.700 14.365 ;
        RECT 34.575 14.195 34.775 14.365 ;
        RECT 35.495 14.235 35.665 14.815 ;
        RECT 35.440 14.195 35.665 14.235 ;
        RECT 32.340 13.735 32.745 13.905 ;
        RECT 32.915 13.735 33.700 13.905 ;
        RECT 33.975 13.455 34.185 13.985 ;
        RECT 34.445 13.670 34.775 14.195 ;
        RECT 35.285 14.110 35.665 14.195 ;
        RECT 34.945 13.455 35.115 14.065 ;
        RECT 35.285 13.675 35.615 14.110 ;
        RECT 35.840 13.455 36.100 14.295 ;
        RECT 36.275 14.200 36.445 14.930 ;
        RECT 36.700 14.905 37.415 15.075 ;
        RECT 36.700 14.695 36.870 14.905 ;
        RECT 38.595 14.840 38.885 16.005 ;
        RECT 40.065 15.075 40.235 15.835 ;
        RECT 40.450 15.245 40.780 16.005 ;
        RECT 40.065 14.905 40.780 15.075 ;
        RECT 40.950 14.930 41.205 15.835 ;
        RECT 36.615 14.365 36.870 14.695 ;
        RECT 36.275 13.625 36.530 14.200 ;
        RECT 36.700 14.175 36.870 14.365 ;
        RECT 37.150 14.355 37.505 14.725 ;
        RECT 39.975 14.355 40.330 14.725 ;
        RECT 40.610 14.695 40.780 14.905 ;
        RECT 40.610 14.365 40.865 14.695 ;
        RECT 36.700 14.005 37.415 14.175 ;
        RECT 36.700 13.455 37.030 13.835 ;
        RECT 37.245 13.625 37.415 14.005 ;
        RECT 38.595 13.455 38.885 14.180 ;
        RECT 40.610 14.175 40.780 14.365 ;
        RECT 41.035 14.200 41.205 14.930 ;
        RECT 41.380 14.855 41.640 16.005 ;
        RECT 41.815 14.930 42.085 15.835 ;
        RECT 42.255 15.245 42.585 16.005 ;
        RECT 42.765 15.075 42.945 15.835 ;
        RECT 44.205 15.385 44.375 15.815 ;
        RECT 44.545 15.555 44.875 16.005 ;
        RECT 44.205 15.155 44.880 15.385 ;
        RECT 40.065 14.005 40.780 14.175 ;
        RECT 40.065 13.625 40.235 14.005 ;
        RECT 40.450 13.455 40.780 13.835 ;
        RECT 40.950 13.625 41.205 14.200 ;
        RECT 41.380 13.455 41.640 14.295 ;
        RECT 41.815 14.130 41.995 14.930 ;
        RECT 42.270 14.905 42.945 15.075 ;
        RECT 42.270 14.760 42.440 14.905 ;
        RECT 42.165 14.430 42.440 14.760 ;
        RECT 42.270 14.175 42.440 14.430 ;
        RECT 42.665 14.355 43.005 14.725 ;
        RECT 41.815 13.625 42.075 14.130 ;
        RECT 42.270 14.005 42.935 14.175 ;
        RECT 44.175 14.135 44.475 14.985 ;
        RECT 44.645 14.505 44.880 15.155 ;
        RECT 45.050 14.845 45.335 15.790 ;
        RECT 45.515 15.535 46.200 16.005 ;
        RECT 45.510 15.015 46.205 15.325 ;
        RECT 46.380 14.950 46.685 15.735 ;
        RECT 45.050 14.695 45.910 14.845 ;
        RECT 45.050 14.675 46.335 14.695 ;
        RECT 44.645 14.175 45.180 14.505 ;
        RECT 45.350 14.315 46.335 14.675 ;
        RECT 44.645 14.025 44.865 14.175 ;
        RECT 42.255 13.455 42.585 13.835 ;
        RECT 42.765 13.625 42.935 14.005 ;
        RECT 44.120 13.455 44.455 13.960 ;
        RECT 44.625 13.650 44.865 14.025 ;
        RECT 45.350 13.980 45.520 14.315 ;
        RECT 46.510 14.145 46.685 14.950 ;
        RECT 47.335 14.915 48.545 16.005 ;
        RECT 47.335 14.375 47.855 14.915 ;
        RECT 48.025 14.205 48.545 14.745 ;
        RECT 45.145 13.785 45.520 13.980 ;
        RECT 45.145 13.640 45.315 13.785 ;
        RECT 45.880 13.455 46.275 13.950 ;
        RECT 46.445 13.625 46.685 14.145 ;
        RECT 47.335 13.455 48.545 14.205 ;
        RECT 12.750 13.285 48.630 13.455 ;
      LAYER met1 ;
        RECT 17.430 204.390 143.010 204.870 ;
        RECT 76.380 204.190 76.700 204.250 ;
        RECT 77.315 204.190 77.605 204.235 ;
        RECT 76.380 204.050 77.605 204.190 ;
        RECT 76.380 203.990 76.700 204.050 ;
        RECT 77.315 204.005 77.605 204.050 ;
        RECT 77.760 203.510 78.080 203.570 ;
        RECT 78.235 203.510 78.525 203.555 ;
        RECT 77.760 203.370 78.525 203.510 ;
        RECT 77.760 203.310 78.080 203.370 ;
        RECT 78.235 203.325 78.525 203.370 ;
        RECT 17.430 201.670 143.010 202.150 ;
        RECT 17.430 198.950 143.010 199.430 ;
        RECT 17.430 196.230 143.010 196.710 ;
        RECT 17.430 193.510 143.010 193.990 ;
        RECT 58.900 192.630 59.220 192.690 ;
        RECT 68.115 192.630 68.405 192.675 ;
        RECT 58.900 192.490 68.405 192.630 ;
        RECT 58.900 192.430 59.220 192.490 ;
        RECT 68.115 192.445 68.405 192.490 ;
        RECT 70.415 192.630 70.705 192.675 ;
        RECT 71.320 192.630 71.640 192.690 ;
        RECT 72.240 192.675 72.560 192.690 ;
        RECT 70.415 192.490 71.640 192.630 ;
        RECT 70.415 192.445 70.705 192.490 ;
        RECT 71.320 192.430 71.640 192.490 ;
        RECT 72.210 192.445 72.560 192.675 ;
        RECT 72.240 192.430 72.560 192.445 ;
        RECT 81.440 192.630 81.760 192.690 ;
        RECT 83.755 192.630 84.045 192.675 ;
        RECT 81.440 192.490 84.045 192.630 ;
        RECT 81.440 192.430 81.760 192.490 ;
        RECT 83.755 192.445 84.045 192.490 ;
        RECT 118.715 192.630 119.005 192.675 ;
        RECT 120.540 192.630 120.860 192.690 ;
        RECT 118.715 192.490 120.860 192.630 ;
        RECT 118.715 192.445 119.005 192.490 ;
        RECT 120.540 192.430 120.860 192.490 ;
        RECT 70.860 192.090 71.180 192.350 ;
        RECT 71.755 192.290 72.045 192.335 ;
        RECT 72.945 192.290 73.235 192.335 ;
        RECT 75.465 192.290 75.755 192.335 ;
        RECT 71.755 192.150 75.755 192.290 ;
        RECT 71.755 192.105 72.045 192.150 ;
        RECT 72.945 192.105 73.235 192.150 ;
        RECT 75.465 192.105 75.755 192.150 ;
        RECT 78.680 192.290 79.000 192.350 ;
        RECT 80.995 192.290 81.285 192.335 ;
        RECT 78.680 192.150 81.285 192.290 ;
        RECT 78.680 192.090 79.000 192.150 ;
        RECT 80.995 192.105 81.285 192.150 ;
        RECT 66.260 191.950 66.580 192.010 ;
        RECT 69.955 191.950 70.245 191.995 ;
        RECT 66.260 191.810 70.245 191.950 ;
        RECT 66.260 191.750 66.580 191.810 ;
        RECT 69.955 191.765 70.245 191.810 ;
        RECT 71.360 191.950 71.650 191.995 ;
        RECT 73.460 191.950 73.750 191.995 ;
        RECT 75.030 191.950 75.320 191.995 ;
        RECT 71.360 191.810 75.320 191.950 ;
        RECT 71.360 191.765 71.650 191.810 ;
        RECT 73.460 191.765 73.750 191.810 ;
        RECT 75.030 191.765 75.320 191.810 ;
        RECT 77.760 191.750 78.080 192.010 ;
        RECT 67.180 191.410 67.500 191.670 ;
        RECT 78.220 191.410 78.540 191.670 ;
        RECT 83.280 191.410 83.600 191.670 ;
        RECT 117.780 191.410 118.100 191.670 ;
        RECT 17.430 190.790 143.010 191.270 ;
        RECT 78.220 190.590 78.540 190.650 ;
        RECT 103.995 190.590 104.285 190.635 ;
        RECT 72.330 190.450 78.540 190.590 ;
        RECT 68.575 189.570 68.865 189.615 ;
        RECT 69.020 189.570 69.340 189.630 ;
        RECT 68.575 189.430 69.340 189.570 ;
        RECT 68.575 189.385 68.865 189.430 ;
        RECT 69.020 189.370 69.340 189.430 ;
        RECT 69.955 189.385 70.245 189.615 ;
        RECT 70.400 189.570 70.720 189.630 ;
        RECT 72.330 189.615 72.470 190.450 ;
        RECT 78.220 190.390 78.540 190.450 ;
        RECT 102.690 190.450 104.285 190.590 ;
        RECT 74.540 190.250 74.860 190.310 ;
        RECT 72.790 190.110 74.860 190.250 ;
        RECT 72.790 189.955 72.930 190.110 ;
        RECT 74.540 190.050 74.860 190.110 ;
        RECT 75.040 190.250 75.330 190.295 ;
        RECT 77.140 190.250 77.430 190.295 ;
        RECT 78.710 190.250 79.000 190.295 ;
        RECT 75.040 190.110 79.000 190.250 ;
        RECT 75.040 190.065 75.330 190.110 ;
        RECT 77.140 190.065 77.430 190.110 ;
        RECT 78.710 190.065 79.000 190.110 ;
        RECT 98.460 190.250 98.750 190.295 ;
        RECT 100.030 190.250 100.320 190.295 ;
        RECT 102.130 190.250 102.420 190.295 ;
        RECT 98.460 190.110 102.420 190.250 ;
        RECT 98.460 190.065 98.750 190.110 ;
        RECT 100.030 190.065 100.320 190.110 ;
        RECT 102.130 190.065 102.420 190.110 ;
        RECT 72.715 189.725 73.005 189.955 ;
        RECT 75.435 189.910 75.725 189.955 ;
        RECT 76.625 189.910 76.915 189.955 ;
        RECT 79.145 189.910 79.435 189.955 ;
        RECT 73.250 189.770 75.275 189.910 ;
        RECT 70.875 189.570 71.165 189.615 ;
        RECT 70.400 189.430 71.165 189.570 ;
        RECT 70.030 189.230 70.170 189.385 ;
        RECT 70.400 189.370 70.720 189.430 ;
        RECT 70.875 189.385 71.165 189.430 ;
        RECT 72.255 189.385 72.545 189.615 ;
        RECT 71.320 189.230 71.640 189.290 ;
        RECT 70.030 189.090 71.640 189.230 ;
        RECT 71.320 189.030 71.640 189.090 ;
        RECT 73.250 188.950 73.390 189.770 ;
        RECT 73.620 189.570 73.940 189.630 ;
        RECT 74.555 189.570 74.845 189.615 ;
        RECT 73.620 189.430 74.845 189.570 ;
        RECT 75.135 189.570 75.275 189.770 ;
        RECT 75.435 189.770 79.435 189.910 ;
        RECT 75.435 189.725 75.725 189.770 ;
        RECT 76.625 189.725 76.915 189.770 ;
        RECT 79.145 189.725 79.435 189.770 ;
        RECT 98.025 189.910 98.315 189.955 ;
        RECT 100.545 189.910 100.835 189.955 ;
        RECT 101.735 189.910 102.025 189.955 ;
        RECT 102.690 189.910 102.830 190.450 ;
        RECT 103.995 190.405 104.285 190.450 ;
        RECT 115.480 190.250 115.770 190.295 ;
        RECT 117.050 190.250 117.340 190.295 ;
        RECT 119.150 190.250 119.440 190.295 ;
        RECT 115.480 190.110 119.440 190.250 ;
        RECT 115.480 190.065 115.770 190.110 ;
        RECT 117.050 190.065 117.340 190.110 ;
        RECT 119.150 190.065 119.440 190.110 ;
        RECT 122.840 190.250 123.130 190.295 ;
        RECT 124.410 190.250 124.700 190.295 ;
        RECT 126.510 190.250 126.800 190.295 ;
        RECT 122.840 190.110 126.800 190.250 ;
        RECT 122.840 190.065 123.130 190.110 ;
        RECT 124.410 190.065 124.700 190.110 ;
        RECT 126.510 190.065 126.800 190.110 ;
        RECT 98.025 189.770 102.025 189.910 ;
        RECT 98.025 189.725 98.315 189.770 ;
        RECT 100.545 189.725 100.835 189.770 ;
        RECT 101.735 189.725 102.025 189.770 ;
        RECT 102.230 189.770 102.830 189.910 ;
        RECT 82.375 189.570 82.665 189.615 ;
        RECT 75.135 189.430 82.665 189.570 ;
        RECT 73.620 189.370 73.940 189.430 ;
        RECT 74.555 189.385 74.845 189.430 ;
        RECT 82.375 189.385 82.665 189.430 ;
        RECT 93.415 189.385 93.705 189.615 ;
        RECT 94.335 189.570 94.625 189.615 ;
        RECT 99.840 189.570 100.160 189.630 ;
        RECT 94.335 189.430 100.160 189.570 ;
        RECT 94.335 189.385 94.625 189.430 ;
        RECT 75.780 189.230 76.070 189.275 ;
        RECT 74.170 189.090 76.070 189.230 ;
        RECT 65.355 188.890 65.645 188.935 ;
        RECT 66.720 188.890 67.040 188.950 ;
        RECT 65.355 188.750 67.040 188.890 ;
        RECT 65.355 188.705 65.645 188.750 ;
        RECT 66.720 188.690 67.040 188.750 ;
        RECT 70.415 188.890 70.705 188.935 ;
        RECT 73.160 188.890 73.480 188.950 ;
        RECT 74.170 188.935 74.310 189.090 ;
        RECT 75.780 189.045 76.070 189.090 ;
        RECT 77.760 189.230 78.080 189.290 ;
        RECT 83.295 189.230 83.585 189.275 ;
        RECT 77.760 189.090 83.585 189.230 ;
        RECT 93.490 189.230 93.630 189.385 ;
        RECT 99.840 189.370 100.160 189.430 ;
        RECT 101.335 189.570 101.625 189.615 ;
        RECT 102.230 189.570 102.370 189.770 ;
        RECT 103.995 189.725 104.285 189.955 ;
        RECT 104.455 189.910 104.745 189.955 ;
        RECT 106.755 189.910 107.045 189.955 ;
        RECT 108.120 189.910 108.440 189.970 ;
        RECT 104.455 189.770 106.050 189.910 ;
        RECT 104.455 189.725 104.745 189.770 ;
        RECT 101.335 189.430 102.370 189.570 ;
        RECT 101.335 189.385 101.625 189.430 ;
        RECT 102.600 189.370 102.920 189.630 ;
        RECT 103.075 189.230 103.365 189.275 ;
        RECT 103.520 189.230 103.840 189.290 ;
        RECT 93.490 189.090 103.840 189.230 ;
        RECT 77.760 189.030 78.080 189.090 ;
        RECT 83.295 189.045 83.585 189.090 ;
        RECT 103.075 189.045 103.365 189.090 ;
        RECT 103.520 189.030 103.840 189.090 ;
        RECT 70.415 188.750 73.480 188.890 ;
        RECT 70.415 188.705 70.705 188.750 ;
        RECT 73.160 188.690 73.480 188.750 ;
        RECT 74.095 188.705 74.385 188.935 ;
        RECT 78.680 188.890 79.000 188.950 ;
        RECT 81.455 188.890 81.745 188.935 ;
        RECT 78.680 188.750 81.745 188.890 ;
        RECT 78.680 188.690 79.000 188.750 ;
        RECT 81.455 188.705 81.745 188.750 ;
        RECT 84.200 188.690 84.520 188.950 ;
        RECT 93.875 188.890 94.165 188.935 ;
        RECT 94.780 188.890 95.100 188.950 ;
        RECT 93.875 188.750 95.100 188.890 ;
        RECT 93.875 188.705 94.165 188.750 ;
        RECT 94.780 188.690 95.100 188.750 ;
        RECT 95.700 188.690 96.020 188.950 ;
        RECT 101.220 188.890 101.540 188.950 ;
        RECT 104.070 188.890 104.210 189.725 ;
        RECT 104.915 189.385 105.205 189.615 ;
        RECT 101.220 188.750 104.210 188.890 ;
        RECT 104.990 188.890 105.130 189.385 ;
        RECT 105.360 189.370 105.680 189.630 ;
        RECT 105.910 189.615 106.050 189.770 ;
        RECT 106.755 189.770 108.440 189.910 ;
        RECT 106.755 189.725 107.045 189.770 ;
        RECT 108.120 189.710 108.440 189.770 ;
        RECT 115.045 189.910 115.335 189.955 ;
        RECT 117.565 189.910 117.855 189.955 ;
        RECT 118.755 189.910 119.045 189.955 ;
        RECT 115.045 189.770 119.045 189.910 ;
        RECT 115.045 189.725 115.335 189.770 ;
        RECT 117.565 189.725 117.855 189.770 ;
        RECT 118.755 189.725 119.045 189.770 ;
        RECT 122.405 189.910 122.695 189.955 ;
        RECT 124.925 189.910 125.215 189.955 ;
        RECT 126.115 189.910 126.405 189.955 ;
        RECT 122.405 189.770 126.405 189.910 ;
        RECT 122.405 189.725 122.695 189.770 ;
        RECT 124.925 189.725 125.215 189.770 ;
        RECT 126.115 189.725 126.405 189.770 ;
        RECT 105.835 189.570 106.125 189.615 ;
        RECT 110.420 189.570 110.740 189.630 ;
        RECT 105.835 189.430 110.740 189.570 ;
        RECT 105.835 189.385 106.125 189.430 ;
        RECT 110.420 189.370 110.740 189.430 ;
        RECT 119.635 189.570 119.925 189.615 ;
        RECT 126.995 189.570 127.285 189.615 ;
        RECT 128.820 189.570 129.140 189.630 ;
        RECT 119.635 189.430 129.140 189.570 ;
        RECT 119.635 189.385 119.925 189.430 ;
        RECT 126.995 189.385 127.285 189.430 ;
        RECT 128.820 189.370 129.140 189.430 ;
        RECT 109.960 189.230 110.280 189.290 ;
        RECT 106.370 189.090 110.280 189.230 ;
        RECT 106.370 188.890 106.510 189.090 ;
        RECT 109.960 189.030 110.280 189.090 ;
        RECT 117.320 189.230 117.640 189.290 ;
        RECT 118.300 189.230 118.590 189.275 ;
        RECT 117.320 189.090 118.590 189.230 ;
        RECT 117.320 189.030 117.640 189.090 ;
        RECT 118.300 189.045 118.590 189.090 ;
        RECT 119.160 189.230 119.480 189.290 ;
        RECT 125.660 189.230 125.950 189.275 ;
        RECT 119.160 189.090 125.950 189.230 ;
        RECT 119.160 189.030 119.480 189.090 ;
        RECT 125.660 189.045 125.950 189.090 ;
        RECT 104.990 188.750 106.510 188.890 ;
        RECT 106.755 188.890 107.045 188.935 ;
        RECT 109.040 188.890 109.360 188.950 ;
        RECT 106.755 188.750 109.360 188.890 ;
        RECT 101.220 188.690 101.540 188.750 ;
        RECT 106.755 188.705 107.045 188.750 ;
        RECT 109.040 188.690 109.360 188.750 ;
        RECT 112.720 188.690 113.040 188.950 ;
        RECT 120.095 188.890 120.385 188.935 ;
        RECT 120.540 188.890 120.860 188.950 ;
        RECT 120.095 188.750 120.860 188.890 ;
        RECT 120.095 188.705 120.385 188.750 ;
        RECT 120.540 188.690 120.860 188.750 ;
        RECT 17.430 188.070 143.010 188.550 ;
        RECT 58.900 187.870 59.220 187.930 ;
        RECT 55.770 187.730 59.220 187.870 ;
        RECT 55.770 187.575 55.910 187.730 ;
        RECT 58.900 187.670 59.220 187.730 ;
        RECT 70.860 187.670 71.180 187.930 ;
        RECT 71.320 187.870 71.640 187.930 ;
        RECT 74.080 187.870 74.400 187.930 ;
        RECT 76.395 187.870 76.685 187.915 ;
        RECT 71.320 187.730 76.685 187.870 ;
        RECT 71.320 187.670 71.640 187.730 ;
        RECT 74.080 187.670 74.400 187.730 ;
        RECT 76.395 187.685 76.685 187.730 ;
        RECT 118.715 187.870 119.005 187.915 ;
        RECT 119.160 187.870 119.480 187.930 ;
        RECT 118.715 187.730 119.480 187.870 ;
        RECT 118.715 187.685 119.005 187.730 ;
        RECT 119.160 187.670 119.480 187.730 ;
        RECT 55.695 187.345 55.985 187.575 ;
        RECT 70.950 187.530 71.090 187.670 ;
        RECT 73.620 187.530 73.940 187.590 ;
        RECT 65.890 187.390 73.940 187.530 ;
        RECT 64.420 187.235 64.740 187.250 ;
        RECT 65.890 187.235 66.030 187.390 ;
        RECT 64.420 187.005 64.770 187.235 ;
        RECT 65.815 187.005 66.105 187.235 ;
        RECT 64.420 186.990 64.740 187.005 ;
        RECT 66.260 186.990 66.580 187.250 ;
        RECT 66.720 186.990 67.040 187.250 ;
        RECT 69.570 187.235 69.710 187.390 ;
        RECT 73.620 187.330 73.940 187.390 ;
        RECT 80.075 187.530 80.365 187.575 ;
        RECT 84.200 187.530 84.520 187.590 ;
        RECT 80.075 187.390 84.520 187.530 ;
        RECT 80.075 187.345 80.365 187.390 ;
        RECT 84.200 187.330 84.520 187.390 ;
        RECT 94.320 187.530 94.640 187.590 ;
        RECT 102.600 187.530 102.920 187.590 ;
        RECT 94.320 187.390 102.920 187.530 ;
        RECT 94.320 187.330 94.640 187.390 ;
        RECT 69.495 187.005 69.785 187.235 ;
        RECT 70.830 187.190 71.120 187.235 ;
        RECT 72.700 187.190 73.020 187.250 ;
        RECT 70.830 187.050 73.020 187.190 ;
        RECT 70.830 187.005 71.120 187.050 ;
        RECT 72.700 186.990 73.020 187.050 ;
        RECT 74.540 187.190 74.860 187.250 ;
        RECT 78.235 187.190 78.525 187.235 ;
        RECT 81.900 187.190 82.220 187.250 ;
        RECT 74.540 187.050 82.220 187.190 ;
        RECT 74.540 186.990 74.860 187.050 ;
        RECT 78.235 187.005 78.525 187.050 ;
        RECT 81.900 186.990 82.220 187.050 ;
        RECT 84.660 186.990 84.980 187.250 ;
        RECT 85.580 186.990 85.900 187.250 ;
        RECT 100.875 187.190 101.165 187.235 ;
        RECT 101.680 187.190 102.000 187.250 ;
        RECT 102.230 187.235 102.370 187.390 ;
        RECT 102.600 187.330 102.920 187.390 ;
        RECT 100.875 187.050 102.000 187.190 ;
        RECT 100.875 187.005 101.165 187.050 ;
        RECT 101.680 186.990 102.000 187.050 ;
        RECT 102.155 187.190 102.445 187.235 ;
        RECT 107.215 187.190 107.505 187.235 ;
        RECT 102.155 187.050 107.505 187.190 ;
        RECT 102.155 187.005 102.445 187.050 ;
        RECT 107.215 187.005 107.505 187.050 ;
        RECT 107.660 187.190 107.980 187.250 ;
        RECT 108.495 187.190 108.785 187.235 ;
        RECT 107.660 187.050 108.785 187.190 ;
        RECT 107.660 186.990 107.980 187.050 ;
        RECT 108.495 187.005 108.785 187.050 ;
        RECT 115.020 187.190 115.340 187.250 ;
        RECT 116.415 187.190 116.705 187.235 ;
        RECT 115.020 187.050 116.705 187.190 ;
        RECT 115.020 186.990 115.340 187.050 ;
        RECT 116.415 187.005 116.705 187.050 ;
        RECT 116.860 186.990 117.180 187.250 ;
        RECT 36.375 186.665 36.665 186.895 ;
        RECT 34.980 186.510 35.300 186.570 ;
        RECT 36.450 186.510 36.590 186.665 ;
        RECT 37.740 186.650 38.060 186.910 ;
        RECT 38.200 186.650 38.520 186.910 ;
        RECT 38.800 186.850 39.090 186.895 ;
        RECT 41.880 186.850 42.200 186.910 ;
        RECT 38.800 186.710 42.200 186.850 ;
        RECT 38.800 186.665 39.090 186.710 ;
        RECT 41.880 186.650 42.200 186.710 ;
        RECT 61.225 186.850 61.515 186.895 ;
        RECT 63.745 186.850 64.035 186.895 ;
        RECT 64.935 186.850 65.225 186.895 ;
        RECT 61.225 186.710 65.225 186.850 ;
        RECT 61.225 186.665 61.515 186.710 ;
        RECT 63.745 186.665 64.035 186.710 ;
        RECT 64.935 186.665 65.225 186.710 ;
        RECT 67.640 186.650 67.960 186.910 ;
        RECT 68.100 186.650 68.420 186.910 ;
        RECT 70.375 186.850 70.665 186.895 ;
        RECT 71.565 186.850 71.855 186.895 ;
        RECT 74.085 186.850 74.375 186.895 ;
        RECT 70.375 186.710 74.375 186.850 ;
        RECT 70.375 186.665 70.665 186.710 ;
        RECT 71.565 186.665 71.855 186.710 ;
        RECT 74.085 186.665 74.375 186.710 ;
        RECT 77.775 186.850 78.065 186.895 ;
        RECT 78.680 186.850 79.000 186.910 ;
        RECT 77.775 186.710 79.000 186.850 ;
        RECT 77.775 186.665 78.065 186.710 ;
        RECT 78.680 186.650 79.000 186.710 ;
        RECT 79.600 186.650 79.920 186.910 ;
        RECT 83.295 186.665 83.585 186.895 ;
        RECT 61.660 186.510 61.950 186.555 ;
        RECT 63.230 186.510 63.520 186.555 ;
        RECT 65.330 186.510 65.620 186.555 ;
        RECT 34.980 186.370 39.350 186.510 ;
        RECT 34.980 186.310 35.300 186.370 ;
        RECT 39.210 186.230 39.350 186.370 ;
        RECT 61.660 186.370 65.620 186.510 ;
        RECT 61.660 186.325 61.950 186.370 ;
        RECT 63.230 186.325 63.520 186.370 ;
        RECT 65.330 186.325 65.620 186.370 ;
        RECT 69.980 186.510 70.270 186.555 ;
        RECT 72.080 186.510 72.370 186.555 ;
        RECT 73.650 186.510 73.940 186.555 ;
        RECT 69.980 186.370 73.940 186.510 ;
        RECT 78.770 186.510 78.910 186.650 ;
        RECT 83.370 186.510 83.510 186.665 ;
        RECT 92.940 186.650 93.260 186.910 ;
        RECT 97.565 186.850 97.855 186.895 ;
        RECT 100.085 186.850 100.375 186.895 ;
        RECT 101.275 186.850 101.565 186.895 ;
        RECT 97.565 186.710 101.565 186.850 ;
        RECT 97.565 186.665 97.855 186.710 ;
        RECT 100.085 186.665 100.375 186.710 ;
        RECT 101.275 186.665 101.565 186.710 ;
        RECT 102.615 186.665 102.905 186.895 ;
        RECT 108.095 186.850 108.385 186.895 ;
        RECT 109.285 186.850 109.575 186.895 ;
        RECT 111.805 186.850 112.095 186.895 ;
        RECT 108.095 186.710 112.095 186.850 ;
        RECT 108.095 186.665 108.385 186.710 ;
        RECT 109.285 186.665 109.575 186.710 ;
        RECT 111.805 186.665 112.095 186.710 ;
        RECT 115.955 186.850 116.245 186.895 ;
        RECT 117.780 186.850 118.100 186.910 ;
        RECT 115.955 186.710 118.100 186.850 ;
        RECT 115.955 186.665 116.245 186.710 ;
        RECT 78.770 186.370 83.510 186.510 ;
        RECT 98.000 186.510 98.290 186.555 ;
        RECT 99.570 186.510 99.860 186.555 ;
        RECT 101.670 186.510 101.960 186.555 ;
        RECT 98.000 186.370 101.960 186.510 ;
        RECT 69.980 186.325 70.270 186.370 ;
        RECT 72.080 186.325 72.370 186.370 ;
        RECT 73.650 186.325 73.940 186.370 ;
        RECT 98.000 186.325 98.290 186.370 ;
        RECT 99.570 186.325 99.860 186.370 ;
        RECT 101.670 186.325 101.960 186.370 ;
        RECT 39.120 185.970 39.440 186.230 ;
        RECT 39.580 185.970 39.900 186.230 ;
        RECT 55.220 185.970 55.540 186.230 ;
        RECT 68.560 185.970 68.880 186.230 ;
        RECT 76.840 185.970 77.160 186.230 ;
        RECT 77.300 186.170 77.620 186.230 ;
        RECT 80.535 186.170 80.825 186.215 ;
        RECT 77.300 186.030 80.825 186.170 ;
        RECT 77.300 185.970 77.620 186.030 ;
        RECT 80.535 185.985 80.825 186.030 ;
        RECT 80.980 186.170 81.300 186.230 ;
        RECT 85.595 186.170 85.885 186.215 ;
        RECT 80.980 186.030 85.885 186.170 ;
        RECT 80.980 185.970 81.300 186.030 ;
        RECT 85.595 185.985 85.885 186.030 ;
        RECT 89.720 186.170 90.040 186.230 ;
        RECT 90.195 186.170 90.485 186.215 ;
        RECT 89.720 186.030 90.485 186.170 ;
        RECT 89.720 185.970 90.040 186.030 ;
        RECT 90.195 185.985 90.485 186.030 ;
        RECT 95.240 186.170 95.560 186.230 ;
        RECT 100.760 186.170 101.080 186.230 ;
        RECT 102.690 186.170 102.830 186.665 ;
        RECT 117.780 186.650 118.100 186.710 ;
        RECT 107.700 186.510 107.990 186.555 ;
        RECT 109.800 186.510 110.090 186.555 ;
        RECT 111.370 186.510 111.660 186.555 ;
        RECT 107.700 186.370 111.660 186.510 ;
        RECT 107.700 186.325 107.990 186.370 ;
        RECT 109.800 186.325 110.090 186.370 ;
        RECT 111.370 186.325 111.660 186.370 ;
        RECT 95.240 186.030 102.830 186.170 ;
        RECT 105.360 186.170 105.680 186.230 ;
        RECT 105.835 186.170 106.125 186.215 ;
        RECT 105.360 186.030 106.125 186.170 ;
        RECT 95.240 185.970 95.560 186.030 ;
        RECT 100.760 185.970 101.080 186.030 ;
        RECT 105.360 185.970 105.680 186.030 ;
        RECT 105.835 185.985 106.125 186.030 ;
        RECT 113.180 186.170 113.500 186.230 ;
        RECT 114.115 186.170 114.405 186.215 ;
        RECT 113.180 186.030 114.405 186.170 ;
        RECT 113.180 185.970 113.500 186.030 ;
        RECT 114.115 185.985 114.405 186.030 ;
        RECT 17.430 185.350 143.010 185.830 ;
        RECT 38.200 185.150 38.520 185.210 ;
        RECT 54.300 185.150 54.620 185.210 ;
        RECT 36.940 185.010 54.620 185.150 ;
        RECT 23.520 184.810 23.810 184.855 ;
        RECT 25.620 184.810 25.910 184.855 ;
        RECT 27.190 184.810 27.480 184.855 ;
        RECT 23.520 184.670 27.480 184.810 ;
        RECT 23.520 184.625 23.810 184.670 ;
        RECT 25.620 184.625 25.910 184.670 ;
        RECT 27.190 184.625 27.480 184.670 ;
        RECT 29.920 184.610 30.240 184.870 ;
        RECT 30.380 184.810 30.700 184.870 ;
        RECT 36.940 184.810 37.080 185.010 ;
        RECT 38.200 184.950 38.520 185.010 ;
        RECT 54.300 184.950 54.620 185.010 ;
        RECT 64.420 184.950 64.740 185.210 ;
        RECT 68.575 185.150 68.865 185.195 ;
        RECT 70.400 185.150 70.720 185.210 ;
        RECT 71.780 185.150 72.100 185.210 ;
        RECT 67.270 185.010 72.100 185.150 ;
        RECT 30.380 184.670 37.080 184.810 ;
        RECT 37.320 184.810 37.610 184.855 ;
        RECT 39.420 184.810 39.710 184.855 ;
        RECT 40.990 184.810 41.280 184.855 ;
        RECT 37.320 184.670 41.280 184.810 ;
        RECT 30.380 184.610 30.700 184.670 ;
        RECT 23.915 184.470 24.205 184.515 ;
        RECT 25.105 184.470 25.395 184.515 ;
        RECT 27.625 184.470 27.915 184.515 ;
        RECT 23.915 184.330 27.915 184.470 ;
        RECT 23.915 184.285 24.205 184.330 ;
        RECT 25.105 184.285 25.395 184.330 ;
        RECT 27.625 184.285 27.915 184.330 ;
        RECT 28.080 184.470 28.400 184.530 ;
        RECT 33.155 184.470 33.445 184.515 ;
        RECT 34.060 184.470 34.380 184.530 ;
        RECT 35.070 184.515 35.210 184.670 ;
        RECT 37.320 184.625 37.610 184.670 ;
        RECT 39.420 184.625 39.710 184.670 ;
        RECT 40.990 184.625 41.280 184.670 ;
        RECT 48.360 184.810 48.650 184.855 ;
        RECT 50.460 184.810 50.750 184.855 ;
        RECT 52.030 184.810 52.320 184.855 ;
        RECT 48.360 184.670 52.320 184.810 ;
        RECT 48.360 184.625 48.650 184.670 ;
        RECT 50.460 184.625 50.750 184.670 ;
        RECT 52.030 184.625 52.320 184.670 ;
        RECT 57.100 184.810 57.390 184.855 ;
        RECT 59.200 184.810 59.490 184.855 ;
        RECT 60.770 184.810 61.060 184.855 ;
        RECT 57.100 184.670 61.060 184.810 ;
        RECT 57.100 184.625 57.390 184.670 ;
        RECT 59.200 184.625 59.490 184.670 ;
        RECT 60.770 184.625 61.060 184.670 ;
        RECT 35.440 184.515 35.760 184.530 ;
        RECT 28.080 184.330 34.380 184.470 ;
        RECT 28.080 184.270 28.400 184.330 ;
        RECT 33.155 184.285 33.445 184.330 ;
        RECT 34.060 184.270 34.380 184.330 ;
        RECT 34.995 184.285 35.285 184.515 ;
        RECT 35.440 184.285 35.870 184.515 ;
        RECT 37.715 184.470 38.005 184.515 ;
        RECT 38.905 184.470 39.195 184.515 ;
        RECT 41.425 184.470 41.715 184.515 ;
        RECT 37.715 184.330 41.715 184.470 ;
        RECT 37.715 184.285 38.005 184.330 ;
        RECT 38.905 184.285 39.195 184.330 ;
        RECT 41.425 184.285 41.715 184.330 ;
        RECT 48.755 184.470 49.045 184.515 ;
        RECT 49.945 184.470 50.235 184.515 ;
        RECT 52.465 184.470 52.755 184.515 ;
        RECT 48.755 184.330 52.755 184.470 ;
        RECT 48.755 184.285 49.045 184.330 ;
        RECT 49.945 184.285 50.235 184.330 ;
        RECT 52.465 184.285 52.755 184.330 ;
        RECT 57.495 184.470 57.785 184.515 ;
        RECT 58.685 184.470 58.975 184.515 ;
        RECT 61.205 184.470 61.495 184.515 ;
        RECT 57.495 184.330 61.495 184.470 ;
        RECT 57.495 184.285 57.785 184.330 ;
        RECT 58.685 184.285 58.975 184.330 ;
        RECT 61.205 184.285 61.495 184.330 ;
        RECT 65.355 184.470 65.645 184.515 ;
        RECT 66.260 184.470 66.580 184.530 ;
        RECT 65.355 184.330 66.580 184.470 ;
        RECT 65.355 184.285 65.645 184.330 ;
        RECT 35.440 184.270 35.760 184.285 ;
        RECT 66.260 184.270 66.580 184.330 ;
        RECT 21.640 184.130 21.960 184.190 ;
        RECT 23.035 184.130 23.325 184.175 ;
        RECT 36.835 184.130 37.125 184.175 ;
        RECT 21.640 183.990 23.325 184.130 ;
        RECT 21.640 183.930 21.960 183.990 ;
        RECT 23.035 183.945 23.325 183.990 ;
        RECT 35.070 183.990 37.125 184.130 ;
        RECT 35.070 183.850 35.210 183.990 ;
        RECT 36.835 183.945 37.125 183.990 ;
        RECT 38.170 184.130 38.460 184.175 ;
        RECT 39.580 184.130 39.900 184.190 ;
        RECT 38.170 183.990 39.900 184.130 ;
        RECT 38.170 183.945 38.460 183.990 ;
        RECT 39.580 183.930 39.900 183.990 ;
        RECT 47.875 184.130 48.165 184.175 ;
        RECT 53.380 184.130 53.700 184.190 ;
        RECT 56.615 184.130 56.905 184.175 ;
        RECT 47.875 183.990 56.905 184.130 ;
        RECT 47.875 183.945 48.165 183.990 ;
        RECT 53.380 183.930 53.700 183.990 ;
        RECT 56.615 183.945 56.905 183.990 ;
        RECT 65.815 184.130 66.105 184.175 ;
        RECT 67.270 184.130 67.410 185.010 ;
        RECT 68.575 184.965 68.865 185.010 ;
        RECT 70.400 184.950 70.720 185.010 ;
        RECT 71.780 184.950 72.100 185.010 ;
        RECT 72.700 184.950 73.020 185.210 ;
        RECT 74.080 185.150 74.400 185.210 ;
        RECT 78.235 185.150 78.525 185.195 ;
        RECT 80.520 185.150 80.840 185.210 ;
        RECT 74.080 185.010 80.840 185.150 ;
        RECT 74.080 184.950 74.400 185.010 ;
        RECT 78.235 184.965 78.525 185.010 ;
        RECT 80.520 184.950 80.840 185.010 ;
        RECT 80.995 185.150 81.285 185.195 ;
        RECT 81.900 185.150 82.220 185.210 ;
        RECT 80.995 185.010 82.220 185.150 ;
        RECT 80.995 184.965 81.285 185.010 ;
        RECT 81.900 184.950 82.220 185.010 ;
        RECT 95.700 185.150 96.020 185.210 ;
        RECT 105.375 185.150 105.665 185.195 ;
        RECT 95.700 185.010 100.990 185.150 ;
        RECT 95.700 184.950 96.020 185.010 ;
        RECT 69.020 184.810 69.340 184.870 ;
        RECT 69.940 184.810 70.260 184.870 ;
        RECT 68.190 184.670 70.260 184.810 ;
        RECT 68.190 184.175 68.330 184.670 ;
        RECT 69.020 184.610 69.340 184.670 ;
        RECT 69.940 184.610 70.260 184.670 ;
        RECT 72.240 184.810 72.560 184.870 ;
        RECT 73.175 184.810 73.465 184.855 ;
        RECT 72.240 184.670 73.465 184.810 ;
        RECT 72.240 184.610 72.560 184.670 ;
        RECT 73.175 184.625 73.465 184.670 ;
        RECT 74.555 184.810 74.845 184.855 ;
        RECT 85.120 184.810 85.440 184.870 ;
        RECT 74.555 184.670 85.440 184.810 ;
        RECT 74.555 184.625 74.845 184.670 ;
        RECT 85.120 184.610 85.440 184.670 ;
        RECT 86.040 184.810 86.330 184.855 ;
        RECT 87.610 184.810 87.900 184.855 ;
        RECT 89.710 184.810 90.000 184.855 ;
        RECT 86.040 184.670 90.000 184.810 ;
        RECT 86.040 184.625 86.330 184.670 ;
        RECT 87.610 184.625 87.900 184.670 ;
        RECT 89.710 184.625 90.000 184.670 ;
        RECT 94.820 184.810 95.110 184.855 ;
        RECT 96.920 184.810 97.210 184.855 ;
        RECT 98.490 184.810 98.780 184.855 ;
        RECT 94.820 184.670 98.780 184.810 ;
        RECT 94.820 184.625 95.110 184.670 ;
        RECT 96.920 184.625 97.210 184.670 ;
        RECT 98.490 184.625 98.780 184.670 ;
        RECT 68.560 184.470 68.880 184.530 ;
        RECT 69.495 184.470 69.785 184.515 ;
        RECT 77.300 184.470 77.620 184.530 ;
        RECT 80.980 184.470 81.300 184.530 ;
        RECT 68.560 184.330 69.785 184.470 ;
        RECT 68.560 184.270 68.880 184.330 ;
        RECT 69.495 184.285 69.785 184.330 ;
        RECT 74.170 184.330 77.620 184.470 ;
        RECT 65.815 183.990 67.410 184.130 ;
        RECT 65.815 183.945 66.105 183.990 ;
        RECT 68.115 183.945 68.405 184.175 ;
        RECT 69.075 184.100 69.365 184.145 ;
        RECT 72.240 184.130 72.560 184.190 ;
        RECT 73.620 184.130 73.940 184.190 ;
        RECT 74.170 184.175 74.310 184.330 ;
        RECT 77.300 184.270 77.620 184.330 ;
        RECT 78.310 184.330 81.300 184.470 ;
        RECT 69.075 183.960 69.710 184.100 ;
        RECT 24.400 183.835 24.720 183.850 ;
        RECT 24.370 183.605 24.720 183.835 ;
        RECT 24.400 183.590 24.720 183.605 ;
        RECT 34.980 183.590 35.300 183.850 ;
        RECT 37.740 183.790 38.060 183.850 ;
        RECT 35.990 183.650 38.060 183.790 ;
        RECT 24.860 183.450 25.180 183.510 ;
        RECT 34.535 183.450 34.825 183.495 ;
        RECT 35.990 183.450 36.130 183.650 ;
        RECT 37.740 183.590 38.060 183.650 ;
        RECT 46.940 183.790 47.260 183.850 ;
        RECT 49.100 183.790 49.390 183.835 ;
        RECT 46.940 183.650 49.390 183.790 ;
        RECT 46.940 183.590 47.260 183.650 ;
        RECT 49.100 183.605 49.390 183.650 ;
        RECT 55.680 183.790 56.000 183.850 ;
        RECT 57.840 183.790 58.130 183.835 ;
        RECT 55.680 183.650 58.130 183.790 ;
        RECT 55.680 183.590 56.000 183.650 ;
        RECT 57.840 183.605 58.130 183.650 ;
        RECT 67.180 183.590 67.500 183.850 ;
        RECT 67.640 183.590 67.960 183.850 ;
        RECT 24.860 183.310 36.130 183.450 ;
        RECT 24.860 183.250 25.180 183.310 ;
        RECT 34.535 183.265 34.825 183.310 ;
        RECT 36.360 183.250 36.680 183.510 ;
        RECT 43.720 183.250 44.040 183.510 ;
        RECT 45.100 183.450 45.420 183.510 ;
        RECT 54.775 183.450 55.065 183.495 ;
        RECT 57.060 183.450 57.380 183.510 ;
        RECT 45.100 183.310 57.380 183.450 ;
        RECT 45.100 183.250 45.420 183.310 ;
        RECT 54.775 183.265 55.065 183.310 ;
        RECT 57.060 183.250 57.380 183.310 ;
        RECT 63.515 183.450 63.805 183.495 ;
        RECT 68.190 183.450 68.330 183.945 ;
        RECT 69.075 183.915 69.365 183.960 ;
        RECT 63.515 183.310 68.330 183.450 ;
        RECT 69.570 183.450 69.710 183.960 ;
        RECT 72.240 183.990 73.940 184.130 ;
        RECT 72.240 183.930 72.560 183.990 ;
        RECT 73.620 183.930 73.940 183.990 ;
        RECT 74.095 183.945 74.385 184.175 ;
        RECT 74.540 184.130 74.860 184.190 ;
        RECT 75.015 184.130 75.305 184.175 ;
        RECT 74.540 183.990 75.305 184.130 ;
        RECT 74.540 183.930 74.860 183.990 ;
        RECT 75.015 183.945 75.305 183.990 ;
        RECT 75.460 183.930 75.780 184.190 ;
        RECT 76.395 184.130 76.685 184.175 ;
        RECT 76.840 184.130 77.160 184.190 ;
        RECT 78.310 184.175 78.450 184.330 ;
        RECT 80.980 184.270 81.300 184.330 ;
        RECT 85.605 184.470 85.895 184.515 ;
        RECT 88.125 184.470 88.415 184.515 ;
        RECT 89.315 184.470 89.605 184.515 ;
        RECT 94.320 184.470 94.640 184.530 ;
        RECT 85.605 184.330 89.605 184.470 ;
        RECT 85.605 184.285 85.895 184.330 ;
        RECT 88.125 184.285 88.415 184.330 ;
        RECT 89.315 184.285 89.605 184.330 ;
        RECT 90.270 184.330 94.640 184.470 ;
        RECT 90.270 184.190 90.410 184.330 ;
        RECT 94.320 184.270 94.640 184.330 ;
        RECT 95.215 184.470 95.505 184.515 ;
        RECT 96.405 184.470 96.695 184.515 ;
        RECT 98.925 184.470 99.215 184.515 ;
        RECT 95.215 184.330 99.215 184.470 ;
        RECT 100.850 184.470 100.990 185.010 ;
        RECT 104.530 185.010 105.665 185.150 ;
        RECT 104.530 184.515 104.670 185.010 ;
        RECT 105.375 184.965 105.665 185.010 ;
        RECT 107.660 185.150 107.980 185.210 ;
        RECT 108.135 185.150 108.425 185.195 ;
        RECT 107.660 185.010 108.425 185.150 ;
        RECT 107.660 184.950 107.980 185.010 ;
        RECT 108.135 184.965 108.425 185.010 ;
        RECT 109.960 185.150 110.280 185.210 ;
        RECT 109.960 185.010 113.870 185.150 ;
        RECT 109.960 184.950 110.280 185.010 ;
        RECT 110.420 184.810 110.740 184.870 ;
        RECT 111.815 184.810 112.105 184.855 ;
        RECT 110.420 184.670 112.105 184.810 ;
        RECT 113.730 184.810 113.870 185.010 ;
        RECT 117.320 184.950 117.640 185.210 ;
        RECT 119.620 185.150 119.940 185.210 ;
        RECT 117.870 185.010 119.940 185.150 ;
        RECT 117.870 184.810 118.010 185.010 ;
        RECT 119.620 184.950 119.940 185.010 ;
        RECT 113.730 184.670 118.010 184.810 ;
        RECT 118.240 184.810 118.560 184.870 ;
        RECT 122.840 184.810 123.160 184.870 ;
        RECT 140.335 184.810 140.625 184.855 ;
        RECT 118.240 184.670 122.610 184.810 ;
        RECT 110.420 184.610 110.740 184.670 ;
        RECT 111.815 184.625 112.105 184.670 ;
        RECT 118.240 184.610 118.560 184.670 ;
        RECT 104.455 184.470 104.745 184.515 ;
        RECT 105.835 184.470 106.125 184.515 ;
        RECT 107.660 184.470 107.980 184.530 ;
        RECT 114.560 184.470 114.880 184.530 ;
        RECT 116.860 184.470 117.180 184.530 ;
        RECT 120.555 184.470 120.845 184.515 ;
        RECT 100.850 184.330 104.745 184.470 ;
        RECT 95.215 184.285 95.505 184.330 ;
        RECT 96.405 184.285 96.695 184.330 ;
        RECT 98.925 184.285 99.215 184.330 ;
        RECT 104.455 184.285 104.745 184.330 ;
        RECT 104.990 184.330 107.980 184.470 ;
        RECT 76.395 183.990 77.160 184.130 ;
        RECT 76.395 183.945 76.685 183.990 ;
        RECT 76.840 183.930 77.160 183.990 ;
        RECT 78.235 183.945 78.525 184.175 ;
        RECT 78.680 183.930 79.000 184.190 ;
        RECT 80.520 183.930 80.840 184.190 ;
        RECT 81.455 183.945 81.745 184.175 ;
        RECT 88.915 184.130 89.205 184.175 ;
        RECT 89.720 184.130 90.040 184.190 ;
        RECT 88.915 183.990 90.040 184.130 ;
        RECT 88.915 183.945 89.205 183.990 ;
        RECT 77.760 183.790 78.080 183.850 ;
        RECT 81.530 183.790 81.670 183.945 ;
        RECT 89.720 183.930 90.040 183.990 ;
        RECT 90.180 183.930 90.500 184.190 ;
        RECT 90.655 183.945 90.945 184.175 ;
        RECT 94.780 184.130 95.100 184.190 ;
        RECT 95.615 184.130 95.905 184.175 ;
        RECT 94.780 183.990 95.905 184.130 ;
        RECT 77.760 183.650 81.670 183.790 ;
        RECT 77.760 183.590 78.080 183.650 ;
        RECT 78.680 183.450 79.000 183.510 ;
        RECT 69.570 183.310 79.000 183.450 ;
        RECT 63.515 183.265 63.805 183.310 ;
        RECT 78.680 183.250 79.000 183.310 ;
        RECT 80.075 183.450 80.365 183.495 ;
        RECT 80.520 183.450 80.840 183.510 ;
        RECT 80.075 183.310 80.840 183.450 ;
        RECT 80.075 183.265 80.365 183.310 ;
        RECT 80.520 183.250 80.840 183.310 ;
        RECT 83.295 183.450 83.585 183.495 ;
        RECT 84.660 183.450 84.980 183.510 ;
        RECT 90.730 183.450 90.870 183.945 ;
        RECT 94.780 183.930 95.100 183.990 ;
        RECT 95.615 183.945 95.905 183.990 ;
        RECT 100.760 184.130 101.080 184.190 ;
        RECT 104.990 184.130 105.130 184.330 ;
        RECT 105.835 184.285 106.125 184.330 ;
        RECT 107.660 184.270 107.980 184.330 ;
        RECT 110.510 184.330 114.880 184.470 ;
        RECT 100.760 183.990 105.130 184.130 ;
        RECT 105.375 184.130 105.665 184.175 ;
        RECT 106.740 184.130 107.060 184.190 ;
        RECT 105.375 183.990 107.060 184.130 ;
        RECT 100.760 183.930 101.080 183.990 ;
        RECT 105.375 183.945 105.665 183.990 ;
        RECT 106.740 183.930 107.060 183.990 ;
        RECT 109.040 183.930 109.360 184.190 ;
        RECT 110.510 184.175 110.650 184.330 ;
        RECT 114.560 184.270 114.880 184.330 ;
        RECT 116.490 184.330 120.845 184.470 ;
        RECT 109.515 183.945 109.805 184.175 ;
        RECT 110.435 183.945 110.725 184.175 ;
        RECT 104.900 183.790 105.220 183.850 ;
        RECT 101.310 183.650 105.220 183.790 ;
        RECT 83.295 183.310 90.870 183.450 ;
        RECT 92.020 183.450 92.340 183.510 ;
        RECT 93.875 183.450 94.165 183.495 ;
        RECT 92.020 183.310 94.165 183.450 ;
        RECT 83.295 183.265 83.585 183.310 ;
        RECT 84.660 183.250 84.980 183.310 ;
        RECT 92.020 183.250 92.340 183.310 ;
        RECT 93.875 183.265 94.165 183.310 ;
        RECT 97.080 183.450 97.400 183.510 ;
        RECT 101.310 183.495 101.450 183.650 ;
        RECT 104.900 183.590 105.220 183.650 ;
        RECT 101.235 183.450 101.525 183.495 ;
        RECT 97.080 183.310 101.525 183.450 ;
        RECT 97.080 183.250 97.400 183.310 ;
        RECT 101.235 183.265 101.525 183.310 ;
        RECT 101.680 183.250 102.000 183.510 ;
        RECT 107.200 183.250 107.520 183.510 ;
        RECT 109.130 183.450 109.270 183.930 ;
        RECT 109.590 183.790 109.730 183.945 ;
        RECT 110.880 183.930 111.200 184.190 ;
        RECT 111.815 183.945 112.105 184.175 ;
        RECT 112.720 184.130 113.040 184.190 ;
        RECT 116.490 184.175 116.630 184.330 ;
        RECT 116.860 184.270 117.180 184.330 ;
        RECT 120.555 184.285 120.845 184.330 ;
        RECT 114.115 184.130 114.405 184.175 ;
        RECT 112.720 183.990 114.405 184.130 ;
        RECT 111.890 183.790 112.030 183.945 ;
        RECT 112.720 183.930 113.040 183.990 ;
        RECT 114.115 183.945 114.405 183.990 ;
        RECT 116.415 183.945 116.705 184.175 ;
        RECT 117.780 183.930 118.100 184.190 ;
        RECT 118.240 184.130 118.560 184.190 ;
        RECT 119.635 184.130 119.925 184.175 ;
        RECT 118.240 183.990 119.925 184.130 ;
        RECT 118.240 183.930 118.560 183.990 ;
        RECT 119.635 183.945 119.925 183.990 ;
        RECT 120.080 183.930 120.400 184.190 ;
        RECT 121.000 183.930 121.320 184.190 ;
        RECT 122.470 184.175 122.610 184.670 ;
        RECT 122.840 184.670 140.625 184.810 ;
        RECT 122.840 184.610 123.160 184.670 ;
        RECT 140.335 184.625 140.625 184.670 ;
        RECT 121.475 183.945 121.765 184.175 ;
        RECT 122.395 183.945 122.685 184.175 ;
        RECT 113.180 183.790 113.500 183.850 ;
        RECT 115.020 183.835 115.340 183.850 ;
        RECT 114.805 183.790 115.340 183.835 ;
        RECT 109.590 183.650 113.500 183.790 ;
        RECT 113.180 183.590 113.500 183.650 ;
        RECT 113.730 183.650 115.340 183.790 ;
        RECT 113.730 183.450 113.870 183.650 ;
        RECT 114.805 183.605 115.340 183.650 ;
        RECT 115.495 183.605 115.785 183.835 ;
        RECT 115.020 183.590 115.340 183.605 ;
        RECT 109.130 183.310 113.870 183.450 ;
        RECT 115.570 183.450 115.710 183.605 ;
        RECT 115.940 183.590 116.260 183.850 ;
        RECT 117.870 183.790 118.010 183.930 ;
        RECT 118.715 183.790 119.005 183.835 ;
        RECT 117.870 183.650 119.005 183.790 ;
        RECT 118.715 183.605 119.005 183.650 ;
        RECT 120.540 183.790 120.860 183.850 ;
        RECT 121.550 183.790 121.690 183.945 ;
        RECT 138.020 183.930 138.340 184.190 ;
        RECT 141.240 183.930 141.560 184.190 ;
        RECT 120.540 183.650 121.690 183.790 ;
        RECT 120.540 183.590 120.860 183.650 ;
        RECT 117.780 183.450 118.100 183.510 ;
        RECT 115.570 183.310 118.100 183.450 ;
        RECT 117.780 183.250 118.100 183.310 ;
        RECT 121.460 183.250 121.780 183.510 ;
        RECT 138.955 183.450 139.245 183.495 ;
        RECT 139.860 183.450 140.180 183.510 ;
        RECT 138.955 183.310 140.180 183.450 ;
        RECT 138.955 183.265 139.245 183.310 ;
        RECT 139.860 183.250 140.180 183.310 ;
        RECT 17.430 182.630 143.010 183.110 ;
        RECT 24.400 182.230 24.720 182.490 ;
        RECT 24.860 182.430 25.180 182.490 ;
        RECT 26.255 182.430 26.545 182.475 ;
        RECT 36.820 182.430 37.140 182.490 ;
        RECT 24.860 182.290 26.545 182.430 ;
        RECT 24.860 182.230 25.180 182.290 ;
        RECT 26.255 182.245 26.545 182.290 ;
        RECT 32.770 182.290 37.140 182.430 ;
        RECT 32.770 182.135 32.910 182.290 ;
        RECT 36.820 182.230 37.140 182.290 ;
        RECT 38.200 182.430 38.520 182.490 ;
        RECT 38.200 182.290 45.790 182.430 ;
        RECT 38.200 182.230 38.520 182.290 ;
        RECT 32.695 181.905 32.985 182.135 ;
        RECT 33.695 182.090 33.985 182.135 ;
        RECT 33.230 181.950 33.985 182.090 ;
        RECT 25.210 181.750 25.500 181.795 ;
        RECT 25.210 181.610 28.310 181.750 ;
        RECT 25.210 181.565 25.500 181.610 ;
        RECT 25.780 181.210 26.100 181.470 ;
        RECT 27.620 181.210 27.940 181.470 ;
        RECT 28.170 181.455 28.310 181.610 ;
        RECT 29.920 181.550 30.240 181.810 ;
        RECT 33.230 181.750 33.370 181.950 ;
        RECT 33.695 181.905 33.985 181.950 ;
        RECT 35.900 181.890 36.220 182.150 ;
        RECT 45.100 182.090 45.420 182.150 ;
        RECT 44.730 181.950 45.420 182.090 ;
        RECT 45.650 182.090 45.790 182.290 ;
        RECT 46.940 182.230 47.260 182.490 ;
        RECT 69.940 182.430 70.260 182.490 ;
        RECT 77.760 182.430 78.080 182.490 ;
        RECT 47.490 182.290 54.990 182.430 ;
        RECT 47.490 182.090 47.630 182.290 ;
        RECT 45.650 181.950 47.630 182.090 ;
        RECT 48.335 182.090 48.625 182.135 ;
        RECT 51.540 182.090 51.860 182.150 ;
        RECT 48.335 181.950 51.860 182.090 ;
        RECT 30.930 181.610 33.370 181.750 ;
        RECT 35.990 181.740 36.130 181.890 ;
        RECT 44.730 181.795 44.870 181.950 ;
        RECT 45.100 181.890 45.420 181.950 ;
        RECT 48.335 181.905 48.625 181.950 ;
        RECT 51.540 181.890 51.860 181.950 ;
        RECT 54.850 181.810 54.990 182.290 ;
        RECT 69.940 182.290 78.080 182.430 ;
        RECT 69.940 182.230 70.260 182.290 ;
        RECT 77.760 182.230 78.080 182.290 ;
        RECT 85.580 182.430 85.900 182.490 ;
        RECT 86.515 182.430 86.805 182.475 ;
        RECT 85.580 182.290 86.805 182.430 ;
        RECT 85.580 182.230 85.900 182.290 ;
        RECT 86.515 182.245 86.805 182.290 ;
        RECT 90.655 182.430 90.945 182.475 ;
        RECT 92.940 182.430 93.260 182.490 ;
        RECT 101.235 182.430 101.525 182.475 ;
        RECT 90.655 182.290 93.260 182.430 ;
        RECT 90.655 182.245 90.945 182.290 ;
        RECT 92.940 182.230 93.260 182.290 ;
        RECT 97.630 182.290 101.525 182.430 ;
        RECT 55.220 182.090 55.540 182.150 ;
        RECT 55.695 182.090 55.985 182.135 ;
        RECT 55.220 181.950 55.985 182.090 ;
        RECT 55.220 181.890 55.540 181.950 ;
        RECT 55.695 181.905 55.985 181.950 ;
        RECT 72.715 182.090 73.005 182.135 ;
        RECT 74.080 182.090 74.400 182.150 ;
        RECT 72.715 181.950 74.400 182.090 ;
        RECT 72.715 181.905 73.005 181.950 ;
        RECT 74.080 181.890 74.400 181.950 ;
        RECT 80.950 182.090 81.240 182.135 ;
        RECT 81.440 182.090 81.760 182.150 ;
        RECT 97.630 182.135 97.770 182.290 ;
        RECT 101.235 182.245 101.525 182.290 ;
        RECT 102.140 182.430 102.460 182.490 ;
        RECT 102.615 182.430 102.905 182.475 ;
        RECT 115.165 182.430 115.455 182.475 ;
        RECT 115.940 182.430 116.260 182.490 ;
        RECT 118.255 182.430 118.545 182.475 ;
        RECT 121.460 182.430 121.780 182.490 ;
        RECT 102.140 182.290 102.905 182.430 ;
        RECT 102.140 182.230 102.460 182.290 ;
        RECT 102.615 182.245 102.905 182.290 ;
        RECT 109.590 182.290 112.950 182.430 ;
        RECT 98.000 182.135 98.320 182.150 ;
        RECT 97.555 182.090 97.845 182.135 ;
        RECT 80.950 181.950 81.760 182.090 ;
        RECT 80.950 181.905 81.240 181.950 ;
        RECT 81.440 181.890 81.760 181.950 ;
        RECT 93.030 181.950 97.845 182.090 ;
        RECT 36.330 181.740 36.620 181.795 ;
        RECT 30.930 181.470 31.070 181.610 ;
        RECT 35.990 181.600 36.620 181.740 ;
        RECT 36.330 181.565 36.620 181.600 ;
        RECT 44.655 181.565 44.945 181.795 ;
        RECT 48.795 181.750 49.085 181.795 ;
        RECT 51.080 181.750 51.400 181.810 ;
        RECT 48.795 181.610 51.400 181.750 ;
        RECT 48.795 181.565 49.085 181.610 ;
        RECT 51.080 181.550 51.400 181.610 ;
        RECT 54.300 181.550 54.620 181.810 ;
        RECT 54.760 181.550 55.080 181.810 ;
        RECT 68.575 181.565 68.865 181.795 ;
        RECT 71.335 181.565 71.625 181.795 ;
        RECT 28.095 181.225 28.385 181.455 ;
        RECT 30.395 181.410 30.685 181.455 ;
        RECT 30.840 181.410 31.160 181.470 ;
        RECT 30.395 181.270 31.160 181.410 ;
        RECT 30.395 181.225 30.685 181.270 ;
        RECT 30.840 181.210 31.160 181.270 ;
        RECT 34.980 181.210 35.300 181.470 ;
        RECT 35.875 181.410 36.165 181.455 ;
        RECT 37.065 181.410 37.355 181.455 ;
        RECT 39.585 181.410 39.875 181.455 ;
        RECT 35.875 181.270 39.875 181.410 ;
        RECT 35.875 181.225 36.165 181.270 ;
        RECT 37.065 181.225 37.355 181.270 ;
        RECT 39.585 181.225 39.875 181.270 ;
        RECT 45.115 181.410 45.405 181.455 ;
        RECT 46.020 181.410 46.340 181.470 ;
        RECT 45.115 181.270 46.340 181.410 ;
        RECT 45.115 181.225 45.405 181.270 ;
        RECT 46.020 181.210 46.340 181.270 ;
        RECT 46.495 181.410 46.785 181.455 ;
        RECT 47.750 181.410 48.040 181.455 ;
        RECT 46.495 181.270 48.040 181.410 ;
        RECT 46.495 181.225 46.785 181.270 ;
        RECT 47.750 181.225 48.040 181.270 ;
        RECT 50.175 181.410 50.465 181.455 ;
        RECT 50.620 181.410 50.940 181.470 ;
        RECT 67.180 181.410 67.500 181.470 ;
        RECT 50.175 181.270 67.500 181.410 ;
        RECT 50.175 181.225 50.465 181.270 ;
        RECT 50.620 181.210 50.940 181.270 ;
        RECT 67.180 181.210 67.500 181.270 ;
        RECT 21.640 181.070 21.960 181.130 ;
        RECT 35.070 181.070 35.210 181.210 ;
        RECT 21.640 180.930 35.210 181.070 ;
        RECT 35.480 181.070 35.770 181.115 ;
        RECT 37.580 181.070 37.870 181.115 ;
        RECT 39.150 181.070 39.440 181.115 ;
        RECT 35.480 180.930 39.440 181.070 ;
        RECT 21.640 180.870 21.960 180.930 ;
        RECT 35.480 180.885 35.770 180.930 ;
        RECT 37.580 180.885 37.870 180.930 ;
        RECT 39.150 180.885 39.440 180.930 ;
        RECT 55.680 180.870 56.000 181.130 ;
        RECT 68.650 181.070 68.790 181.565 ;
        RECT 69.020 181.410 69.340 181.470 ;
        RECT 70.875 181.410 71.165 181.455 ;
        RECT 69.020 181.270 71.165 181.410 ;
        RECT 71.410 181.410 71.550 181.565 ;
        RECT 71.780 181.550 72.100 181.810 ;
        RECT 92.020 181.550 92.340 181.810 ;
        RECT 92.480 181.550 92.800 181.810 ;
        RECT 93.030 181.795 93.170 181.950 ;
        RECT 97.555 181.905 97.845 181.950 ;
        RECT 98.000 181.905 98.430 182.135 ;
        RECT 101.680 182.090 102.000 182.150 ;
        RECT 103.995 182.090 104.285 182.135 ;
        RECT 101.680 181.950 104.285 182.090 ;
        RECT 98.000 181.890 98.320 181.905 ;
        RECT 101.680 181.890 102.000 181.950 ;
        RECT 103.995 181.905 104.285 181.950 ;
        RECT 104.900 182.090 105.220 182.150 ;
        RECT 109.590 182.090 109.730 182.290 ;
        RECT 104.900 181.950 109.730 182.090 ;
        RECT 104.900 181.890 105.220 181.950 ;
        RECT 92.955 181.565 93.245 181.795 ;
        RECT 93.875 181.750 94.165 181.795 ;
        RECT 103.520 181.750 103.840 181.810 ;
        RECT 93.875 181.610 95.470 181.750 ;
        RECT 93.875 181.565 94.165 181.610 ;
        RECT 72.240 181.410 72.560 181.470 ;
        RECT 79.615 181.410 79.905 181.455 ;
        RECT 71.410 181.270 72.010 181.410 ;
        RECT 69.020 181.210 69.340 181.270 ;
        RECT 70.875 181.225 71.165 181.270 ;
        RECT 69.495 181.070 69.785 181.115 ;
        RECT 68.650 180.930 69.785 181.070 ;
        RECT 71.870 181.070 72.010 181.270 ;
        RECT 72.240 181.270 79.905 181.410 ;
        RECT 72.240 181.210 72.560 181.270 ;
        RECT 79.615 181.225 79.905 181.270 ;
        RECT 80.495 181.410 80.785 181.455 ;
        RECT 81.685 181.410 81.975 181.455 ;
        RECT 84.205 181.410 84.495 181.455 ;
        RECT 80.495 181.270 84.495 181.410 ;
        RECT 80.495 181.225 80.785 181.270 ;
        RECT 81.685 181.225 81.975 181.270 ;
        RECT 84.205 181.225 84.495 181.270 ;
        RECT 89.720 181.410 90.040 181.470 ;
        RECT 93.030 181.410 93.170 181.565 ;
        RECT 95.330 181.470 95.470 181.610 ;
        RECT 99.010 181.610 103.840 181.750 ;
        RECT 89.720 181.270 93.170 181.410 ;
        RECT 95.240 181.410 95.560 181.470 ;
        RECT 95.715 181.410 96.005 181.455 ;
        RECT 95.240 181.270 96.005 181.410 ;
        RECT 89.720 181.210 90.040 181.270 ;
        RECT 95.240 181.210 95.560 181.270 ;
        RECT 95.715 181.225 96.005 181.270 ;
        RECT 73.160 181.070 73.480 181.130 ;
        RECT 71.870 180.930 73.480 181.070 ;
        RECT 69.495 180.885 69.785 180.930 ;
        RECT 73.160 180.870 73.480 180.930 ;
        RECT 80.100 181.070 80.390 181.115 ;
        RECT 82.200 181.070 82.490 181.115 ;
        RECT 83.770 181.070 84.060 181.115 ;
        RECT 80.100 180.930 84.060 181.070 ;
        RECT 80.100 180.885 80.390 180.930 ;
        RECT 82.200 180.885 82.490 180.930 ;
        RECT 83.770 180.885 84.060 180.930 ;
        RECT 29.920 180.730 30.240 180.790 ;
        RECT 33.615 180.730 33.905 180.775 ;
        RECT 29.920 180.590 33.905 180.730 ;
        RECT 29.920 180.530 30.240 180.590 ;
        RECT 33.615 180.545 33.905 180.590 ;
        RECT 34.535 180.730 34.825 180.775 ;
        RECT 34.980 180.730 35.300 180.790 ;
        RECT 34.535 180.590 35.300 180.730 ;
        RECT 34.535 180.545 34.825 180.590 ;
        RECT 34.980 180.530 35.300 180.590 ;
        RECT 36.360 180.730 36.680 180.790 ;
        RECT 38.660 180.730 38.980 180.790 ;
        RECT 41.895 180.730 42.185 180.775 ;
        RECT 36.360 180.590 42.185 180.730 ;
        RECT 36.360 180.530 36.680 180.590 ;
        RECT 38.660 180.530 38.980 180.590 ;
        RECT 41.895 180.545 42.185 180.590 ;
        RECT 68.115 180.730 68.405 180.775 ;
        RECT 70.400 180.730 70.720 180.790 ;
        RECT 68.115 180.590 70.720 180.730 ;
        RECT 68.115 180.545 68.405 180.590 ;
        RECT 70.400 180.530 70.720 180.590 ;
        RECT 71.320 180.530 71.640 180.790 ;
        RECT 71.780 180.730 72.100 180.790 ;
        RECT 73.635 180.730 73.925 180.775 ;
        RECT 71.780 180.590 73.925 180.730 ;
        RECT 71.780 180.530 72.100 180.590 ;
        RECT 73.635 180.545 73.925 180.590 ;
        RECT 80.980 180.730 81.300 180.790 ;
        RECT 89.260 180.730 89.580 180.790 ;
        RECT 80.980 180.590 89.580 180.730 ;
        RECT 95.790 180.730 95.930 181.225 ;
        RECT 97.080 181.210 97.400 181.470 ;
        RECT 99.010 181.115 99.150 181.610 ;
        RECT 103.520 181.550 103.840 181.610 ;
        RECT 104.455 181.565 104.745 181.795 ;
        RECT 99.840 181.410 100.160 181.470 ;
        RECT 104.530 181.410 104.670 181.565 ;
        RECT 105.360 181.550 105.680 181.810 ;
        RECT 106.740 181.550 107.060 181.810 ;
        RECT 107.660 181.750 107.980 181.810 ;
        RECT 108.135 181.750 108.425 181.795 ;
        RECT 107.660 181.610 108.425 181.750 ;
        RECT 107.660 181.550 107.980 181.610 ;
        RECT 108.135 181.565 108.425 181.610 ;
        RECT 108.580 181.550 108.900 181.810 ;
        RECT 109.590 181.795 109.730 181.950 ;
        RECT 109.960 182.090 110.280 182.150 ;
        RECT 112.810 182.135 112.950 182.290 ;
        RECT 115.165 182.290 121.780 182.430 ;
        RECT 115.165 182.245 115.455 182.290 ;
        RECT 115.940 182.230 116.260 182.290 ;
        RECT 118.255 182.245 118.545 182.290 ;
        RECT 121.460 182.230 121.780 182.290 ;
        RECT 135.735 182.245 136.025 182.475 ;
        RECT 110.435 182.090 110.725 182.135 ;
        RECT 109.960 181.950 110.725 182.090 ;
        RECT 109.960 181.890 110.280 181.950 ;
        RECT 110.435 181.905 110.725 181.950 ;
        RECT 111.585 181.920 111.875 181.965 ;
        RECT 109.515 181.565 109.805 181.795 ;
        RECT 111.585 181.750 111.950 181.920 ;
        RECT 112.735 181.905 113.025 182.135 ;
        RECT 113.640 182.090 113.960 182.150 ;
        RECT 114.115 182.090 114.405 182.135 ;
        RECT 113.640 181.950 114.405 182.090 ;
        RECT 113.640 181.890 113.960 181.950 ;
        RECT 114.115 181.905 114.405 181.950 ;
        RECT 115.940 181.750 116.260 181.810 ;
        RECT 111.585 181.735 116.260 181.750 ;
        RECT 111.810 181.610 116.260 181.735 ;
        RECT 115.940 181.550 116.260 181.610 ;
        RECT 128.835 181.750 129.125 181.795 ;
        RECT 129.280 181.750 129.600 181.810 ;
        RECT 128.835 181.610 129.600 181.750 ;
        RECT 128.835 181.565 129.125 181.610 ;
        RECT 129.280 181.550 129.600 181.610 ;
        RECT 130.170 181.750 130.460 181.795 ;
        RECT 133.880 181.750 134.200 181.810 ;
        RECT 130.170 181.610 134.200 181.750 ;
        RECT 135.810 181.750 135.950 182.245 ;
        RECT 138.020 181.750 138.340 181.810 ;
        RECT 138.955 181.750 139.245 181.795 ;
        RECT 135.810 181.610 139.245 181.750 ;
        RECT 130.170 181.565 130.460 181.610 ;
        RECT 133.880 181.550 134.200 181.610 ;
        RECT 138.020 181.550 138.340 181.610 ;
        RECT 138.955 181.565 139.245 181.610 ;
        RECT 139.860 181.550 140.180 181.810 ;
        RECT 99.840 181.270 104.670 181.410 ;
        RECT 99.840 181.210 100.160 181.270 ;
        RECT 98.935 180.885 99.225 181.115 ;
        RECT 99.395 180.885 99.685 181.115 ;
        RECT 100.300 181.070 100.620 181.130 ;
        RECT 105.835 181.070 106.125 181.115 ;
        RECT 108.670 181.070 108.810 181.550 ;
        RECT 109.040 181.410 109.360 181.470 ;
        RECT 120.080 181.410 120.400 181.470 ;
        RECT 109.040 181.270 120.400 181.410 ;
        RECT 109.040 181.210 109.360 181.270 ;
        RECT 120.080 181.210 120.400 181.270 ;
        RECT 129.715 181.410 130.005 181.455 ;
        RECT 130.905 181.410 131.195 181.455 ;
        RECT 133.425 181.410 133.715 181.455 ;
        RECT 129.715 181.270 133.715 181.410 ;
        RECT 129.715 181.225 130.005 181.270 ;
        RECT 130.905 181.225 131.195 181.270 ;
        RECT 133.425 181.225 133.715 181.270 ;
        RECT 135.720 181.410 136.040 181.470 ;
        RECT 136.195 181.410 136.485 181.455 ;
        RECT 135.720 181.270 136.485 181.410 ;
        RECT 135.720 181.210 136.040 181.270 ;
        RECT 136.195 181.225 136.485 181.270 ;
        RECT 113.640 181.070 113.960 181.130 ;
        RECT 116.415 181.070 116.705 181.115 ;
        RECT 117.320 181.070 117.640 181.130 ;
        RECT 100.300 180.930 106.125 181.070 ;
        RECT 99.470 180.730 99.610 180.885 ;
        RECT 100.300 180.870 100.620 180.930 ;
        RECT 105.835 180.885 106.125 180.930 ;
        RECT 107.290 180.930 112.030 181.070 ;
        RECT 95.790 180.590 99.610 180.730 ;
        RECT 80.980 180.530 81.300 180.590 ;
        RECT 89.260 180.530 89.580 180.590 ;
        RECT 101.220 180.530 101.540 180.790 ;
        RECT 102.155 180.730 102.445 180.775 ;
        RECT 107.290 180.730 107.430 180.930 ;
        RECT 111.890 180.790 112.030 180.930 ;
        RECT 113.640 180.930 117.640 181.070 ;
        RECT 113.640 180.870 113.960 180.930 ;
        RECT 116.415 180.885 116.705 180.930 ;
        RECT 117.320 180.870 117.640 180.930 ;
        RECT 129.320 181.070 129.610 181.115 ;
        RECT 131.420 181.070 131.710 181.115 ;
        RECT 132.990 181.070 133.280 181.115 ;
        RECT 129.320 180.930 133.280 181.070 ;
        RECT 129.320 180.885 129.610 180.930 ;
        RECT 131.420 180.885 131.710 180.930 ;
        RECT 132.990 180.885 133.280 180.930 ;
        RECT 102.155 180.590 107.430 180.730 ;
        RECT 102.155 180.545 102.445 180.590 ;
        RECT 107.660 180.530 107.980 180.790 ;
        RECT 109.500 180.730 109.820 180.790 ;
        RECT 110.880 180.730 111.200 180.790 ;
        RECT 109.500 180.590 111.200 180.730 ;
        RECT 109.500 180.530 109.820 180.590 ;
        RECT 110.880 180.530 111.200 180.590 ;
        RECT 111.800 180.530 112.120 180.790 ;
        RECT 115.035 180.730 115.325 180.775 ;
        RECT 115.480 180.730 115.800 180.790 ;
        RECT 115.035 180.590 115.800 180.730 ;
        RECT 115.035 180.545 115.325 180.590 ;
        RECT 115.480 180.530 115.800 180.590 ;
        RECT 115.955 180.730 116.245 180.775 ;
        RECT 116.860 180.730 117.180 180.790 ;
        RECT 115.955 180.590 117.180 180.730 ;
        RECT 115.955 180.545 116.245 180.590 ;
        RECT 116.860 180.530 117.180 180.590 ;
        RECT 117.780 180.730 118.100 180.790 ;
        RECT 118.255 180.730 118.545 180.775 ;
        RECT 118.700 180.730 119.020 180.790 ;
        RECT 117.780 180.590 119.020 180.730 ;
        RECT 117.780 180.530 118.100 180.590 ;
        RECT 118.255 180.545 118.545 180.590 ;
        RECT 118.700 180.530 119.020 180.590 ;
        RECT 119.160 180.530 119.480 180.790 ;
        RECT 140.780 180.530 141.100 180.790 ;
        RECT 17.430 179.910 143.010 180.390 ;
        RECT 29.920 179.710 30.240 179.770 ;
        RECT 34.520 179.710 34.840 179.770 ;
        RECT 29.920 179.570 34.840 179.710 ;
        RECT 29.920 179.510 30.240 179.570 ;
        RECT 34.520 179.510 34.840 179.570 ;
        RECT 35.440 179.710 35.760 179.770 ;
        RECT 35.915 179.710 36.205 179.755 ;
        RECT 35.440 179.570 36.205 179.710 ;
        RECT 35.440 179.510 35.760 179.570 ;
        RECT 35.915 179.525 36.205 179.570 ;
        RECT 39.120 179.710 39.440 179.770 ;
        RECT 99.855 179.710 100.145 179.755 ;
        RECT 101.220 179.710 101.540 179.770 ;
        RECT 39.120 179.570 49.930 179.710 ;
        RECT 39.120 179.510 39.440 179.570 ;
        RECT 25.780 179.370 26.100 179.430 ;
        RECT 30.380 179.370 30.700 179.430 ;
        RECT 25.780 179.230 30.700 179.370 ;
        RECT 25.780 179.170 26.100 179.230 ;
        RECT 30.380 179.170 30.700 179.230 ;
        RECT 30.840 179.370 31.160 179.430 ;
        RECT 37.740 179.370 38.060 179.430 ;
        RECT 30.840 179.230 38.060 179.370 ;
        RECT 30.840 179.170 31.160 179.230 ;
        RECT 37.740 179.170 38.060 179.230 ;
        RECT 38.215 179.370 38.505 179.415 ;
        RECT 43.720 179.370 44.040 179.430 ;
        RECT 38.215 179.230 44.040 179.370 ;
        RECT 38.215 179.185 38.505 179.230 ;
        RECT 43.720 179.170 44.040 179.230 ;
        RECT 49.790 179.370 49.930 179.570 ;
        RECT 99.855 179.570 101.540 179.710 ;
        RECT 99.855 179.525 100.145 179.570 ;
        RECT 101.220 179.510 101.540 179.570 ;
        RECT 101.695 179.710 101.985 179.755 ;
        RECT 106.740 179.710 107.060 179.770 ;
        RECT 101.695 179.570 107.060 179.710 ;
        RECT 101.695 179.525 101.985 179.570 ;
        RECT 106.740 179.510 107.060 179.570 ;
        RECT 108.580 179.710 108.900 179.770 ;
        RECT 109.960 179.710 110.280 179.770 ;
        RECT 108.580 179.570 110.280 179.710 ;
        RECT 108.580 179.510 108.900 179.570 ;
        RECT 109.960 179.510 110.280 179.570 ;
        RECT 112.275 179.710 112.565 179.755 ;
        RECT 112.720 179.710 113.040 179.770 ;
        RECT 118.700 179.710 119.020 179.770 ;
        RECT 112.275 179.570 115.250 179.710 ;
        RECT 112.275 179.525 112.565 179.570 ;
        RECT 112.720 179.510 113.040 179.570 ;
        RECT 55.220 179.370 55.540 179.430 ;
        RECT 73.160 179.370 73.480 179.430 ;
        RECT 94.335 179.370 94.625 179.415 ;
        RECT 98.015 179.370 98.305 179.415 ;
        RECT 49.790 179.230 55.540 179.370 ;
        RECT 24.400 178.830 24.720 179.090 ;
        RECT 25.870 179.030 26.010 179.170 ;
        RECT 24.950 178.890 26.010 179.030 ;
        RECT 35.530 178.890 40.730 179.030 ;
        RECT 23.940 178.690 24.260 178.750 ;
        RECT 24.950 178.690 25.090 178.890 ;
        RECT 23.940 178.550 25.090 178.690 ;
        RECT 25.320 178.690 25.640 178.750 ;
        RECT 25.795 178.690 26.085 178.735 ;
        RECT 27.620 178.690 27.940 178.750 ;
        RECT 25.320 178.550 27.940 178.690 ;
        RECT 23.940 178.490 24.260 178.550 ;
        RECT 25.320 178.490 25.640 178.550 ;
        RECT 25.795 178.505 26.085 178.550 ;
        RECT 27.620 178.490 27.940 178.550 ;
        RECT 34.980 178.690 35.300 178.750 ;
        RECT 35.530 178.690 35.670 178.890 ;
        RECT 34.980 178.550 35.670 178.690 ;
        RECT 34.980 178.490 35.300 178.550 ;
        RECT 35.915 178.505 36.205 178.735 ;
        RECT 23.370 178.350 23.660 178.395 ;
        RECT 29.920 178.350 30.240 178.410 ;
        RECT 23.370 178.210 30.240 178.350 ;
        RECT 23.370 178.165 23.660 178.210 ;
        RECT 29.920 178.150 30.240 178.210 ;
        RECT 22.560 177.810 22.880 178.070 ;
        RECT 35.990 178.010 36.130 178.505 ;
        RECT 36.360 178.490 36.680 178.750 ;
        RECT 37.280 178.490 37.600 178.750 ;
        RECT 37.740 178.690 38.060 178.750 ;
        RECT 40.055 178.690 40.345 178.735 ;
        RECT 37.740 178.550 40.345 178.690 ;
        RECT 37.740 178.490 38.060 178.550 ;
        RECT 40.055 178.505 40.345 178.550 ;
        RECT 37.370 178.350 37.510 178.490 ;
        RECT 39.595 178.350 39.885 178.395 ;
        RECT 37.370 178.210 39.885 178.350 ;
        RECT 40.590 178.350 40.730 178.890 ;
        RECT 41.880 178.830 42.200 179.090 ;
        RECT 49.790 179.075 49.930 179.230 ;
        RECT 55.220 179.170 55.540 179.230 ;
        RECT 64.510 179.230 73.480 179.370 ;
        RECT 43.275 179.030 43.565 179.075 ;
        RECT 49.715 179.030 50.005 179.075 ;
        RECT 42.430 178.890 43.565 179.030 ;
        RECT 49.605 178.890 50.005 179.030 ;
        RECT 41.420 178.490 41.740 178.750 ;
        RECT 42.430 178.735 42.570 178.890 ;
        RECT 43.275 178.845 43.565 178.890 ;
        RECT 49.715 178.845 50.005 178.890 ;
        RECT 63.975 179.030 64.265 179.075 ;
        RECT 64.510 179.030 64.650 179.230 ;
        RECT 73.160 179.170 73.480 179.230 ;
        RECT 92.570 179.230 98.305 179.370 ;
        RECT 92.570 179.090 92.710 179.230 ;
        RECT 94.335 179.185 94.625 179.230 ;
        RECT 98.015 179.185 98.305 179.230 ;
        RECT 98.460 179.370 98.780 179.430 ;
        RECT 103.995 179.370 104.285 179.415 ;
        RECT 109.040 179.370 109.360 179.430 ;
        RECT 115.110 179.415 115.250 179.570 ;
        RECT 116.490 179.570 119.020 179.710 ;
        RECT 98.460 179.230 109.360 179.370 ;
        RECT 98.460 179.170 98.780 179.230 ;
        RECT 103.995 179.185 104.285 179.230 ;
        RECT 109.040 179.170 109.360 179.230 ;
        RECT 115.035 179.185 115.325 179.415 ;
        RECT 115.480 179.370 115.800 179.430 ;
        RECT 116.490 179.370 116.630 179.570 ;
        RECT 118.700 179.510 119.020 179.570 ;
        RECT 119.620 179.710 119.940 179.770 ;
        RECT 121.460 179.710 121.780 179.770 ;
        RECT 119.620 179.570 121.780 179.710 ;
        RECT 119.620 179.510 119.940 179.570 ;
        RECT 121.460 179.510 121.780 179.570 ;
        RECT 124.235 179.525 124.525 179.755 ;
        RECT 115.480 179.230 116.630 179.370 ;
        RECT 117.335 179.370 117.625 179.415 ;
        RECT 117.780 179.370 118.100 179.430 ;
        RECT 117.335 179.230 118.100 179.370 ;
        RECT 118.790 179.370 118.930 179.510 ;
        RECT 121.935 179.370 122.225 179.415 ;
        RECT 118.790 179.230 122.225 179.370 ;
        RECT 63.975 178.890 64.650 179.030 ;
        RECT 64.895 179.030 65.185 179.075 ;
        RECT 66.275 179.030 66.565 179.075 ;
        RECT 64.895 178.890 66.565 179.030 ;
        RECT 63.975 178.845 64.265 178.890 ;
        RECT 64.895 178.845 65.185 178.890 ;
        RECT 66.275 178.845 66.565 178.890 ;
        RECT 67.640 179.030 67.960 179.090 ;
        RECT 67.640 178.890 71.090 179.030 ;
        RECT 67.640 178.830 67.960 178.890 ;
        RECT 42.355 178.505 42.645 178.735 ;
        RECT 42.815 178.505 43.105 178.735 ;
        RECT 42.890 178.350 43.030 178.505 ;
        RECT 43.720 178.490 44.040 178.750 ;
        RECT 47.400 178.690 47.720 178.750 ;
        RECT 53.395 178.690 53.685 178.735 ;
        RECT 47.400 178.550 53.685 178.690 ;
        RECT 47.400 178.490 47.720 178.550 ;
        RECT 53.395 178.505 53.685 178.550 ;
        RECT 54.315 178.690 54.605 178.735 ;
        RECT 57.520 178.690 57.840 178.750 ;
        RECT 54.315 178.550 57.840 178.690 ;
        RECT 54.315 178.505 54.605 178.550 ;
        RECT 57.520 178.490 57.840 178.550 ;
        RECT 64.435 178.505 64.725 178.735 ;
        RECT 65.355 178.505 65.645 178.735 ;
        RECT 68.100 178.690 68.420 178.750 ;
        RECT 69.020 178.690 69.340 178.750 ;
        RECT 68.100 178.550 69.340 178.690 ;
        RECT 40.590 178.210 43.030 178.350 ;
        RECT 52.140 178.350 52.430 178.395 ;
        RECT 53.855 178.350 54.145 178.395 ;
        RECT 52.140 178.210 54.145 178.350 ;
        RECT 39.595 178.165 39.885 178.210 ;
        RECT 52.140 178.165 52.430 178.210 ;
        RECT 53.855 178.165 54.145 178.210 ;
        RECT 36.865 178.010 37.155 178.055 ;
        RECT 35.990 177.870 37.155 178.010 ;
        RECT 36.865 177.825 37.155 177.870 ;
        RECT 38.660 178.010 38.980 178.070 ;
        RECT 39.135 178.010 39.425 178.055 ;
        RECT 38.660 177.870 39.425 178.010 ;
        RECT 38.660 177.810 38.980 177.870 ;
        RECT 39.135 177.825 39.425 177.870 ;
        RECT 40.975 178.010 41.265 178.055 ;
        RECT 41.420 178.010 41.740 178.070 ;
        RECT 46.020 178.010 46.340 178.070 ;
        RECT 40.975 177.870 46.340 178.010 ;
        RECT 40.975 177.825 41.265 177.870 ;
        RECT 41.420 177.810 41.740 177.870 ;
        RECT 46.020 177.810 46.340 177.870 ;
        RECT 51.080 177.810 51.400 178.070 ;
        RECT 51.540 177.810 51.860 178.070 ;
        RECT 52.920 177.810 53.240 178.070 ;
        RECT 62.580 178.010 62.900 178.070 ;
        RECT 63.055 178.010 63.345 178.055 ;
        RECT 62.580 177.870 63.345 178.010 ;
        RECT 64.510 178.010 64.650 178.505 ;
        RECT 65.430 178.350 65.570 178.505 ;
        RECT 68.100 178.490 68.420 178.550 ;
        RECT 69.020 178.490 69.340 178.550 ;
        RECT 70.400 178.350 70.720 178.410 ;
        RECT 65.430 178.210 70.720 178.350 ;
        RECT 70.950 178.350 71.090 178.890 ;
        RECT 72.790 178.890 74.770 179.030 ;
        RECT 71.320 178.690 71.640 178.750 ;
        RECT 72.790 178.735 72.930 178.890 ;
        RECT 74.630 178.750 74.770 178.890 ;
        RECT 92.480 178.830 92.800 179.090 ;
        RECT 95.240 179.030 95.560 179.090 ;
        RECT 96.635 179.030 96.925 179.075 ;
        RECT 102.140 179.030 102.460 179.090 ;
        RECT 113.640 179.030 113.960 179.090 ;
        RECT 95.240 178.890 96.925 179.030 ;
        RECT 95.240 178.830 95.560 178.890 ;
        RECT 96.635 178.845 96.925 178.890 ;
        RECT 100.390 178.890 102.460 179.030 ;
        RECT 72.715 178.690 73.005 178.735 ;
        RECT 71.320 178.550 73.005 178.690 ;
        RECT 71.320 178.490 71.640 178.550 ;
        RECT 72.715 178.505 73.005 178.550 ;
        RECT 73.620 178.490 73.940 178.750 ;
        RECT 74.540 178.490 74.860 178.750 ;
        RECT 75.015 178.505 75.305 178.735 ;
        RECT 74.095 178.350 74.385 178.395 ;
        RECT 75.090 178.350 75.230 178.505 ;
        RECT 75.920 178.490 76.240 178.750 ;
        RECT 79.600 178.690 79.920 178.750 ;
        RECT 82.375 178.690 82.665 178.735 ;
        RECT 79.600 178.550 82.665 178.690 ;
        RECT 79.600 178.490 79.920 178.550 ;
        RECT 82.375 178.505 82.665 178.550 ;
        RECT 89.720 178.690 90.040 178.750 ;
        RECT 92.035 178.690 92.325 178.735 ;
        RECT 89.720 178.550 92.325 178.690 ;
        RECT 92.570 178.690 92.710 178.830 ;
        RECT 92.955 178.690 93.245 178.735 ;
        RECT 92.570 178.550 93.245 178.690 ;
        RECT 89.720 178.490 90.040 178.550 ;
        RECT 92.035 178.505 92.325 178.550 ;
        RECT 92.955 178.505 93.245 178.550 ;
        RECT 93.415 178.505 93.705 178.735 ;
        RECT 94.335 178.690 94.625 178.735 ;
        RECT 97.080 178.690 97.400 178.750 ;
        RECT 98.000 178.690 98.320 178.750 ;
        RECT 99.840 178.690 100.160 178.750 ;
        RECT 100.390 178.735 100.530 178.890 ;
        RECT 102.140 178.830 102.460 178.890 ;
        RECT 112.270 178.890 113.960 179.030 ;
        RECT 115.110 179.030 115.250 179.185 ;
        RECT 115.480 179.170 115.800 179.230 ;
        RECT 117.335 179.185 117.625 179.230 ;
        RECT 117.780 179.170 118.100 179.230 ;
        RECT 121.935 179.185 122.225 179.230 ;
        RECT 118.240 179.030 118.560 179.090 ;
        RECT 118.715 179.030 119.005 179.075 ;
        RECT 115.110 178.890 119.005 179.030 ;
        RECT 94.335 178.550 97.770 178.690 ;
        RECT 94.335 178.505 94.625 178.550 ;
        RECT 70.950 178.210 75.230 178.350 ;
        RECT 93.490 178.350 93.630 178.505 ;
        RECT 97.080 178.490 97.400 178.550 ;
        RECT 95.700 178.350 96.020 178.410 ;
        RECT 93.490 178.210 96.020 178.350 ;
        RECT 97.630 178.350 97.770 178.550 ;
        RECT 98.000 178.550 100.160 178.690 ;
        RECT 98.000 178.490 98.320 178.550 ;
        RECT 99.840 178.490 100.160 178.550 ;
        RECT 100.315 178.505 100.605 178.735 ;
        RECT 101.235 178.505 101.525 178.735 ;
        RECT 105.370 178.505 105.660 178.735 ;
        RECT 105.835 178.690 106.125 178.735 ;
        RECT 107.200 178.690 107.520 178.750 ;
        RECT 105.835 178.550 107.520 178.690 ;
        RECT 112.270 178.565 112.410 178.890 ;
        RECT 113.640 178.830 113.960 178.890 ;
        RECT 118.240 178.830 118.560 178.890 ;
        RECT 118.715 178.845 119.005 178.890 ;
        RECT 119.635 179.030 119.925 179.075 ;
        RECT 122.380 179.030 122.700 179.090 ;
        RECT 119.635 178.890 122.700 179.030 ;
        RECT 119.635 178.845 119.925 178.890 ;
        RECT 122.380 178.830 122.700 178.890 ;
        RECT 122.855 179.030 123.145 179.075 ;
        RECT 124.310 179.030 124.450 179.525 ;
        RECT 133.880 179.510 134.200 179.770 ;
        RECT 125.600 179.030 125.920 179.090 ;
        RECT 122.855 178.890 125.920 179.030 ;
        RECT 122.855 178.845 123.145 178.890 ;
        RECT 125.600 178.830 125.920 178.890 ;
        RECT 129.280 179.030 129.600 179.090 ;
        RECT 136.655 179.030 136.945 179.075 ;
        RECT 129.280 178.890 136.945 179.030 ;
        RECT 129.280 178.830 129.600 178.890 ;
        RECT 136.655 178.845 136.945 178.890 ;
        RECT 115.020 178.690 115.340 178.750 ;
        RECT 105.835 178.505 106.125 178.550 ;
        RECT 101.310 178.350 101.450 178.505 ;
        RECT 97.630 178.210 101.450 178.350 ;
        RECT 105.450 178.350 105.590 178.505 ;
        RECT 107.200 178.490 107.520 178.550 ;
        RECT 110.420 178.350 110.740 178.410 ;
        RECT 105.450 178.210 110.740 178.350 ;
        RECT 112.045 178.380 112.410 178.565 ;
        RECT 113.270 178.550 115.340 178.690 ;
        RECT 113.270 178.395 113.410 178.550 ;
        RECT 115.020 178.490 115.340 178.550 ;
        RECT 115.940 178.690 116.260 178.750 ;
        RECT 115.940 178.550 118.930 178.690 ;
        RECT 115.940 178.490 116.260 178.550 ;
        RECT 112.045 178.335 112.335 178.380 ;
        RECT 70.400 178.150 70.720 178.210 ;
        RECT 74.095 178.165 74.385 178.210 ;
        RECT 95.700 178.150 96.020 178.210 ;
        RECT 110.420 178.150 110.740 178.210 ;
        RECT 113.195 178.165 113.485 178.395 ;
        RECT 67.640 178.010 67.960 178.070 ;
        RECT 64.510 177.870 67.960 178.010 ;
        RECT 62.580 177.810 62.900 177.870 ;
        RECT 63.055 177.825 63.345 177.870 ;
        RECT 67.640 177.810 67.960 177.870 ;
        RECT 69.955 178.010 70.245 178.055 ;
        RECT 71.320 178.010 71.640 178.070 ;
        RECT 69.955 177.870 71.640 178.010 ;
        RECT 69.955 177.825 70.245 177.870 ;
        RECT 71.320 177.810 71.640 177.870 ;
        RECT 75.475 178.010 75.765 178.055 ;
        RECT 77.760 178.010 78.080 178.070 ;
        RECT 75.475 177.870 78.080 178.010 ;
        RECT 75.475 177.825 75.765 177.870 ;
        RECT 77.760 177.810 78.080 177.870 ;
        RECT 84.200 178.010 84.520 178.070 ;
        RECT 85.120 178.010 85.440 178.070 ;
        RECT 85.595 178.010 85.885 178.055 ;
        RECT 84.200 177.870 85.885 178.010 ;
        RECT 84.200 177.810 84.520 177.870 ;
        RECT 85.120 177.810 85.440 177.870 ;
        RECT 85.595 177.825 85.885 177.870 ;
        RECT 92.495 178.010 92.785 178.055 ;
        RECT 98.000 178.010 98.320 178.070 ;
        RECT 92.495 177.870 98.320 178.010 ;
        RECT 92.495 177.825 92.785 177.870 ;
        RECT 98.000 177.810 98.320 177.870 ;
        RECT 98.935 178.010 99.225 178.055 ;
        RECT 110.880 178.010 111.200 178.070 ;
        RECT 98.935 177.870 111.200 178.010 ;
        RECT 98.935 177.825 99.225 177.870 ;
        RECT 110.880 177.810 111.200 177.870 ;
        RECT 111.340 177.810 111.660 178.070 ;
        RECT 115.940 177.810 116.260 178.070 ;
        RECT 116.490 178.055 116.630 178.550 ;
        RECT 118.790 178.410 118.930 178.550 ;
        RECT 119.175 178.660 119.465 178.735 ;
        RECT 119.175 178.640 119.850 178.660 ;
        RECT 119.175 178.520 119.940 178.640 ;
        RECT 119.175 178.505 119.465 178.520 ;
        RECT 118.700 178.150 119.020 178.410 ;
        RECT 119.620 178.380 119.940 178.520 ;
        RECT 121.475 178.505 121.765 178.735 ;
        RECT 122.470 178.690 122.610 178.830 ;
        RECT 123.315 178.690 123.605 178.735 ;
        RECT 122.470 178.550 123.605 178.690 ;
        RECT 123.315 178.505 123.605 178.550 ;
        RECT 121.550 178.350 121.690 178.505 ;
        RECT 135.720 178.490 136.040 178.750 ;
        RECT 138.035 178.505 138.325 178.735 ;
        RECT 120.170 178.210 121.690 178.350 ;
        RECT 130.200 178.350 130.520 178.410 ;
        RECT 138.110 178.350 138.250 178.505 ;
        RECT 139.860 178.490 140.180 178.750 ;
        RECT 130.200 178.210 138.250 178.350 ;
        RECT 116.415 177.825 116.705 178.055 ;
        RECT 117.780 178.010 118.100 178.070 ;
        RECT 120.170 178.010 120.310 178.210 ;
        RECT 130.200 178.150 130.520 178.210 ;
        RECT 117.780 177.870 120.310 178.010 ;
        RECT 121.015 178.010 121.305 178.055 ;
        RECT 121.920 178.010 122.240 178.070 ;
        RECT 121.015 177.870 122.240 178.010 ;
        RECT 117.780 177.810 118.100 177.870 ;
        RECT 121.015 177.825 121.305 177.870 ;
        RECT 121.920 177.810 122.240 177.870 ;
        RECT 122.855 178.010 123.145 178.055 ;
        RECT 123.760 178.010 124.080 178.070 ;
        RECT 122.855 177.870 124.080 178.010 ;
        RECT 122.855 177.825 123.145 177.870 ;
        RECT 123.760 177.810 124.080 177.870 ;
        RECT 131.580 178.010 131.900 178.070 ;
        RECT 136.195 178.010 136.485 178.055 ;
        RECT 131.580 177.870 136.485 178.010 ;
        RECT 131.580 177.810 131.900 177.870 ;
        RECT 136.195 177.825 136.485 177.870 ;
        RECT 138.940 177.810 139.260 178.070 ;
        RECT 140.795 178.010 141.085 178.055 ;
        RECT 141.700 178.010 142.020 178.070 ;
        RECT 140.795 177.870 142.020 178.010 ;
        RECT 140.795 177.825 141.085 177.870 ;
        RECT 141.700 177.810 142.020 177.870 ;
        RECT 17.430 177.190 143.010 177.670 ;
        RECT 29.920 176.790 30.240 177.050 ;
        RECT 46.480 176.990 46.800 177.050 ;
        RECT 48.875 176.990 49.165 177.035 ;
        RECT 46.110 176.850 49.165 176.990 ;
        RECT 22.560 176.650 22.880 176.710 ;
        RECT 23.340 176.650 23.630 176.695 ;
        RECT 22.560 176.510 23.630 176.650 ;
        RECT 22.560 176.450 22.880 176.510 ;
        RECT 23.340 176.465 23.630 176.510 ;
        RECT 16.120 176.310 16.440 176.370 ;
        RECT 18.895 176.310 19.185 176.355 ;
        RECT 16.120 176.170 19.185 176.310 ;
        RECT 16.120 176.110 16.440 176.170 ;
        RECT 18.895 176.125 19.185 176.170 ;
        RECT 28.540 176.310 28.860 176.370 ;
        RECT 29.475 176.310 29.765 176.355 ;
        RECT 28.540 176.170 29.765 176.310 ;
        RECT 28.540 176.110 28.860 176.170 ;
        RECT 29.475 176.125 29.765 176.170 ;
        RECT 30.395 176.310 30.685 176.355 ;
        RECT 30.840 176.310 31.160 176.370 ;
        RECT 46.110 176.355 46.250 176.850 ;
        RECT 46.480 176.790 46.800 176.850 ;
        RECT 48.875 176.805 49.165 176.850 ;
        RECT 49.715 176.990 50.005 177.035 ;
        RECT 57.520 176.990 57.840 177.050 ;
        RECT 49.715 176.850 57.840 176.990 ;
        RECT 49.715 176.805 50.005 176.850 ;
        RECT 57.520 176.790 57.840 176.850 ;
        RECT 68.575 176.990 68.865 177.035 ;
        RECT 70.860 176.990 71.180 177.050 ;
        RECT 68.575 176.850 71.180 176.990 ;
        RECT 68.575 176.805 68.865 176.850 ;
        RECT 70.860 176.790 71.180 176.850 ;
        RECT 71.320 176.790 71.640 177.050 ;
        RECT 73.160 176.990 73.480 177.050 ;
        RECT 75.920 176.990 76.240 177.050 ;
        RECT 73.160 176.850 76.240 176.990 ;
        RECT 73.160 176.790 73.480 176.850 ;
        RECT 75.920 176.790 76.240 176.850 ;
        RECT 79.600 176.790 79.920 177.050 ;
        RECT 122.840 176.990 123.160 177.050 ;
        RECT 114.190 176.850 123.160 176.990 ;
        RECT 47.875 176.465 48.165 176.695 ;
        RECT 53.380 176.650 53.700 176.710 ;
        RECT 50.250 176.510 53.700 176.650 ;
        RECT 30.395 176.170 31.160 176.310 ;
        RECT 30.395 176.125 30.685 176.170 ;
        RECT 30.840 176.110 31.160 176.170 ;
        RECT 46.035 176.125 46.325 176.355 ;
        RECT 46.495 176.125 46.785 176.355 ;
        RECT 46.940 176.310 47.260 176.370 ;
        RECT 47.415 176.310 47.705 176.355 ;
        RECT 47.950 176.310 48.090 176.465 ;
        RECT 50.250 176.355 50.390 176.510 ;
        RECT 53.380 176.450 53.700 176.510 ;
        RECT 75.460 176.650 75.780 176.710 ;
        RECT 79.140 176.650 79.460 176.710 ;
        RECT 75.460 176.510 79.460 176.650 ;
        RECT 75.460 176.450 75.780 176.510 ;
        RECT 79.140 176.450 79.460 176.510 ;
        RECT 46.940 176.170 48.090 176.310 ;
        RECT 21.640 175.970 21.960 176.030 ;
        RECT 22.115 175.970 22.405 176.015 ;
        RECT 21.640 175.830 22.405 175.970 ;
        RECT 21.640 175.770 21.960 175.830 ;
        RECT 22.115 175.785 22.405 175.830 ;
        RECT 22.995 175.970 23.285 176.015 ;
        RECT 24.185 175.970 24.475 176.015 ;
        RECT 26.705 175.970 26.995 176.015 ;
        RECT 22.995 175.830 26.995 175.970 ;
        RECT 22.995 175.785 23.285 175.830 ;
        RECT 24.185 175.785 24.475 175.830 ;
        RECT 26.705 175.785 26.995 175.830 ;
        RECT 45.560 175.970 45.880 176.030 ;
        RECT 46.110 175.970 46.250 176.125 ;
        RECT 45.560 175.830 46.250 175.970 ;
        RECT 45.560 175.770 45.880 175.830 ;
        RECT 22.600 175.630 22.890 175.675 ;
        RECT 24.700 175.630 24.990 175.675 ;
        RECT 26.270 175.630 26.560 175.675 ;
        RECT 22.600 175.490 26.560 175.630 ;
        RECT 22.600 175.445 22.890 175.490 ;
        RECT 24.700 175.445 24.990 175.490 ;
        RECT 26.270 175.445 26.560 175.490 ;
        RECT 19.815 175.290 20.105 175.335 ;
        RECT 28.080 175.290 28.400 175.350 ;
        RECT 19.815 175.150 28.400 175.290 ;
        RECT 19.815 175.105 20.105 175.150 ;
        RECT 28.080 175.090 28.400 175.150 ;
        RECT 29.000 175.090 29.320 175.350 ;
        RECT 44.180 175.290 44.500 175.350 ;
        RECT 45.100 175.290 45.420 175.350 ;
        RECT 46.570 175.290 46.710 176.125 ;
        RECT 46.940 176.110 47.260 176.170 ;
        RECT 47.415 176.125 47.705 176.170 ;
        RECT 47.400 175.430 47.720 175.690 ;
        RECT 47.950 175.630 48.090 176.170 ;
        RECT 50.175 176.125 50.465 176.355 ;
        RECT 51.510 176.310 51.800 176.355 ;
        RECT 52.920 176.310 53.240 176.370 ;
        RECT 51.510 176.170 53.240 176.310 ;
        RECT 51.510 176.125 51.800 176.170 ;
        RECT 52.920 176.110 53.240 176.170 ;
        RECT 63.010 176.310 63.300 176.355 ;
        RECT 69.495 176.310 69.785 176.355 ;
        RECT 63.010 176.170 69.785 176.310 ;
        RECT 63.010 176.125 63.300 176.170 ;
        RECT 69.495 176.125 69.785 176.170 ;
        RECT 70.400 176.110 70.720 176.370 ;
        RECT 71.780 176.110 72.100 176.370 ;
        RECT 72.240 176.110 72.560 176.370 ;
        RECT 73.590 176.310 73.880 176.355 ;
        RECT 76.380 176.310 76.700 176.370 ;
        RECT 73.590 176.170 76.700 176.310 ;
        RECT 73.590 176.125 73.880 176.170 ;
        RECT 76.380 176.110 76.700 176.170 ;
        RECT 51.055 175.970 51.345 176.015 ;
        RECT 52.245 175.970 52.535 176.015 ;
        RECT 54.765 175.970 55.055 176.015 ;
        RECT 51.055 175.830 55.055 175.970 ;
        RECT 51.055 175.785 51.345 175.830 ;
        RECT 52.245 175.785 52.535 175.830 ;
        RECT 54.765 175.785 55.055 175.830 ;
        RECT 59.820 175.970 60.140 176.030 ;
        RECT 61.675 175.970 61.965 176.015 ;
        RECT 59.820 175.830 61.965 175.970 ;
        RECT 59.820 175.770 60.140 175.830 ;
        RECT 61.675 175.785 61.965 175.830 ;
        RECT 62.555 175.970 62.845 176.015 ;
        RECT 63.745 175.970 64.035 176.015 ;
        RECT 66.265 175.970 66.555 176.015 ;
        RECT 62.555 175.830 66.555 175.970 ;
        RECT 62.555 175.785 62.845 175.830 ;
        RECT 63.745 175.785 64.035 175.830 ;
        RECT 66.265 175.785 66.555 175.830 ;
        RECT 73.135 175.970 73.425 176.015 ;
        RECT 74.325 175.970 74.615 176.015 ;
        RECT 76.845 175.970 77.135 176.015 ;
        RECT 73.135 175.830 77.135 175.970 ;
        RECT 73.135 175.785 73.425 175.830 ;
        RECT 74.325 175.785 74.615 175.830 ;
        RECT 76.845 175.785 77.135 175.830 ;
        RECT 50.660 175.630 50.950 175.675 ;
        RECT 52.760 175.630 53.050 175.675 ;
        RECT 54.330 175.630 54.620 175.675 ;
        RECT 47.950 175.490 50.390 175.630 ;
        RECT 48.795 175.290 49.085 175.335 ;
        RECT 44.180 175.150 49.085 175.290 ;
        RECT 50.250 175.290 50.390 175.490 ;
        RECT 50.660 175.490 54.620 175.630 ;
        RECT 50.660 175.445 50.950 175.490 ;
        RECT 52.760 175.445 53.050 175.490 ;
        RECT 54.330 175.445 54.620 175.490 ;
        RECT 62.160 175.630 62.450 175.675 ;
        RECT 64.260 175.630 64.550 175.675 ;
        RECT 65.830 175.630 66.120 175.675 ;
        RECT 62.160 175.490 66.120 175.630 ;
        RECT 62.160 175.445 62.450 175.490 ;
        RECT 64.260 175.445 64.550 175.490 ;
        RECT 65.830 175.445 66.120 175.490 ;
        RECT 72.740 175.630 73.030 175.675 ;
        RECT 74.840 175.630 75.130 175.675 ;
        RECT 76.410 175.630 76.700 175.675 ;
        RECT 79.690 175.630 79.830 176.790 ;
        RECT 113.655 176.650 113.945 176.695 ;
        RECT 72.740 175.490 76.700 175.630 ;
        RECT 72.740 175.445 73.030 175.490 ;
        RECT 74.840 175.445 75.130 175.490 ;
        RECT 76.410 175.445 76.700 175.490 ;
        RECT 78.770 175.490 79.830 175.630 ;
        RECT 80.150 176.510 90.870 176.650 ;
        RECT 57.075 175.290 57.365 175.335 ;
        RECT 59.360 175.290 59.680 175.350 ;
        RECT 50.250 175.150 59.680 175.290 ;
        RECT 44.180 175.090 44.500 175.150 ;
        RECT 45.100 175.090 45.420 175.150 ;
        RECT 48.795 175.105 49.085 175.150 ;
        RECT 57.075 175.105 57.365 175.150 ;
        RECT 59.360 175.090 59.680 175.150 ;
        RECT 73.160 175.290 73.480 175.350 ;
        RECT 78.770 175.290 78.910 175.490 ;
        RECT 80.150 175.350 80.290 176.510 ;
        RECT 85.235 176.310 85.525 176.355 ;
        RECT 86.040 176.310 86.360 176.370 ;
        RECT 85.235 176.170 86.360 176.310 ;
        RECT 85.235 176.125 85.525 176.170 ;
        RECT 86.040 176.110 86.360 176.170 ;
        RECT 86.515 176.310 86.805 176.355 ;
        RECT 90.180 176.310 90.500 176.370 ;
        RECT 86.515 176.170 90.500 176.310 ;
        RECT 86.515 176.125 86.805 176.170 ;
        RECT 90.180 176.110 90.500 176.170 ;
        RECT 81.925 175.970 82.215 176.015 ;
        RECT 84.445 175.970 84.735 176.015 ;
        RECT 85.635 175.970 85.925 176.015 ;
        RECT 81.925 175.830 85.925 175.970 ;
        RECT 81.925 175.785 82.215 175.830 ;
        RECT 84.445 175.785 84.735 175.830 ;
        RECT 85.635 175.785 85.925 175.830 ;
        RECT 89.735 175.970 90.025 176.015 ;
        RECT 90.730 175.970 90.870 176.510 ;
        RECT 111.890 176.510 113.945 176.650 ;
        RECT 111.890 176.370 112.030 176.510 ;
        RECT 113.655 176.465 113.945 176.510 ;
        RECT 110.895 176.310 111.185 176.355 ;
        RECT 111.800 176.310 112.120 176.370 ;
        RECT 110.895 176.170 112.120 176.310 ;
        RECT 110.895 176.125 111.185 176.170 ;
        RECT 111.800 176.110 112.120 176.170 ;
        RECT 112.275 176.310 112.565 176.355 ;
        RECT 114.190 176.310 114.330 176.850 ;
        RECT 122.840 176.790 123.160 176.850 ;
        RECT 124.235 176.990 124.525 177.035 ;
        RECT 128.820 176.990 129.140 177.050 ;
        RECT 137.575 176.990 137.865 177.035 ;
        RECT 124.235 176.850 129.140 176.990 ;
        RECT 124.235 176.805 124.525 176.850 ;
        RECT 128.820 176.790 129.140 176.850 ;
        RECT 129.370 176.850 137.865 176.990 ;
        RECT 116.860 176.650 117.180 176.710 ;
        RECT 119.635 176.650 119.925 176.695 ;
        RECT 123.300 176.650 123.620 176.710 ;
        RECT 116.860 176.510 124.910 176.650 ;
        RECT 116.860 176.450 117.180 176.510 ;
        RECT 119.635 176.465 119.925 176.510 ;
        RECT 123.300 176.450 123.620 176.510 ;
        RECT 112.275 176.170 114.330 176.310 ;
        RECT 112.275 176.125 112.565 176.170 ;
        RECT 114.560 176.110 114.880 176.370 ;
        RECT 115.955 176.310 116.245 176.355 ;
        RECT 117.780 176.310 118.100 176.370 ;
        RECT 115.955 176.170 118.100 176.310 ;
        RECT 115.955 176.125 116.245 176.170 ;
        RECT 117.780 176.110 118.100 176.170 ;
        RECT 118.240 176.310 118.560 176.370 ;
        RECT 118.715 176.310 119.005 176.355 ;
        RECT 120.540 176.310 120.860 176.370 ;
        RECT 118.240 176.170 120.860 176.310 ;
        RECT 118.240 176.110 118.560 176.170 ;
        RECT 118.715 176.125 119.005 176.170 ;
        RECT 120.540 176.110 120.860 176.170 ;
        RECT 121.015 176.310 121.305 176.355 ;
        RECT 121.460 176.310 121.780 176.370 ;
        RECT 121.015 176.170 121.780 176.310 ;
        RECT 121.015 176.125 121.305 176.170 ;
        RECT 121.460 176.110 121.780 176.170 ;
        RECT 121.920 176.110 122.240 176.370 ;
        RECT 124.770 176.355 124.910 176.510 ;
        RECT 122.395 176.125 122.685 176.355 ;
        RECT 122.855 176.125 123.145 176.355 ;
        RECT 124.695 176.125 124.985 176.355 ;
        RECT 126.075 176.310 126.365 176.355 ;
        RECT 127.900 176.310 128.220 176.370 ;
        RECT 129.370 176.355 129.510 176.850 ;
        RECT 137.575 176.805 137.865 176.850 ;
        RECT 126.075 176.170 128.220 176.310 ;
        RECT 126.075 176.125 126.365 176.170 ;
        RECT 89.735 175.830 90.870 175.970 ;
        RECT 111.340 175.970 111.660 176.030 ;
        RECT 113.640 175.970 113.960 176.030 ;
        RECT 111.340 175.830 113.960 175.970 ;
        RECT 89.735 175.785 90.025 175.830 ;
        RECT 111.340 175.770 111.660 175.830 ;
        RECT 113.640 175.770 113.960 175.830 ;
        RECT 115.480 175.970 115.800 176.030 ;
        RECT 116.415 175.970 116.705 176.015 ;
        RECT 115.480 175.830 116.705 175.970 ;
        RECT 115.480 175.770 115.800 175.830 ;
        RECT 116.415 175.785 116.705 175.830 ;
        RECT 117.335 175.970 117.625 176.015 ;
        RECT 120.080 175.970 120.400 176.030 ;
        RECT 122.470 175.970 122.610 176.125 ;
        RECT 117.335 175.830 118.470 175.970 ;
        RECT 117.335 175.785 117.625 175.830 ;
        RECT 82.360 175.630 82.650 175.675 ;
        RECT 83.930 175.630 84.220 175.675 ;
        RECT 86.030 175.630 86.320 175.675 ;
        RECT 82.360 175.490 86.320 175.630 ;
        RECT 82.360 175.445 82.650 175.490 ;
        RECT 83.930 175.445 84.220 175.490 ;
        RECT 86.030 175.445 86.320 175.490 ;
        RECT 111.800 175.430 112.120 175.690 ;
        RECT 117.780 175.630 118.100 175.690 ;
        RECT 112.350 175.490 118.100 175.630 ;
        RECT 118.330 175.630 118.470 175.830 ;
        RECT 120.080 175.830 122.610 175.970 ;
        RECT 120.080 175.770 120.400 175.830 ;
        RECT 121.000 175.630 121.320 175.690 ;
        RECT 122.930 175.630 123.070 176.125 ;
        RECT 127.900 176.110 128.220 176.170 ;
        RECT 129.295 176.125 129.585 176.355 ;
        RECT 129.740 176.310 130.060 176.370 ;
        RECT 130.660 176.310 130.980 176.370 ;
        RECT 132.040 176.355 132.360 176.370 ;
        RECT 129.740 176.170 130.980 176.310 ;
        RECT 129.740 176.110 130.060 176.170 ;
        RECT 130.660 176.110 130.980 176.170 ;
        RECT 132.010 176.125 132.360 176.355 ;
        RECT 137.650 176.310 137.790 176.805 ;
        RECT 140.795 176.310 141.085 176.355 ;
        RECT 137.650 176.170 141.085 176.310 ;
        RECT 140.795 176.125 141.085 176.170 ;
        RECT 132.040 176.110 132.360 176.125 ;
        RECT 126.520 175.770 126.840 176.030 ;
        RECT 131.555 175.970 131.845 176.015 ;
        RECT 132.745 175.970 133.035 176.015 ;
        RECT 135.265 175.970 135.555 176.015 ;
        RECT 131.555 175.830 135.555 175.970 ;
        RECT 131.555 175.785 131.845 175.830 ;
        RECT 132.745 175.785 133.035 175.830 ;
        RECT 135.265 175.785 135.555 175.830 ;
        RECT 118.330 175.490 119.850 175.630 ;
        RECT 73.160 175.150 78.910 175.290 ;
        RECT 79.155 175.290 79.445 175.335 ;
        RECT 80.060 175.290 80.380 175.350 ;
        RECT 79.155 175.150 80.380 175.290 ;
        RECT 73.160 175.090 73.480 175.150 ;
        RECT 79.155 175.105 79.445 175.150 ;
        RECT 80.060 175.090 80.380 175.150 ;
        RECT 80.980 175.290 81.300 175.350 ;
        RECT 86.975 175.290 87.265 175.335 ;
        RECT 80.980 175.150 87.265 175.290 ;
        RECT 80.980 175.090 81.300 175.150 ;
        RECT 86.975 175.105 87.265 175.150 ;
        RECT 107.660 175.290 107.980 175.350 ;
        RECT 112.350 175.290 112.490 175.490 ;
        RECT 117.780 175.430 118.100 175.490 ;
        RECT 107.660 175.150 112.490 175.290 ;
        RECT 112.720 175.290 113.040 175.350 ;
        RECT 113.195 175.290 113.485 175.335 ;
        RECT 112.720 175.150 113.485 175.290 ;
        RECT 107.660 175.090 107.980 175.150 ;
        RECT 112.720 175.090 113.040 175.150 ;
        RECT 113.195 175.105 113.485 175.150 ;
        RECT 115.035 175.290 115.325 175.335 ;
        RECT 115.940 175.290 116.260 175.350 ;
        RECT 115.035 175.150 116.260 175.290 ;
        RECT 115.035 175.105 115.325 175.150 ;
        RECT 115.940 175.090 116.260 175.150 ;
        RECT 116.875 175.290 117.165 175.335 ;
        RECT 117.320 175.290 117.640 175.350 ;
        RECT 116.875 175.150 117.640 175.290 ;
        RECT 116.875 175.105 117.165 175.150 ;
        RECT 117.320 175.090 117.640 175.150 ;
        RECT 118.240 175.090 118.560 175.350 ;
        RECT 119.710 175.290 119.850 175.490 ;
        RECT 121.000 175.490 123.070 175.630 ;
        RECT 121.000 175.430 121.320 175.490 ;
        RECT 130.200 175.430 130.520 175.690 ;
        RECT 131.160 175.630 131.450 175.675 ;
        RECT 133.260 175.630 133.550 175.675 ;
        RECT 134.830 175.630 135.120 175.675 ;
        RECT 131.160 175.490 135.120 175.630 ;
        RECT 131.160 175.445 131.450 175.490 ;
        RECT 133.260 175.445 133.550 175.490 ;
        RECT 134.830 175.445 135.120 175.490 ;
        RECT 124.680 175.290 125.000 175.350 ;
        RECT 119.710 175.150 125.000 175.290 ;
        RECT 124.680 175.090 125.000 175.150 ;
        RECT 138.020 175.090 138.340 175.350 ;
        RECT 17.430 174.470 143.010 174.950 ;
        RECT 28.540 174.070 28.860 174.330 ;
        RECT 37.755 174.270 38.045 174.315 ;
        RECT 38.660 174.270 38.980 174.330 ;
        RECT 37.755 174.130 38.980 174.270 ;
        RECT 37.755 174.085 38.045 174.130 ;
        RECT 21.680 173.930 21.970 173.975 ;
        RECT 23.780 173.930 24.070 173.975 ;
        RECT 25.350 173.930 25.640 173.975 ;
        RECT 21.680 173.790 25.640 173.930 ;
        RECT 21.680 173.745 21.970 173.790 ;
        RECT 23.780 173.745 24.070 173.790 ;
        RECT 25.350 173.745 25.640 173.790 ;
        RECT 22.075 173.590 22.365 173.635 ;
        RECT 23.265 173.590 23.555 173.635 ;
        RECT 25.785 173.590 26.075 173.635 ;
        RECT 22.075 173.450 26.075 173.590 ;
        RECT 22.075 173.405 22.365 173.450 ;
        RECT 23.265 173.405 23.555 173.450 ;
        RECT 25.785 173.405 26.075 173.450 ;
        RECT 28.080 173.590 28.400 173.650 ;
        RECT 37.830 173.590 37.970 174.085 ;
        RECT 38.660 174.070 38.980 174.130 ;
        RECT 68.100 174.070 68.420 174.330 ;
        RECT 71.780 174.270 72.100 174.330 ;
        RECT 75.460 174.270 75.780 174.330 ;
        RECT 71.780 174.130 75.780 174.270 ;
        RECT 71.780 174.070 72.100 174.130 ;
        RECT 75.460 174.070 75.780 174.130 ;
        RECT 75.920 174.270 76.240 174.330 ;
        RECT 78.695 174.270 78.985 174.315 ;
        RECT 75.920 174.130 78.985 174.270 ;
        RECT 75.920 174.070 76.240 174.130 ;
        RECT 78.695 174.085 78.985 174.130 ;
        RECT 79.140 174.270 79.460 174.330 ;
        RECT 79.615 174.270 79.905 174.315 ;
        RECT 82.360 174.270 82.680 174.330 ;
        RECT 79.140 174.130 82.680 174.270 ;
        RECT 79.140 174.070 79.460 174.130 ;
        RECT 79.615 174.085 79.905 174.130 ;
        RECT 82.360 174.070 82.680 174.130 ;
        RECT 86.040 174.270 86.360 174.330 ;
        RECT 86.515 174.270 86.805 174.315 ;
        RECT 86.040 174.130 86.805 174.270 ;
        RECT 86.040 174.070 86.360 174.130 ;
        RECT 86.515 174.085 86.805 174.130 ;
        RECT 111.800 174.270 112.120 174.330 ;
        RECT 113.655 174.270 113.945 174.315 ;
        RECT 111.800 174.130 113.945 174.270 ;
        RECT 111.800 174.070 112.120 174.130 ;
        RECT 39.595 173.930 39.885 173.975 ;
        RECT 40.500 173.930 40.820 173.990 ;
        RECT 39.595 173.790 40.820 173.930 ;
        RECT 39.595 173.745 39.885 173.790 ;
        RECT 40.500 173.730 40.820 173.790 ;
        RECT 40.960 173.930 41.280 173.990 ;
        RECT 45.100 173.930 45.420 173.990 ;
        RECT 51.540 173.930 51.830 173.975 ;
        RECT 53.110 173.930 53.400 173.975 ;
        RECT 55.210 173.930 55.500 173.975 ;
        RECT 40.960 173.790 48.550 173.930 ;
        RECT 40.960 173.730 41.280 173.790 ;
        RECT 45.100 173.730 45.420 173.790 ;
        RECT 42.355 173.590 42.645 173.635 ;
        RECT 43.720 173.590 44.040 173.650 ;
        RECT 28.080 173.450 33.370 173.590 ;
        RECT 28.080 173.390 28.400 173.450 ;
        RECT 21.195 173.250 21.485 173.295 ;
        RECT 21.640 173.250 21.960 173.310 ;
        RECT 23.940 173.250 24.260 173.310 ;
        RECT 21.195 173.110 24.260 173.250 ;
        RECT 21.195 173.065 21.485 173.110 ;
        RECT 21.640 173.050 21.960 173.110 ;
        RECT 23.940 173.050 24.260 173.110 ;
        RECT 26.240 173.250 26.560 173.310 ;
        RECT 28.555 173.250 28.845 173.295 ;
        RECT 26.240 173.110 28.845 173.250 ;
        RECT 26.240 173.050 26.560 173.110 ;
        RECT 28.555 173.065 28.845 173.110 ;
        RECT 29.000 173.250 29.320 173.310 ;
        RECT 29.475 173.250 29.765 173.295 ;
        RECT 32.220 173.250 32.540 173.310 ;
        RECT 33.230 173.295 33.370 173.450 ;
        RECT 36.910 173.450 37.970 173.590 ;
        RECT 38.750 173.450 44.040 173.590 ;
        RECT 36.910 173.295 37.050 173.450 ;
        RECT 38.750 173.295 38.890 173.450 ;
        RECT 42.355 173.405 42.645 173.450 ;
        RECT 43.720 173.390 44.040 173.450 ;
        RECT 44.180 173.590 44.500 173.650 ;
        RECT 47.875 173.590 48.165 173.635 ;
        RECT 44.180 173.450 48.165 173.590 ;
        RECT 44.180 173.390 44.500 173.450 ;
        RECT 47.875 173.405 48.165 173.450 ;
        RECT 29.000 173.110 32.540 173.250 ;
        RECT 29.000 173.050 29.320 173.110 ;
        RECT 29.475 173.065 29.765 173.110 ;
        RECT 32.220 173.050 32.540 173.110 ;
        RECT 33.155 173.065 33.445 173.295 ;
        RECT 36.370 173.065 36.660 173.295 ;
        RECT 36.835 173.065 37.125 173.295 ;
        RECT 37.295 173.065 37.585 173.295 ;
        RECT 38.675 173.065 38.965 173.295 ;
        RECT 22.560 172.955 22.880 172.970 ;
        RECT 22.530 172.725 22.880 172.955 ;
        RECT 35.900 172.910 36.220 172.970 ;
        RECT 36.405 172.910 36.545 173.065 ;
        RECT 37.370 172.910 37.510 173.065 ;
        RECT 40.960 173.050 41.280 173.310 ;
        RECT 41.435 173.250 41.725 173.295 ;
        RECT 41.880 173.250 42.200 173.310 ;
        RECT 41.435 173.110 42.200 173.250 ;
        RECT 41.435 173.065 41.725 173.110 ;
        RECT 41.880 173.050 42.200 173.110 ;
        RECT 42.815 173.250 43.105 173.295 ;
        RECT 43.275 173.250 43.565 173.295 ;
        RECT 44.640 173.250 44.960 173.310 ;
        RECT 42.815 173.110 44.960 173.250 ;
        RECT 42.815 173.065 43.105 173.110 ;
        RECT 43.275 173.065 43.565 173.110 ;
        RECT 44.640 173.050 44.960 173.110 ;
        RECT 46.955 173.250 47.245 173.295 ;
        RECT 48.410 173.250 48.550 173.790 ;
        RECT 51.540 173.790 55.500 173.930 ;
        RECT 51.540 173.745 51.830 173.790 ;
        RECT 53.110 173.745 53.400 173.790 ;
        RECT 55.210 173.745 55.500 173.790 ;
        RECT 59.360 173.730 59.680 173.990 ;
        RECT 61.700 173.930 61.990 173.975 ;
        RECT 63.800 173.930 64.090 173.975 ;
        RECT 65.370 173.930 65.660 173.975 ;
        RECT 61.700 173.790 65.660 173.930 ;
        RECT 61.700 173.745 61.990 173.790 ;
        RECT 63.800 173.745 64.090 173.790 ;
        RECT 65.370 173.745 65.660 173.790 ;
        RECT 72.790 173.790 74.770 173.930 ;
        RECT 51.105 173.590 51.395 173.635 ;
        RECT 53.625 173.590 53.915 173.635 ;
        RECT 54.815 173.590 55.105 173.635 ;
        RECT 51.105 173.450 55.105 173.590 ;
        RECT 51.105 173.405 51.395 173.450 ;
        RECT 53.625 173.405 53.915 173.450 ;
        RECT 54.815 173.405 55.105 173.450 ;
        RECT 62.095 173.590 62.385 173.635 ;
        RECT 63.285 173.590 63.575 173.635 ;
        RECT 65.805 173.590 66.095 173.635 ;
        RECT 72.790 173.590 72.930 173.790 ;
        RECT 62.095 173.450 66.095 173.590 ;
        RECT 62.095 173.405 62.385 173.450 ;
        RECT 63.285 173.405 63.575 173.450 ;
        RECT 65.805 173.405 66.095 173.450 ;
        RECT 68.650 173.450 72.930 173.590 ;
        RECT 74.630 173.590 74.770 173.790 ;
        RECT 75.000 173.730 75.320 173.990 ;
        RECT 83.740 173.930 84.060 173.990 ;
        RECT 112.275 173.930 112.565 173.975 ;
        RECT 83.740 173.790 88.110 173.930 ;
        RECT 83.740 173.730 84.060 173.790 ;
        RECT 75.460 173.590 75.780 173.650 ;
        RECT 76.395 173.590 76.685 173.635 ;
        RECT 74.630 173.450 76.685 173.590 ;
        RECT 55.695 173.250 55.985 173.295 ;
        RECT 59.820 173.250 60.140 173.310 ;
        RECT 62.580 173.295 62.900 173.310 ;
        RECT 68.650 173.295 68.790 173.450 ;
        RECT 75.460 173.390 75.780 173.450 ;
        RECT 76.395 173.405 76.685 173.450 ;
        RECT 76.840 173.390 77.160 173.650 ;
        RECT 77.315 173.590 77.605 173.635 ;
        RECT 79.140 173.590 79.460 173.650 ;
        RECT 77.315 173.450 79.460 173.590 ;
        RECT 77.315 173.405 77.605 173.450 ;
        RECT 79.140 173.390 79.460 173.450 ;
        RECT 80.060 173.390 80.380 173.650 ;
        RECT 83.280 173.390 83.600 173.650 ;
        RECT 84.200 173.390 84.520 173.650 ;
        RECT 87.435 173.590 87.725 173.635 ;
        RECT 84.750 173.450 87.725 173.590 ;
        RECT 61.215 173.250 61.505 173.295 ;
        RECT 62.550 173.250 62.900 173.295 ;
        RECT 46.955 173.110 48.550 173.250 ;
        RECT 53.470 173.110 61.505 173.250 ;
        RECT 62.385 173.110 62.900 173.250 ;
        RECT 46.955 173.065 47.245 173.110 ;
        RECT 53.470 172.970 53.610 173.110 ;
        RECT 55.695 173.065 55.985 173.110 ;
        RECT 59.820 173.050 60.140 173.110 ;
        RECT 61.215 173.065 61.505 173.110 ;
        RECT 62.550 173.065 62.900 173.110 ;
        RECT 68.575 173.065 68.865 173.295 ;
        RECT 69.495 173.250 69.785 173.295 ;
        RECT 72.700 173.250 73.020 173.310 ;
        RECT 69.495 173.110 73.020 173.250 ;
        RECT 69.495 173.065 69.785 173.110 ;
        RECT 62.580 173.050 62.900 173.065 ;
        RECT 72.700 173.050 73.020 173.110 ;
        RECT 74.080 173.050 74.400 173.310 ;
        RECT 75.920 173.050 76.240 173.310 ;
        RECT 78.190 173.250 78.480 173.295 ;
        RECT 77.850 173.110 78.480 173.250 ;
        RECT 45.115 172.910 45.405 172.955 ;
        RECT 22.560 172.710 22.880 172.725 ;
        RECT 34.150 172.770 45.405 172.910 ;
        RECT 28.080 172.370 28.400 172.630 ;
        RECT 34.150 172.615 34.290 172.770 ;
        RECT 35.900 172.710 36.220 172.770 ;
        RECT 45.115 172.725 45.405 172.770 ;
        RECT 45.560 172.910 45.880 172.970 ;
        RECT 45.560 172.770 49.470 172.910 ;
        RECT 45.560 172.710 45.880 172.770 ;
        RECT 34.075 172.385 34.365 172.615 ;
        RECT 34.980 172.370 35.300 172.630 ;
        RECT 40.040 172.370 40.360 172.630 ;
        RECT 46.020 172.370 46.340 172.630 ;
        RECT 48.780 172.370 49.100 172.630 ;
        RECT 49.330 172.570 49.470 172.770 ;
        RECT 53.380 172.710 53.700 172.970 ;
        RECT 53.840 172.910 54.160 172.970 ;
        RECT 54.360 172.910 54.650 172.955 ;
        RECT 53.840 172.770 54.650 172.910 ;
        RECT 53.840 172.710 54.160 172.770 ;
        RECT 54.360 172.725 54.650 172.770 ;
        RECT 56.600 172.710 56.920 172.970 ;
        RECT 57.060 172.910 57.380 172.970 ;
        RECT 57.995 172.910 58.285 172.955 ;
        RECT 57.060 172.770 58.285 172.910 ;
        RECT 57.060 172.710 57.380 172.770 ;
        RECT 57.995 172.725 58.285 172.770 ;
        RECT 57.535 172.570 57.825 172.615 ;
        RECT 49.330 172.430 57.825 172.570 ;
        RECT 57.535 172.385 57.825 172.430 ;
        RECT 58.440 172.370 58.760 172.630 ;
        RECT 69.480 172.370 69.800 172.630 ;
        RECT 71.320 172.370 71.640 172.630 ;
        RECT 72.790 172.570 72.930 173.050 ;
        RECT 77.850 172.570 77.990 173.110 ;
        RECT 78.190 173.065 78.480 173.110 ;
        RECT 80.520 173.250 80.840 173.310 ;
        RECT 81.455 173.250 81.745 173.295 ;
        RECT 84.750 173.250 84.890 173.450 ;
        RECT 87.435 173.405 87.725 173.450 ;
        RECT 80.520 173.110 84.890 173.250 ;
        RECT 80.520 173.050 80.840 173.110 ;
        RECT 81.455 173.065 81.745 173.110 ;
        RECT 86.960 173.050 87.280 173.310 ;
        RECT 87.970 173.295 88.110 173.790 ;
        RECT 98.090 173.790 112.565 173.930 ;
        RECT 98.090 173.635 98.230 173.790 ;
        RECT 112.275 173.745 112.565 173.790 ;
        RECT 98.015 173.405 98.305 173.635 ;
        RECT 98.920 173.590 99.240 173.650 ;
        RECT 103.075 173.590 103.365 173.635 ;
        RECT 98.920 173.450 103.365 173.590 ;
        RECT 98.920 173.390 99.240 173.450 ;
        RECT 103.075 173.405 103.365 173.450 ;
        RECT 107.200 173.590 107.520 173.650 ;
        RECT 112.810 173.590 112.950 174.130 ;
        RECT 113.655 174.085 113.945 174.130 ;
        RECT 115.480 174.070 115.800 174.330 ;
        RECT 117.780 174.270 118.100 174.330 ;
        RECT 116.950 174.130 118.100 174.270 ;
        RECT 115.020 173.930 115.340 173.990 ;
        RECT 116.950 173.930 117.090 174.130 ;
        RECT 117.780 174.070 118.100 174.130 ;
        RECT 121.015 174.270 121.305 174.315 ;
        RECT 123.300 174.270 123.620 174.330 ;
        RECT 121.015 174.130 123.620 174.270 ;
        RECT 121.015 174.085 121.305 174.130 ;
        RECT 123.300 174.070 123.620 174.130 ;
        RECT 128.835 174.270 129.125 174.315 ;
        RECT 131.580 174.270 131.900 174.330 ;
        RECT 128.835 174.130 131.900 174.270 ;
        RECT 128.835 174.085 129.125 174.130 ;
        RECT 131.580 174.070 131.900 174.130 ;
        RECT 132.040 174.270 132.360 174.330 ;
        RECT 132.975 174.270 133.265 174.315 ;
        RECT 132.040 174.130 133.265 174.270 ;
        RECT 132.040 174.070 132.360 174.130 ;
        RECT 132.975 174.085 133.265 174.130 ;
        RECT 114.190 173.790 115.340 173.930 ;
        RECT 114.190 173.635 114.330 173.790 ;
        RECT 115.020 173.730 115.340 173.790 ;
        RECT 115.570 173.790 117.090 173.930 ;
        RECT 107.200 173.450 112.950 173.590 ;
        RECT 107.200 173.390 107.520 173.450 ;
        RECT 87.895 173.065 88.185 173.295 ;
        RECT 97.095 173.250 97.385 173.295 ;
        RECT 98.460 173.250 98.780 173.310 ;
        RECT 97.095 173.110 98.780 173.250 ;
        RECT 97.095 173.065 97.385 173.110 ;
        RECT 98.460 173.050 98.780 173.110 ;
        RECT 99.380 173.250 99.700 173.310 ;
        RECT 109.130 173.295 109.270 173.450 ;
        RECT 114.115 173.405 114.405 173.635 ;
        RECT 102.155 173.250 102.445 173.295 ;
        RECT 99.380 173.110 102.445 173.250 ;
        RECT 99.380 173.050 99.700 173.110 ;
        RECT 102.155 173.065 102.445 173.110 ;
        RECT 109.055 173.065 109.345 173.295 ;
        RECT 109.515 173.065 109.805 173.295 ;
        RECT 84.675 172.910 84.965 172.955 ;
        RECT 107.660 172.910 107.980 172.970 ;
        RECT 109.590 172.910 109.730 173.065 ;
        RECT 110.420 173.050 110.740 173.310 ;
        RECT 111.340 173.050 111.660 173.310 ;
        RECT 111.815 173.065 112.105 173.295 ;
        RECT 84.675 172.770 88.110 172.910 ;
        RECT 84.675 172.725 84.965 172.770 ;
        RECT 87.970 172.630 88.110 172.770 ;
        RECT 107.660 172.770 109.730 172.910 ;
        RECT 111.890 172.910 112.030 173.065 ;
        RECT 112.720 173.050 113.040 173.310 ;
        RECT 113.640 173.050 113.960 173.310 ;
        RECT 115.020 173.250 115.340 173.310 ;
        RECT 115.570 173.250 115.710 173.790 ;
        RECT 116.950 173.590 117.090 173.790 ;
        RECT 118.700 173.930 119.020 173.990 ;
        RECT 120.080 173.930 120.400 173.990 ;
        RECT 118.700 173.790 120.400 173.930 ;
        RECT 118.700 173.730 119.020 173.790 ;
        RECT 120.080 173.730 120.400 173.790 ;
        RECT 134.380 173.930 134.670 173.975 ;
        RECT 136.480 173.930 136.770 173.975 ;
        RECT 138.050 173.930 138.340 173.975 ;
        RECT 134.380 173.790 138.340 173.930 ;
        RECT 134.380 173.745 134.670 173.790 ;
        RECT 136.480 173.745 136.770 173.790 ;
        RECT 138.050 173.745 138.340 173.790 ;
        RECT 117.795 173.590 118.085 173.635 ;
        RECT 116.950 173.450 118.085 173.590 ;
        RECT 117.795 173.405 118.085 173.450 ;
        RECT 119.635 173.590 119.925 173.635 ;
        RECT 129.755 173.590 130.045 173.635 ;
        RECT 119.635 173.450 130.045 173.590 ;
        RECT 119.635 173.405 119.925 173.450 ;
        RECT 129.755 173.405 130.045 173.450 ;
        RECT 130.660 173.590 130.980 173.650 ;
        RECT 133.895 173.590 134.185 173.635 ;
        RECT 130.660 173.450 134.185 173.590 ;
        RECT 130.660 173.390 130.980 173.450 ;
        RECT 133.895 173.405 134.185 173.450 ;
        RECT 134.775 173.590 135.065 173.635 ;
        RECT 135.965 173.590 136.255 173.635 ;
        RECT 138.485 173.590 138.775 173.635 ;
        RECT 134.775 173.450 138.775 173.590 ;
        RECT 134.775 173.405 135.065 173.450 ;
        RECT 135.965 173.405 136.255 173.450 ;
        RECT 138.485 173.405 138.775 173.450 ;
        RECT 115.020 173.110 115.710 173.250 ;
        RECT 115.020 173.050 115.340 173.110 ;
        RECT 115.940 173.050 116.260 173.310 ;
        RECT 116.860 173.050 117.180 173.310 ;
        RECT 117.335 173.260 117.625 173.295 ;
        RECT 118.240 173.260 118.560 173.310 ;
        RECT 117.335 173.120 118.560 173.260 ;
        RECT 117.335 173.065 117.625 173.120 ;
        RECT 118.240 173.050 118.560 173.120 ;
        RECT 118.700 173.050 119.020 173.310 ;
        RECT 120.095 173.250 120.385 173.295 ;
        RECT 120.540 173.250 120.860 173.310 ;
        RECT 120.095 173.110 120.860 173.250 ;
        RECT 120.095 173.065 120.385 173.110 ;
        RECT 120.540 173.050 120.860 173.110 ;
        RECT 121.015 173.250 121.305 173.295 ;
        RECT 124.235 173.250 124.525 173.295 ;
        RECT 126.075 173.250 126.365 173.295 ;
        RECT 121.015 173.110 123.530 173.250 ;
        RECT 121.015 173.065 121.305 173.110 ;
        RECT 123.390 172.970 123.530 173.110 ;
        RECT 124.235 173.110 126.365 173.250 ;
        RECT 124.235 173.065 124.525 173.110 ;
        RECT 126.075 173.065 126.365 173.110 ;
        RECT 126.520 173.250 126.840 173.310 ;
        RECT 126.995 173.250 127.285 173.295 ;
        RECT 126.520 173.110 127.285 173.250 ;
        RECT 126.520 173.050 126.840 173.110 ;
        RECT 126.995 173.065 127.285 173.110 ;
        RECT 127.900 173.050 128.220 173.310 ;
        RECT 131.135 173.250 131.425 173.295 ;
        RECT 138.020 173.250 138.340 173.310 ;
        RECT 131.135 173.110 138.340 173.250 ;
        RECT 131.135 173.065 131.425 173.110 ;
        RECT 138.020 173.050 138.340 173.110 ;
        RECT 115.480 172.910 115.800 172.970 ;
        RECT 119.620 172.910 119.940 172.970 ;
        RECT 122.395 172.910 122.685 172.955 ;
        RECT 111.890 172.770 115.800 172.910 ;
        RECT 107.660 172.710 107.980 172.770 ;
        RECT 115.480 172.710 115.800 172.770 ;
        RECT 119.275 172.770 122.685 172.910 ;
        RECT 72.790 172.430 77.990 172.570 ;
        RECT 87.880 172.370 88.200 172.630 ;
        RECT 95.240 172.370 95.560 172.630 ;
        RECT 97.555 172.570 97.845 172.615 ;
        RECT 99.395 172.570 99.685 172.615 ;
        RECT 97.555 172.430 99.685 172.570 ;
        RECT 97.555 172.385 97.845 172.430 ;
        RECT 99.395 172.385 99.685 172.430 ;
        RECT 105.360 172.570 105.680 172.630 ;
        RECT 106.295 172.570 106.585 172.615 ;
        RECT 105.360 172.430 106.585 172.570 ;
        RECT 105.360 172.370 105.680 172.430 ;
        RECT 106.295 172.385 106.585 172.430 ;
        RECT 109.040 172.570 109.360 172.630 ;
        RECT 109.515 172.570 109.805 172.615 ;
        RECT 109.040 172.430 109.805 172.570 ;
        RECT 109.040 172.370 109.360 172.430 ;
        RECT 109.515 172.385 109.805 172.430 ;
        RECT 110.880 172.570 111.200 172.630 ;
        RECT 119.275 172.570 119.415 172.770 ;
        RECT 119.620 172.710 119.940 172.770 ;
        RECT 122.395 172.725 122.685 172.770 ;
        RECT 123.300 172.910 123.620 172.970 ;
        RECT 124.680 172.910 125.000 172.970 ;
        RECT 135.260 172.955 135.580 172.970 ;
        RECT 123.300 172.770 125.000 172.910 ;
        RECT 123.300 172.710 123.620 172.770 ;
        RECT 124.680 172.710 125.000 172.770 ;
        RECT 127.455 172.725 127.745 172.955 ;
        RECT 135.230 172.725 135.580 172.955 ;
        RECT 110.880 172.430 119.415 172.570 ;
        RECT 110.880 172.370 111.200 172.430 ;
        RECT 121.920 172.370 122.240 172.630 ;
        RECT 125.140 172.570 125.460 172.630 ;
        RECT 127.530 172.570 127.670 172.725 ;
        RECT 135.260 172.710 135.580 172.725 ;
        RECT 125.140 172.430 127.670 172.570 ;
        RECT 130.200 172.570 130.520 172.630 ;
        RECT 130.675 172.570 130.965 172.615 ;
        RECT 130.200 172.430 130.965 172.570 ;
        RECT 125.140 172.370 125.460 172.430 ;
        RECT 130.200 172.370 130.520 172.430 ;
        RECT 130.675 172.385 130.965 172.430 ;
        RECT 140.780 172.370 141.100 172.630 ;
        RECT 17.430 171.750 143.010 172.230 ;
        RECT 22.115 171.550 22.405 171.595 ;
        RECT 22.560 171.550 22.880 171.610 ;
        RECT 22.115 171.410 22.880 171.550 ;
        RECT 22.115 171.365 22.405 171.410 ;
        RECT 22.560 171.350 22.880 171.410 ;
        RECT 23.480 171.350 23.800 171.610 ;
        RECT 23.940 171.550 24.260 171.610 ;
        RECT 48.780 171.550 49.100 171.610 ;
        RECT 58.440 171.550 58.760 171.610 ;
        RECT 74.540 171.550 74.860 171.610 ;
        RECT 76.380 171.550 76.700 171.610 ;
        RECT 76.855 171.550 77.145 171.595 ;
        RECT 23.940 171.410 38.890 171.550 ;
        RECT 23.940 171.350 24.260 171.410 ;
        RECT 25.780 171.210 26.100 171.270 ;
        RECT 26.555 171.210 26.845 171.255 ;
        RECT 25.780 171.070 26.845 171.210 ;
        RECT 25.780 171.010 26.100 171.070 ;
        RECT 26.555 171.025 26.845 171.070 ;
        RECT 27.635 171.210 27.925 171.255 ;
        RECT 28.080 171.210 28.400 171.270 ;
        RECT 29.015 171.210 29.305 171.255 ;
        RECT 27.635 171.070 29.305 171.210 ;
        RECT 27.635 171.025 27.925 171.070 ;
        RECT 28.080 171.010 28.400 171.070 ;
        RECT 29.015 171.025 29.305 171.070 ;
        RECT 30.840 171.010 31.160 171.270 ;
        RECT 32.220 171.210 32.540 171.270 ;
        RECT 38.750 171.255 38.890 171.410 ;
        RECT 48.780 171.410 60.970 171.550 ;
        RECT 48.780 171.350 49.100 171.410 ;
        RECT 58.440 171.350 58.760 171.410 ;
        RECT 38.675 171.210 38.965 171.255 ;
        RECT 53.380 171.210 53.700 171.270 ;
        RECT 55.235 171.210 55.525 171.255 ;
        RECT 57.060 171.210 57.380 171.270 ;
        RECT 32.220 171.070 36.130 171.210 ;
        RECT 32.220 171.010 32.540 171.070 ;
        RECT 20.735 170.685 21.025 170.915 ;
        RECT 20.810 170.190 20.950 170.685 ;
        RECT 21.640 170.670 21.960 170.930 ;
        RECT 23.955 170.870 24.245 170.915 ;
        RECT 24.400 170.870 24.720 170.930 ;
        RECT 23.955 170.730 24.720 170.870 ;
        RECT 23.955 170.685 24.245 170.730 ;
        RECT 24.400 170.670 24.720 170.730 ;
        RECT 25.320 170.670 25.640 170.930 ;
        RECT 29.475 170.685 29.765 170.915 ;
        RECT 21.195 170.530 21.485 170.575 ;
        RECT 22.910 170.530 23.200 170.575 ;
        RECT 21.195 170.390 23.200 170.530 ;
        RECT 21.195 170.345 21.485 170.390 ;
        RECT 22.910 170.345 23.200 170.390 ;
        RECT 28.095 170.530 28.385 170.575 ;
        RECT 29.000 170.530 29.320 170.590 ;
        RECT 28.095 170.390 29.320 170.530 ;
        RECT 28.095 170.345 28.385 170.390 ;
        RECT 29.000 170.330 29.320 170.390 ;
        RECT 25.795 170.190 26.085 170.235 ;
        RECT 26.240 170.190 26.560 170.250 ;
        RECT 20.810 170.050 26.560 170.190 ;
        RECT 25.795 170.005 26.085 170.050 ;
        RECT 26.240 169.990 26.560 170.050 ;
        RECT 23.020 169.850 23.340 169.910 ;
        RECT 26.715 169.850 27.005 169.895 ;
        RECT 29.550 169.850 29.690 170.685 ;
        RECT 29.920 170.670 30.240 170.930 ;
        RECT 34.075 170.870 34.365 170.915 ;
        RECT 34.520 170.870 34.840 170.930 ;
        RECT 34.075 170.730 34.840 170.870 ;
        RECT 34.075 170.685 34.365 170.730 ;
        RECT 34.520 170.670 34.840 170.730 ;
        RECT 34.980 170.670 35.300 170.930 ;
        RECT 35.440 170.670 35.760 170.930 ;
        RECT 35.990 170.915 36.130 171.070 ;
        RECT 38.675 171.070 43.950 171.210 ;
        RECT 38.675 171.025 38.965 171.070 ;
        RECT 43.810 170.915 43.950 171.070 ;
        RECT 53.380 171.070 57.380 171.210 ;
        RECT 53.380 171.010 53.700 171.070 ;
        RECT 55.235 171.025 55.525 171.070 ;
        RECT 57.060 171.010 57.380 171.070 ;
        RECT 57.520 171.210 57.840 171.270 ;
        RECT 57.520 171.070 60.050 171.210 ;
        RECT 57.520 171.010 57.840 171.070 ;
        RECT 59.910 170.915 60.050 171.070 ;
        RECT 60.830 170.915 60.970 171.410 ;
        RECT 74.540 171.410 76.150 171.550 ;
        RECT 74.540 171.350 74.860 171.410 ;
        RECT 74.080 171.210 74.400 171.270 ;
        RECT 75.000 171.255 75.320 171.270 ;
        RECT 75.000 171.210 75.350 171.255 ;
        RECT 76.010 171.210 76.150 171.410 ;
        RECT 76.380 171.410 77.145 171.550 ;
        RECT 76.380 171.350 76.700 171.410 ;
        RECT 76.855 171.365 77.145 171.410 ;
        RECT 78.695 171.550 78.985 171.595 ;
        RECT 80.980 171.550 81.300 171.610 ;
        RECT 78.695 171.410 81.300 171.550 ;
        RECT 78.695 171.365 78.985 171.410 ;
        RECT 80.980 171.350 81.300 171.410 ;
        RECT 81.900 171.350 82.220 171.610 ;
        RECT 87.880 171.350 88.200 171.610 ;
        RECT 90.195 171.550 90.485 171.595 ;
        RECT 95.255 171.550 95.545 171.595 ;
        RECT 98.920 171.550 99.240 171.610 ;
        RECT 90.195 171.410 99.240 171.550 ;
        RECT 90.195 171.365 90.485 171.410 ;
        RECT 95.255 171.365 95.545 171.410 ;
        RECT 98.920 171.350 99.240 171.410 ;
        RECT 102.615 171.365 102.905 171.595 ;
        RECT 110.880 171.550 111.200 171.610 ;
        RECT 103.610 171.410 111.200 171.550 ;
        RECT 80.535 171.210 80.825 171.255 ;
        RECT 74.080 171.070 74.770 171.210 ;
        RECT 74.080 171.010 74.400 171.070 ;
        RECT 35.915 170.685 36.205 170.915 ;
        RECT 42.815 170.685 43.105 170.915 ;
        RECT 43.735 170.685 44.025 170.915 ;
        RECT 59.375 170.685 59.665 170.915 ;
        RECT 59.835 170.685 60.125 170.915 ;
        RECT 60.755 170.685 61.045 170.915 ;
        RECT 74.630 170.870 74.770 171.070 ;
        RECT 75.000 171.070 75.515 171.210 ;
        RECT 76.010 171.070 80.825 171.210 ;
        RECT 75.000 171.025 75.350 171.070 ;
        RECT 80.535 171.025 80.825 171.070 ;
        RECT 81.455 171.210 81.745 171.255 ;
        RECT 82.360 171.210 82.680 171.270 ;
        RECT 86.960 171.210 87.280 171.270 ;
        RECT 81.455 171.070 82.680 171.210 ;
        RECT 81.455 171.025 81.745 171.070 ;
        RECT 75.000 171.010 75.320 171.025 ;
        RECT 82.360 171.010 82.680 171.070 ;
        RECT 82.910 171.070 87.280 171.210 ;
        RECT 74.630 170.730 77.070 170.870 ;
        RECT 34.610 170.530 34.750 170.670 ;
        RECT 37.280 170.530 37.600 170.590 ;
        RECT 34.610 170.390 37.600 170.530 ;
        RECT 42.890 170.530 43.030 170.685 ;
        RECT 59.450 170.530 59.590 170.685 ;
        RECT 64.420 170.530 64.740 170.590 ;
        RECT 42.890 170.390 64.740 170.530 ;
        RECT 37.280 170.330 37.600 170.390 ;
        RECT 64.420 170.330 64.740 170.390 ;
        RECT 71.805 170.530 72.095 170.575 ;
        RECT 74.325 170.530 74.615 170.575 ;
        RECT 75.515 170.530 75.805 170.575 ;
        RECT 71.805 170.390 75.805 170.530 ;
        RECT 71.805 170.345 72.095 170.390 ;
        RECT 74.325 170.345 74.615 170.390 ;
        RECT 75.515 170.345 75.805 170.390 ;
        RECT 76.380 170.330 76.700 170.590 ;
        RECT 76.930 170.530 77.070 170.730 ;
        RECT 77.760 170.670 78.080 170.930 ;
        RECT 79.140 170.670 79.460 170.930 ;
        RECT 79.600 170.870 79.920 170.930 ;
        RECT 82.910 170.915 83.050 171.070 ;
        RECT 86.960 171.010 87.280 171.070 ;
        RECT 100.930 171.210 101.220 171.255 ;
        RECT 102.690 171.210 102.830 171.365 ;
        RECT 100.930 171.070 102.830 171.210 ;
        RECT 100.930 171.025 101.220 171.070 ;
        RECT 82.835 170.870 83.125 170.915 ;
        RECT 79.600 170.730 83.125 170.870 ;
        RECT 79.600 170.670 79.920 170.730 ;
        RECT 82.835 170.685 83.125 170.730 ;
        RECT 83.740 170.670 84.060 170.930 ;
        RECT 88.800 170.870 89.120 170.930 ;
        RECT 89.735 170.870 90.025 170.915 ;
        RECT 98.460 170.870 98.780 170.930 ;
        RECT 103.610 170.915 103.750 171.410 ;
        RECT 110.880 171.350 111.200 171.410 ;
        RECT 115.020 171.550 115.340 171.610 ;
        RECT 116.875 171.550 117.165 171.595 ;
        RECT 115.020 171.410 117.165 171.550 ;
        RECT 115.020 171.350 115.340 171.410 ;
        RECT 116.875 171.365 117.165 171.410 ;
        RECT 118.700 171.350 119.020 171.610 ;
        RECT 126.520 171.550 126.840 171.610 ;
        RECT 126.150 171.410 126.840 171.550 ;
        RECT 104.455 171.210 104.745 171.255 ;
        RECT 105.835 171.210 106.125 171.255 ;
        RECT 109.040 171.210 109.360 171.270 ;
        RECT 122.840 171.210 123.160 171.270 ;
        RECT 126.150 171.255 126.290 171.410 ;
        RECT 126.520 171.350 126.840 171.410 ;
        RECT 127.440 171.550 127.760 171.610 ;
        RECT 130.200 171.550 130.520 171.610 ;
        RECT 131.135 171.550 131.425 171.595 ;
        RECT 127.440 171.410 129.970 171.550 ;
        RECT 127.440 171.350 127.760 171.410 ;
        RECT 104.455 171.070 106.125 171.210 ;
        RECT 104.455 171.025 104.745 171.070 ;
        RECT 105.835 171.025 106.125 171.070 ;
        RECT 106.370 171.070 109.360 171.210 ;
        RECT 88.800 170.730 90.025 170.870 ;
        RECT 88.800 170.670 89.120 170.730 ;
        RECT 89.735 170.685 90.025 170.730 ;
        RECT 91.190 170.730 98.780 170.870 ;
        RECT 83.830 170.530 83.970 170.670 ;
        RECT 76.930 170.390 83.970 170.530 ;
        RECT 84.200 170.330 84.520 170.590 ;
        RECT 91.190 170.575 91.330 170.730 ;
        RECT 98.460 170.670 98.780 170.730 ;
        RECT 103.535 170.685 103.825 170.915 ;
        RECT 103.995 170.685 104.285 170.915 ;
        RECT 91.115 170.345 91.405 170.575 ;
        RECT 97.565 170.530 97.855 170.575 ;
        RECT 100.085 170.530 100.375 170.575 ;
        RECT 101.275 170.530 101.565 170.575 ;
        RECT 97.565 170.390 101.565 170.530 ;
        RECT 97.565 170.345 97.855 170.390 ;
        RECT 100.085 170.345 100.375 170.390 ;
        RECT 101.275 170.345 101.565 170.390 ;
        RECT 102.140 170.330 102.460 170.590 ;
        RECT 104.070 170.530 104.210 170.685 ;
        RECT 105.360 170.670 105.680 170.930 ;
        RECT 106.370 170.530 106.510 171.070 ;
        RECT 109.040 171.010 109.360 171.070 ;
        RECT 118.790 171.070 123.160 171.210 ;
        RECT 106.755 170.685 107.045 170.915 ;
        RECT 107.215 170.685 107.505 170.915 ;
        RECT 104.070 170.390 106.510 170.530 ;
        RECT 72.240 170.190 72.530 170.235 ;
        RECT 73.810 170.190 74.100 170.235 ;
        RECT 75.910 170.190 76.200 170.235 ;
        RECT 78.680 170.190 79.000 170.250 ;
        RECT 72.240 170.050 76.200 170.190 ;
        RECT 72.240 170.005 72.530 170.050 ;
        RECT 73.810 170.005 74.100 170.050 ;
        RECT 75.910 170.005 76.200 170.050 ;
        RECT 76.470 170.050 79.000 170.190 ;
        RECT 23.020 169.710 29.690 169.850 ;
        RECT 37.295 169.850 37.585 169.895 ;
        RECT 37.740 169.850 38.060 169.910 ;
        RECT 37.295 169.710 38.060 169.850 ;
        RECT 23.020 169.650 23.340 169.710 ;
        RECT 26.715 169.665 27.005 169.710 ;
        RECT 37.295 169.665 37.585 169.710 ;
        RECT 37.740 169.650 38.060 169.710 ;
        RECT 55.220 169.850 55.540 169.910 ;
        RECT 59.835 169.850 60.125 169.895 ;
        RECT 55.220 169.710 60.125 169.850 ;
        RECT 55.220 169.650 55.540 169.710 ;
        RECT 59.835 169.665 60.125 169.710 ;
        RECT 69.495 169.850 69.785 169.895 ;
        RECT 74.540 169.850 74.860 169.910 ;
        RECT 76.470 169.850 76.610 170.050 ;
        RECT 78.680 169.990 79.000 170.050 ;
        RECT 87.435 170.190 87.725 170.235 ;
        RECT 88.340 170.190 88.660 170.250 ;
        RECT 87.435 170.050 88.660 170.190 ;
        RECT 87.435 170.005 87.725 170.050 ;
        RECT 88.340 169.990 88.660 170.050 ;
        RECT 98.000 170.190 98.290 170.235 ;
        RECT 99.570 170.190 99.860 170.235 ;
        RECT 101.670 170.190 101.960 170.235 ;
        RECT 98.000 170.050 101.960 170.190 ;
        RECT 106.830 170.190 106.970 170.685 ;
        RECT 107.290 170.530 107.430 170.685 ;
        RECT 108.120 170.670 108.440 170.930 ;
        RECT 108.580 170.870 108.900 170.930 ;
        RECT 110.420 170.870 110.740 170.930 ;
        RECT 108.580 170.730 110.740 170.870 ;
        RECT 108.580 170.670 108.900 170.730 ;
        RECT 110.420 170.670 110.740 170.730 ;
        RECT 112.720 170.870 113.040 170.930 ;
        RECT 114.575 170.870 114.865 170.915 ;
        RECT 112.720 170.730 114.865 170.870 ;
        RECT 112.720 170.670 113.040 170.730 ;
        RECT 114.575 170.685 114.865 170.730 ;
        RECT 115.035 170.685 115.325 170.915 ;
        RECT 116.415 170.870 116.705 170.915 ;
        RECT 116.415 170.730 117.090 170.870 ;
        RECT 116.415 170.685 116.705 170.730 ;
        RECT 111.340 170.530 111.660 170.590 ;
        RECT 107.290 170.390 111.660 170.530 ;
        RECT 111.340 170.330 111.660 170.390 ;
        RECT 110.880 170.190 111.200 170.250 ;
        RECT 106.830 170.050 111.200 170.190 ;
        RECT 98.000 170.005 98.290 170.050 ;
        RECT 99.570 170.005 99.860 170.050 ;
        RECT 101.670 170.005 101.960 170.050 ;
        RECT 110.880 169.990 111.200 170.050 ;
        RECT 114.560 170.190 114.880 170.250 ;
        RECT 115.110 170.190 115.250 170.685 ;
        RECT 115.480 170.530 115.800 170.590 ;
        RECT 115.955 170.530 116.245 170.575 ;
        RECT 115.480 170.390 116.245 170.530 ;
        RECT 115.480 170.330 115.800 170.390 ;
        RECT 115.955 170.345 116.245 170.390 ;
        RECT 114.560 170.050 115.250 170.190 ;
        RECT 116.950 170.190 117.090 170.730 ;
        RECT 117.795 170.860 118.085 170.915 ;
        RECT 118.790 170.870 118.930 171.070 ;
        RECT 122.840 171.010 123.160 171.070 ;
        RECT 126.075 171.210 126.365 171.255 ;
        RECT 129.295 171.210 129.585 171.255 ;
        RECT 126.075 171.070 129.585 171.210 ;
        RECT 129.830 171.210 129.970 171.410 ;
        RECT 130.200 171.410 131.425 171.550 ;
        RECT 130.200 171.350 130.520 171.410 ;
        RECT 131.135 171.365 131.425 171.410 ;
        RECT 135.260 171.350 135.580 171.610 ;
        RECT 136.655 171.550 136.945 171.595 ;
        RECT 139.860 171.550 140.180 171.610 ;
        RECT 136.655 171.410 140.180 171.550 ;
        RECT 136.655 171.365 136.945 171.410 ;
        RECT 139.860 171.350 140.180 171.410 ;
        RECT 133.435 171.210 133.725 171.255 ;
        RECT 137.115 171.210 137.405 171.255 ;
        RECT 129.830 171.070 130.430 171.210 ;
        RECT 126.075 171.025 126.365 171.070 ;
        RECT 129.295 171.025 129.585 171.070 ;
        RECT 118.330 170.860 118.930 170.870 ;
        RECT 117.795 170.730 118.930 170.860 ;
        RECT 119.175 170.870 119.465 170.915 ;
        RECT 120.080 170.870 120.400 170.930 ;
        RECT 119.175 170.730 120.400 170.870 ;
        RECT 117.795 170.720 118.470 170.730 ;
        RECT 117.795 170.685 118.085 170.720 ;
        RECT 119.175 170.685 119.465 170.730 ;
        RECT 120.080 170.670 120.400 170.730 ;
        RECT 121.015 170.870 121.305 170.915 ;
        RECT 121.460 170.870 121.780 170.930 ;
        RECT 121.015 170.730 121.780 170.870 ;
        RECT 121.015 170.685 121.305 170.730 ;
        RECT 121.460 170.670 121.780 170.730 ;
        RECT 121.935 170.685 122.225 170.915 ;
        RECT 117.320 170.530 117.640 170.590 ;
        RECT 122.010 170.530 122.150 170.685 ;
        RECT 122.380 170.670 122.700 170.930 ;
        RECT 123.775 170.685 124.065 170.915 ;
        RECT 124.220 170.870 124.540 170.930 ;
        RECT 125.155 170.870 125.445 170.915 ;
        RECT 126.535 170.870 126.825 170.915 ;
        RECT 124.220 170.730 125.445 170.870 ;
        RECT 117.320 170.390 122.150 170.530 ;
        RECT 117.320 170.330 117.640 170.390 ;
        RECT 122.840 170.330 123.160 170.590 ;
        RECT 118.240 170.190 118.560 170.250 ;
        RECT 121.920 170.190 122.240 170.250 ;
        RECT 123.850 170.190 123.990 170.685 ;
        RECT 124.220 170.670 124.540 170.730 ;
        RECT 125.155 170.685 125.445 170.730 ;
        RECT 126.150 170.730 126.825 170.870 ;
        RECT 126.150 170.590 126.290 170.730 ;
        RECT 126.535 170.685 126.825 170.730 ;
        RECT 126.995 170.870 127.285 170.915 ;
        RECT 127.440 170.870 127.760 170.930 ;
        RECT 126.995 170.730 127.760 170.870 ;
        RECT 126.995 170.685 127.285 170.730 ;
        RECT 127.440 170.670 127.760 170.730 ;
        RECT 128.360 170.670 128.680 170.930 ;
        RECT 129.740 170.670 130.060 170.930 ;
        RECT 130.290 170.915 130.430 171.070 ;
        RECT 133.435 171.070 137.405 171.210 ;
        RECT 133.435 171.025 133.725 171.070 ;
        RECT 137.115 171.025 137.405 171.070 ;
        RECT 130.215 170.685 130.505 170.915 ;
        RECT 135.735 170.870 136.025 170.915 ;
        RECT 140.335 170.870 140.625 170.915 ;
        RECT 140.780 170.870 141.100 170.930 ;
        RECT 135.735 170.730 141.100 170.870 ;
        RECT 135.735 170.685 136.025 170.730 ;
        RECT 140.335 170.685 140.625 170.730 ;
        RECT 140.780 170.670 141.100 170.730 ;
        RECT 126.060 170.330 126.380 170.590 ;
        RECT 132.055 170.530 132.345 170.575 ;
        RECT 127.530 170.390 132.345 170.530 ;
        RECT 116.950 170.050 123.990 170.190 ;
        RECT 124.695 170.190 124.985 170.235 ;
        RECT 127.530 170.190 127.670 170.390 ;
        RECT 132.055 170.345 132.345 170.390 ;
        RECT 132.975 170.345 133.265 170.575 ;
        RECT 124.695 170.050 127.670 170.190 ;
        RECT 127.915 170.190 128.205 170.235 ;
        RECT 133.050 170.190 133.190 170.345 ;
        RECT 127.915 170.050 133.190 170.190 ;
        RECT 114.560 169.990 114.880 170.050 ;
        RECT 69.495 169.710 76.610 169.850 ;
        RECT 76.840 169.850 77.160 169.910 ;
        RECT 79.140 169.850 79.460 169.910 ;
        RECT 79.615 169.850 79.905 169.895 ;
        RECT 76.840 169.710 79.905 169.850 ;
        RECT 69.495 169.665 69.785 169.710 ;
        RECT 74.540 169.650 74.860 169.710 ;
        RECT 76.840 169.650 77.160 169.710 ;
        RECT 79.140 169.650 79.460 169.710 ;
        RECT 79.615 169.665 79.905 169.710 ;
        RECT 83.280 169.850 83.600 169.910 ;
        RECT 87.880 169.850 88.200 169.910 ;
        RECT 83.280 169.710 88.200 169.850 ;
        RECT 83.280 169.650 83.600 169.710 ;
        RECT 87.880 169.650 88.200 169.710 ;
        RECT 113.640 169.650 113.960 169.910 ;
        RECT 115.110 169.850 115.250 170.050 ;
        RECT 118.240 169.990 118.560 170.050 ;
        RECT 121.920 169.990 122.240 170.050 ;
        RECT 124.695 170.005 124.985 170.050 ;
        RECT 127.915 170.005 128.205 170.050 ;
        RECT 127.440 169.850 127.760 169.910 ;
        RECT 115.110 169.710 127.760 169.850 ;
        RECT 127.440 169.650 127.760 169.710 ;
        RECT 17.430 169.030 143.010 169.510 ;
        RECT 21.640 168.830 21.960 168.890 ;
        RECT 26.715 168.830 27.005 168.875 ;
        RECT 21.640 168.690 27.005 168.830 ;
        RECT 21.640 168.630 21.960 168.690 ;
        RECT 26.715 168.645 27.005 168.690 ;
        RECT 28.080 168.830 28.400 168.890 ;
        RECT 30.840 168.830 31.160 168.890 ;
        RECT 33.155 168.830 33.445 168.875 ;
        RECT 28.080 168.690 33.445 168.830 ;
        RECT 28.080 168.630 28.400 168.690 ;
        RECT 30.840 168.630 31.160 168.690 ;
        RECT 33.155 168.645 33.445 168.690 ;
        RECT 43.735 168.830 44.025 168.875 ;
        RECT 46.020 168.830 46.340 168.890 ;
        RECT 43.735 168.690 46.340 168.830 ;
        RECT 43.735 168.645 44.025 168.690 ;
        RECT 46.020 168.630 46.340 168.690 ;
        RECT 53.840 168.630 54.160 168.890 ;
        RECT 82.835 168.830 83.125 168.875 ;
        RECT 84.200 168.830 84.520 168.890 ;
        RECT 82.835 168.690 84.520 168.830 ;
        RECT 82.835 168.645 83.125 168.690 ;
        RECT 84.200 168.630 84.520 168.690 ;
        RECT 97.095 168.830 97.385 168.875 ;
        RECT 97.540 168.830 97.860 168.890 ;
        RECT 99.380 168.830 99.700 168.890 ;
        RECT 97.095 168.690 99.700 168.830 ;
        RECT 97.095 168.645 97.385 168.690 ;
        RECT 97.540 168.630 97.860 168.690 ;
        RECT 99.380 168.630 99.700 168.690 ;
        RECT 109.040 168.830 109.360 168.890 ;
        RECT 115.940 168.830 116.260 168.890 ;
        RECT 121.460 168.830 121.780 168.890 ;
        RECT 109.040 168.690 115.710 168.830 ;
        RECT 109.040 168.630 109.360 168.690 ;
        RECT 34.995 168.305 35.285 168.535 ;
        RECT 53.380 168.490 53.700 168.550 ;
        RECT 54.300 168.490 54.620 168.550 ;
        RECT 52.550 168.350 54.620 168.490 ;
        RECT 29.920 168.150 30.240 168.210 ;
        RECT 25.870 168.010 30.240 168.150 ;
        RECT 25.870 167.870 26.010 168.010 ;
        RECT 29.920 167.950 30.240 168.010 ;
        RECT 32.220 168.150 32.540 168.210 ;
        RECT 33.615 168.150 33.905 168.195 ;
        RECT 32.220 168.010 33.905 168.150 ;
        RECT 35.070 168.150 35.210 168.305 ;
        RECT 35.070 168.010 38.890 168.150 ;
        RECT 32.220 167.950 32.540 168.010 ;
        RECT 33.615 167.965 33.905 168.010 ;
        RECT 25.335 167.810 25.625 167.855 ;
        RECT 25.780 167.810 26.100 167.870 ;
        RECT 25.335 167.670 26.100 167.810 ;
        RECT 25.335 167.625 25.625 167.670 ;
        RECT 25.780 167.610 26.100 167.670 ;
        RECT 26.715 167.810 27.005 167.855 ;
        RECT 28.080 167.810 28.400 167.870 ;
        RECT 26.715 167.670 28.400 167.810 ;
        RECT 26.715 167.625 27.005 167.670 ;
        RECT 28.080 167.610 28.400 167.670 ;
        RECT 31.300 167.810 31.620 167.870 ;
        RECT 33.155 167.810 33.445 167.855 ;
        RECT 31.300 167.670 33.445 167.810 ;
        RECT 31.300 167.610 31.620 167.670 ;
        RECT 33.155 167.625 33.445 167.670 ;
        RECT 34.980 167.810 35.300 167.870 ;
        RECT 36.375 167.810 36.665 167.855 ;
        RECT 34.980 167.670 36.665 167.810 ;
        RECT 34.980 167.610 35.300 167.670 ;
        RECT 36.375 167.625 36.665 167.670 ;
        RECT 37.280 167.610 37.600 167.870 ;
        RECT 37.740 167.610 38.060 167.870 ;
        RECT 38.750 167.855 38.890 168.010 ;
        RECT 40.130 168.010 44.410 168.150 ;
        RECT 40.130 167.870 40.270 168.010 ;
        RECT 38.675 167.625 38.965 167.855 ;
        RECT 39.135 167.625 39.425 167.855 ;
        RECT 39.595 167.810 39.885 167.855 ;
        RECT 40.040 167.810 40.360 167.870 ;
        RECT 39.595 167.670 40.360 167.810 ;
        RECT 39.595 167.625 39.885 167.670 ;
        RECT 39.210 167.470 39.350 167.625 ;
        RECT 40.040 167.610 40.360 167.670 ;
        RECT 40.500 167.810 40.820 167.870 ;
        RECT 44.270 167.855 44.410 168.010 ;
        RECT 50.620 167.950 50.940 168.210 ;
        RECT 52.550 168.195 52.690 168.350 ;
        RECT 53.380 168.290 53.700 168.350 ;
        RECT 54.300 168.290 54.620 168.350 ;
        RECT 85.580 168.490 85.870 168.535 ;
        RECT 87.150 168.490 87.440 168.535 ;
        RECT 89.250 168.490 89.540 168.535 ;
        RECT 85.580 168.350 89.540 168.490 ;
        RECT 85.580 168.305 85.870 168.350 ;
        RECT 87.150 168.305 87.440 168.350 ;
        RECT 89.250 168.305 89.540 168.350 ;
        RECT 90.680 168.490 90.970 168.535 ;
        RECT 92.780 168.490 93.070 168.535 ;
        RECT 94.350 168.490 94.640 168.535 ;
        RECT 90.680 168.350 94.640 168.490 ;
        RECT 90.680 168.305 90.970 168.350 ;
        RECT 92.780 168.305 93.070 168.350 ;
        RECT 94.350 168.305 94.640 168.350 ;
        RECT 102.140 168.490 102.430 168.535 ;
        RECT 103.710 168.490 104.000 168.535 ;
        RECT 105.810 168.490 106.100 168.535 ;
        RECT 102.140 168.350 106.100 168.490 ;
        RECT 102.140 168.305 102.430 168.350 ;
        RECT 103.710 168.305 104.000 168.350 ;
        RECT 105.810 168.305 106.100 168.350 ;
        RECT 108.580 168.490 108.900 168.550 ;
        RECT 113.195 168.490 113.485 168.535 ;
        RECT 108.580 168.350 113.485 168.490 ;
        RECT 108.580 168.290 108.900 168.350 ;
        RECT 113.195 168.305 113.485 168.350 ;
        RECT 52.475 167.965 52.765 168.195 ;
        RECT 56.600 168.150 56.920 168.210 ;
        RECT 54.390 168.010 56.920 168.150 ;
        RECT 54.390 167.870 54.530 168.010 ;
        RECT 56.600 167.950 56.920 168.010 ;
        RECT 85.145 168.150 85.435 168.195 ;
        RECT 87.665 168.150 87.955 168.195 ;
        RECT 88.855 168.150 89.145 168.195 ;
        RECT 85.145 168.010 89.145 168.150 ;
        RECT 85.145 167.965 85.435 168.010 ;
        RECT 87.665 167.965 87.955 168.010 ;
        RECT 88.855 167.965 89.145 168.010 ;
        RECT 89.735 168.150 90.025 168.195 ;
        RECT 90.180 168.150 90.500 168.210 ;
        RECT 89.735 168.010 90.500 168.150 ;
        RECT 89.735 167.965 90.025 168.010 ;
        RECT 90.180 167.950 90.500 168.010 ;
        RECT 91.075 168.150 91.365 168.195 ;
        RECT 92.265 168.150 92.555 168.195 ;
        RECT 94.785 168.150 95.075 168.195 ;
        RECT 91.075 168.010 95.075 168.150 ;
        RECT 91.075 167.965 91.365 168.010 ;
        RECT 92.265 167.965 92.555 168.010 ;
        RECT 94.785 167.965 95.075 168.010 ;
        RECT 101.705 168.150 101.995 168.195 ;
        RECT 104.225 168.150 104.515 168.195 ;
        RECT 105.415 168.150 105.705 168.195 ;
        RECT 101.705 168.010 105.705 168.150 ;
        RECT 101.705 167.965 101.995 168.010 ;
        RECT 104.225 167.965 104.515 168.010 ;
        RECT 105.415 167.965 105.705 168.010 ;
        RECT 107.200 168.150 107.520 168.210 ;
        RECT 113.655 168.150 113.945 168.195 ;
        RECT 107.200 168.010 113.945 168.150 ;
        RECT 107.200 167.950 107.520 168.010 ;
        RECT 113.655 167.965 113.945 168.010 ;
        RECT 115.035 167.965 115.325 168.195 ;
        RECT 42.355 167.810 42.645 167.855 ;
        RECT 40.500 167.670 42.645 167.810 ;
        RECT 40.500 167.610 40.820 167.670 ;
        RECT 42.355 167.625 42.645 167.670 ;
        RECT 44.195 167.810 44.485 167.855 ;
        RECT 45.575 167.810 45.865 167.855 ;
        RECT 44.195 167.670 45.865 167.810 ;
        RECT 44.195 167.625 44.485 167.670 ;
        RECT 45.575 167.625 45.865 167.670 ;
        RECT 54.300 167.610 54.620 167.870 ;
        RECT 55.220 167.610 55.540 167.870 ;
        RECT 57.060 167.610 57.380 167.870 ;
        RECT 64.420 167.810 64.740 167.870 ;
        RECT 67.180 167.810 67.500 167.870 ;
        RECT 64.420 167.670 67.500 167.810 ;
        RECT 64.420 167.610 64.740 167.670 ;
        RECT 67.180 167.610 67.500 167.670 ;
        RECT 68.575 167.810 68.865 167.855 ;
        RECT 69.480 167.810 69.800 167.870 ;
        RECT 70.415 167.810 70.705 167.855 ;
        RECT 72.240 167.810 72.560 167.870 ;
        RECT 76.380 167.810 76.700 167.870 ;
        RECT 68.575 167.670 76.700 167.810 ;
        RECT 68.575 167.625 68.865 167.670 ;
        RECT 69.480 167.610 69.800 167.670 ;
        RECT 70.415 167.625 70.705 167.670 ;
        RECT 72.240 167.610 72.560 167.670 ;
        RECT 76.380 167.610 76.700 167.670 ;
        RECT 80.535 167.625 80.825 167.855 ;
        RECT 81.455 167.810 81.745 167.855 ;
        RECT 82.360 167.810 82.680 167.870 ;
        RECT 81.455 167.670 82.680 167.810 ;
        RECT 81.455 167.625 81.745 167.670 ;
        RECT 44.655 167.470 44.945 167.515 ;
        RECT 46.020 167.470 46.340 167.530 ;
        RECT 39.210 167.330 46.340 167.470 ;
        RECT 44.655 167.285 44.945 167.330 ;
        RECT 46.020 167.270 46.340 167.330 ;
        RECT 53.060 167.470 53.350 167.515 ;
        RECT 54.775 167.470 55.065 167.515 ;
        RECT 53.060 167.330 55.065 167.470 ;
        RECT 53.060 167.285 53.350 167.330 ;
        RECT 54.775 167.285 55.065 167.330 ;
        RECT 69.020 167.470 69.340 167.530 ;
        RECT 71.320 167.470 71.640 167.530 ;
        RECT 80.610 167.470 80.750 167.625 ;
        RECT 82.360 167.610 82.680 167.670 ;
        RECT 91.530 167.810 91.820 167.855 ;
        RECT 95.240 167.810 95.560 167.870 ;
        RECT 91.530 167.670 95.560 167.810 ;
        RECT 91.530 167.625 91.820 167.670 ;
        RECT 95.240 167.610 95.560 167.670 ;
        RECT 102.140 167.810 102.460 167.870 ;
        RECT 106.295 167.810 106.585 167.855 ;
        RECT 102.140 167.670 106.585 167.810 ;
        RECT 102.140 167.610 102.460 167.670 ;
        RECT 106.295 167.625 106.585 167.670 ;
        RECT 108.120 167.610 108.440 167.870 ;
        RECT 111.340 167.810 111.660 167.870 ;
        RECT 112.735 167.810 113.025 167.855 ;
        RECT 111.340 167.670 113.025 167.810 ;
        RECT 111.340 167.610 111.660 167.670 ;
        RECT 112.735 167.625 113.025 167.670 ;
        RECT 114.115 167.810 114.405 167.855 ;
        RECT 115.110 167.810 115.250 167.965 ;
        RECT 114.115 167.670 115.250 167.810 ;
        RECT 115.570 167.810 115.710 168.690 ;
        RECT 115.940 168.690 121.780 168.830 ;
        RECT 115.940 168.630 116.260 168.690 ;
        RECT 121.460 168.630 121.780 168.690 ;
        RECT 122.840 168.630 123.160 168.890 ;
        RECT 116.860 168.490 117.180 168.550 ;
        RECT 116.030 168.350 117.180 168.490 ;
        RECT 116.030 168.195 116.170 168.350 ;
        RECT 116.860 168.290 117.180 168.350 ;
        RECT 118.700 168.490 119.020 168.550 ;
        RECT 122.395 168.490 122.685 168.535 ;
        RECT 128.360 168.490 128.680 168.550 ;
        RECT 118.700 168.350 120.770 168.490 ;
        RECT 118.700 168.290 119.020 168.350 ;
        RECT 115.955 167.965 116.245 168.195 ;
        RECT 116.415 168.150 116.705 168.195 ;
        RECT 117.780 168.150 118.100 168.210 ;
        RECT 116.415 168.010 118.100 168.150 ;
        RECT 116.415 167.965 116.705 168.010 ;
        RECT 117.780 167.950 118.100 168.010 ;
        RECT 116.860 167.810 117.180 167.870 ;
        RECT 115.570 167.670 117.180 167.810 ;
        RECT 114.115 167.625 114.405 167.670 ;
        RECT 116.860 167.610 117.180 167.670 ;
        RECT 117.335 167.810 117.625 167.855 ;
        RECT 118.700 167.810 119.020 167.870 ;
        RECT 120.080 167.810 120.400 167.870 ;
        RECT 120.630 167.855 120.770 168.350 ;
        RECT 122.395 168.350 128.680 168.490 ;
        RECT 122.395 168.305 122.685 168.350 ;
        RECT 128.360 168.290 128.680 168.350 ;
        RECT 124.220 168.150 124.540 168.210 ;
        RECT 136.655 168.150 136.945 168.195 ;
        RECT 124.220 168.010 136.945 168.150 ;
        RECT 124.220 167.950 124.540 168.010 ;
        RECT 136.655 167.965 136.945 168.010 ;
        RECT 117.335 167.670 118.010 167.810 ;
        RECT 117.335 167.625 117.625 167.670 ;
        RECT 69.020 167.330 80.750 167.470 ;
        RECT 86.040 167.470 86.360 167.530 ;
        RECT 88.400 167.470 88.690 167.515 ;
        RECT 86.040 167.330 88.690 167.470 ;
        RECT 69.020 167.270 69.340 167.330 ;
        RECT 71.320 167.270 71.640 167.330 ;
        RECT 86.040 167.270 86.360 167.330 ;
        RECT 88.400 167.285 88.690 167.330 ;
        RECT 105.070 167.470 105.360 167.515 ;
        RECT 111.815 167.470 112.105 167.515 ;
        RECT 105.070 167.330 112.105 167.470 ;
        RECT 105.070 167.285 105.360 167.330 ;
        RECT 111.815 167.285 112.105 167.330 ;
        RECT 23.020 167.130 23.340 167.190 ;
        RECT 25.795 167.130 26.085 167.175 ;
        RECT 23.020 166.990 26.085 167.130 ;
        RECT 23.020 166.930 23.340 166.990 ;
        RECT 25.795 166.945 26.085 166.990 ;
        RECT 37.295 167.130 37.585 167.175 ;
        RECT 40.040 167.130 40.360 167.190 ;
        RECT 37.295 166.990 40.360 167.130 ;
        RECT 37.295 166.945 37.585 166.990 ;
        RECT 40.040 166.930 40.360 166.990 ;
        RECT 40.960 166.930 41.280 167.190 ;
        RECT 41.420 166.930 41.740 167.190 ;
        RECT 46.480 166.930 46.800 167.190 ;
        RECT 52.015 167.130 52.305 167.175 ;
        RECT 55.220 167.130 55.540 167.190 ;
        RECT 52.015 166.990 55.540 167.130 ;
        RECT 52.015 166.945 52.305 166.990 ;
        RECT 55.220 166.930 55.540 166.990 ;
        RECT 80.980 166.930 81.300 167.190 ;
        RECT 99.395 167.130 99.685 167.175 ;
        RECT 103.520 167.130 103.840 167.190 ;
        RECT 108.120 167.130 108.440 167.190 ;
        RECT 99.395 166.990 108.440 167.130 ;
        RECT 99.395 166.945 99.685 166.990 ;
        RECT 103.520 166.930 103.840 166.990 ;
        RECT 108.120 166.930 108.440 166.990 ;
        RECT 111.355 167.130 111.645 167.175 ;
        RECT 117.870 167.130 118.010 167.670 ;
        RECT 118.700 167.670 120.400 167.810 ;
        RECT 118.700 167.610 119.020 167.670 ;
        RECT 120.080 167.610 120.400 167.670 ;
        RECT 120.555 167.625 120.845 167.855 ;
        RECT 121.475 167.810 121.765 167.855 ;
        RECT 122.380 167.810 122.700 167.870 ;
        RECT 123.300 167.810 123.620 167.870 ;
        RECT 121.475 167.670 123.620 167.810 ;
        RECT 121.475 167.625 121.765 167.670 ;
        RECT 122.380 167.610 122.700 167.670 ;
        RECT 123.300 167.610 123.620 167.670 ;
        RECT 124.680 167.610 125.000 167.870 ;
        RECT 131.580 167.610 131.900 167.870 ;
        RECT 138.480 167.810 138.800 167.870 ;
        RECT 140.795 167.810 141.085 167.855 ;
        RECT 138.480 167.670 141.085 167.810 ;
        RECT 138.480 167.610 138.800 167.670 ;
        RECT 140.795 167.625 141.085 167.670 ;
        RECT 123.760 167.270 124.080 167.530 ;
        RECT 135.735 167.470 136.025 167.515 ;
        RECT 138.035 167.470 138.325 167.515 ;
        RECT 135.735 167.330 138.325 167.470 ;
        RECT 135.735 167.285 136.025 167.330 ;
        RECT 138.035 167.285 138.325 167.330 ;
        RECT 111.355 166.990 118.010 167.130 ;
        RECT 118.240 167.130 118.560 167.190 ;
        RECT 121.000 167.130 121.320 167.190 ;
        RECT 118.240 166.990 121.320 167.130 ;
        RECT 111.355 166.945 111.645 166.990 ;
        RECT 118.240 166.930 118.560 166.990 ;
        RECT 121.000 166.930 121.320 166.990 ;
        RECT 129.740 167.130 130.060 167.190 ;
        RECT 131.120 167.130 131.440 167.190 ;
        RECT 129.740 166.990 131.440 167.130 ;
        RECT 129.740 166.930 130.060 166.990 ;
        RECT 131.120 166.930 131.440 166.990 ;
        RECT 132.500 166.930 132.820 167.190 ;
        RECT 133.880 166.930 134.200 167.190 ;
        RECT 134.340 167.130 134.660 167.190 ;
        RECT 136.195 167.130 136.485 167.175 ;
        RECT 134.340 166.990 136.485 167.130 ;
        RECT 134.340 166.930 134.660 166.990 ;
        RECT 136.195 166.945 136.485 166.990 ;
        RECT 17.430 166.310 143.010 166.790 ;
        RECT 74.080 166.110 74.400 166.170 ;
        RECT 76.395 166.110 76.685 166.155 ;
        RECT 74.080 165.970 76.685 166.110 ;
        RECT 74.080 165.910 74.400 165.970 ;
        RECT 76.395 165.925 76.685 165.970 ;
        RECT 81.440 165.910 81.760 166.170 ;
        RECT 83.755 166.110 84.045 166.155 ;
        RECT 84.200 166.110 84.520 166.170 ;
        RECT 83.755 165.970 84.520 166.110 ;
        RECT 83.755 165.925 84.045 165.970 ;
        RECT 84.200 165.910 84.520 165.970 ;
        RECT 86.040 165.910 86.360 166.170 ;
        RECT 107.200 165.910 107.520 166.170 ;
        RECT 116.860 166.110 117.180 166.170 ;
        RECT 118.125 166.110 118.415 166.155 ;
        RECT 122.840 166.110 123.160 166.170 ;
        RECT 116.860 165.970 118.415 166.110 ;
        RECT 116.860 165.910 117.180 165.970 ;
        RECT 118.125 165.925 118.415 165.970 ;
        RECT 119.250 165.970 123.160 166.110 ;
        RECT 23.480 165.770 23.800 165.830 ;
        RECT 27.620 165.770 27.940 165.830 ;
        RECT 40.960 165.770 41.280 165.830 ;
        RECT 51.080 165.770 51.400 165.830 ;
        RECT 52.920 165.770 53.240 165.830 ;
        RECT 57.075 165.770 57.365 165.815 ;
        RECT 23.480 165.630 25.550 165.770 ;
        RECT 23.480 165.570 23.800 165.630 ;
        RECT 23.020 165.230 23.340 165.490 ;
        RECT 25.410 165.475 25.550 165.630 ;
        RECT 25.870 165.630 27.940 165.770 ;
        RECT 25.335 165.430 25.625 165.475 ;
        RECT 25.870 165.430 26.010 165.630 ;
        RECT 27.620 165.570 27.940 165.630 ;
        RECT 28.170 165.630 40.270 165.770 ;
        RECT 25.335 165.290 26.010 165.430 ;
        RECT 26.255 165.430 26.545 165.475 ;
        RECT 28.170 165.430 28.310 165.630 ;
        RECT 26.255 165.290 28.310 165.430 ;
        RECT 25.335 165.245 25.625 165.290 ;
        RECT 26.255 165.245 26.545 165.290 ;
        RECT 30.840 165.230 31.160 165.490 ;
        RECT 32.220 165.430 32.540 165.490 ;
        RECT 34.075 165.430 34.365 165.475 ;
        RECT 32.220 165.290 34.365 165.430 ;
        RECT 32.220 165.230 32.540 165.290 ;
        RECT 34.075 165.245 34.365 165.290 ;
        RECT 35.440 165.430 35.760 165.490 ;
        RECT 39.595 165.430 39.885 165.475 ;
        RECT 35.440 165.290 39.885 165.430 ;
        RECT 35.440 165.230 35.760 165.290 ;
        RECT 39.595 165.245 39.885 165.290 ;
        RECT 23.495 165.090 23.785 165.135 ;
        RECT 25.780 165.090 26.100 165.150 ;
        RECT 23.495 164.950 26.100 165.090 ;
        RECT 23.495 164.905 23.785 164.950 ;
        RECT 25.780 164.890 26.100 164.950 ;
        RECT 31.300 164.890 31.620 165.150 ;
        RECT 34.535 165.090 34.825 165.135 ;
        RECT 34.980 165.090 35.300 165.150 ;
        RECT 34.535 164.950 35.300 165.090 ;
        RECT 34.535 164.905 34.825 164.950 ;
        RECT 34.980 164.890 35.300 164.950 ;
        RECT 32.695 164.750 32.985 164.795 ;
        RECT 35.530 164.750 35.670 165.230 ;
        RECT 32.695 164.610 35.670 164.750 ;
        RECT 40.130 164.750 40.270 165.630 ;
        RECT 40.960 165.630 44.410 165.770 ;
        RECT 40.960 165.570 41.280 165.630 ;
        RECT 40.515 165.430 40.805 165.475 ;
        RECT 41.420 165.430 41.740 165.490 ;
        RECT 40.515 165.290 41.740 165.430 ;
        RECT 40.515 165.245 40.805 165.290 ;
        RECT 41.420 165.230 41.740 165.290 ;
        RECT 41.880 165.430 42.200 165.490 ;
        RECT 44.270 165.475 44.410 165.630 ;
        RECT 51.080 165.630 57.365 165.770 ;
        RECT 51.080 165.570 51.400 165.630 ;
        RECT 52.920 165.570 53.240 165.630 ;
        RECT 57.075 165.585 57.365 165.630 ;
        RECT 66.735 165.770 67.025 165.815 ;
        RECT 70.720 165.770 71.010 165.815 ;
        RECT 109.040 165.770 109.360 165.830 ;
        RECT 119.250 165.815 119.390 165.970 ;
        RECT 122.840 165.910 123.160 165.970 ;
        RECT 124.220 165.910 124.540 166.170 ;
        RECT 130.675 166.110 130.965 166.155 ;
        RECT 131.580 166.110 131.900 166.170 ;
        RECT 138.035 166.110 138.325 166.155 ;
        RECT 138.480 166.110 138.800 166.170 ;
        RECT 130.675 165.970 131.900 166.110 ;
        RECT 130.675 165.925 130.965 165.970 ;
        RECT 131.580 165.910 131.900 165.970 ;
        RECT 132.130 165.970 138.800 166.110 ;
        RECT 66.735 165.630 71.010 165.770 ;
        RECT 66.735 165.585 67.025 165.630 ;
        RECT 70.720 165.585 71.010 165.630 ;
        RECT 106.370 165.630 109.360 165.770 ;
        RECT 43.735 165.430 44.025 165.475 ;
        RECT 41.880 165.290 44.025 165.430 ;
        RECT 41.880 165.230 42.200 165.290 ;
        RECT 43.735 165.245 44.025 165.290 ;
        RECT 44.200 165.245 44.490 165.475 ;
        RECT 44.640 165.430 44.960 165.490 ;
        RECT 46.480 165.475 46.800 165.490 ;
        RECT 45.115 165.430 45.405 165.475 ;
        RECT 44.640 165.290 45.405 165.430 ;
        RECT 44.640 165.230 44.960 165.290 ;
        RECT 45.115 165.245 45.405 165.290 ;
        RECT 45.575 165.245 45.865 165.475 ;
        RECT 46.265 165.245 46.800 165.475 ;
        RECT 41.510 165.090 41.650 165.230 ;
        RECT 45.650 165.090 45.790 165.245 ;
        RECT 46.480 165.230 46.800 165.245 ;
        RECT 53.840 165.230 54.160 165.490 ;
        RECT 65.355 165.430 65.645 165.475 ;
        RECT 69.020 165.430 69.340 165.490 ;
        RECT 65.355 165.290 69.340 165.430 ;
        RECT 65.355 165.245 65.645 165.290 ;
        RECT 69.020 165.230 69.340 165.290 ;
        RECT 69.480 165.230 69.800 165.490 ;
        RECT 82.360 165.430 82.680 165.490 ;
        RECT 84.215 165.430 84.505 165.475 ;
        RECT 82.360 165.290 84.505 165.430 ;
        RECT 82.360 165.230 82.680 165.290 ;
        RECT 84.215 165.245 84.505 165.290 ;
        RECT 87.895 165.430 88.185 165.475 ;
        RECT 95.240 165.430 95.560 165.490 ;
        RECT 87.895 165.290 95.560 165.430 ;
        RECT 87.895 165.245 88.185 165.290 ;
        RECT 95.240 165.230 95.560 165.290 ;
        RECT 98.000 165.230 98.320 165.490 ;
        RECT 106.370 165.475 106.510 165.630 ;
        RECT 109.040 165.570 109.360 165.630 ;
        RECT 119.175 165.585 119.465 165.815 ;
        RECT 120.080 165.770 120.400 165.830 ;
        RECT 132.130 165.770 132.270 165.970 ;
        RECT 138.035 165.925 138.325 165.970 ;
        RECT 138.480 165.910 138.800 165.970 ;
        RECT 140.780 165.910 141.100 166.170 ;
        RECT 120.080 165.630 122.610 165.770 ;
        RECT 120.080 165.570 120.400 165.630 ;
        RECT 106.295 165.245 106.585 165.475 ;
        RECT 107.215 165.430 107.505 165.475 ;
        RECT 108.120 165.430 108.440 165.490 ;
        RECT 107.215 165.290 108.440 165.430 ;
        RECT 107.215 165.245 107.505 165.290 ;
        RECT 108.120 165.230 108.440 165.290 ;
        RECT 121.015 165.430 121.305 165.475 ;
        RECT 121.460 165.430 121.780 165.490 ;
        RECT 122.470 165.475 122.610 165.630 ;
        RECT 129.830 165.630 132.270 165.770 ;
        RECT 132.470 165.770 132.760 165.815 ;
        RECT 133.880 165.770 134.200 165.830 ;
        RECT 132.470 165.630 134.200 165.770 ;
        RECT 129.830 165.475 129.970 165.630 ;
        RECT 132.470 165.585 132.760 165.630 ;
        RECT 133.880 165.570 134.200 165.630 ;
        RECT 136.180 165.770 136.500 165.830 ;
        RECT 136.180 165.630 140.090 165.770 ;
        RECT 136.180 165.570 136.500 165.630 ;
        RECT 121.015 165.290 121.780 165.430 ;
        RECT 121.015 165.245 121.305 165.290 ;
        RECT 121.460 165.230 121.780 165.290 ;
        RECT 121.935 165.245 122.225 165.475 ;
        RECT 122.395 165.245 122.685 165.475 ;
        RECT 122.855 165.245 123.145 165.475 ;
        RECT 129.755 165.245 130.045 165.475 ;
        RECT 130.660 165.430 130.980 165.490 ;
        RECT 131.135 165.430 131.425 165.475 ;
        RECT 130.660 165.290 131.425 165.430 ;
        RECT 41.510 164.950 45.790 165.090 ;
        RECT 54.300 164.890 54.620 165.150 ;
        RECT 55.220 165.090 55.540 165.150 ;
        RECT 56.155 165.090 56.445 165.135 ;
        RECT 55.220 164.950 56.445 165.090 ;
        RECT 55.220 164.890 55.540 164.950 ;
        RECT 56.155 164.905 56.445 164.950 ;
        RECT 66.735 164.905 67.025 165.135 ;
        RECT 70.375 165.090 70.665 165.135 ;
        RECT 71.565 165.090 71.855 165.135 ;
        RECT 74.085 165.090 74.375 165.135 ;
        RECT 70.375 164.950 74.375 165.090 ;
        RECT 70.375 164.905 70.665 164.950 ;
        RECT 71.565 164.905 71.855 164.950 ;
        RECT 74.085 164.905 74.375 164.950 ;
        RECT 49.240 164.750 49.560 164.810 ;
        RECT 51.540 164.750 51.860 164.810 ;
        RECT 52.460 164.750 52.780 164.810 ;
        RECT 63.960 164.750 64.280 164.810 ;
        RECT 40.130 164.610 64.280 164.750 ;
        RECT 32.695 164.565 32.985 164.610 ;
        RECT 49.240 164.550 49.560 164.610 ;
        RECT 51.540 164.550 51.860 164.610 ;
        RECT 52.460 164.550 52.780 164.610 ;
        RECT 63.960 164.550 64.280 164.610 ;
        RECT 24.860 164.210 25.180 164.470 ;
        RECT 35.455 164.410 35.745 164.455 ;
        RECT 35.900 164.410 36.220 164.470 ;
        RECT 39.595 164.410 39.885 164.455 ;
        RECT 35.455 164.270 39.885 164.410 ;
        RECT 35.455 164.225 35.745 164.270 ;
        RECT 35.900 164.210 36.220 164.270 ;
        RECT 39.595 164.225 39.885 164.270 ;
        RECT 41.435 164.410 41.725 164.455 ;
        RECT 41.880 164.410 42.200 164.470 ;
        RECT 41.435 164.270 42.200 164.410 ;
        RECT 41.435 164.225 41.725 164.270 ;
        RECT 41.880 164.210 42.200 164.270 ;
        RECT 46.940 164.210 47.260 164.470 ;
        RECT 55.695 164.410 55.985 164.455 ;
        RECT 63.500 164.410 63.820 164.470 ;
        RECT 55.695 164.270 63.820 164.410 ;
        RECT 55.695 164.225 55.985 164.270 ;
        RECT 63.500 164.210 63.820 164.270 ;
        RECT 65.800 164.210 66.120 164.470 ;
        RECT 66.810 164.410 66.950 164.905 ;
        RECT 78.220 164.890 78.540 165.150 ;
        RECT 80.060 165.090 80.380 165.150 ;
        RECT 84.675 165.090 84.965 165.135 ;
        RECT 80.060 164.950 84.965 165.090 ;
        RECT 80.060 164.890 80.380 164.950 ;
        RECT 84.675 164.905 84.965 164.950 ;
        RECT 88.340 164.890 88.660 165.150 ;
        RECT 89.260 164.890 89.580 165.150 ;
        RECT 90.180 165.090 90.500 165.150 ;
        RECT 101.695 165.090 101.985 165.135 ;
        RECT 102.140 165.090 102.460 165.150 ;
        RECT 90.180 164.950 102.460 165.090 ;
        RECT 122.010 165.090 122.150 165.245 ;
        RECT 122.010 164.950 122.380 165.090 ;
        RECT 90.180 164.890 90.500 164.950 ;
        RECT 101.695 164.905 101.985 164.950 ;
        RECT 102.140 164.890 102.460 164.950 ;
        RECT 122.240 164.810 122.380 164.950 ;
        RECT 69.980 164.750 70.270 164.795 ;
        RECT 72.080 164.750 72.370 164.795 ;
        RECT 73.650 164.750 73.940 164.795 ;
        RECT 80.980 164.750 81.300 164.810 ;
        RECT 69.980 164.610 73.940 164.750 ;
        RECT 69.980 164.565 70.270 164.610 ;
        RECT 72.080 164.565 72.370 164.610 ;
        RECT 73.650 164.565 73.940 164.610 ;
        RECT 76.010 164.610 81.300 164.750 ;
        RECT 122.240 164.610 122.700 164.810 ;
        RECT 76.010 164.410 76.150 164.610 ;
        RECT 80.980 164.550 81.300 164.610 ;
        RECT 122.380 164.550 122.700 164.610 ;
        RECT 66.810 164.270 76.150 164.410 ;
        RECT 81.900 164.210 82.220 164.470 ;
        RECT 117.320 164.210 117.640 164.470 ;
        RECT 117.780 164.410 118.100 164.470 ;
        RECT 118.255 164.410 118.545 164.455 ;
        RECT 117.780 164.270 118.545 164.410 ;
        RECT 117.780 164.210 118.100 164.270 ;
        RECT 118.255 164.225 118.545 164.270 ;
        RECT 119.620 164.410 119.940 164.470 ;
        RECT 121.920 164.410 122.240 164.470 ;
        RECT 122.930 164.410 123.070 165.245 ;
        RECT 130.660 165.230 130.980 165.290 ;
        RECT 131.135 165.245 131.425 165.290 ;
        RECT 139.400 165.230 139.720 165.490 ;
        RECT 139.950 165.475 140.090 165.630 ;
        RECT 139.875 165.245 140.165 165.475 ;
        RECT 132.015 165.090 132.305 165.135 ;
        RECT 133.205 165.090 133.495 165.135 ;
        RECT 135.725 165.090 136.015 165.135 ;
        RECT 132.015 164.950 136.015 165.090 ;
        RECT 132.015 164.905 132.305 164.950 ;
        RECT 133.205 164.905 133.495 164.950 ;
        RECT 135.725 164.905 136.015 164.950 ;
        RECT 131.620 164.750 131.910 164.795 ;
        RECT 133.720 164.750 134.010 164.795 ;
        RECT 135.290 164.750 135.580 164.795 ;
        RECT 131.620 164.610 135.580 164.750 ;
        RECT 131.620 164.565 131.910 164.610 ;
        RECT 133.720 164.565 134.010 164.610 ;
        RECT 135.290 164.565 135.580 164.610 ;
        RECT 124.680 164.410 125.000 164.470 ;
        RECT 119.620 164.270 125.000 164.410 ;
        RECT 119.620 164.210 119.940 164.270 ;
        RECT 121.920 164.210 122.240 164.270 ;
        RECT 124.680 164.210 125.000 164.270 ;
        RECT 138.480 164.210 138.800 164.470 ;
        RECT 17.430 163.590 143.010 164.070 ;
        RECT 19.815 163.390 20.105 163.435 ;
        RECT 32.680 163.390 33.000 163.450 ;
        RECT 19.815 163.250 33.000 163.390 ;
        RECT 19.815 163.205 20.105 163.250 ;
        RECT 32.680 163.190 33.000 163.250 ;
        RECT 37.280 163.390 37.600 163.450 ;
        RECT 39.135 163.390 39.425 163.435 ;
        RECT 64.420 163.390 64.740 163.450 ;
        RECT 37.280 163.250 39.425 163.390 ;
        RECT 37.280 163.190 37.600 163.250 ;
        RECT 39.135 163.205 39.425 163.250 ;
        RECT 39.655 163.250 64.740 163.390 ;
        RECT 25.320 163.050 25.640 163.110 ;
        RECT 39.655 163.050 39.795 163.250 ;
        RECT 64.420 163.190 64.740 163.250 ;
        RECT 70.415 163.390 70.705 163.435 ;
        RECT 73.175 163.390 73.465 163.435 ;
        RECT 74.540 163.390 74.860 163.450 ;
        RECT 70.415 163.250 74.860 163.390 ;
        RECT 70.415 163.205 70.705 163.250 ;
        RECT 73.175 163.205 73.465 163.250 ;
        RECT 74.540 163.190 74.860 163.250 ;
        RECT 80.980 163.190 81.300 163.450 ;
        RECT 95.240 163.190 95.560 163.450 ;
        RECT 119.635 163.390 119.925 163.435 ;
        RECT 124.220 163.390 124.540 163.450 ;
        RECT 119.635 163.250 124.540 163.390 ;
        RECT 119.635 163.205 119.925 163.250 ;
        RECT 124.220 163.190 124.540 163.250 ;
        RECT 130.215 163.390 130.505 163.435 ;
        RECT 134.340 163.390 134.660 163.450 ;
        RECT 130.215 163.250 134.660 163.390 ;
        RECT 130.215 163.205 130.505 163.250 ;
        RECT 134.340 163.190 134.660 163.250 ;
        RECT 25.320 162.910 39.795 163.050 ;
        RECT 51.080 163.050 51.400 163.110 ;
        RECT 54.300 163.050 54.620 163.110 ;
        RECT 59.360 163.050 59.650 163.095 ;
        RECT 60.930 163.050 61.220 163.095 ;
        RECT 63.030 163.050 63.320 163.095 ;
        RECT 51.080 162.910 54.990 163.050 ;
        RECT 25.320 162.850 25.640 162.910 ;
        RECT 23.035 162.710 23.325 162.755 ;
        RECT 24.400 162.710 24.720 162.770 ;
        RECT 23.035 162.570 24.720 162.710 ;
        RECT 23.035 162.525 23.325 162.570 ;
        RECT 24.400 162.510 24.720 162.570 ;
        RECT 24.860 162.710 25.180 162.770 ;
        RECT 27.050 162.710 27.340 162.755 ;
        RECT 24.860 162.570 27.340 162.710 ;
        RECT 24.860 162.510 25.180 162.570 ;
        RECT 27.050 162.525 27.340 162.570 ;
        RECT 27.620 162.510 27.940 162.770 ;
        RECT 29.550 162.755 29.690 162.910 ;
        RECT 51.080 162.850 51.400 162.910 ;
        RECT 54.300 162.850 54.620 162.910 ;
        RECT 29.475 162.525 29.765 162.755 ;
        RECT 40.040 162.510 40.360 162.770 ;
        RECT 40.500 162.710 40.820 162.770 ;
        RECT 45.560 162.710 45.880 162.770 ;
        RECT 40.500 162.570 52.230 162.710 ;
        RECT 40.500 162.510 40.820 162.570 ;
        RECT 16.120 162.370 16.440 162.430 ;
        RECT 18.895 162.370 19.185 162.415 ;
        RECT 16.120 162.230 19.185 162.370 ;
        RECT 16.120 162.170 16.440 162.230 ;
        RECT 18.895 162.185 19.185 162.230 ;
        RECT 22.575 162.370 22.865 162.415 ;
        RECT 23.480 162.370 23.800 162.430 ;
        RECT 22.575 162.230 23.800 162.370 ;
        RECT 24.490 162.370 24.630 162.510 ;
        RECT 28.095 162.370 28.385 162.415 ;
        RECT 24.490 162.230 28.385 162.370 ;
        RECT 22.575 162.185 22.865 162.230 ;
        RECT 23.480 162.170 23.800 162.230 ;
        RECT 28.095 162.185 28.385 162.230 ;
        RECT 30.840 162.370 31.160 162.430 ;
        RECT 31.315 162.370 31.605 162.415 ;
        RECT 30.840 162.230 31.605 162.370 ;
        RECT 30.840 162.170 31.160 162.230 ;
        RECT 31.315 162.185 31.605 162.230 ;
        RECT 32.220 162.170 32.540 162.430 ;
        RECT 35.440 162.170 35.760 162.430 ;
        RECT 35.900 162.170 36.220 162.430 ;
        RECT 36.835 162.185 37.125 162.415 ;
        RECT 25.335 162.030 25.625 162.075 ;
        RECT 25.780 162.030 26.100 162.090 ;
        RECT 25.335 161.890 26.100 162.030 ;
        RECT 36.910 162.030 37.050 162.185 ;
        RECT 37.280 162.170 37.600 162.430 ;
        RECT 38.660 162.415 38.980 162.430 ;
        RECT 38.615 162.185 38.980 162.415 ;
        RECT 38.660 162.170 38.980 162.185 ;
        RECT 40.960 162.170 41.280 162.430 ;
        RECT 44.640 162.370 44.960 162.430 ;
        RECT 45.190 162.415 45.330 162.570 ;
        RECT 45.560 162.510 45.880 162.570 ;
        RECT 41.510 162.230 44.960 162.370 ;
        RECT 39.580 162.030 39.900 162.090 ;
        RECT 41.510 162.030 41.650 162.230 ;
        RECT 44.640 162.170 44.960 162.230 ;
        RECT 45.115 162.185 45.405 162.415 ;
        RECT 48.780 162.370 49.100 162.430 ;
        RECT 52.090 162.415 52.230 162.570 ;
        RECT 53.840 162.510 54.160 162.770 ;
        RECT 54.850 162.755 54.990 162.910 ;
        RECT 59.360 162.910 63.320 163.050 ;
        RECT 59.360 162.865 59.650 162.910 ;
        RECT 60.930 162.865 61.220 162.910 ;
        RECT 63.030 162.865 63.320 162.910 ;
        RECT 65.800 163.050 66.120 163.110 ;
        RECT 74.080 163.050 74.400 163.110 ;
        RECT 65.800 162.910 74.400 163.050 ;
        RECT 65.800 162.850 66.120 162.910 ;
        RECT 74.080 162.850 74.400 162.910 ;
        RECT 54.775 162.525 55.065 162.755 ;
        RECT 58.925 162.710 59.215 162.755 ;
        RECT 61.445 162.710 61.735 162.755 ;
        RECT 62.635 162.710 62.925 162.755 ;
        RECT 58.925 162.570 62.925 162.710 ;
        RECT 58.925 162.525 59.215 162.570 ;
        RECT 61.445 162.525 61.735 162.570 ;
        RECT 62.635 162.525 62.925 162.570 ;
        RECT 73.620 162.710 73.940 162.770 ;
        RECT 74.630 162.710 74.770 163.190 ;
        RECT 78.235 162.865 78.525 163.095 ;
        RECT 124.680 163.050 125.000 163.110 ;
        RECT 124.680 162.910 125.830 163.050 ;
        RECT 73.620 162.510 74.080 162.710 ;
        RECT 74.630 162.570 76.610 162.710 ;
        RECT 50.635 162.370 50.925 162.415 ;
        RECT 48.780 162.230 50.925 162.370 ;
        RECT 48.780 162.170 49.100 162.230 ;
        RECT 50.635 162.185 50.925 162.230 ;
        RECT 52.015 162.185 52.305 162.415 ;
        RECT 53.395 162.185 53.685 162.415 ;
        RECT 54.315 162.370 54.605 162.415 ;
        RECT 56.600 162.370 56.920 162.430 ;
        RECT 54.315 162.230 56.920 162.370 ;
        RECT 54.315 162.185 54.605 162.230 ;
        RECT 36.910 161.890 39.900 162.030 ;
        RECT 25.335 161.845 25.625 161.890 ;
        RECT 25.780 161.830 26.100 161.890 ;
        RECT 39.580 161.830 39.900 161.890 ;
        RECT 41.050 161.890 41.650 162.030 ;
        RECT 21.640 161.490 21.960 161.750 ;
        RECT 26.240 161.490 26.560 161.750 ;
        RECT 31.775 161.690 32.065 161.735 ;
        RECT 34.060 161.690 34.380 161.750 ;
        RECT 31.775 161.550 34.380 161.690 ;
        RECT 31.775 161.505 32.065 161.550 ;
        RECT 34.060 161.490 34.380 161.550 ;
        RECT 38.215 161.690 38.505 161.735 ;
        RECT 41.050 161.690 41.190 161.890 ;
        RECT 44.180 161.830 44.500 162.090 ;
        RECT 53.470 162.030 53.610 162.185 ;
        RECT 56.600 162.170 56.920 162.230 ;
        RECT 63.040 162.370 63.360 162.430 ;
        RECT 63.515 162.370 63.805 162.415 ;
        RECT 73.940 162.370 74.080 162.510 ;
        RECT 76.470 162.415 76.610 162.570 ;
        RECT 75.935 162.370 76.225 162.415 ;
        RECT 63.040 162.230 63.805 162.370 ;
        RECT 63.040 162.170 63.360 162.230 ;
        RECT 63.515 162.185 63.805 162.230 ;
        RECT 72.330 162.230 76.225 162.370 ;
        RECT 72.330 162.090 72.470 162.230 ;
        RECT 75.935 162.185 76.225 162.230 ;
        RECT 76.395 162.185 76.685 162.415 ;
        RECT 76.855 162.370 77.145 162.415 ;
        RECT 77.300 162.370 77.620 162.430 ;
        RECT 76.855 162.230 77.620 162.370 ;
        RECT 76.855 162.185 77.145 162.230 ;
        RECT 77.300 162.170 77.620 162.230 ;
        RECT 77.775 162.370 78.065 162.415 ;
        RECT 78.310 162.370 78.450 162.865 ;
        RECT 124.680 162.850 125.000 162.910 ;
        RECT 78.680 162.710 79.000 162.770 ;
        RECT 79.615 162.710 79.905 162.755 ;
        RECT 78.680 162.570 79.905 162.710 ;
        RECT 78.680 162.510 79.000 162.570 ;
        RECT 79.615 162.525 79.905 162.570 ;
        RECT 87.880 162.510 88.200 162.770 ;
        RECT 97.540 162.510 97.860 162.770 ;
        RECT 98.460 162.510 98.780 162.770 ;
        RECT 121.920 162.710 122.240 162.770 ;
        RECT 121.920 162.570 125.370 162.710 ;
        RECT 121.920 162.510 122.240 162.570 ;
        RECT 77.775 162.230 78.450 162.370 ;
        RECT 77.775 162.185 78.065 162.230 ;
        RECT 79.155 162.185 79.445 162.415 ;
        RECT 80.060 162.370 80.380 162.430 ;
        RECT 81.455 162.370 81.745 162.415 ;
        RECT 80.060 162.230 81.745 162.370 ;
        RECT 60.280 162.030 60.600 162.090 ;
        RECT 62.180 162.030 62.470 162.075 ;
        RECT 49.330 161.890 56.830 162.030 ;
        RECT 38.215 161.550 41.190 161.690 ;
        RECT 41.420 161.690 41.740 161.750 ;
        RECT 41.895 161.690 42.185 161.735 ;
        RECT 41.420 161.550 42.185 161.690 ;
        RECT 38.215 161.505 38.505 161.550 ;
        RECT 41.420 161.490 41.740 161.550 ;
        RECT 41.895 161.505 42.185 161.550 ;
        RECT 43.260 161.490 43.580 161.750 ;
        RECT 44.270 161.690 44.410 161.830 ;
        RECT 49.330 161.690 49.470 161.890 ;
        RECT 44.270 161.550 49.470 161.690 ;
        RECT 49.700 161.490 50.020 161.750 ;
        RECT 51.555 161.690 51.845 161.735 ;
        RECT 53.840 161.690 54.160 161.750 ;
        RECT 51.555 161.550 54.160 161.690 ;
        RECT 51.555 161.505 51.845 161.550 ;
        RECT 53.840 161.490 54.160 161.550 ;
        RECT 55.680 161.490 56.000 161.750 ;
        RECT 56.690 161.735 56.830 161.890 ;
        RECT 60.280 161.890 62.470 162.030 ;
        RECT 60.280 161.830 60.600 161.890 ;
        RECT 62.180 161.845 62.470 161.890 ;
        RECT 69.495 162.030 69.785 162.075 ;
        RECT 72.240 162.030 72.560 162.090 ;
        RECT 69.495 161.890 72.560 162.030 ;
        RECT 69.495 161.845 69.785 161.890 ;
        RECT 72.240 161.830 72.560 161.890 ;
        RECT 73.160 162.075 73.480 162.090 ;
        RECT 73.160 161.845 73.545 162.075 ;
        RECT 79.230 162.030 79.370 162.185 ;
        RECT 80.060 162.170 80.380 162.230 ;
        RECT 81.455 162.185 81.745 162.230 ;
        RECT 83.755 162.370 84.045 162.415 ;
        RECT 84.200 162.370 84.520 162.430 ;
        RECT 83.755 162.230 84.520 162.370 ;
        RECT 83.755 162.185 84.045 162.230 ;
        RECT 84.200 162.170 84.520 162.230 ;
        RECT 84.660 162.370 84.980 162.430 ;
        RECT 91.115 162.370 91.405 162.415 ;
        RECT 84.660 162.230 91.405 162.370 ;
        RECT 84.660 162.170 84.980 162.230 ;
        RECT 91.115 162.185 91.405 162.230 ;
        RECT 96.160 162.370 96.480 162.430 ;
        RECT 100.775 162.370 101.065 162.415 ;
        RECT 96.160 162.230 101.065 162.370 ;
        RECT 96.160 162.170 96.480 162.230 ;
        RECT 100.775 162.185 101.065 162.230 ;
        RECT 115.480 162.370 115.800 162.430 ;
        RECT 117.795 162.370 118.085 162.415 ;
        RECT 115.480 162.230 118.085 162.370 ;
        RECT 115.480 162.170 115.800 162.230 ;
        RECT 117.795 162.185 118.085 162.230 ;
        RECT 118.715 162.370 119.005 162.415 ;
        RECT 119.160 162.370 119.480 162.430 ;
        RECT 118.715 162.230 119.480 162.370 ;
        RECT 118.715 162.185 119.005 162.230 ;
        RECT 119.160 162.170 119.480 162.230 ;
        RECT 119.620 162.370 119.940 162.430 ;
        RECT 119.620 162.365 120.770 162.370 ;
        RECT 121.015 162.365 121.305 162.415 ;
        RECT 119.620 162.230 121.305 162.365 ;
        RECT 119.620 162.170 119.940 162.230 ;
        RECT 120.630 162.225 121.305 162.230 ;
        RECT 121.015 162.185 121.305 162.225 ;
        RECT 74.170 161.890 79.370 162.030 ;
        RECT 88.815 162.030 89.105 162.075 ;
        RECT 101.220 162.030 101.540 162.090 ;
        RECT 121.475 162.075 121.765 162.305 ;
        RECT 123.300 162.170 123.620 162.430 ;
        RECT 123.760 162.170 124.080 162.430 ;
        RECT 125.230 162.415 125.370 162.570 ;
        RECT 125.690 162.415 125.830 162.910 ;
        RECT 129.740 162.710 130.060 162.770 ;
        RECT 136.655 162.710 136.945 162.755 ;
        RECT 129.740 162.570 136.945 162.710 ;
        RECT 129.740 162.510 130.060 162.570 ;
        RECT 136.655 162.525 136.945 162.570 ;
        RECT 124.695 162.370 124.985 162.415 ;
        RECT 124.310 162.230 124.985 162.370 ;
        RECT 88.815 161.890 101.540 162.030 ;
        RECT 73.160 161.830 73.480 161.845 ;
        RECT 70.400 161.735 70.720 161.750 ;
        RECT 56.615 161.505 56.905 161.735 ;
        RECT 70.400 161.505 70.785 161.735 ;
        RECT 70.400 161.490 70.720 161.505 ;
        RECT 71.320 161.490 71.640 161.750 ;
        RECT 74.170 161.735 74.310 161.890 ;
        RECT 88.815 161.845 89.105 161.890 ;
        RECT 101.220 161.830 101.540 161.890 ;
        RECT 74.095 161.505 74.385 161.735 ;
        RECT 74.555 161.690 74.845 161.735 ;
        RECT 76.840 161.690 77.160 161.750 ;
        RECT 74.555 161.550 77.160 161.690 ;
        RECT 74.555 161.505 74.845 161.550 ;
        RECT 76.840 161.490 77.160 161.550 ;
        RECT 86.515 161.690 86.805 161.735 ;
        RECT 88.355 161.690 88.645 161.735 ;
        RECT 86.515 161.550 88.645 161.690 ;
        RECT 86.515 161.505 86.805 161.550 ;
        RECT 88.355 161.505 88.645 161.550 ;
        RECT 89.720 161.690 90.040 161.750 ;
        RECT 90.655 161.690 90.945 161.735 ;
        RECT 89.720 161.550 90.945 161.690 ;
        RECT 89.720 161.490 90.040 161.550 ;
        RECT 90.655 161.505 90.945 161.550 ;
        RECT 92.020 161.690 92.340 161.750 ;
        RECT 94.335 161.690 94.625 161.735 ;
        RECT 92.020 161.550 94.625 161.690 ;
        RECT 92.020 161.490 92.340 161.550 ;
        RECT 94.335 161.505 94.625 161.550 ;
        RECT 97.095 161.690 97.385 161.735 ;
        RECT 97.540 161.690 97.860 161.750 ;
        RECT 97.095 161.550 97.860 161.690 ;
        RECT 97.095 161.505 97.385 161.550 ;
        RECT 97.540 161.490 97.860 161.550 ;
        RECT 103.995 161.690 104.285 161.735 ;
        RECT 104.900 161.690 105.220 161.750 ;
        RECT 103.995 161.550 105.220 161.690 ;
        RECT 103.995 161.505 104.285 161.550 ;
        RECT 104.900 161.490 105.220 161.550 ;
        RECT 109.960 161.690 110.280 161.750 ;
        RECT 113.180 161.690 113.500 161.750 ;
        RECT 118.700 161.690 119.020 161.750 ;
        RECT 109.960 161.550 119.020 161.690 ;
        RECT 109.960 161.490 110.280 161.550 ;
        RECT 113.180 161.490 113.500 161.550 ;
        RECT 118.700 161.490 119.020 161.550 ;
        RECT 120.080 161.490 120.400 161.750 ;
        RECT 121.000 161.690 121.320 161.750 ;
        RECT 121.550 161.690 121.690 162.075 ;
        RECT 122.840 161.830 123.160 162.090 ;
        RECT 121.000 161.550 121.690 161.690 ;
        RECT 121.920 161.690 122.240 161.750 ;
        RECT 124.310 161.690 124.450 162.230 ;
        RECT 124.695 162.185 124.985 162.230 ;
        RECT 125.155 162.185 125.445 162.415 ;
        RECT 125.615 162.185 125.905 162.415 ;
        RECT 127.455 162.370 127.745 162.415 ;
        RECT 127.900 162.370 128.220 162.430 ;
        RECT 127.455 162.230 128.220 162.370 ;
        RECT 127.455 162.185 127.745 162.230 ;
        RECT 127.900 162.170 128.220 162.230 ;
        RECT 129.295 162.370 129.585 162.415 ;
        RECT 130.200 162.370 130.520 162.430 ;
        RECT 129.295 162.230 130.520 162.370 ;
        RECT 129.295 162.185 129.585 162.230 ;
        RECT 130.200 162.170 130.520 162.230 ;
        RECT 137.560 162.370 137.880 162.430 ;
        RECT 139.400 162.370 139.720 162.430 ;
        RECT 140.795 162.370 141.085 162.415 ;
        RECT 137.560 162.230 141.085 162.370 ;
        RECT 137.560 162.170 137.880 162.230 ;
        RECT 139.400 162.170 139.720 162.230 ;
        RECT 140.795 162.185 141.085 162.230 ;
        RECT 126.520 162.030 126.840 162.090 ;
        RECT 128.375 162.030 128.665 162.075 ;
        RECT 126.520 161.890 128.665 162.030 ;
        RECT 126.520 161.830 126.840 161.890 ;
        RECT 128.375 161.845 128.665 161.890 ;
        RECT 128.835 162.030 129.125 162.075 ;
        RECT 132.960 162.030 133.280 162.090 ;
        RECT 128.835 161.890 133.280 162.030 ;
        RECT 128.835 161.845 129.125 161.890 ;
        RECT 132.960 161.830 133.280 161.890 ;
        RECT 135.735 162.030 136.025 162.075 ;
        RECT 138.035 162.030 138.325 162.075 ;
        RECT 135.735 161.890 138.325 162.030 ;
        RECT 135.735 161.845 136.025 161.890 ;
        RECT 138.035 161.845 138.325 161.890 ;
        RECT 121.920 161.550 124.450 161.690 ;
        RECT 126.995 161.690 127.285 161.735 ;
        RECT 133.420 161.690 133.740 161.750 ;
        RECT 126.995 161.550 133.740 161.690 ;
        RECT 121.000 161.490 121.320 161.550 ;
        RECT 121.920 161.490 122.240 161.550 ;
        RECT 126.995 161.505 127.285 161.550 ;
        RECT 133.420 161.490 133.740 161.550 ;
        RECT 133.880 161.490 134.200 161.750 ;
        RECT 134.800 161.690 135.120 161.750 ;
        RECT 136.195 161.690 136.485 161.735 ;
        RECT 134.800 161.550 136.485 161.690 ;
        RECT 134.800 161.490 135.120 161.550 ;
        RECT 136.195 161.505 136.485 161.550 ;
        RECT 17.430 160.870 143.010 161.350 ;
        RECT 21.195 160.670 21.485 160.715 ;
        RECT 23.020 160.670 23.340 160.730 ;
        RECT 32.220 160.670 32.540 160.730 ;
        RECT 36.835 160.670 37.125 160.715 ;
        RECT 38.200 160.670 38.520 160.730 ;
        RECT 21.195 160.530 35.670 160.670 ;
        RECT 21.195 160.485 21.485 160.530 ;
        RECT 23.020 160.470 23.340 160.530 ;
        RECT 32.220 160.470 32.540 160.530 ;
        RECT 35.530 160.375 35.670 160.530 ;
        RECT 36.835 160.530 38.520 160.670 ;
        RECT 36.835 160.485 37.125 160.530 ;
        RECT 38.200 160.470 38.520 160.530 ;
        RECT 39.580 160.670 39.900 160.730 ;
        RECT 48.780 160.670 49.100 160.730 ;
        RECT 39.580 160.530 49.100 160.670 ;
        RECT 39.580 160.470 39.900 160.530 ;
        RECT 48.780 160.470 49.100 160.530 ;
        RECT 52.460 160.670 52.780 160.730 ;
        RECT 53.395 160.670 53.685 160.715 ;
        RECT 52.460 160.530 53.685 160.670 ;
        RECT 52.460 160.470 52.780 160.530 ;
        RECT 53.395 160.485 53.685 160.530 ;
        RECT 53.840 160.670 54.160 160.730 ;
        RECT 55.235 160.670 55.525 160.715 ;
        RECT 53.840 160.530 55.525 160.670 ;
        RECT 53.840 160.470 54.160 160.530 ;
        RECT 55.235 160.485 55.525 160.530 ;
        RECT 56.140 160.670 56.460 160.730 ;
        RECT 64.435 160.670 64.725 160.715 ;
        RECT 56.140 160.530 64.725 160.670 ;
        RECT 56.140 160.470 56.460 160.530 ;
        RECT 64.435 160.485 64.725 160.530 ;
        RECT 73.160 160.670 73.480 160.730 ;
        RECT 73.635 160.670 73.925 160.715 ;
        RECT 73.160 160.530 73.925 160.670 ;
        RECT 73.160 160.470 73.480 160.530 ;
        RECT 73.635 160.485 73.925 160.530 ;
        RECT 74.080 160.470 74.400 160.730 ;
        RECT 76.395 160.670 76.685 160.715 ;
        RECT 77.300 160.670 77.620 160.730 ;
        RECT 76.395 160.530 77.620 160.670 ;
        RECT 76.395 160.485 76.685 160.530 ;
        RECT 77.300 160.470 77.620 160.530 ;
        RECT 79.600 160.470 79.920 160.730 ;
        RECT 80.980 160.470 81.300 160.730 ;
        RECT 81.915 160.670 82.205 160.715 ;
        RECT 84.200 160.670 84.520 160.730 ;
        RECT 81.915 160.530 84.520 160.670 ;
        RECT 81.915 160.485 82.205 160.530 ;
        RECT 84.200 160.470 84.520 160.530 ;
        RECT 108.580 160.670 108.900 160.730 ;
        RECT 110.895 160.670 111.185 160.715 ;
        RECT 115.020 160.670 115.340 160.730 ;
        RECT 121.000 160.670 121.320 160.730 ;
        RECT 108.580 160.530 121.320 160.670 ;
        RECT 108.580 160.470 108.900 160.530 ;
        RECT 110.895 160.485 111.185 160.530 ;
        RECT 115.020 160.470 115.340 160.530 ;
        RECT 121.000 160.470 121.320 160.530 ;
        RECT 127.900 160.670 128.220 160.730 ;
        RECT 128.375 160.670 128.665 160.715 ;
        RECT 127.900 160.530 128.665 160.670 ;
        RECT 127.900 160.470 128.220 160.530 ;
        RECT 128.375 160.485 128.665 160.530 ;
        RECT 137.560 160.470 137.880 160.730 ;
        RECT 138.940 160.470 139.260 160.730 ;
        RECT 33.615 160.330 33.905 160.375 ;
        RECT 34.995 160.330 35.285 160.375 ;
        RECT 25.640 160.190 28.310 160.330 ;
        RECT 23.940 159.990 24.260 160.050 ;
        RECT 25.640 159.990 25.780 160.190 ;
        RECT 23.940 159.850 25.780 159.990 ;
        RECT 26.700 160.035 27.020 160.050 ;
        RECT 28.170 160.035 28.310 160.190 ;
        RECT 33.615 160.190 35.285 160.330 ;
        RECT 33.615 160.145 33.905 160.190 ;
        RECT 34.995 160.145 35.285 160.190 ;
        RECT 35.455 160.145 35.745 160.375 ;
        RECT 40.500 160.330 40.820 160.390 ;
        RECT 44.180 160.330 44.500 160.390 ;
        RECT 35.990 160.190 40.820 160.330 ;
        RECT 26.700 159.990 27.050 160.035 ;
        RECT 26.700 159.850 27.215 159.990 ;
        RECT 23.940 159.790 24.260 159.850 ;
        RECT 26.700 159.805 27.050 159.850 ;
        RECT 28.095 159.805 28.385 160.035 ;
        RECT 26.700 159.790 27.020 159.805 ;
        RECT 31.760 159.790 32.080 160.050 ;
        RECT 32.220 159.990 32.540 160.050 ;
        RECT 32.220 159.850 32.735 159.990 ;
        RECT 32.220 159.790 32.540 159.850 ;
        RECT 34.060 159.790 34.380 160.050 ;
        RECT 35.990 160.035 36.130 160.190 ;
        RECT 40.500 160.130 40.820 160.190 ;
        RECT 41.050 160.190 44.500 160.330 ;
        RECT 35.915 159.805 36.205 160.035 ;
        RECT 39.580 159.990 39.870 160.035 ;
        RECT 41.050 159.990 41.190 160.190 ;
        RECT 44.180 160.130 44.500 160.190 ;
        RECT 48.320 160.330 48.640 160.390 ;
        RECT 51.540 160.330 51.860 160.390 ;
        RECT 53.930 160.330 54.070 160.470 ;
        RECT 63.500 160.375 63.820 160.390 ;
        RECT 48.320 160.190 54.070 160.330 ;
        RECT 48.320 160.130 48.640 160.190 ;
        RECT 39.580 159.850 41.190 159.990 ;
        RECT 39.580 159.805 39.870 159.850 ;
        RECT 41.420 159.790 41.740 160.050 ;
        RECT 41.880 159.790 42.200 160.050 ;
        RECT 46.480 159.790 46.800 160.050 ;
        RECT 47.860 159.790 48.180 160.050 ;
        RECT 50.250 160.035 50.390 160.190 ;
        RECT 51.540 160.130 51.860 160.190 ;
        RECT 63.390 160.145 63.820 160.375 ;
        RECT 63.500 160.130 63.820 160.145 ;
        RECT 63.960 160.130 64.280 160.390 ;
        RECT 74.170 160.330 74.310 160.470 ;
        RECT 79.140 160.330 79.460 160.390 ;
        RECT 74.170 160.190 79.460 160.330 ;
        RECT 49.255 159.805 49.545 160.035 ;
        RECT 50.175 159.805 50.465 160.035 ;
        RECT 23.505 159.650 23.795 159.695 ;
        RECT 26.025 159.650 26.315 159.695 ;
        RECT 27.215 159.650 27.505 159.695 ;
        RECT 23.505 159.510 27.505 159.650 ;
        RECT 23.505 159.465 23.795 159.510 ;
        RECT 26.025 159.465 26.315 159.510 ;
        RECT 27.215 159.465 27.505 159.510 ;
        RECT 45.575 159.650 45.865 159.695 ;
        RECT 46.940 159.650 47.260 159.710 ;
        RECT 45.575 159.510 47.260 159.650 ;
        RECT 45.575 159.465 45.865 159.510 ;
        RECT 46.940 159.450 47.260 159.510 ;
        RECT 47.400 159.650 47.720 159.710 ;
        RECT 49.330 159.650 49.470 159.805 ;
        RECT 51.080 159.790 51.400 160.050 ;
        RECT 53.980 159.990 54.270 160.035 ;
        RECT 54.760 159.990 55.080 160.050 ;
        RECT 53.980 159.850 55.080 159.990 ;
        RECT 53.980 159.805 54.270 159.850 ;
        RECT 54.760 159.790 55.080 159.850 ;
        RECT 60.855 159.990 61.145 160.035 ;
        RECT 73.160 159.990 73.480 160.050 ;
        RECT 74.095 159.990 74.385 160.035 ;
        RECT 60.855 159.850 63.270 159.990 ;
        RECT 60.855 159.805 61.145 159.850 ;
        RECT 47.400 159.510 49.470 159.650 ;
        RECT 50.620 159.650 50.940 159.710 ;
        RECT 51.555 159.650 51.845 159.695 ;
        RECT 50.620 159.510 51.845 159.650 ;
        RECT 47.400 159.450 47.720 159.510 ;
        RECT 50.620 159.450 50.940 159.510 ;
        RECT 51.555 159.465 51.845 159.510 ;
        RECT 52.920 159.450 53.240 159.710 ;
        RECT 57.545 159.650 57.835 159.695 ;
        RECT 60.065 159.650 60.355 159.695 ;
        RECT 61.255 159.650 61.545 159.695 ;
        RECT 57.545 159.510 61.545 159.650 ;
        RECT 57.545 159.465 57.835 159.510 ;
        RECT 60.065 159.465 60.355 159.510 ;
        RECT 61.255 159.465 61.545 159.510 ;
        RECT 62.135 159.650 62.425 159.695 ;
        RECT 62.580 159.650 62.900 159.710 ;
        RECT 62.135 159.510 62.900 159.650 ;
        RECT 62.135 159.465 62.425 159.510 ;
        RECT 62.580 159.450 62.900 159.510 ;
        RECT 23.940 159.310 24.230 159.355 ;
        RECT 25.510 159.310 25.800 159.355 ;
        RECT 27.610 159.310 27.900 159.355 ;
        RECT 23.940 159.170 27.900 159.310 ;
        RECT 23.940 159.125 24.230 159.170 ;
        RECT 25.510 159.125 25.800 159.170 ;
        RECT 27.610 159.125 27.900 159.170 ;
        RECT 48.335 159.310 48.625 159.355 ;
        RECT 53.010 159.310 53.150 159.450 ;
        RECT 48.335 159.170 53.150 159.310 ;
        RECT 54.775 159.310 55.065 159.355 ;
        RECT 57.980 159.310 58.270 159.355 ;
        RECT 59.550 159.310 59.840 159.355 ;
        RECT 61.650 159.310 61.940 159.355 ;
        RECT 63.130 159.310 63.270 159.850 ;
        RECT 73.160 159.850 74.385 159.990 ;
        RECT 73.160 159.790 73.480 159.850 ;
        RECT 74.095 159.805 74.385 159.850 ;
        RECT 75.475 159.805 75.765 160.035 ;
        RECT 64.420 159.650 64.740 159.710 ;
        RECT 65.815 159.650 66.105 159.695 ;
        RECT 64.420 159.510 66.105 159.650 ;
        RECT 64.420 159.450 64.740 159.510 ;
        RECT 65.815 159.465 66.105 159.510 ;
        RECT 71.335 159.650 71.625 159.695 ;
        RECT 73.620 159.650 73.940 159.710 ;
        RECT 71.335 159.510 73.940 159.650 ;
        RECT 71.335 159.465 71.625 159.510 ;
        RECT 73.620 159.450 73.940 159.510 ;
        RECT 75.000 159.450 75.320 159.710 ;
        RECT 75.550 159.650 75.690 159.805 ;
        RECT 76.840 159.790 77.160 160.050 ;
        RECT 77.390 160.035 77.530 160.190 ;
        RECT 79.140 160.130 79.460 160.190 ;
        RECT 89.720 160.375 90.040 160.390 ;
        RECT 89.720 160.330 90.070 160.375 ;
        RECT 101.850 160.330 102.140 160.375 ;
        RECT 103.535 160.330 103.825 160.375 ;
        RECT 113.195 160.330 113.485 160.375 ;
        RECT 127.455 160.330 127.745 160.375 ;
        RECT 132.010 160.330 132.300 160.375 ;
        RECT 133.880 160.330 134.200 160.390 ;
        RECT 89.720 160.190 90.235 160.330 ;
        RECT 101.850 160.190 103.825 160.330 ;
        RECT 89.720 160.145 90.070 160.190 ;
        RECT 101.850 160.145 102.140 160.190 ;
        RECT 103.535 160.145 103.825 160.190 ;
        RECT 105.910 160.190 122.150 160.330 ;
        RECT 89.720 160.130 90.040 160.145 ;
        RECT 77.315 159.805 77.605 160.035 ;
        RECT 77.760 159.990 78.080 160.050 ;
        RECT 78.235 159.990 78.525 160.035 ;
        RECT 77.760 159.850 78.525 159.990 ;
        RECT 77.760 159.790 78.080 159.850 ;
        RECT 78.235 159.805 78.525 159.850 ;
        RECT 78.695 159.990 78.985 160.035 ;
        RECT 81.900 159.990 82.220 160.050 ;
        RECT 78.695 159.850 82.220 159.990 ;
        RECT 78.695 159.805 78.985 159.850 ;
        RECT 81.900 159.790 82.220 159.850 ;
        RECT 83.740 159.790 84.060 160.050 ;
        RECT 90.640 159.990 90.960 160.050 ;
        RECT 91.115 159.990 91.405 160.035 ;
        RECT 90.640 159.850 91.405 159.990 ;
        RECT 90.640 159.790 90.960 159.850 ;
        RECT 91.115 159.805 91.405 159.850 ;
        RECT 102.600 159.990 102.920 160.050 ;
        RECT 103.075 159.990 103.365 160.035 ;
        RECT 102.600 159.850 103.365 159.990 ;
        RECT 102.600 159.790 102.920 159.850 ;
        RECT 103.075 159.805 103.365 159.850 ;
        RECT 104.455 159.805 104.745 160.035 ;
        RECT 80.060 159.650 80.380 159.710 ;
        RECT 75.550 159.510 80.380 159.650 ;
        RECT 80.060 159.450 80.380 159.510 ;
        RECT 86.525 159.650 86.815 159.695 ;
        RECT 89.045 159.650 89.335 159.695 ;
        RECT 90.235 159.650 90.525 159.695 ;
        RECT 86.525 159.510 90.525 159.650 ;
        RECT 86.525 159.465 86.815 159.510 ;
        RECT 89.045 159.465 89.335 159.510 ;
        RECT 90.235 159.465 90.525 159.510 ;
        RECT 98.485 159.650 98.775 159.695 ;
        RECT 101.005 159.650 101.295 159.695 ;
        RECT 102.195 159.650 102.485 159.695 ;
        RECT 98.485 159.510 102.485 159.650 ;
        RECT 104.530 159.650 104.670 159.805 ;
        RECT 104.900 159.790 105.220 160.050 ;
        RECT 105.910 159.695 106.050 160.190 ;
        RECT 113.195 160.145 113.485 160.190 ;
        RECT 106.295 159.990 106.585 160.035 ;
        RECT 107.200 159.990 107.520 160.050 ;
        RECT 106.295 159.850 107.520 159.990 ;
        RECT 106.295 159.805 106.585 159.850 ;
        RECT 107.200 159.790 107.520 159.850 ;
        RECT 109.960 159.790 110.280 160.050 ;
        RECT 111.340 159.990 111.660 160.050 ;
        RECT 112.275 159.990 112.565 160.035 ;
        RECT 111.340 159.850 112.565 159.990 ;
        RECT 111.340 159.790 111.660 159.850 ;
        RECT 112.275 159.805 112.565 159.850 ;
        RECT 112.720 159.790 113.040 160.050 ;
        RECT 113.655 159.805 113.945 160.035 ;
        RECT 114.115 159.805 114.405 160.035 ;
        RECT 104.530 159.510 105.130 159.650 ;
        RECT 98.485 159.465 98.775 159.510 ;
        RECT 101.005 159.465 101.295 159.510 ;
        RECT 102.195 159.465 102.485 159.510 ;
        RECT 54.775 159.170 57.750 159.310 ;
        RECT 48.335 159.125 48.625 159.170 ;
        RECT 54.775 159.125 55.065 159.170 ;
        RECT 38.675 158.970 38.965 159.015 ;
        RECT 49.240 158.970 49.560 159.030 ;
        RECT 38.675 158.830 49.560 158.970 ;
        RECT 38.675 158.785 38.965 158.830 ;
        RECT 49.240 158.770 49.560 158.830 ;
        RECT 50.635 158.970 50.925 159.015 ;
        RECT 54.300 158.970 54.620 159.030 ;
        RECT 50.635 158.830 54.620 158.970 ;
        RECT 57.610 158.970 57.750 159.170 ;
        RECT 57.980 159.170 61.940 159.310 ;
        RECT 57.980 159.125 58.270 159.170 ;
        RECT 59.550 159.125 59.840 159.170 ;
        RECT 61.650 159.125 61.940 159.170 ;
        RECT 62.670 159.170 63.270 159.310 ;
        RECT 73.175 159.310 73.465 159.355 ;
        RECT 76.380 159.310 76.700 159.370 ;
        RECT 73.175 159.170 76.700 159.310 ;
        RECT 62.120 158.970 62.440 159.030 ;
        RECT 62.670 159.015 62.810 159.170 ;
        RECT 73.175 159.125 73.465 159.170 ;
        RECT 76.380 159.110 76.700 159.170 ;
        RECT 86.960 159.310 87.250 159.355 ;
        RECT 88.530 159.310 88.820 159.355 ;
        RECT 90.630 159.310 90.920 159.355 ;
        RECT 86.960 159.170 90.920 159.310 ;
        RECT 86.960 159.125 87.250 159.170 ;
        RECT 88.530 159.125 88.820 159.170 ;
        RECT 90.630 159.125 90.920 159.170 ;
        RECT 98.920 159.310 99.210 159.355 ;
        RECT 100.490 159.310 100.780 159.355 ;
        RECT 102.590 159.310 102.880 159.355 ;
        RECT 98.920 159.170 102.880 159.310 ;
        RECT 98.920 159.125 99.210 159.170 ;
        RECT 100.490 159.125 100.780 159.170 ;
        RECT 102.590 159.125 102.880 159.170 ;
        RECT 57.610 158.830 62.440 158.970 ;
        RECT 50.635 158.785 50.925 158.830 ;
        RECT 54.300 158.770 54.620 158.830 ;
        RECT 62.120 158.770 62.440 158.830 ;
        RECT 62.595 158.785 62.885 159.015 ;
        RECT 71.320 158.970 71.640 159.030 ;
        RECT 74.095 158.970 74.385 159.015 ;
        RECT 71.320 158.830 74.385 158.970 ;
        RECT 71.320 158.770 71.640 158.830 ;
        RECT 74.095 158.785 74.385 158.830 ;
        RECT 74.540 158.970 74.860 159.030 ;
        RECT 81.915 158.970 82.205 159.015 ;
        RECT 74.540 158.830 82.205 158.970 ;
        RECT 74.540 158.770 74.860 158.830 ;
        RECT 81.915 158.785 82.205 158.830 ;
        RECT 96.160 158.770 96.480 159.030 ;
        RECT 104.990 158.970 105.130 159.510 ;
        RECT 105.835 159.465 106.125 159.695 ;
        RECT 109.040 159.650 109.360 159.710 ;
        RECT 111.815 159.650 112.105 159.695 ;
        RECT 112.810 159.650 112.950 159.790 ;
        RECT 109.040 159.510 112.950 159.650 ;
        RECT 113.180 159.650 113.500 159.710 ;
        RECT 113.730 159.650 113.870 159.805 ;
        RECT 113.180 159.510 113.870 159.650 ;
        RECT 114.190 159.650 114.330 159.805 ;
        RECT 114.560 159.790 114.880 160.050 ;
        RECT 115.035 159.805 115.325 160.035 ;
        RECT 115.110 159.650 115.250 159.805 ;
        RECT 115.480 159.790 115.800 160.050 ;
        RECT 116.400 159.790 116.720 160.050 ;
        RECT 119.160 159.990 119.480 160.050 ;
        RECT 119.635 159.990 119.925 160.035 ;
        RECT 117.410 159.850 119.925 159.990 ;
        RECT 115.955 159.650 116.245 159.695 ;
        RECT 117.410 159.650 117.550 159.850 ;
        RECT 119.160 159.790 119.480 159.850 ;
        RECT 119.635 159.805 119.925 159.850 ;
        RECT 120.080 159.790 120.400 160.050 ;
        RECT 121.000 159.790 121.320 160.050 ;
        RECT 121.475 159.805 121.765 160.035 ;
        RECT 114.190 159.510 114.790 159.650 ;
        RECT 115.110 159.510 117.550 159.650 ;
        RECT 109.040 159.450 109.360 159.510 ;
        RECT 111.815 159.465 112.105 159.510 ;
        RECT 113.180 159.450 113.500 159.510 ;
        RECT 112.260 159.310 112.580 159.370 ;
        RECT 114.650 159.310 114.790 159.510 ;
        RECT 115.955 159.465 116.245 159.510 ;
        RECT 117.780 159.450 118.100 159.710 ;
        RECT 121.550 159.650 121.690 159.805 ;
        RECT 121.090 159.510 121.690 159.650 ;
        RECT 122.010 159.650 122.150 160.190 ;
        RECT 127.455 160.190 130.890 160.330 ;
        RECT 127.455 160.145 127.745 160.190 ;
        RECT 130.750 160.050 130.890 160.190 ;
        RECT 132.010 160.190 134.200 160.330 ;
        RECT 132.010 160.145 132.300 160.190 ;
        RECT 133.880 160.130 134.200 160.190 ;
        RECT 123.300 159.790 123.620 160.050 ;
        RECT 125.600 159.990 125.920 160.050 ;
        RECT 128.375 159.990 128.665 160.035 ;
        RECT 125.600 159.850 128.665 159.990 ;
        RECT 125.600 159.790 125.920 159.850 ;
        RECT 128.375 159.805 128.665 159.850 ;
        RECT 129.295 159.805 129.585 160.035 ;
        RECT 129.370 159.650 129.510 159.805 ;
        RECT 130.660 159.790 130.980 160.050 ;
        RECT 138.035 159.990 138.325 160.035 ;
        RECT 138.480 159.990 138.800 160.050 ;
        RECT 138.035 159.850 138.800 159.990 ;
        RECT 138.035 159.805 138.325 159.850 ;
        RECT 138.480 159.790 138.800 159.850 ;
        RECT 139.860 159.790 140.180 160.050 ;
        RECT 122.010 159.510 129.510 159.650 ;
        RECT 131.555 159.650 131.845 159.695 ;
        RECT 132.745 159.650 133.035 159.695 ;
        RECT 135.265 159.650 135.555 159.695 ;
        RECT 131.555 159.510 135.555 159.650 ;
        RECT 112.260 159.170 118.470 159.310 ;
        RECT 112.260 159.110 112.580 159.170 ;
        RECT 118.330 159.030 118.470 159.170 ;
        RECT 118.700 159.110 119.020 159.370 ;
        RECT 121.090 159.310 121.230 159.510 ;
        RECT 131.555 159.465 131.845 159.510 ;
        RECT 132.745 159.465 133.035 159.510 ;
        RECT 135.265 159.465 135.555 159.510 ;
        RECT 121.460 159.310 121.780 159.370 ;
        RECT 125.600 159.310 125.920 159.370 ;
        RECT 121.090 159.170 125.920 159.310 ;
        RECT 121.460 159.110 121.780 159.170 ;
        RECT 125.600 159.110 125.920 159.170 ;
        RECT 131.160 159.310 131.450 159.355 ;
        RECT 133.260 159.310 133.550 159.355 ;
        RECT 134.830 159.310 135.120 159.355 ;
        RECT 131.160 159.170 135.120 159.310 ;
        RECT 131.160 159.125 131.450 159.170 ;
        RECT 133.260 159.125 133.550 159.170 ;
        RECT 134.830 159.125 135.120 159.170 ;
        RECT 114.100 158.970 114.420 159.030 ;
        RECT 104.990 158.830 114.420 158.970 ;
        RECT 114.100 158.770 114.420 158.830 ;
        RECT 118.240 158.970 118.560 159.030 ;
        RECT 120.080 158.970 120.400 159.030 ;
        RECT 121.015 158.970 121.305 159.015 ;
        RECT 118.240 158.830 121.305 158.970 ;
        RECT 118.240 158.770 118.560 158.830 ;
        RECT 120.080 158.770 120.400 158.830 ;
        RECT 121.015 158.785 121.305 158.830 ;
        RECT 122.380 158.970 122.700 159.030 ;
        RECT 122.855 158.970 123.145 159.015 ;
        RECT 122.380 158.830 123.145 158.970 ;
        RECT 122.380 158.770 122.700 158.830 ;
        RECT 122.855 158.785 123.145 158.830 ;
        RECT 140.780 158.770 141.100 159.030 ;
        RECT 17.430 158.150 143.010 158.630 ;
        RECT 25.780 157.950 26.100 158.010 ;
        RECT 26.715 157.950 27.005 157.995 ;
        RECT 31.760 157.950 32.080 158.010 ;
        RECT 25.780 157.810 32.080 157.950 ;
        RECT 25.780 157.750 26.100 157.810 ;
        RECT 26.715 157.765 27.005 157.810 ;
        RECT 31.760 157.750 32.080 157.810 ;
        RECT 38.660 157.950 38.980 158.010 ;
        RECT 39.135 157.950 39.425 157.995 ;
        RECT 46.020 157.950 46.340 158.010 ;
        RECT 38.660 157.810 39.425 157.950 ;
        RECT 38.660 157.750 38.980 157.810 ;
        RECT 39.135 157.765 39.425 157.810 ;
        RECT 39.655 157.810 46.340 157.950 ;
        RECT 20.300 157.610 20.590 157.655 ;
        RECT 22.400 157.610 22.690 157.655 ;
        RECT 23.970 157.610 24.260 157.655 ;
        RECT 20.300 157.470 24.260 157.610 ;
        RECT 20.300 157.425 20.590 157.470 ;
        RECT 22.400 157.425 22.690 157.470 ;
        RECT 23.970 157.425 24.260 157.470 ;
        RECT 32.680 157.610 33.000 157.670 ;
        RECT 39.655 157.610 39.795 157.810 ;
        RECT 46.020 157.750 46.340 157.810 ;
        RECT 46.480 157.950 46.800 158.010 ;
        RECT 49.255 157.950 49.545 157.995 ;
        RECT 46.480 157.810 49.545 157.950 ;
        RECT 46.480 157.750 46.800 157.810 ;
        RECT 49.255 157.765 49.545 157.810 ;
        RECT 55.235 157.950 55.525 157.995 ;
        RECT 60.280 157.950 60.600 158.010 ;
        RECT 55.235 157.810 60.600 157.950 ;
        RECT 55.235 157.765 55.525 157.810 ;
        RECT 60.280 157.750 60.600 157.810 ;
        RECT 74.095 157.950 74.385 157.995 ;
        RECT 74.540 157.950 74.860 158.010 ;
        RECT 74.095 157.810 74.860 157.950 ;
        RECT 74.095 157.765 74.385 157.810 ;
        RECT 74.540 157.750 74.860 157.810 ;
        RECT 75.000 157.750 75.320 158.010 ;
        RECT 77.775 157.950 78.065 157.995 ;
        RECT 78.680 157.950 79.000 158.010 ;
        RECT 77.775 157.810 79.000 157.950 ;
        RECT 77.775 157.765 78.065 157.810 ;
        RECT 78.680 157.750 79.000 157.810 ;
        RECT 82.360 157.750 82.680 158.010 ;
        RECT 87.880 157.950 88.200 158.010 ;
        RECT 87.880 157.810 92.250 157.950 ;
        RECT 87.880 157.750 88.200 157.810 ;
        RECT 32.680 157.470 39.795 157.610 ;
        RECT 43.735 157.610 44.025 157.655 ;
        RECT 47.860 157.610 48.180 157.670 ;
        RECT 43.735 157.470 48.180 157.610 ;
        RECT 32.680 157.410 33.000 157.470 ;
        RECT 43.735 157.425 44.025 157.470 ;
        RECT 47.860 157.410 48.180 157.470 ;
        RECT 50.620 157.610 50.940 157.670 ;
        RECT 50.620 157.470 52.230 157.610 ;
        RECT 50.620 157.410 50.940 157.470 ;
        RECT 20.695 157.270 20.985 157.315 ;
        RECT 21.885 157.270 22.175 157.315 ;
        RECT 24.405 157.270 24.695 157.315 ;
        RECT 43.260 157.270 43.580 157.330 ;
        RECT 47.415 157.270 47.705 157.315 ;
        RECT 48.780 157.270 49.100 157.330 ;
        RECT 52.090 157.315 52.230 157.470 ;
        RECT 56.600 157.410 56.920 157.670 ;
        RECT 59.360 157.610 59.650 157.655 ;
        RECT 60.930 157.610 61.220 157.655 ;
        RECT 63.030 157.610 63.320 157.655 ;
        RECT 59.360 157.470 63.320 157.610 ;
        RECT 59.360 157.425 59.650 157.470 ;
        RECT 60.930 157.425 61.220 157.470 ;
        RECT 63.030 157.425 63.320 157.470 ;
        RECT 72.240 157.410 72.560 157.670 ;
        RECT 20.695 157.130 24.695 157.270 ;
        RECT 20.695 157.085 20.985 157.130 ;
        RECT 21.885 157.085 22.175 157.130 ;
        RECT 24.405 157.085 24.695 157.130 ;
        RECT 40.130 157.130 46.250 157.270 ;
        RECT 19.815 156.930 20.105 156.975 ;
        RECT 23.480 156.930 23.800 156.990 ;
        RECT 19.815 156.790 23.800 156.930 ;
        RECT 19.815 156.745 20.105 156.790 ;
        RECT 23.480 156.730 23.800 156.790 ;
        RECT 31.760 156.930 32.080 156.990 ;
        RECT 40.130 156.975 40.270 157.130 ;
        RECT 43.260 157.070 43.580 157.130 ;
        RECT 31.760 156.790 33.370 156.930 ;
        RECT 31.760 156.730 32.080 156.790 ;
        RECT 21.150 156.590 21.440 156.635 ;
        RECT 21.640 156.590 21.960 156.650 ;
        RECT 21.150 156.450 21.960 156.590 ;
        RECT 21.150 156.405 21.440 156.450 ;
        RECT 21.640 156.390 21.960 156.450 ;
        RECT 32.680 156.390 33.000 156.650 ;
        RECT 33.230 156.590 33.370 156.790 ;
        RECT 40.055 156.745 40.345 156.975 ;
        RECT 40.960 156.730 41.280 156.990 ;
        RECT 41.435 156.745 41.725 156.975 ;
        RECT 41.510 156.590 41.650 156.745 ;
        RECT 44.640 156.730 44.960 156.990 ;
        RECT 45.115 156.930 45.405 156.975 ;
        RECT 46.110 156.930 46.250 157.130 ;
        RECT 47.415 157.130 50.265 157.270 ;
        RECT 47.415 157.085 47.705 157.130 ;
        RECT 48.780 157.070 49.100 157.130 ;
        RECT 46.955 156.930 47.245 156.975 ;
        RECT 45.115 156.790 45.790 156.930 ;
        RECT 46.110 156.790 47.245 156.930 ;
        RECT 45.115 156.745 45.405 156.790 ;
        RECT 33.230 156.450 41.650 156.590 ;
        RECT 32.235 156.250 32.525 156.295 ;
        RECT 34.060 156.250 34.380 156.310 ;
        RECT 32.235 156.110 34.380 156.250 ;
        RECT 45.650 156.250 45.790 156.790 ;
        RECT 46.955 156.745 47.245 156.790 ;
        RECT 47.860 156.730 48.180 156.990 ;
        RECT 48.320 156.730 48.640 156.990 ;
        RECT 50.125 156.975 50.265 157.130 ;
        RECT 52.015 157.085 52.305 157.315 ;
        RECT 53.380 157.270 53.700 157.330 ;
        RECT 53.855 157.270 54.145 157.315 ;
        RECT 53.380 157.130 54.145 157.270 ;
        RECT 53.380 157.070 53.700 157.130 ;
        RECT 53.855 157.085 54.145 157.130 ;
        RECT 54.440 157.270 54.730 157.315 ;
        RECT 55.680 157.270 56.000 157.330 ;
        RECT 54.440 157.130 56.000 157.270 ;
        RECT 54.440 157.085 54.730 157.130 ;
        RECT 55.680 157.070 56.000 157.130 ;
        RECT 58.925 157.270 59.215 157.315 ;
        RECT 61.445 157.270 61.735 157.315 ;
        RECT 62.635 157.270 62.925 157.315 ;
        RECT 58.925 157.130 62.925 157.270 ;
        RECT 74.630 157.270 74.770 157.750 ;
        RECT 77.315 157.425 77.605 157.655 ;
        RECT 75.475 157.270 75.765 157.315 ;
        RECT 74.630 157.130 75.765 157.270 ;
        RECT 58.925 157.085 59.215 157.130 ;
        RECT 61.445 157.085 61.735 157.130 ;
        RECT 62.635 157.085 62.925 157.130 ;
        RECT 75.475 157.085 75.765 157.130 ;
        RECT 49.835 156.790 50.265 156.975 ;
        RECT 50.635 156.930 50.925 156.975 ;
        RECT 51.540 156.930 51.860 156.990 ;
        RECT 50.635 156.790 51.860 156.930 ;
        RECT 49.835 156.745 50.125 156.790 ;
        RECT 50.635 156.745 50.925 156.790 ;
        RECT 51.540 156.730 51.860 156.790 ;
        RECT 62.120 156.975 62.440 156.990 ;
        RECT 62.120 156.930 62.470 156.975 ;
        RECT 63.040 156.930 63.360 156.990 ;
        RECT 63.515 156.930 63.805 156.975 ;
        RECT 70.875 156.930 71.165 156.975 ;
        RECT 62.120 156.790 62.635 156.930 ;
        RECT 63.040 156.790 63.805 156.930 ;
        RECT 62.120 156.745 62.470 156.790 ;
        RECT 62.120 156.730 62.440 156.745 ;
        RECT 63.040 156.730 63.360 156.790 ;
        RECT 63.515 156.745 63.805 156.790 ;
        RECT 66.810 156.790 71.165 156.930 ;
        RECT 46.035 156.590 46.325 156.635 ;
        RECT 53.395 156.590 53.685 156.635 ;
        RECT 55.220 156.590 55.540 156.650 ;
        RECT 46.035 156.450 49.930 156.590 ;
        RECT 46.035 156.405 46.325 156.450 ;
        RECT 49.790 156.310 49.930 156.450 ;
        RECT 53.395 156.450 55.540 156.590 ;
        RECT 63.590 156.590 63.730 156.745 ;
        RECT 66.810 156.650 66.950 156.790 ;
        RECT 70.875 156.745 71.165 156.790 ;
        RECT 64.895 156.590 65.185 156.635 ;
        RECT 66.720 156.590 67.040 156.650 ;
        RECT 63.590 156.450 67.040 156.590 ;
        RECT 53.395 156.405 53.685 156.450 ;
        RECT 55.220 156.390 55.540 156.450 ;
        RECT 64.895 156.405 65.185 156.450 ;
        RECT 66.720 156.390 67.040 156.450 ;
        RECT 67.180 156.390 67.500 156.650 ;
        RECT 77.390 156.590 77.530 157.425 ;
        RECT 78.695 157.270 78.985 157.315 ;
        RECT 82.450 157.270 82.590 157.750 ;
        RECT 85.120 157.610 85.410 157.655 ;
        RECT 86.690 157.610 86.980 157.655 ;
        RECT 88.790 157.610 89.080 157.655 ;
        RECT 85.120 157.470 89.080 157.610 ;
        RECT 92.110 157.610 92.250 157.810 ;
        RECT 101.220 157.750 101.540 158.010 ;
        RECT 108.580 157.750 108.900 158.010 ;
        RECT 110.880 157.950 111.200 158.010 ;
        RECT 114.560 157.950 114.880 158.010 ;
        RECT 110.880 157.810 114.880 157.950 ;
        RECT 110.880 157.750 111.200 157.810 ;
        RECT 114.560 157.750 114.880 157.810 ;
        RECT 116.860 157.950 117.180 158.010 ;
        RECT 118.240 157.950 118.560 158.010 ;
        RECT 116.860 157.810 118.560 157.950 ;
        RECT 116.860 157.750 117.180 157.810 ;
        RECT 118.240 157.750 118.560 157.810 ;
        RECT 119.635 157.950 119.925 157.995 ;
        RECT 129.740 157.950 130.060 158.010 ;
        RECT 119.635 157.810 130.060 157.950 ;
        RECT 119.635 157.765 119.925 157.810 ;
        RECT 129.740 157.750 130.060 157.810 ;
        RECT 98.000 157.610 98.320 157.670 ;
        RECT 123.300 157.610 123.620 157.670 ;
        RECT 92.110 157.470 92.710 157.610 ;
        RECT 85.120 157.425 85.410 157.470 ;
        RECT 86.690 157.425 86.980 157.470 ;
        RECT 88.790 157.425 89.080 157.470 ;
        RECT 92.570 157.330 92.710 157.470 ;
        RECT 96.710 157.470 123.620 157.610 ;
        RECT 78.695 157.130 82.590 157.270 ;
        RECT 84.685 157.270 84.975 157.315 ;
        RECT 87.205 157.270 87.495 157.315 ;
        RECT 88.395 157.270 88.685 157.315 ;
        RECT 92.035 157.270 92.325 157.315 ;
        RECT 84.685 157.130 88.685 157.270 ;
        RECT 78.695 157.085 78.985 157.130 ;
        RECT 84.685 157.085 84.975 157.130 ;
        RECT 87.205 157.085 87.495 157.130 ;
        RECT 88.395 157.085 88.685 157.130 ;
        RECT 88.890 157.130 92.325 157.270 ;
        RECT 81.455 156.930 81.745 156.975 ;
        RECT 88.890 156.930 89.030 157.130 ;
        RECT 92.035 157.085 92.325 157.130 ;
        RECT 92.480 157.070 92.800 157.330 ;
        RECT 81.455 156.790 89.030 156.930 ;
        RECT 81.455 156.745 81.745 156.790 ;
        RECT 89.260 156.730 89.580 156.990 ;
        RECT 94.780 156.930 95.100 156.990 ;
        RECT 96.175 156.930 96.465 156.975 ;
        RECT 96.710 156.930 96.850 157.470 ;
        RECT 98.000 157.410 98.320 157.470 ;
        RECT 123.300 157.410 123.620 157.470 ;
        RECT 103.520 157.070 103.840 157.330 ;
        RECT 103.995 157.085 104.285 157.315 ;
        RECT 94.780 156.790 96.850 156.930 ;
        RECT 98.460 156.930 98.780 156.990 ;
        RECT 101.220 156.930 101.540 156.990 ;
        RECT 104.070 156.930 104.210 157.085 ;
        RECT 109.500 157.070 109.820 157.330 ;
        RECT 116.400 157.270 116.720 157.330 ;
        RECT 117.795 157.270 118.085 157.315 ;
        RECT 120.080 157.270 120.400 157.330 ;
        RECT 116.400 157.130 118.085 157.270 ;
        RECT 116.400 157.070 116.720 157.130 ;
        RECT 117.795 157.085 118.085 157.130 ;
        RECT 118.330 157.130 120.400 157.270 ;
        RECT 98.460 156.790 104.210 156.930 ;
        RECT 108.120 156.930 108.440 156.990 ;
        RECT 110.435 156.930 110.725 156.975 ;
        RECT 108.120 156.790 115.710 156.930 ;
        RECT 94.780 156.730 95.100 156.790 ;
        RECT 96.175 156.745 96.465 156.790 ;
        RECT 98.460 156.730 98.780 156.790 ;
        RECT 101.220 156.730 101.540 156.790 ;
        RECT 108.120 156.730 108.440 156.790 ;
        RECT 110.435 156.745 110.725 156.790 ;
        RECT 84.660 156.590 84.980 156.650 ;
        RECT 77.390 156.450 84.980 156.590 ;
        RECT 84.660 156.390 84.980 156.450 ;
        RECT 88.050 156.590 88.340 156.635 ;
        RECT 88.050 156.450 89.950 156.590 ;
        RECT 88.050 156.405 88.340 156.450 ;
        RECT 47.860 156.250 48.180 156.310 ;
        RECT 45.650 156.110 48.180 156.250 ;
        RECT 32.235 156.065 32.525 156.110 ;
        RECT 34.060 156.050 34.380 156.110 ;
        RECT 47.860 156.050 48.180 156.110 ;
        RECT 49.700 156.050 50.020 156.310 ;
        RECT 50.160 156.050 50.480 156.310 ;
        RECT 74.080 156.050 74.400 156.310 ;
        RECT 89.810 156.295 89.950 156.450 ;
        RECT 99.840 156.390 100.160 156.650 ;
        RECT 89.735 156.065 90.025 156.295 ;
        RECT 91.560 156.050 91.880 156.310 ;
        RECT 103.060 156.050 103.380 156.310 ;
        RECT 109.515 156.250 109.805 156.295 ;
        RECT 110.420 156.250 110.740 156.310 ;
        RECT 109.515 156.110 110.740 156.250 ;
        RECT 115.570 156.250 115.710 156.790 ;
        RECT 115.955 156.745 116.245 156.975 ;
        RECT 116.030 156.590 116.170 156.745 ;
        RECT 116.860 156.730 117.180 156.990 ;
        RECT 117.335 156.940 117.625 156.975 ;
        RECT 118.330 156.940 118.470 157.130 ;
        RECT 120.080 157.070 120.400 157.130 ;
        RECT 133.420 157.270 133.740 157.330 ;
        RECT 136.655 157.270 136.945 157.315 ;
        RECT 133.420 157.130 136.945 157.270 ;
        RECT 133.420 157.070 133.740 157.130 ;
        RECT 136.655 157.085 136.945 157.130 ;
        RECT 117.335 156.800 118.470 156.940 ;
        RECT 118.715 156.930 119.005 156.975 ;
        RECT 119.620 156.930 119.940 156.990 ;
        RECT 117.335 156.745 117.625 156.800 ;
        RECT 118.715 156.790 119.940 156.930 ;
        RECT 118.715 156.745 119.005 156.790 ;
        RECT 119.620 156.730 119.940 156.790 ;
        RECT 120.540 156.930 120.860 156.990 ;
        RECT 121.015 156.930 121.305 156.975 ;
        RECT 120.540 156.790 121.305 156.930 ;
        RECT 120.540 156.730 120.860 156.790 ;
        RECT 121.015 156.745 121.305 156.790 ;
        RECT 121.460 156.730 121.780 156.990 ;
        RECT 123.315 156.930 123.605 156.975 ;
        RECT 130.660 156.930 130.980 156.990 ;
        RECT 123.315 156.790 130.980 156.930 ;
        RECT 123.315 156.745 123.605 156.790 ;
        RECT 130.660 156.730 130.980 156.790 ;
        RECT 137.560 156.930 137.880 156.990 ;
        RECT 140.795 156.930 141.085 156.975 ;
        RECT 137.560 156.790 141.085 156.930 ;
        RECT 137.560 156.730 137.880 156.790 ;
        RECT 140.795 156.745 141.085 156.790 ;
        RECT 117.780 156.590 118.100 156.650 ;
        RECT 116.030 156.450 118.100 156.590 ;
        RECT 117.780 156.390 118.100 156.450 ;
        RECT 118.240 156.590 118.560 156.650 ;
        RECT 120.095 156.590 120.385 156.635 ;
        RECT 121.550 156.590 121.690 156.730 ;
        RECT 118.240 156.450 120.385 156.590 ;
        RECT 118.240 156.390 118.560 156.450 ;
        RECT 120.095 156.405 120.385 156.450 ;
        RECT 120.630 156.450 121.690 156.590 ;
        RECT 135.735 156.590 136.025 156.635 ;
        RECT 138.035 156.590 138.325 156.635 ;
        RECT 135.735 156.450 138.325 156.590 ;
        RECT 120.630 156.250 120.770 156.450 ;
        RECT 135.735 156.405 136.025 156.450 ;
        RECT 138.035 156.405 138.325 156.450 ;
        RECT 115.570 156.110 120.770 156.250 ;
        RECT 109.515 156.065 109.805 156.110 ;
        RECT 110.420 156.050 110.740 156.110 ;
        RECT 121.460 156.050 121.780 156.310 ;
        RECT 132.040 156.250 132.360 156.310 ;
        RECT 133.895 156.250 134.185 156.295 ;
        RECT 132.040 156.110 134.185 156.250 ;
        RECT 132.040 156.050 132.360 156.110 ;
        RECT 133.895 156.065 134.185 156.110 ;
        RECT 134.340 156.250 134.660 156.310 ;
        RECT 136.195 156.250 136.485 156.295 ;
        RECT 134.340 156.110 136.485 156.250 ;
        RECT 134.340 156.050 134.660 156.110 ;
        RECT 136.195 156.065 136.485 156.110 ;
        RECT 17.430 155.430 143.010 155.910 ;
        RECT 30.840 155.230 31.160 155.290 ;
        RECT 27.710 155.090 31.160 155.230 ;
        RECT 27.710 154.595 27.850 155.090 ;
        RECT 30.840 155.030 31.160 155.090 ;
        RECT 34.980 155.030 35.300 155.290 ;
        RECT 48.335 155.045 48.625 155.275 ;
        RECT 53.395 155.230 53.685 155.275 ;
        RECT 54.760 155.230 55.080 155.290 ;
        RECT 53.395 155.090 55.080 155.230 ;
        RECT 53.395 155.045 53.685 155.090 ;
        RECT 48.410 154.890 48.550 155.045 ;
        RECT 54.760 155.030 55.080 155.090 ;
        RECT 67.180 155.230 67.500 155.290 ;
        RECT 85.580 155.230 85.900 155.290 ;
        RECT 94.780 155.230 95.100 155.290 ;
        RECT 117.320 155.230 117.640 155.290 ;
        RECT 67.180 155.090 95.100 155.230 ;
        RECT 67.180 155.030 67.500 155.090 ;
        RECT 85.580 155.030 85.900 155.090 ;
        RECT 94.780 155.030 95.100 155.090 ;
        RECT 110.050 155.090 117.640 155.230 ;
        RECT 48.795 154.890 49.085 154.935 ;
        RECT 96.175 154.890 96.465 154.935 ;
        RECT 96.620 154.890 96.940 154.950 ;
        RECT 99.840 154.890 100.160 154.950 ;
        RECT 28.170 154.750 34.140 154.890 ;
        RECT 48.410 154.750 49.085 154.890 ;
        RECT 27.635 154.365 27.925 154.595 ;
        RECT 28.170 154.255 28.310 154.750 ;
        RECT 34.000 154.610 34.140 154.750 ;
        RECT 48.795 154.705 49.085 154.750 ;
        RECT 49.330 154.750 50.390 154.890 ;
        RECT 30.840 154.550 31.160 154.610 ;
        RECT 34.000 154.595 34.380 154.610 ;
        RECT 33.155 154.550 33.445 154.595 ;
        RECT 30.840 154.410 33.445 154.550 ;
        RECT 30.840 154.350 31.160 154.410 ;
        RECT 33.155 154.365 33.445 154.410 ;
        RECT 33.925 154.550 34.380 154.595 ;
        RECT 43.260 154.550 43.580 154.610 ;
        RECT 33.925 154.410 43.580 154.550 ;
        RECT 33.925 154.365 34.380 154.410 ;
        RECT 28.095 154.025 28.385 154.255 ;
        RECT 29.475 154.210 29.765 154.255 ;
        RECT 31.300 154.210 31.620 154.270 ;
        RECT 29.475 154.070 31.620 154.210 ;
        RECT 33.230 154.210 33.370 154.365 ;
        RECT 34.060 154.350 34.380 154.365 ;
        RECT 43.260 154.350 43.580 154.410 ;
        RECT 43.720 154.350 44.040 154.610 ;
        RECT 46.495 154.550 46.785 154.595 ;
        RECT 47.400 154.550 47.720 154.610 ;
        RECT 46.495 154.410 47.720 154.550 ;
        RECT 46.495 154.365 46.785 154.410 ;
        RECT 47.400 154.350 47.720 154.410 ;
        RECT 47.860 154.550 48.180 154.610 ;
        RECT 49.330 154.550 49.470 154.750 ;
        RECT 47.860 154.410 49.470 154.550 ;
        RECT 47.860 154.350 48.180 154.410 ;
        RECT 49.700 154.350 50.020 154.610 ;
        RECT 50.250 154.595 50.390 154.750 ;
        RECT 91.190 154.750 100.160 154.890 ;
        RECT 50.175 154.550 50.465 154.595 ;
        RECT 55.235 154.550 55.525 154.595 ;
        RECT 56.600 154.550 56.920 154.610 ;
        RECT 70.860 154.595 71.180 154.610 ;
        RECT 50.175 154.410 56.920 154.550 ;
        RECT 50.175 154.365 50.465 154.410 ;
        RECT 55.235 154.365 55.525 154.410 ;
        RECT 56.600 154.350 56.920 154.410 ;
        RECT 70.830 154.365 71.180 154.595 ;
        RECT 70.860 154.350 71.180 154.365 ;
        RECT 76.380 154.550 76.700 154.610 ;
        RECT 79.615 154.550 79.905 154.595 ;
        RECT 76.380 154.410 79.905 154.550 ;
        RECT 76.380 154.350 76.700 154.410 ;
        RECT 79.615 154.365 79.905 154.410 ;
        RECT 87.995 154.550 88.285 154.595 ;
        RECT 89.260 154.550 89.580 154.610 ;
        RECT 91.190 154.550 91.330 154.750 ;
        RECT 96.175 154.705 96.465 154.750 ;
        RECT 96.620 154.690 96.940 154.750 ;
        RECT 99.840 154.690 100.160 154.750 ;
        RECT 103.075 154.890 103.365 154.935 ;
        RECT 103.980 154.890 104.300 154.950 ;
        RECT 103.075 154.750 104.300 154.890 ;
        RECT 103.075 154.705 103.365 154.750 ;
        RECT 103.980 154.690 104.300 154.750 ;
        RECT 107.675 154.890 107.965 154.935 ;
        RECT 109.040 154.890 109.360 154.950 ;
        RECT 107.675 154.750 109.360 154.890 ;
        RECT 107.675 154.705 107.965 154.750 ;
        RECT 109.040 154.690 109.360 154.750 ;
        RECT 87.995 154.410 89.030 154.550 ;
        RECT 87.995 154.365 88.285 154.410 ;
        RECT 42.800 154.210 43.120 154.270 ;
        RECT 43.810 154.210 43.950 154.350 ;
        RECT 33.230 154.070 43.950 154.210 ;
        RECT 46.955 154.210 47.245 154.255 ;
        RECT 51.540 154.210 51.860 154.270 ;
        RECT 46.955 154.070 51.860 154.210 ;
        RECT 29.475 154.025 29.765 154.070 ;
        RECT 31.300 154.010 31.620 154.070 ;
        RECT 42.800 154.010 43.120 154.070 ;
        RECT 46.955 154.025 47.245 154.070 ;
        RECT 51.540 154.010 51.860 154.070 ;
        RECT 54.300 154.210 54.620 154.270 ;
        RECT 54.775 154.210 55.065 154.255 ;
        RECT 54.300 154.070 55.065 154.210 ;
        RECT 54.300 154.010 54.620 154.070 ;
        RECT 54.775 154.025 55.065 154.070 ;
        RECT 66.720 154.210 67.040 154.270 ;
        RECT 69.495 154.210 69.785 154.255 ;
        RECT 66.720 154.070 69.785 154.210 ;
        RECT 66.720 154.010 67.040 154.070 ;
        RECT 69.495 154.025 69.785 154.070 ;
        RECT 70.375 154.210 70.665 154.255 ;
        RECT 71.565 154.210 71.855 154.255 ;
        RECT 74.085 154.210 74.375 154.255 ;
        RECT 70.375 154.070 74.375 154.210 ;
        RECT 70.375 154.025 70.665 154.070 ;
        RECT 71.565 154.025 71.855 154.070 ;
        RECT 74.085 154.025 74.375 154.070 ;
        RECT 84.685 154.210 84.975 154.255 ;
        RECT 87.205 154.210 87.495 154.255 ;
        RECT 88.395 154.210 88.685 154.255 ;
        RECT 84.685 154.070 88.685 154.210 ;
        RECT 88.890 154.210 89.030 154.410 ;
        RECT 89.260 154.410 91.330 154.550 ;
        RECT 89.260 154.350 89.580 154.410 ;
        RECT 91.575 154.365 91.865 154.595 ;
        RECT 88.890 154.070 89.950 154.210 ;
        RECT 84.685 154.025 84.975 154.070 ;
        RECT 87.205 154.025 87.495 154.070 ;
        RECT 88.395 154.025 88.685 154.070 ;
        RECT 41.420 153.870 41.740 153.930 ;
        RECT 89.810 153.915 89.950 154.070 ;
        RECT 51.095 153.870 51.385 153.915 ;
        RECT 41.420 153.730 51.385 153.870 ;
        RECT 41.420 153.670 41.740 153.730 ;
        RECT 51.095 153.685 51.385 153.730 ;
        RECT 69.980 153.870 70.270 153.915 ;
        RECT 72.080 153.870 72.370 153.915 ;
        RECT 73.650 153.870 73.940 153.915 ;
        RECT 76.855 153.870 77.145 153.915 ;
        RECT 69.980 153.730 73.940 153.870 ;
        RECT 69.980 153.685 70.270 153.730 ;
        RECT 72.080 153.685 72.370 153.730 ;
        RECT 73.650 153.685 73.940 153.730 ;
        RECT 75.550 153.730 77.145 153.870 ;
        RECT 44.195 153.530 44.485 153.575 ;
        RECT 44.640 153.530 44.960 153.590 ;
        RECT 46.020 153.530 46.340 153.590 ;
        RECT 44.195 153.390 46.340 153.530 ;
        RECT 44.195 153.345 44.485 153.390 ;
        RECT 44.640 153.330 44.960 153.390 ;
        RECT 46.020 153.330 46.340 153.390 ;
        RECT 50.160 153.330 50.480 153.590 ;
        RECT 73.160 153.530 73.480 153.590 ;
        RECT 75.550 153.530 75.690 153.730 ;
        RECT 76.855 153.685 77.145 153.730 ;
        RECT 85.120 153.870 85.410 153.915 ;
        RECT 86.690 153.870 86.980 153.915 ;
        RECT 88.790 153.870 89.080 153.915 ;
        RECT 85.120 153.730 89.080 153.870 ;
        RECT 85.120 153.685 85.410 153.730 ;
        RECT 86.690 153.685 86.980 153.730 ;
        RECT 88.790 153.685 89.080 153.730 ;
        RECT 89.735 153.685 90.025 153.915 ;
        RECT 91.650 153.870 91.790 154.365 ;
        RECT 92.020 154.350 92.340 154.610 ;
        RECT 101.220 154.550 101.540 154.610 ;
        RECT 107.215 154.550 107.505 154.595 ;
        RECT 109.515 154.550 109.805 154.595 ;
        RECT 101.220 154.410 104.210 154.550 ;
        RECT 101.220 154.350 101.540 154.410 ;
        RECT 92.480 154.010 92.800 154.270 ;
        RECT 103.520 154.010 103.840 154.270 ;
        RECT 104.070 154.255 104.210 154.410 ;
        RECT 107.215 154.410 109.805 154.550 ;
        RECT 107.215 154.365 107.505 154.410 ;
        RECT 109.515 154.365 109.805 154.410 ;
        RECT 103.995 154.025 104.285 154.255 ;
        RECT 108.135 154.210 108.425 154.255 ;
        RECT 110.050 154.210 110.190 155.090 ;
        RECT 117.320 155.030 117.640 155.090 ;
        RECT 118.700 155.230 119.020 155.290 ;
        RECT 122.380 155.230 122.700 155.290 ;
        RECT 118.700 155.090 122.700 155.230 ;
        RECT 118.700 155.030 119.020 155.090 ;
        RECT 122.380 155.030 122.700 155.090 ;
        RECT 122.855 155.230 123.145 155.275 ;
        RECT 123.760 155.230 124.080 155.290 ;
        RECT 122.855 155.090 124.080 155.230 ;
        RECT 122.855 155.045 123.145 155.090 ;
        RECT 123.760 155.030 124.080 155.090 ;
        RECT 137.560 155.030 137.880 155.290 ;
        RECT 138.955 155.230 139.245 155.275 ;
        RECT 139.860 155.230 140.180 155.290 ;
        RECT 138.955 155.090 140.180 155.230 ;
        RECT 138.955 155.045 139.245 155.090 ;
        RECT 139.860 155.030 140.180 155.090 ;
        RECT 110.420 154.890 110.740 154.950 ;
        RECT 114.115 154.890 114.405 154.935 ;
        RECT 110.420 154.750 114.405 154.890 ;
        RECT 110.420 154.690 110.740 154.750 ;
        RECT 114.115 154.705 114.405 154.750 ;
        RECT 114.575 154.890 114.865 154.935 ;
        RECT 114.575 154.750 118.930 154.890 ;
        RECT 114.575 154.705 114.865 154.750 ;
        RECT 113.180 154.350 113.500 154.610 ;
        RECT 115.020 154.350 115.340 154.610 ;
        RECT 115.480 154.550 115.800 154.610 ;
        RECT 116.400 154.550 116.720 154.610 ;
        RECT 117.795 154.550 118.085 154.595 ;
        RECT 115.480 154.410 118.085 154.550 ;
        RECT 115.480 154.350 115.800 154.410 ;
        RECT 116.400 154.350 116.720 154.410 ;
        RECT 117.795 154.365 118.085 154.410 ;
        RECT 118.240 154.550 118.560 154.610 ;
        RECT 118.790 154.550 118.930 154.750 ;
        RECT 123.300 154.690 123.620 154.950 ;
        RECT 118.240 154.410 118.930 154.550 ;
        RECT 120.080 154.550 120.400 154.610 ;
        RECT 121.015 154.550 121.305 154.595 ;
        RECT 120.080 154.410 121.305 154.550 ;
        RECT 118.240 154.350 118.560 154.410 ;
        RECT 120.080 154.350 120.400 154.410 ;
        RECT 121.015 154.365 121.305 154.410 ;
        RECT 121.920 154.350 122.240 154.610 ;
        RECT 128.360 154.350 128.680 154.610 ;
        RECT 129.295 154.365 129.585 154.595 ;
        RECT 108.135 154.070 110.190 154.210 ;
        RECT 108.135 154.025 108.425 154.070 ;
        RECT 112.275 154.025 112.565 154.255 ;
        RECT 101.235 153.870 101.525 153.915 ;
        RECT 91.650 153.730 101.525 153.870 ;
        RECT 101.235 153.685 101.525 153.730 ;
        RECT 104.440 153.870 104.760 153.930 ;
        RECT 112.350 153.870 112.490 154.025 ;
        RECT 117.320 154.010 117.640 154.270 ;
        RECT 118.700 154.010 119.020 154.270 ;
        RECT 126.980 154.010 127.300 154.270 ;
        RECT 104.440 153.730 112.490 153.870 ;
        RECT 114.560 153.870 114.880 153.930 ;
        RECT 122.840 153.870 123.160 153.930 ;
        RECT 129.370 153.870 129.510 154.365 ;
        RECT 130.660 154.350 130.980 154.610 ;
        RECT 132.040 154.595 132.360 154.610 ;
        RECT 132.010 154.550 132.360 154.595 ;
        RECT 131.845 154.410 132.360 154.550 ;
        RECT 137.650 154.550 137.790 155.030 ;
        RECT 138.035 154.550 138.325 154.595 ;
        RECT 137.650 154.410 138.325 154.550 ;
        RECT 132.010 154.365 132.360 154.410 ;
        RECT 138.035 154.365 138.325 154.410 ;
        RECT 139.875 154.365 140.165 154.595 ;
        RECT 132.040 154.350 132.360 154.365 ;
        RECT 131.555 154.210 131.845 154.255 ;
        RECT 132.745 154.210 133.035 154.255 ;
        RECT 135.265 154.210 135.555 154.255 ;
        RECT 131.555 154.070 135.555 154.210 ;
        RECT 131.555 154.025 131.845 154.070 ;
        RECT 132.745 154.025 133.035 154.070 ;
        RECT 135.265 154.025 135.555 154.070 ;
        RECT 135.720 154.210 136.040 154.270 ;
        RECT 139.950 154.210 140.090 154.365 ;
        RECT 135.720 154.070 140.090 154.210 ;
        RECT 135.720 154.010 136.040 154.070 ;
        RECT 114.560 153.730 129.510 153.870 ;
        RECT 131.160 153.870 131.450 153.915 ;
        RECT 133.260 153.870 133.550 153.915 ;
        RECT 134.830 153.870 135.120 153.915 ;
        RECT 131.160 153.730 135.120 153.870 ;
        RECT 104.440 153.670 104.760 153.730 ;
        RECT 114.560 153.670 114.880 153.730 ;
        RECT 122.840 153.670 123.160 153.730 ;
        RECT 131.160 153.685 131.450 153.730 ;
        RECT 133.260 153.685 133.550 153.730 ;
        RECT 134.830 153.685 135.120 153.730 ;
        RECT 140.780 153.670 141.100 153.930 ;
        RECT 73.160 153.390 75.690 153.530 ;
        RECT 73.160 153.330 73.480 153.390 ;
        RECT 76.380 153.330 76.700 153.590 ;
        RECT 82.375 153.530 82.665 153.575 ;
        RECT 84.660 153.530 84.980 153.590 ;
        RECT 82.375 153.390 84.980 153.530 ;
        RECT 82.375 153.345 82.665 153.390 ;
        RECT 84.660 153.330 84.980 153.390 ;
        RECT 105.360 153.330 105.680 153.590 ;
        RECT 115.940 153.330 116.260 153.590 ;
        RECT 116.400 153.330 116.720 153.590 ;
        RECT 121.000 153.530 121.320 153.590 ;
        RECT 121.935 153.530 122.225 153.575 ;
        RECT 124.220 153.530 124.540 153.590 ;
        RECT 128.360 153.530 128.680 153.590 ;
        RECT 121.000 153.390 128.680 153.530 ;
        RECT 121.000 153.330 121.320 153.390 ;
        RECT 121.935 153.345 122.225 153.390 ;
        RECT 124.220 153.330 124.540 153.390 ;
        RECT 128.360 153.330 128.680 153.390 ;
        RECT 129.740 153.530 130.060 153.590 ;
        RECT 130.215 153.530 130.505 153.575 ;
        RECT 129.740 153.390 130.505 153.530 ;
        RECT 129.740 153.330 130.060 153.390 ;
        RECT 130.215 153.345 130.505 153.390 ;
        RECT 17.430 152.710 143.010 153.190 ;
        RECT 70.860 152.310 71.180 152.570 ;
        RECT 91.560 152.510 91.880 152.570 ;
        RECT 92.955 152.510 93.245 152.555 ;
        RECT 91.560 152.370 93.245 152.510 ;
        RECT 91.560 152.310 91.880 152.370 ;
        RECT 92.955 152.325 93.245 152.370 ;
        RECT 103.535 152.510 103.825 152.555 ;
        RECT 104.440 152.510 104.760 152.570 ;
        RECT 103.535 152.370 104.760 152.510 ;
        RECT 103.535 152.325 103.825 152.370 ;
        RECT 104.440 152.310 104.760 152.370 ;
        RECT 111.355 152.510 111.645 152.555 ;
        RECT 113.180 152.510 113.500 152.570 ;
        RECT 111.355 152.370 113.500 152.510 ;
        RECT 111.355 152.325 111.645 152.370 ;
        RECT 113.180 152.310 113.500 152.370 ;
        RECT 40.040 152.170 40.360 152.230 ;
        RECT 45.100 152.170 45.420 152.230 ;
        RECT 40.040 152.030 45.420 152.170 ;
        RECT 40.040 151.970 40.360 152.030 ;
        RECT 45.100 151.970 45.420 152.030 ;
        RECT 97.120 152.170 97.410 152.215 ;
        RECT 99.220 152.170 99.510 152.215 ;
        RECT 100.790 152.170 101.080 152.215 ;
        RECT 97.120 152.030 101.080 152.170 ;
        RECT 97.120 151.985 97.410 152.030 ;
        RECT 99.220 151.985 99.510 152.030 ;
        RECT 100.790 151.985 101.080 152.030 ;
        RECT 122.380 152.170 122.700 152.230 ;
        RECT 134.380 152.170 134.670 152.215 ;
        RECT 136.480 152.170 136.770 152.215 ;
        RECT 138.050 152.170 138.340 152.215 ;
        RECT 122.380 152.030 129.970 152.170 ;
        RECT 122.380 151.970 122.700 152.030 ;
        RECT 39.135 151.830 39.425 151.875 ;
        RECT 44.195 151.830 44.485 151.875 ;
        RECT 39.135 151.690 44.485 151.830 ;
        RECT 39.135 151.645 39.425 151.690 ;
        RECT 44.195 151.645 44.485 151.690 ;
        RECT 73.160 151.630 73.480 151.890 ;
        RECT 73.635 151.645 73.925 151.875 ;
        RECT 74.080 151.830 74.400 151.890 ;
        RECT 79.155 151.830 79.445 151.875 ;
        RECT 74.080 151.690 79.445 151.830 ;
        RECT 42.800 151.290 43.120 151.550 ;
        RECT 43.720 151.290 44.040 151.550 ;
        RECT 73.710 151.490 73.850 151.645 ;
        RECT 74.080 151.630 74.400 151.690 ;
        RECT 79.155 151.645 79.445 151.690 ;
        RECT 80.060 151.830 80.380 151.890 ;
        RECT 87.880 151.830 88.200 151.890 ;
        RECT 80.060 151.690 88.200 151.830 ;
        RECT 80.060 151.630 80.380 151.690 ;
        RECT 87.880 151.630 88.200 151.690 ;
        RECT 88.340 151.830 88.660 151.890 ;
        RECT 89.735 151.830 90.025 151.875 ;
        RECT 88.340 151.690 90.025 151.830 ;
        RECT 88.340 151.630 88.660 151.690 ;
        RECT 89.735 151.645 90.025 151.690 ;
        RECT 90.655 151.830 90.945 151.875 ;
        RECT 96.160 151.830 96.480 151.890 ;
        RECT 90.655 151.690 96.480 151.830 ;
        RECT 90.655 151.645 90.945 151.690 ;
        RECT 96.160 151.630 96.480 151.690 ;
        RECT 96.620 151.630 96.940 151.890 ;
        RECT 97.515 151.830 97.805 151.875 ;
        RECT 98.705 151.830 98.995 151.875 ;
        RECT 101.225 151.830 101.515 151.875 ;
        RECT 97.515 151.690 101.515 151.830 ;
        RECT 97.515 151.645 97.805 151.690 ;
        RECT 98.705 151.645 98.995 151.690 ;
        RECT 101.225 151.645 101.515 151.690 ;
        RECT 103.520 151.830 103.840 151.890 ;
        RECT 108.135 151.830 108.425 151.875 ;
        RECT 103.520 151.690 108.425 151.830 ;
        RECT 103.520 151.630 103.840 151.690 ;
        RECT 108.135 151.645 108.425 151.690 ;
        RECT 113.195 151.830 113.485 151.875 ;
        RECT 116.400 151.830 116.720 151.890 ;
        RECT 129.830 151.875 129.970 152.030 ;
        RECT 134.380 152.030 138.340 152.170 ;
        RECT 134.380 151.985 134.670 152.030 ;
        RECT 136.480 151.985 136.770 152.030 ;
        RECT 138.050 151.985 138.340 152.030 ;
        RECT 113.195 151.690 116.720 151.830 ;
        RECT 113.195 151.645 113.485 151.690 ;
        RECT 116.400 151.630 116.720 151.690 ;
        RECT 120.170 151.690 121.690 151.830 ;
        RECT 80.150 151.490 80.290 151.630 ;
        RECT 73.710 151.350 80.290 151.490 ;
        RECT 97.970 151.490 98.260 151.535 ;
        RECT 105.360 151.490 105.680 151.550 ;
        RECT 97.970 151.350 105.680 151.490 ;
        RECT 97.970 151.305 98.260 151.350 ;
        RECT 105.360 151.290 105.680 151.350 ;
        RECT 111.800 151.290 112.120 151.550 ;
        RECT 112.275 151.490 112.565 151.535 ;
        RECT 113.640 151.490 113.960 151.550 ;
        RECT 112.275 151.350 113.960 151.490 ;
        RECT 112.275 151.305 112.565 151.350 ;
        RECT 113.640 151.290 113.960 151.350 ;
        RECT 114.560 151.290 114.880 151.550 ;
        RECT 115.955 151.305 116.245 151.535 ;
        RECT 119.175 151.490 119.465 151.535 ;
        RECT 120.170 151.490 120.310 151.690 ;
        RECT 119.175 151.350 120.310 151.490 ;
        RECT 119.175 151.305 119.465 151.350 ;
        RECT 120.555 151.305 120.845 151.535 ;
        RECT 72.715 151.150 73.005 151.195 ;
        RECT 76.840 151.150 77.160 151.210 ;
        RECT 107.660 151.150 107.980 151.210 ;
        RECT 72.715 151.010 74.080 151.150 ;
        RECT 72.715 150.965 73.005 151.010 ;
        RECT 19.800 150.810 20.120 150.870 ;
        RECT 69.940 150.810 70.260 150.870 ;
        RECT 19.800 150.670 70.260 150.810 ;
        RECT 73.940 150.810 74.080 151.010 ;
        RECT 76.840 151.010 107.980 151.150 ;
        RECT 76.840 150.950 77.160 151.010 ;
        RECT 107.660 150.950 107.980 151.010 ;
        RECT 110.420 151.150 110.740 151.210 ;
        RECT 113.195 151.150 113.485 151.195 ;
        RECT 110.420 151.010 113.485 151.150 ;
        RECT 116.030 151.150 116.170 151.305 ;
        RECT 116.400 151.150 116.720 151.210 ;
        RECT 116.030 151.010 116.720 151.150 ;
        RECT 110.420 150.950 110.740 151.010 ;
        RECT 113.195 150.965 113.485 151.010 ;
        RECT 116.400 150.950 116.720 151.010 ;
        RECT 118.240 151.150 118.560 151.210 ;
        RECT 120.630 151.150 120.770 151.305 ;
        RECT 121.000 151.290 121.320 151.550 ;
        RECT 121.550 151.490 121.690 151.690 ;
        RECT 129.755 151.645 130.045 151.875 ;
        RECT 134.775 151.830 135.065 151.875 ;
        RECT 135.965 151.830 136.255 151.875 ;
        RECT 138.485 151.830 138.775 151.875 ;
        RECT 134.775 151.690 138.775 151.830 ;
        RECT 134.775 151.645 135.065 151.690 ;
        RECT 135.965 151.645 136.255 151.690 ;
        RECT 138.485 151.645 138.775 151.690 ;
        RECT 122.395 151.490 122.685 151.535 ;
        RECT 126.980 151.490 127.300 151.550 ;
        RECT 133.895 151.490 134.185 151.535 ;
        RECT 121.550 151.350 122.685 151.490 ;
        RECT 122.395 151.305 122.685 151.350 ;
        RECT 123.390 151.350 134.185 151.490 ;
        RECT 118.240 151.010 120.770 151.150 ;
        RECT 118.240 150.950 118.560 151.010 ;
        RECT 121.460 150.950 121.780 151.210 ;
        RECT 123.390 151.195 123.530 151.350 ;
        RECT 126.980 151.290 127.300 151.350 ;
        RECT 133.895 151.305 134.185 151.350 ;
        RECT 123.315 150.965 123.605 151.195 ;
        RECT 135.120 151.150 135.410 151.195 ;
        RECT 133.050 151.010 135.410 151.150 ;
        RECT 75.920 150.810 76.240 150.870 ;
        RECT 73.940 150.670 76.240 150.810 ;
        RECT 19.800 150.610 20.120 150.670 ;
        RECT 69.940 150.610 70.260 150.670 ;
        RECT 75.920 150.610 76.240 150.670 ;
        RECT 76.380 150.610 76.700 150.870 ;
        RECT 91.100 150.610 91.420 150.870 ;
        RECT 114.575 150.810 114.865 150.855 ;
        RECT 117.320 150.810 117.640 150.870 ;
        RECT 114.575 150.670 117.640 150.810 ;
        RECT 114.575 150.625 114.865 150.670 ;
        RECT 117.320 150.610 117.640 150.670 ;
        RECT 119.620 150.610 119.940 150.870 ;
        RECT 120.540 150.810 120.860 150.870 ;
        RECT 123.390 150.810 123.530 150.965 ;
        RECT 120.540 150.670 123.530 150.810 ;
        RECT 120.540 150.610 120.860 150.670 ;
        RECT 130.660 150.610 130.980 150.870 ;
        RECT 131.120 150.610 131.440 150.870 ;
        RECT 133.050 150.855 133.190 151.010 ;
        RECT 135.120 150.965 135.410 151.010 ;
        RECT 132.975 150.625 133.265 150.855 ;
        RECT 139.400 150.810 139.720 150.870 ;
        RECT 140.795 150.810 141.085 150.855 ;
        RECT 139.400 150.670 141.085 150.810 ;
        RECT 139.400 150.610 139.720 150.670 ;
        RECT 140.795 150.625 141.085 150.670 ;
        RECT 17.430 149.990 143.010 150.470 ;
        RECT 19.800 149.590 20.120 149.850 ;
        RECT 34.075 149.790 34.365 149.835 ;
        RECT 34.980 149.790 35.300 149.850 ;
        RECT 34.075 149.650 35.300 149.790 ;
        RECT 34.075 149.605 34.365 149.650 ;
        RECT 34.980 149.590 35.300 149.650 ;
        RECT 40.960 149.790 41.280 149.850 ;
        RECT 42.355 149.790 42.645 149.835 ;
        RECT 40.960 149.650 42.645 149.790 ;
        RECT 40.960 149.590 41.280 149.650 ;
        RECT 42.355 149.605 42.645 149.650 ;
        RECT 74.080 149.790 74.400 149.850 ;
        RECT 76.395 149.790 76.685 149.835 ;
        RECT 74.080 149.650 76.685 149.790 ;
        RECT 74.080 149.590 74.400 149.650 ;
        RECT 76.395 149.605 76.685 149.650 ;
        RECT 103.520 149.590 103.840 149.850 ;
        RECT 115.940 149.790 116.260 149.850 ;
        RECT 106.830 149.650 116.260 149.790 ;
        RECT 20.720 149.450 21.040 149.510 ;
        RECT 39.580 149.450 39.900 149.510 ;
        RECT 40.055 149.450 40.345 149.495 ;
        RECT 42.800 149.450 43.120 149.510 ;
        RECT 44.655 149.450 44.945 149.495 ;
        RECT 20.720 149.310 39.350 149.450 ;
        RECT 20.720 149.250 21.040 149.310 ;
        RECT 16.120 149.110 16.440 149.170 ;
        RECT 18.895 149.110 19.185 149.155 ;
        RECT 16.120 148.970 19.185 149.110 ;
        RECT 16.120 148.910 16.440 148.970 ;
        RECT 18.895 148.925 19.185 148.970 ;
        RECT 23.480 148.910 23.800 149.170 ;
        RECT 23.940 149.110 24.260 149.170 ;
        RECT 24.775 149.110 25.065 149.155 ;
        RECT 23.940 148.970 25.065 149.110 ;
        RECT 23.940 148.910 24.260 148.970 ;
        RECT 24.775 148.925 25.065 148.970 ;
        RECT 31.300 149.110 31.620 149.170 ;
        RECT 31.775 149.110 32.065 149.155 ;
        RECT 31.300 148.970 32.065 149.110 ;
        RECT 31.300 148.910 31.620 148.970 ;
        RECT 31.775 148.925 32.065 148.970 ;
        RECT 34.370 149.110 34.660 149.155 ;
        RECT 35.900 149.110 36.220 149.170 ;
        RECT 34.370 148.970 36.220 149.110 ;
        RECT 34.370 148.925 34.660 148.970 ;
        RECT 35.900 148.910 36.220 148.970 ;
        RECT 24.375 148.770 24.665 148.815 ;
        RECT 25.565 148.770 25.855 148.815 ;
        RECT 28.085 148.770 28.375 148.815 ;
        RECT 24.375 148.630 28.375 148.770 ;
        RECT 24.375 148.585 24.665 148.630 ;
        RECT 25.565 148.585 25.855 148.630 ;
        RECT 28.085 148.585 28.375 148.630 ;
        RECT 23.980 148.430 24.270 148.475 ;
        RECT 26.080 148.430 26.370 148.475 ;
        RECT 27.650 148.430 27.940 148.475 ;
        RECT 23.980 148.290 27.940 148.430 ;
        RECT 23.980 148.245 24.270 148.290 ;
        RECT 26.080 148.245 26.370 148.290 ;
        RECT 27.650 148.245 27.940 148.290 ;
        RECT 30.395 148.090 30.685 148.135 ;
        RECT 32.220 148.090 32.540 148.150 ;
        RECT 30.395 147.950 32.540 148.090 ;
        RECT 30.395 147.905 30.685 147.950 ;
        RECT 32.220 147.890 32.540 147.950 ;
        RECT 34.995 148.090 35.285 148.135 ;
        RECT 35.440 148.090 35.760 148.150 ;
        RECT 34.995 147.950 35.760 148.090 ;
        RECT 39.210 148.090 39.350 149.310 ;
        RECT 39.580 149.310 44.945 149.450 ;
        RECT 39.580 149.250 39.900 149.310 ;
        RECT 40.055 149.265 40.345 149.310 ;
        RECT 42.800 149.250 43.120 149.310 ;
        RECT 44.655 149.265 44.945 149.310 ;
        RECT 70.400 149.450 70.720 149.510 ;
        RECT 97.970 149.450 98.260 149.495 ;
        RECT 106.830 149.450 106.970 149.650 ;
        RECT 115.940 149.590 116.260 149.650 ;
        RECT 126.075 149.790 126.365 149.835 ;
        RECT 130.660 149.790 130.980 149.850 ;
        RECT 126.075 149.650 130.980 149.790 ;
        RECT 126.075 149.605 126.365 149.650 ;
        RECT 130.660 149.590 130.980 149.650 ;
        RECT 131.120 149.790 131.440 149.850 ;
        RECT 136.195 149.790 136.485 149.835 ;
        RECT 131.120 149.650 136.485 149.790 ;
        RECT 131.120 149.590 131.440 149.650 ;
        RECT 136.195 149.605 136.485 149.650 ;
        RECT 124.235 149.450 124.525 149.495 ;
        RECT 126.980 149.450 127.300 149.510 ;
        RECT 127.455 149.450 127.745 149.495 ;
        RECT 70.400 149.310 83.970 149.450 ;
        RECT 70.400 149.250 70.720 149.310 ;
        RECT 43.720 149.110 44.040 149.170 ;
        RECT 41.510 148.970 44.040 149.110 ;
        RECT 41.510 148.490 41.650 148.970 ;
        RECT 43.720 148.910 44.040 148.970 ;
        RECT 70.830 149.110 71.120 149.155 ;
        RECT 72.240 149.110 72.560 149.170 ;
        RECT 70.830 148.970 72.560 149.110 ;
        RECT 70.830 148.925 71.120 148.970 ;
        RECT 72.240 148.910 72.560 148.970 ;
        RECT 78.680 148.910 79.000 149.170 ;
        RECT 83.830 149.155 83.970 149.310 ;
        RECT 97.970 149.310 106.970 149.450 ;
        RECT 111.890 149.310 120.310 149.450 ;
        RECT 97.970 149.265 98.260 149.310 ;
        RECT 79.155 149.110 79.445 149.155 ;
        RECT 80.995 149.110 81.285 149.155 ;
        RECT 79.155 148.970 81.285 149.110 ;
        RECT 79.155 148.925 79.445 148.970 ;
        RECT 80.995 148.925 81.285 148.970 ;
        RECT 83.755 148.925 84.045 149.155 ;
        RECT 96.620 148.910 96.940 149.170 ;
        RECT 110.420 149.155 110.740 149.170 ;
        RECT 111.890 149.155 112.030 149.310 ;
        RECT 110.420 149.110 110.770 149.155 ;
        RECT 110.420 148.970 110.935 149.110 ;
        RECT 110.420 148.925 110.770 148.970 ;
        RECT 111.815 148.925 112.105 149.155 ;
        RECT 116.400 149.110 116.720 149.170 ;
        RECT 113.270 148.970 116.720 149.110 ;
        RECT 110.420 148.910 110.740 148.925 ;
        RECT 66.720 148.770 67.040 148.830 ;
        RECT 69.495 148.770 69.785 148.815 ;
        RECT 66.720 148.630 69.785 148.770 ;
        RECT 66.720 148.570 67.040 148.630 ;
        RECT 69.495 148.585 69.785 148.630 ;
        RECT 70.375 148.770 70.665 148.815 ;
        RECT 71.565 148.770 71.855 148.815 ;
        RECT 74.085 148.770 74.375 148.815 ;
        RECT 70.375 148.630 74.375 148.770 ;
        RECT 70.375 148.585 70.665 148.630 ;
        RECT 71.565 148.585 71.855 148.630 ;
        RECT 74.085 148.585 74.375 148.630 ;
        RECT 80.060 148.570 80.380 148.830 ;
        RECT 97.515 148.770 97.805 148.815 ;
        RECT 98.705 148.770 98.995 148.815 ;
        RECT 101.225 148.770 101.515 148.815 ;
        RECT 97.515 148.630 101.515 148.770 ;
        RECT 97.515 148.585 97.805 148.630 ;
        RECT 98.705 148.585 98.995 148.630 ;
        RECT 101.225 148.585 101.515 148.630 ;
        RECT 107.225 148.770 107.515 148.815 ;
        RECT 109.745 148.770 110.035 148.815 ;
        RECT 110.935 148.770 111.225 148.815 ;
        RECT 107.225 148.630 111.225 148.770 ;
        RECT 107.225 148.585 107.515 148.630 ;
        RECT 109.745 148.585 110.035 148.630 ;
        RECT 110.935 148.585 111.225 148.630 ;
        RECT 41.420 148.230 41.740 148.490 ;
        RECT 69.980 148.430 70.270 148.475 ;
        RECT 72.080 148.430 72.370 148.475 ;
        RECT 73.650 148.430 73.940 148.475 ;
        RECT 76.855 148.430 77.145 148.475 ;
        RECT 44.270 148.290 69.710 148.430 ;
        RECT 44.270 148.090 44.410 148.290 ;
        RECT 39.210 147.950 44.410 148.090 ;
        RECT 44.640 148.090 44.960 148.150 ;
        RECT 45.575 148.090 45.865 148.135 ;
        RECT 44.640 147.950 45.865 148.090 ;
        RECT 69.570 148.090 69.710 148.290 ;
        RECT 69.980 148.290 73.940 148.430 ;
        RECT 69.980 148.245 70.270 148.290 ;
        RECT 72.080 148.245 72.370 148.290 ;
        RECT 73.650 148.245 73.940 148.290 ;
        RECT 75.550 148.290 77.145 148.430 ;
        RECT 70.860 148.090 71.180 148.150 ;
        RECT 69.570 147.950 71.180 148.090 ;
        RECT 34.995 147.905 35.285 147.950 ;
        RECT 35.440 147.890 35.760 147.950 ;
        RECT 44.640 147.890 44.960 147.950 ;
        RECT 45.575 147.905 45.865 147.950 ;
        RECT 70.860 147.890 71.180 147.950 ;
        RECT 73.160 148.090 73.480 148.150 ;
        RECT 75.550 148.090 75.690 148.290 ;
        RECT 76.855 148.245 77.145 148.290 ;
        RECT 97.120 148.430 97.410 148.475 ;
        RECT 99.220 148.430 99.510 148.475 ;
        RECT 100.790 148.430 101.080 148.475 ;
        RECT 97.120 148.290 101.080 148.430 ;
        RECT 97.120 148.245 97.410 148.290 ;
        RECT 99.220 148.245 99.510 148.290 ;
        RECT 100.790 148.245 101.080 148.290 ;
        RECT 107.660 148.430 107.950 148.475 ;
        RECT 109.230 148.430 109.520 148.475 ;
        RECT 111.330 148.430 111.620 148.475 ;
        RECT 107.660 148.290 111.620 148.430 ;
        RECT 107.660 148.245 107.950 148.290 ;
        RECT 109.230 148.245 109.520 148.290 ;
        RECT 111.330 148.245 111.620 148.290 ;
        RECT 113.270 148.150 113.410 148.970 ;
        RECT 116.400 148.910 116.720 148.970 ;
        RECT 118.815 149.110 119.105 149.155 ;
        RECT 119.620 149.110 119.940 149.170 ;
        RECT 118.815 148.970 119.940 149.110 ;
        RECT 118.815 148.925 119.105 148.970 ;
        RECT 119.620 148.910 119.940 148.970 ;
        RECT 120.170 148.815 120.310 149.310 ;
        RECT 124.235 149.310 130.890 149.450 ;
        RECT 124.235 149.265 124.525 149.310 ;
        RECT 126.980 149.250 127.300 149.310 ;
        RECT 127.455 149.265 127.745 149.310 ;
        RECT 121.015 148.925 121.305 149.155 ;
        RECT 115.505 148.770 115.795 148.815 ;
        RECT 118.025 148.770 118.315 148.815 ;
        RECT 119.215 148.770 119.505 148.815 ;
        RECT 115.505 148.630 119.505 148.770 ;
        RECT 115.505 148.585 115.795 148.630 ;
        RECT 118.025 148.585 118.315 148.630 ;
        RECT 119.215 148.585 119.505 148.630 ;
        RECT 120.095 148.770 120.385 148.815 ;
        RECT 120.540 148.770 120.860 148.830 ;
        RECT 120.095 148.630 120.860 148.770 ;
        RECT 120.095 148.585 120.385 148.630 ;
        RECT 120.540 148.570 120.860 148.630 ;
        RECT 115.940 148.430 116.230 148.475 ;
        RECT 117.510 148.430 117.800 148.475 ;
        RECT 119.610 148.430 119.900 148.475 ;
        RECT 115.940 148.290 119.900 148.430 ;
        RECT 115.940 148.245 116.230 148.290 ;
        RECT 117.510 148.245 117.800 148.290 ;
        RECT 119.610 148.245 119.900 148.290 ;
        RECT 73.160 147.950 75.690 148.090 ;
        RECT 88.340 148.090 88.660 148.150 ;
        RECT 101.220 148.090 101.540 148.150 ;
        RECT 88.340 147.950 101.540 148.090 ;
        RECT 73.160 147.890 73.480 147.950 ;
        RECT 88.340 147.890 88.660 147.950 ;
        RECT 101.220 147.890 101.540 147.950 ;
        RECT 104.915 148.090 105.205 148.135 ;
        RECT 105.360 148.090 105.680 148.150 ;
        RECT 104.915 147.950 105.680 148.090 ;
        RECT 104.915 147.905 105.205 147.950 ;
        RECT 105.360 147.890 105.680 147.950 ;
        RECT 113.180 147.890 113.500 148.150 ;
        RECT 113.640 148.090 113.960 148.150 ;
        RECT 121.090 148.090 121.230 148.925 ;
        RECT 121.920 148.910 122.240 149.170 ;
        RECT 122.380 149.110 122.700 149.170 ;
        RECT 123.315 149.110 123.605 149.155 ;
        RECT 122.380 148.970 123.605 149.110 ;
        RECT 122.380 148.910 122.700 148.970 ;
        RECT 123.315 148.925 123.605 148.970 ;
        RECT 124.680 148.910 125.000 149.170 ;
        RECT 125.140 148.910 125.460 149.170 ;
        RECT 126.535 148.925 126.825 149.155 ;
        RECT 121.475 148.770 121.765 148.815 ;
        RECT 126.610 148.770 126.750 148.925 ;
        RECT 127.900 148.910 128.220 149.170 ;
        RECT 128.375 148.925 128.665 149.155 ;
        RECT 128.450 148.770 128.590 148.925 ;
        RECT 129.740 148.910 130.060 149.170 ;
        RECT 130.750 149.155 130.890 149.310 ;
        RECT 130.675 148.925 130.965 149.155 ;
        RECT 131.120 148.910 131.440 149.170 ;
        RECT 131.595 148.925 131.885 149.155 ;
        RECT 134.815 149.110 135.105 149.155 ;
        RECT 139.400 149.110 139.720 149.170 ;
        RECT 134.815 148.970 139.720 149.110 ;
        RECT 134.815 148.925 135.105 148.970 ;
        RECT 131.670 148.770 131.810 148.925 ;
        RECT 139.400 148.910 139.720 148.970 ;
        RECT 139.875 149.110 140.165 149.155 ;
        RECT 140.320 149.110 140.640 149.170 ;
        RECT 139.875 148.970 140.640 149.110 ;
        RECT 139.875 148.925 140.165 148.970 ;
        RECT 140.320 148.910 140.640 148.970 ;
        RECT 121.475 148.630 126.750 148.770 ;
        RECT 127.990 148.630 131.810 148.770 ;
        RECT 121.475 148.585 121.765 148.630 ;
        RECT 125.140 148.430 125.460 148.490 ;
        RECT 127.440 148.430 127.760 148.490 ;
        RECT 127.990 148.430 128.130 148.630 ;
        RECT 125.140 148.290 128.130 148.430 ;
        RECT 132.515 148.430 132.805 148.475 ;
        RECT 134.340 148.430 134.660 148.490 ;
        RECT 132.515 148.290 134.660 148.430 ;
        RECT 125.140 148.230 125.460 148.290 ;
        RECT 127.440 148.230 127.760 148.290 ;
        RECT 132.515 148.245 132.805 148.290 ;
        RECT 134.340 148.230 134.660 148.290 ;
        RECT 135.720 148.230 136.040 148.490 ;
        RECT 113.640 147.950 121.230 148.090 ;
        RECT 129.295 148.090 129.585 148.135 ;
        RECT 134.800 148.090 135.120 148.150 ;
        RECT 129.295 147.950 135.120 148.090 ;
        RECT 113.640 147.890 113.960 147.950 ;
        RECT 129.295 147.905 129.585 147.950 ;
        RECT 134.800 147.890 135.120 147.950 ;
        RECT 140.780 147.890 141.100 148.150 ;
        RECT 17.430 147.270 143.010 147.750 ;
        RECT 19.815 147.070 20.105 147.115 ;
        RECT 20.720 147.070 21.040 147.130 ;
        RECT 19.815 146.930 21.040 147.070 ;
        RECT 19.815 146.885 20.105 146.930 ;
        RECT 20.720 146.870 21.040 146.930 ;
        RECT 23.940 146.870 24.260 147.130 ;
        RECT 24.860 146.870 25.180 147.130 ;
        RECT 45.560 147.070 45.880 147.130 ;
        RECT 46.495 147.070 46.785 147.115 ;
        RECT 45.560 146.930 46.785 147.070 ;
        RECT 45.560 146.870 45.880 146.930 ;
        RECT 46.495 146.885 46.785 146.930 ;
        RECT 66.735 147.070 67.025 147.115 ;
        RECT 70.400 147.070 70.720 147.130 ;
        RECT 66.735 146.930 70.720 147.070 ;
        RECT 66.735 146.885 67.025 146.930 ;
        RECT 70.400 146.870 70.720 146.930 ;
        RECT 72.240 147.070 72.560 147.130 ;
        RECT 74.095 147.070 74.385 147.115 ;
        RECT 72.240 146.930 74.385 147.070 ;
        RECT 72.240 146.870 72.560 146.930 ;
        RECT 74.095 146.885 74.385 146.930 ;
        RECT 78.680 147.070 79.000 147.130 ;
        RECT 103.075 147.070 103.365 147.115 ;
        RECT 78.680 146.930 103.365 147.070 ;
        RECT 78.680 146.870 79.000 146.930 ;
        RECT 103.075 146.885 103.365 146.930 ;
        RECT 112.735 147.070 113.025 147.115 ;
        RECT 118.700 147.070 119.020 147.130 ;
        RECT 112.735 146.930 119.020 147.070 ;
        RECT 112.735 146.885 113.025 146.930 ;
        RECT 118.700 146.870 119.020 146.930 ;
        RECT 123.315 147.070 123.605 147.115 ;
        RECT 130.660 147.070 130.980 147.130 ;
        RECT 123.315 146.930 130.980 147.070 ;
        RECT 123.315 146.885 123.605 146.930 ;
        RECT 130.660 146.870 130.980 146.930 ;
        RECT 140.795 147.070 141.085 147.115 ;
        RECT 142.160 147.070 142.480 147.130 ;
        RECT 140.795 146.930 142.480 147.070 ;
        RECT 140.795 146.885 141.085 146.930 ;
        RECT 142.160 146.870 142.480 146.930 ;
        RECT 69.480 146.730 69.770 146.775 ;
        RECT 71.050 146.730 71.340 146.775 ;
        RECT 73.150 146.730 73.440 146.775 ;
        RECT 69.480 146.590 73.440 146.730 ;
        RECT 69.480 146.545 69.770 146.590 ;
        RECT 71.050 146.545 71.340 146.590 ;
        RECT 73.150 146.545 73.440 146.590 ;
        RECT 75.920 146.730 76.240 146.790 ;
        RECT 98.935 146.730 99.225 146.775 ;
        RECT 104.440 146.730 104.760 146.790 ;
        RECT 75.920 146.590 99.225 146.730 ;
        RECT 75.920 146.530 76.240 146.590 ;
        RECT 98.935 146.545 99.225 146.590 ;
        RECT 101.310 146.590 104.760 146.730 ;
        RECT 28.080 146.390 28.400 146.450 ;
        RECT 25.640 146.250 28.400 146.390 ;
        RECT 22.575 145.865 22.865 146.095 ;
        RECT 23.495 146.050 23.785 146.095 ;
        RECT 25.640 146.050 25.780 146.250 ;
        RECT 28.080 146.190 28.400 146.250 ;
        RECT 28.540 146.390 28.860 146.450 ;
        RECT 41.420 146.390 41.740 146.450 ;
        RECT 69.045 146.390 69.335 146.435 ;
        RECT 71.565 146.390 71.855 146.435 ;
        RECT 72.755 146.390 73.045 146.435 ;
        RECT 28.540 146.250 33.830 146.390 ;
        RECT 28.540 146.190 28.860 146.250 ;
        RECT 23.495 145.910 25.780 146.050 ;
        RECT 23.495 145.865 23.785 145.910 ;
        RECT 19.340 145.510 19.660 145.770 ;
        RECT 22.650 145.370 22.790 145.865 ;
        RECT 26.240 145.850 26.560 146.110 ;
        RECT 27.175 146.050 27.465 146.095 ;
        RECT 29.920 146.050 30.240 146.110 ;
        RECT 27.175 145.910 30.240 146.050 ;
        RECT 27.175 145.865 27.465 145.910 ;
        RECT 29.920 145.850 30.240 145.910 ;
        RECT 32.220 145.850 32.540 146.110 ;
        RECT 23.035 145.710 23.325 145.755 ;
        RECT 24.715 145.710 25.005 145.755 ;
        RECT 23.035 145.570 25.005 145.710 ;
        RECT 23.035 145.525 23.325 145.570 ;
        RECT 24.715 145.525 25.005 145.570 ;
        RECT 25.320 145.710 25.640 145.770 ;
        RECT 25.795 145.710 26.085 145.755 ;
        RECT 25.320 145.570 26.085 145.710 ;
        RECT 25.320 145.510 25.640 145.570 ;
        RECT 25.795 145.525 26.085 145.570 ;
        RECT 28.540 145.510 28.860 145.770 ;
        RECT 29.475 145.710 29.765 145.755 ;
        RECT 31.760 145.710 32.080 145.770 ;
        RECT 33.690 145.755 33.830 146.250 ;
        RECT 40.125 146.250 41.740 146.390 ;
        RECT 40.125 146.095 40.265 146.250 ;
        RECT 41.420 146.190 41.740 146.250 ;
        RECT 59.450 146.250 63.270 146.390 ;
        RECT 40.050 145.865 40.340 146.095 ;
        RECT 40.500 145.850 40.820 146.110 ;
        RECT 44.640 145.850 44.960 146.110 ;
        RECT 45.575 146.050 45.865 146.095 ;
        RECT 48.780 146.050 49.100 146.110 ;
        RECT 45.575 145.910 49.100 146.050 ;
        RECT 45.575 145.865 45.865 145.910 ;
        RECT 29.475 145.570 32.080 145.710 ;
        RECT 29.475 145.525 29.765 145.570 ;
        RECT 31.760 145.510 32.080 145.570 ;
        RECT 33.615 145.710 33.905 145.755 ;
        RECT 40.590 145.710 40.730 145.850 ;
        RECT 33.615 145.570 40.730 145.710 ;
        RECT 33.615 145.525 33.905 145.570 ;
        RECT 45.650 145.430 45.790 145.865 ;
        RECT 48.780 145.850 49.100 145.910 ;
        RECT 54.760 146.050 55.080 146.110 ;
        RECT 59.450 146.095 59.590 146.250 ;
        RECT 63.130 146.095 63.270 146.250 ;
        RECT 69.045 146.250 73.045 146.390 ;
        RECT 69.045 146.205 69.335 146.250 ;
        RECT 71.565 146.205 71.855 146.250 ;
        RECT 72.755 146.205 73.045 146.250 ;
        RECT 76.380 146.190 76.700 146.450 ;
        RECT 77.315 146.390 77.605 146.435 ;
        RECT 80.060 146.390 80.380 146.450 ;
        RECT 86.975 146.390 87.265 146.435 ;
        RECT 88.340 146.390 88.660 146.450 ;
        RECT 77.315 146.250 80.380 146.390 ;
        RECT 77.315 146.205 77.605 146.250 ;
        RECT 80.060 146.190 80.380 146.250 ;
        RECT 86.130 146.250 88.660 146.390 ;
        RECT 59.375 146.050 59.665 146.095 ;
        RECT 62.135 146.050 62.425 146.095 ;
        RECT 54.760 145.910 59.665 146.050 ;
        RECT 54.760 145.850 55.080 145.910 ;
        RECT 59.375 145.865 59.665 145.910 ;
        RECT 61.290 145.910 62.425 146.050 ;
        RECT 57.060 145.710 57.380 145.770 ;
        RECT 58.455 145.710 58.745 145.755 ;
        RECT 57.060 145.570 58.745 145.710 ;
        RECT 57.060 145.510 57.380 145.570 ;
        RECT 58.455 145.525 58.745 145.570 ;
        RECT 59.820 145.710 60.140 145.770 ;
        RECT 61.290 145.755 61.430 145.910 ;
        RECT 62.135 145.865 62.425 145.910 ;
        RECT 63.055 145.865 63.345 146.095 ;
        RECT 72.355 146.050 72.645 146.095 ;
        RECT 73.160 146.050 73.480 146.110 ;
        RECT 72.355 145.910 73.480 146.050 ;
        RECT 72.355 145.865 72.645 145.910 ;
        RECT 73.160 145.850 73.480 145.910 ;
        RECT 73.620 145.850 73.940 146.110 ;
        RECT 77.760 146.050 78.080 146.110 ;
        RECT 86.130 146.050 86.270 146.250 ;
        RECT 86.975 146.205 87.265 146.250 ;
        RECT 88.340 146.190 88.660 146.250 ;
        RECT 88.800 146.190 89.120 146.450 ;
        RECT 101.310 146.435 101.450 146.590 ;
        RECT 104.440 146.530 104.760 146.590 ;
        RECT 113.640 146.730 113.960 146.790 ;
        RECT 115.035 146.730 115.325 146.775 ;
        RECT 124.235 146.730 124.525 146.775 ;
        RECT 125.140 146.730 125.460 146.790 ;
        RECT 113.640 146.590 115.325 146.730 ;
        RECT 113.640 146.530 113.960 146.590 ;
        RECT 115.035 146.545 115.325 146.590 ;
        RECT 120.170 146.590 125.460 146.730 ;
        RECT 101.235 146.205 101.525 146.435 ;
        RECT 101.680 146.390 102.000 146.450 ;
        RECT 120.170 146.435 120.310 146.590 ;
        RECT 124.235 146.545 124.525 146.590 ;
        RECT 125.140 146.530 125.460 146.590 ;
        RECT 126.560 146.730 126.850 146.775 ;
        RECT 128.660 146.730 128.950 146.775 ;
        RECT 130.230 146.730 130.520 146.775 ;
        RECT 126.560 146.590 130.520 146.730 ;
        RECT 126.560 146.545 126.850 146.590 ;
        RECT 128.660 146.545 128.950 146.590 ;
        RECT 130.230 146.545 130.520 146.590 ;
        RECT 132.975 146.730 133.265 146.775 ;
        RECT 132.975 146.590 136.870 146.730 ;
        RECT 132.975 146.545 133.265 146.590 ;
        RECT 136.730 146.450 136.870 146.590 ;
        RECT 105.835 146.390 106.125 146.435 ;
        RECT 101.680 146.250 106.125 146.390 ;
        RECT 101.680 146.190 102.000 146.250 ;
        RECT 105.835 146.205 106.125 146.250 ;
        RECT 120.095 146.205 120.385 146.435 ;
        RECT 120.540 146.390 120.860 146.450 ;
        RECT 125.600 146.390 125.920 146.450 ;
        RECT 126.075 146.390 126.365 146.435 ;
        RECT 120.540 146.250 126.365 146.390 ;
        RECT 120.540 146.190 120.860 146.250 ;
        RECT 125.600 146.190 125.920 146.250 ;
        RECT 126.075 146.205 126.365 146.250 ;
        RECT 126.955 146.390 127.245 146.435 ;
        RECT 128.145 146.390 128.435 146.435 ;
        RECT 130.665 146.390 130.955 146.435 ;
        RECT 126.955 146.250 130.955 146.390 ;
        RECT 126.955 146.205 127.245 146.250 ;
        RECT 128.145 146.205 128.435 146.250 ;
        RECT 130.665 146.205 130.955 146.250 ;
        RECT 136.640 146.190 136.960 146.450 ;
        RECT 77.760 145.910 86.270 146.050 ;
        RECT 86.515 146.050 86.805 146.095 ;
        RECT 105.360 146.050 105.680 146.110 ;
        RECT 108.595 146.050 108.885 146.095 ;
        RECT 86.515 145.910 105.130 146.050 ;
        RECT 77.760 145.850 78.080 145.910 ;
        RECT 86.515 145.865 86.805 145.910 ;
        RECT 61.215 145.710 61.505 145.755 ;
        RECT 59.820 145.570 61.505 145.710 ;
        RECT 59.820 145.510 60.140 145.570 ;
        RECT 61.215 145.525 61.505 145.570 ;
        RECT 75.935 145.710 76.225 145.755 ;
        RECT 75.935 145.570 79.830 145.710 ;
        RECT 75.935 145.525 76.225 145.570 ;
        RECT 26.700 145.370 27.020 145.430 ;
        RECT 22.650 145.230 27.020 145.370 ;
        RECT 26.700 145.170 27.020 145.230 ;
        RECT 27.620 145.170 27.940 145.430 ;
        RECT 30.840 145.170 31.160 145.430 ;
        RECT 32.695 145.370 32.985 145.415 ;
        RECT 35.900 145.370 36.220 145.430 ;
        RECT 32.695 145.230 36.220 145.370 ;
        RECT 32.695 145.185 32.985 145.230 ;
        RECT 35.900 145.170 36.220 145.230 ;
        RECT 38.660 145.170 38.980 145.430 ;
        RECT 44.195 145.370 44.485 145.415 ;
        RECT 45.560 145.370 45.880 145.430 ;
        RECT 44.195 145.230 45.880 145.370 ;
        RECT 44.195 145.185 44.485 145.230 ;
        RECT 45.560 145.170 45.880 145.230 ;
        RECT 56.600 145.370 56.920 145.430 ;
        RECT 60.755 145.370 61.045 145.415 ;
        RECT 56.600 145.230 61.045 145.370 ;
        RECT 56.600 145.170 56.920 145.230 ;
        RECT 60.755 145.185 61.045 145.230 ;
        RECT 63.040 145.170 63.360 145.430 ;
        RECT 78.680 145.170 79.000 145.430 ;
        RECT 79.690 145.370 79.830 145.570 ;
        RECT 80.060 145.510 80.380 145.770 ;
        RECT 100.775 145.710 101.065 145.755 ;
        RECT 104.440 145.710 104.760 145.770 ;
        RECT 100.775 145.570 104.760 145.710 ;
        RECT 104.990 145.710 105.130 145.910 ;
        RECT 105.360 145.910 108.885 146.050 ;
        RECT 105.360 145.850 105.680 145.910 ;
        RECT 108.595 145.865 108.885 145.910 ;
        RECT 111.815 146.050 112.105 146.095 ;
        RECT 112.275 146.050 112.565 146.095 ;
        RECT 111.815 145.910 112.565 146.050 ;
        RECT 111.815 145.865 112.105 145.910 ;
        RECT 112.275 145.865 112.565 145.910 ;
        RECT 112.720 146.050 113.040 146.110 ;
        RECT 114.575 146.050 114.865 146.095 ;
        RECT 112.720 145.910 114.865 146.050 ;
        RECT 112.720 145.850 113.040 145.910 ;
        RECT 114.575 145.865 114.865 145.910 ;
        RECT 115.480 145.850 115.800 146.110 ;
        RECT 121.460 145.850 121.780 146.110 ;
        RECT 125.140 146.050 125.460 146.110 ;
        RECT 130.200 146.050 130.520 146.110 ;
        RECT 125.140 145.910 130.520 146.050 ;
        RECT 125.140 145.850 125.460 145.910 ;
        RECT 130.200 145.850 130.520 145.910 ;
        RECT 138.020 145.850 138.340 146.110 ;
        RECT 139.875 145.865 140.165 146.095 ;
        RECT 113.180 145.710 113.500 145.770 ;
        RECT 104.990 145.570 113.500 145.710 ;
        RECT 100.775 145.525 101.065 145.570 ;
        RECT 104.440 145.510 104.760 145.570 ;
        RECT 113.180 145.510 113.500 145.570 ;
        RECT 127.410 145.710 127.700 145.755 ;
        RECT 128.360 145.710 128.680 145.770 ;
        RECT 127.410 145.570 128.680 145.710 ;
        RECT 127.410 145.525 127.700 145.570 ;
        RECT 128.360 145.510 128.680 145.570 ;
        RECT 128.820 145.710 129.140 145.770 ;
        RECT 139.950 145.710 140.090 145.865 ;
        RECT 128.820 145.570 140.090 145.710 ;
        RECT 128.820 145.510 129.140 145.570 ;
        RECT 84.215 145.370 84.505 145.415 ;
        RECT 79.690 145.230 84.505 145.370 ;
        RECT 84.215 145.185 84.505 145.230 ;
        RECT 86.040 145.170 86.360 145.430 ;
        RECT 91.560 145.170 91.880 145.430 ;
        RECT 104.900 145.170 105.220 145.430 ;
        RECT 116.860 145.370 117.180 145.430 ;
        RECT 121.015 145.370 121.305 145.415 ;
        RECT 116.860 145.230 121.305 145.370 ;
        RECT 116.860 145.170 117.180 145.230 ;
        RECT 121.015 145.185 121.305 145.230 ;
        RECT 133.420 145.370 133.740 145.430 ;
        RECT 133.895 145.370 134.185 145.415 ;
        RECT 133.420 145.230 134.185 145.370 ;
        RECT 133.420 145.170 133.740 145.230 ;
        RECT 133.895 145.185 134.185 145.230 ;
        RECT 138.940 145.170 139.260 145.430 ;
        RECT 17.430 144.550 143.010 145.030 ;
        RECT 25.795 144.350 26.085 144.395 ;
        RECT 27.620 144.350 27.940 144.410 ;
        RECT 25.795 144.210 27.940 144.350 ;
        RECT 25.795 144.165 26.085 144.210 ;
        RECT 27.620 144.150 27.940 144.210 ;
        RECT 31.760 144.350 32.080 144.410 ;
        RECT 34.075 144.350 34.365 144.395 ;
        RECT 39.580 144.350 39.900 144.410 ;
        RECT 31.760 144.210 34.365 144.350 ;
        RECT 31.760 144.150 32.080 144.210 ;
        RECT 34.075 144.165 34.365 144.210 ;
        RECT 36.910 144.210 39.900 144.350 ;
        RECT 21.655 143.825 21.945 144.055 ;
        RECT 26.715 144.010 27.005 144.055 ;
        RECT 28.400 144.010 28.690 144.055 ;
        RECT 26.715 143.870 28.690 144.010 ;
        RECT 34.150 144.010 34.290 144.165 ;
        RECT 34.150 143.870 35.210 144.010 ;
        RECT 26.715 143.825 27.005 143.870 ;
        RECT 28.400 143.825 28.690 143.870 ;
        RECT 21.730 143.670 21.870 143.825 ;
        RECT 24.860 143.670 25.180 143.730 ;
        RECT 21.730 143.530 25.180 143.670 ;
        RECT 24.860 143.470 25.180 143.530 ;
        RECT 25.335 143.670 25.625 143.715 ;
        RECT 26.240 143.670 26.560 143.730 ;
        RECT 27.620 143.670 27.940 143.730 ;
        RECT 25.335 143.530 27.940 143.670 ;
        RECT 25.335 143.485 25.625 143.530 ;
        RECT 26.240 143.470 26.560 143.530 ;
        RECT 27.620 143.470 27.940 143.530 ;
        RECT 32.680 143.670 33.000 143.730 ;
        RECT 34.535 143.670 34.825 143.715 ;
        RECT 32.680 143.530 34.825 143.670 ;
        RECT 32.680 143.470 33.000 143.530 ;
        RECT 34.535 143.485 34.825 143.530 ;
        RECT 21.730 143.190 24.170 143.330 ;
        RECT 20.735 142.650 21.025 142.695 ;
        RECT 21.180 142.650 21.500 142.710 ;
        RECT 21.730 142.695 21.870 143.190 ;
        RECT 24.030 143.035 24.170 143.190 ;
        RECT 27.160 143.130 27.480 143.390 ;
        RECT 28.055 143.330 28.345 143.375 ;
        RECT 29.245 143.330 29.535 143.375 ;
        RECT 31.765 143.330 32.055 143.375 ;
        RECT 28.055 143.190 32.055 143.330 ;
        RECT 35.070 143.330 35.210 143.870 ;
        RECT 36.910 143.715 37.050 144.210 ;
        RECT 39.580 144.150 39.900 144.210 ;
        RECT 73.175 144.350 73.465 144.395 ;
        RECT 78.220 144.350 78.540 144.410 ;
        RECT 73.175 144.210 78.540 144.350 ;
        RECT 73.175 144.165 73.465 144.210 ;
        RECT 78.220 144.150 78.540 144.210 ;
        RECT 78.680 144.350 79.000 144.410 ;
        RECT 89.735 144.350 90.025 144.395 ;
        RECT 91.560 144.350 91.880 144.410 ;
        RECT 78.680 144.210 89.490 144.350 ;
        RECT 78.680 144.150 79.000 144.210 ;
        RECT 37.295 144.010 37.585 144.055 ;
        RECT 38.660 144.010 38.980 144.070 ;
        RECT 39.135 144.010 39.425 144.055 ;
        RECT 37.295 143.870 38.430 144.010 ;
        RECT 37.295 143.825 37.585 143.870 ;
        RECT 38.290 143.715 38.430 143.870 ;
        RECT 38.660 143.870 39.425 144.010 ;
        RECT 38.660 143.810 38.980 143.870 ;
        RECT 39.135 143.825 39.425 143.870 ;
        RECT 40.960 144.010 41.280 144.070 ;
        RECT 43.735 144.010 44.025 144.055 ;
        RECT 66.720 144.010 67.040 144.070 ;
        RECT 73.620 144.010 73.940 144.070 ;
        RECT 40.960 143.870 44.025 144.010 ;
        RECT 40.960 143.810 41.280 143.870 ;
        RECT 43.735 143.825 44.025 143.870 ;
        RECT 61.750 143.870 80.290 144.010 ;
        RECT 36.835 143.485 37.125 143.715 ;
        RECT 37.755 143.485 38.045 143.715 ;
        RECT 38.215 143.485 38.505 143.715 ;
        RECT 39.595 143.485 39.885 143.715 ;
        RECT 40.055 143.670 40.345 143.715 ;
        RECT 41.880 143.670 42.200 143.730 ;
        RECT 45.100 143.670 45.420 143.730 ;
        RECT 40.055 143.530 45.420 143.670 ;
        RECT 40.055 143.485 40.345 143.530 ;
        RECT 37.830 143.330 37.970 143.485 ;
        RECT 39.670 143.330 39.810 143.485 ;
        RECT 41.880 143.470 42.200 143.530 ;
        RECT 45.100 143.470 45.420 143.530 ;
        RECT 45.575 143.670 45.865 143.715 ;
        RECT 50.160 143.670 50.480 143.730 ;
        RECT 57.520 143.670 57.840 143.730 ;
        RECT 45.575 143.530 57.840 143.670 ;
        RECT 45.575 143.485 45.865 143.530 ;
        RECT 50.160 143.470 50.480 143.530 ;
        RECT 35.070 143.190 39.810 143.330 ;
        RECT 40.500 143.330 40.820 143.390 ;
        RECT 44.655 143.330 44.945 143.375 ;
        RECT 40.500 143.190 44.945 143.330 ;
        RECT 28.055 143.145 28.345 143.190 ;
        RECT 29.245 143.145 29.535 143.190 ;
        RECT 31.765 143.145 32.055 143.190 ;
        RECT 40.500 143.130 40.820 143.190 ;
        RECT 44.655 143.145 44.945 143.190 ;
        RECT 23.495 142.805 23.785 143.035 ;
        RECT 23.955 142.990 24.245 143.035 ;
        RECT 25.320 142.990 25.640 143.050 ;
        RECT 23.955 142.850 25.640 142.990 ;
        RECT 23.955 142.805 24.245 142.850 ;
        RECT 20.735 142.510 21.500 142.650 ;
        RECT 20.735 142.465 21.025 142.510 ;
        RECT 21.180 142.450 21.500 142.510 ;
        RECT 21.655 142.465 21.945 142.695 ;
        RECT 23.570 142.650 23.710 142.805 ;
        RECT 25.320 142.790 25.640 142.850 ;
        RECT 27.660 142.990 27.950 143.035 ;
        RECT 29.760 142.990 30.050 143.035 ;
        RECT 31.330 142.990 31.620 143.035 ;
        RECT 27.660 142.850 31.620 142.990 ;
        RECT 27.660 142.805 27.950 142.850 ;
        RECT 29.760 142.805 30.050 142.850 ;
        RECT 31.330 142.805 31.620 142.850 ;
        RECT 45.100 142.790 45.420 143.050 ;
        RECT 54.390 143.035 54.530 143.530 ;
        RECT 57.520 143.470 57.840 143.530 ;
        RECT 57.980 143.670 58.300 143.730 ;
        RECT 59.880 143.670 60.170 143.715 ;
        RECT 57.980 143.530 60.170 143.670 ;
        RECT 57.980 143.470 58.300 143.530 ;
        RECT 59.880 143.485 60.170 143.530 ;
        RECT 60.740 143.670 61.060 143.730 ;
        RECT 61.750 143.715 61.890 143.870 ;
        RECT 66.720 143.810 67.040 143.870 ;
        RECT 73.620 143.810 73.940 143.870 ;
        RECT 63.040 143.715 63.360 143.730 ;
        RECT 61.215 143.670 61.505 143.715 ;
        RECT 61.675 143.670 61.965 143.715 ;
        RECT 63.010 143.670 63.360 143.715 ;
        RECT 60.740 143.530 61.965 143.670 ;
        RECT 62.845 143.530 63.360 143.670 ;
        RECT 60.740 143.470 61.060 143.530 ;
        RECT 61.215 143.485 61.505 143.530 ;
        RECT 61.675 143.485 61.965 143.530 ;
        RECT 63.010 143.485 63.360 143.530 ;
        RECT 63.040 143.470 63.360 143.485 ;
        RECT 69.940 143.470 70.260 143.730 ;
        RECT 70.860 143.470 71.180 143.730 ;
        RECT 72.715 143.670 73.005 143.715 ;
        RECT 77.300 143.670 77.620 143.730 ;
        RECT 72.715 143.530 77.620 143.670 ;
        RECT 72.715 143.485 73.005 143.530 ;
        RECT 77.300 143.470 77.620 143.530 ;
        RECT 78.680 143.715 79.000 143.730 ;
        RECT 80.150 143.715 80.290 143.870 ;
        RECT 81.900 143.715 82.220 143.730 ;
        RECT 78.680 143.670 79.030 143.715 ;
        RECT 80.075 143.670 80.365 143.715 ;
        RECT 80.535 143.670 80.825 143.715 ;
        RECT 78.680 143.530 79.195 143.670 ;
        RECT 80.075 143.530 80.825 143.670 ;
        RECT 78.680 143.485 79.030 143.530 ;
        RECT 80.075 143.485 80.365 143.530 ;
        RECT 80.535 143.485 80.825 143.530 ;
        RECT 81.870 143.485 82.220 143.715 ;
        RECT 78.680 143.470 79.000 143.485 ;
        RECT 81.900 143.470 82.220 143.485 ;
        RECT 56.625 143.330 56.915 143.375 ;
        RECT 59.145 143.330 59.435 143.375 ;
        RECT 60.335 143.330 60.625 143.375 ;
        RECT 56.625 143.190 60.625 143.330 ;
        RECT 56.625 143.145 56.915 143.190 ;
        RECT 59.145 143.145 59.435 143.190 ;
        RECT 60.335 143.145 60.625 143.190 ;
        RECT 62.555 143.330 62.845 143.375 ;
        RECT 63.745 143.330 64.035 143.375 ;
        RECT 66.265 143.330 66.555 143.375 ;
        RECT 62.555 143.190 66.555 143.330 ;
        RECT 62.555 143.145 62.845 143.190 ;
        RECT 63.745 143.145 64.035 143.190 ;
        RECT 66.265 143.145 66.555 143.190 ;
        RECT 75.485 143.330 75.775 143.375 ;
        RECT 78.005 143.330 78.295 143.375 ;
        RECT 79.195 143.330 79.485 143.375 ;
        RECT 75.485 143.190 79.485 143.330 ;
        RECT 75.485 143.145 75.775 143.190 ;
        RECT 78.005 143.145 78.295 143.190 ;
        RECT 79.195 143.145 79.485 143.190 ;
        RECT 81.415 143.330 81.705 143.375 ;
        RECT 82.605 143.330 82.895 143.375 ;
        RECT 85.125 143.330 85.415 143.375 ;
        RECT 81.415 143.190 85.415 143.330 ;
        RECT 81.415 143.145 81.705 143.190 ;
        RECT 82.605 143.145 82.895 143.190 ;
        RECT 85.125 143.145 85.415 143.190 ;
        RECT 87.880 143.130 88.200 143.390 ;
        RECT 89.350 143.330 89.490 144.210 ;
        RECT 89.735 144.210 91.880 144.350 ;
        RECT 89.735 144.165 90.025 144.210 ;
        RECT 91.560 144.150 91.880 144.210 ;
        RECT 121.920 144.350 122.240 144.410 ;
        RECT 121.920 144.210 123.070 144.350 ;
        RECT 121.920 144.150 122.240 144.210 ;
        RECT 90.195 144.010 90.485 144.055 ;
        RECT 90.640 144.010 90.960 144.070 ;
        RECT 90.195 143.870 90.960 144.010 ;
        RECT 90.195 143.825 90.485 143.870 ;
        RECT 90.640 143.810 90.960 143.870 ;
        RECT 97.540 144.010 97.860 144.070 ;
        RECT 97.540 143.870 102.370 144.010 ;
        RECT 97.540 143.810 97.860 143.870 ;
        RECT 102.230 143.715 102.370 143.870 ;
        RECT 122.380 143.810 122.700 144.070 ;
        RECT 97.095 143.670 97.385 143.715 ;
        RECT 99.395 143.670 99.685 143.715 ;
        RECT 97.095 143.530 99.685 143.670 ;
        RECT 97.095 143.485 97.385 143.530 ;
        RECT 99.395 143.485 99.685 143.530 ;
        RECT 102.155 143.485 102.445 143.715 ;
        RECT 119.160 143.670 119.480 143.730 ;
        RECT 122.930 143.715 123.070 144.210 ;
        RECT 128.360 144.150 128.680 144.410 ;
        RECT 130.215 144.350 130.505 144.395 ;
        RECT 133.420 144.350 133.740 144.410 ;
        RECT 130.215 144.210 133.740 144.350 ;
        RECT 130.215 144.165 130.505 144.210 ;
        RECT 133.420 144.150 133.740 144.210 ;
        RECT 137.575 144.350 137.865 144.395 ;
        RECT 138.020 144.350 138.340 144.410 ;
        RECT 137.575 144.210 138.340 144.350 ;
        RECT 137.575 144.165 137.865 144.210 ;
        RECT 138.020 144.150 138.340 144.210 ;
        RECT 130.660 143.810 130.980 144.070 ;
        RECT 121.935 143.670 122.225 143.715 ;
        RECT 119.160 143.530 122.225 143.670 ;
        RECT 119.160 143.470 119.480 143.530 ;
        RECT 121.935 143.485 122.225 143.530 ;
        RECT 122.855 143.485 123.145 143.715 ;
        RECT 136.640 143.470 136.960 143.730 ;
        RECT 90.655 143.330 90.945 143.375 ;
        RECT 89.350 143.190 90.945 143.330 ;
        RECT 90.655 143.145 90.945 143.190 ;
        RECT 95.700 143.330 96.020 143.390 ;
        RECT 97.555 143.330 97.845 143.375 ;
        RECT 95.700 143.190 97.845 143.330 ;
        RECT 54.315 142.805 54.605 143.035 ;
        RECT 57.060 142.990 57.350 143.035 ;
        RECT 58.630 142.990 58.920 143.035 ;
        RECT 60.730 142.990 61.020 143.035 ;
        RECT 57.060 142.850 61.020 142.990 ;
        RECT 57.060 142.805 57.350 142.850 ;
        RECT 58.630 142.805 58.920 142.850 ;
        RECT 60.730 142.805 61.020 142.850 ;
        RECT 62.160 142.990 62.450 143.035 ;
        RECT 64.260 142.990 64.550 143.035 ;
        RECT 65.830 142.990 66.120 143.035 ;
        RECT 62.160 142.850 66.120 142.990 ;
        RECT 62.160 142.805 62.450 142.850 ;
        RECT 64.260 142.805 64.550 142.850 ;
        RECT 65.830 142.805 66.120 142.850 ;
        RECT 75.920 142.990 76.210 143.035 ;
        RECT 77.490 142.990 77.780 143.035 ;
        RECT 79.590 142.990 79.880 143.035 ;
        RECT 75.920 142.850 79.880 142.990 ;
        RECT 75.920 142.805 76.210 142.850 ;
        RECT 77.490 142.805 77.780 142.850 ;
        RECT 79.590 142.805 79.880 142.850 ;
        RECT 81.020 142.990 81.310 143.035 ;
        RECT 83.120 142.990 83.410 143.035 ;
        RECT 84.690 142.990 84.980 143.035 ;
        RECT 81.020 142.850 84.980 142.990 ;
        RECT 87.970 142.990 88.110 143.130 ;
        RECT 89.720 142.990 90.040 143.050 ;
        RECT 87.970 142.850 90.040 142.990 ;
        RECT 90.730 142.990 90.870 143.145 ;
        RECT 95.700 143.130 96.020 143.190 ;
        RECT 97.555 143.145 97.845 143.190 ;
        RECT 98.015 143.145 98.305 143.375 ;
        RECT 114.100 143.330 114.420 143.390 ;
        RECT 114.100 143.190 126.750 143.330 ;
        RECT 98.090 142.990 98.230 143.145 ;
        RECT 114.100 143.130 114.420 143.190 ;
        RECT 90.730 142.850 98.230 142.990 ;
        RECT 98.460 142.990 98.780 143.050 ;
        RECT 125.140 142.990 125.460 143.050 ;
        RECT 98.460 142.850 125.460 142.990 ;
        RECT 126.610 142.990 126.750 143.190 ;
        RECT 131.135 143.145 131.425 143.375 ;
        RECT 131.210 142.990 131.350 143.145 ;
        RECT 126.610 142.850 131.350 142.990 ;
        RECT 81.020 142.805 81.310 142.850 ;
        RECT 83.120 142.805 83.410 142.850 ;
        RECT 84.690 142.805 84.980 142.850 ;
        RECT 89.720 142.790 90.040 142.850 ;
        RECT 98.460 142.790 98.780 142.850 ;
        RECT 125.140 142.790 125.460 142.850 ;
        RECT 26.240 142.650 26.560 142.710 ;
        RECT 28.540 142.650 28.860 142.710 ;
        RECT 23.570 142.510 28.860 142.650 ;
        RECT 26.240 142.450 26.560 142.510 ;
        RECT 28.540 142.450 28.860 142.510 ;
        RECT 30.380 142.650 30.700 142.710 ;
        RECT 34.995 142.650 35.285 142.695 ;
        RECT 30.380 142.510 35.285 142.650 ;
        RECT 30.380 142.450 30.700 142.510 ;
        RECT 34.995 142.465 35.285 142.510 ;
        RECT 36.820 142.650 37.140 142.710 ;
        RECT 40.040 142.650 40.360 142.710 ;
        RECT 36.820 142.510 40.360 142.650 ;
        RECT 36.820 142.450 37.140 142.510 ;
        RECT 40.040 142.450 40.360 142.510 ;
        RECT 40.975 142.650 41.265 142.695 ;
        RECT 42.340 142.650 42.660 142.710 ;
        RECT 40.975 142.510 42.660 142.650 ;
        RECT 40.975 142.465 41.265 142.510 ;
        RECT 42.340 142.450 42.660 142.510 ;
        RECT 44.640 142.450 44.960 142.710 ;
        RECT 68.560 142.450 68.880 142.710 ;
        RECT 81.440 142.650 81.760 142.710 ;
        RECT 86.040 142.650 86.360 142.710 ;
        RECT 87.435 142.650 87.725 142.695 ;
        RECT 81.440 142.510 87.725 142.650 ;
        RECT 81.440 142.450 81.760 142.510 ;
        RECT 86.040 142.450 86.360 142.510 ;
        RECT 87.435 142.465 87.725 142.510 ;
        RECT 87.895 142.650 88.185 142.695 ;
        RECT 88.800 142.650 89.120 142.710 ;
        RECT 87.895 142.510 89.120 142.650 ;
        RECT 87.895 142.465 88.185 142.510 ;
        RECT 88.800 142.450 89.120 142.510 ;
        RECT 95.240 142.450 95.560 142.710 ;
        RECT 120.540 142.650 120.860 142.710 ;
        RECT 136.180 142.650 136.500 142.710 ;
        RECT 120.540 142.510 136.500 142.650 ;
        RECT 120.540 142.450 120.860 142.510 ;
        RECT 136.180 142.450 136.500 142.510 ;
        RECT 17.430 141.830 143.010 142.310 ;
        RECT 27.635 141.445 27.925 141.675 ;
        RECT 21.220 141.290 21.510 141.335 ;
        RECT 23.320 141.290 23.610 141.335 ;
        RECT 24.890 141.290 25.180 141.335 ;
        RECT 21.220 141.150 25.180 141.290 ;
        RECT 27.710 141.290 27.850 141.445 ;
        RECT 28.080 141.430 28.400 141.690 ;
        RECT 29.000 141.630 29.320 141.690 ;
        RECT 30.380 141.630 30.700 141.690 ;
        RECT 29.000 141.490 30.700 141.630 ;
        RECT 29.000 141.430 29.320 141.490 ;
        RECT 30.380 141.430 30.700 141.490 ;
        RECT 34.075 141.630 34.365 141.675 ;
        RECT 35.900 141.630 36.220 141.690 ;
        RECT 37.280 141.630 37.600 141.690 ;
        RECT 40.055 141.630 40.345 141.675 ;
        RECT 34.075 141.490 37.600 141.630 ;
        RECT 34.075 141.445 34.365 141.490 ;
        RECT 28.540 141.290 28.860 141.350 ;
        RECT 34.150 141.290 34.290 141.445 ;
        RECT 35.900 141.430 36.220 141.490 ;
        RECT 37.280 141.430 37.600 141.490 ;
        RECT 37.830 141.490 40.345 141.630 ;
        RECT 27.710 141.150 34.290 141.290 ;
        RECT 21.220 141.105 21.510 141.150 ;
        RECT 23.320 141.105 23.610 141.150 ;
        RECT 24.890 141.105 25.180 141.150 ;
        RECT 28.540 141.090 28.860 141.150 ;
        RECT 34.995 141.105 35.285 141.335 ;
        RECT 21.615 140.950 21.905 140.995 ;
        RECT 22.805 140.950 23.095 140.995 ;
        RECT 25.325 140.950 25.615 140.995 ;
        RECT 21.615 140.810 25.615 140.950 ;
        RECT 21.615 140.765 21.905 140.810 ;
        RECT 22.805 140.765 23.095 140.810 ;
        RECT 25.325 140.765 25.615 140.810 ;
        RECT 27.620 140.950 27.940 141.010 ;
        RECT 31.315 140.950 31.605 140.995 ;
        RECT 35.070 140.950 35.210 141.105 ;
        RECT 37.830 140.950 37.970 141.490 ;
        RECT 40.055 141.445 40.345 141.490 ;
        RECT 52.460 141.630 52.780 141.690 ;
        RECT 54.775 141.630 55.065 141.675 ;
        RECT 59.820 141.630 60.140 141.690 ;
        RECT 52.460 141.490 60.140 141.630 ;
        RECT 52.460 141.430 52.780 141.490 ;
        RECT 54.775 141.445 55.065 141.490 ;
        RECT 59.820 141.430 60.140 141.490 ;
        RECT 69.495 141.630 69.785 141.675 ;
        RECT 69.940 141.630 70.260 141.690 ;
        RECT 69.495 141.490 70.260 141.630 ;
        RECT 69.495 141.445 69.785 141.490 ;
        RECT 69.940 141.430 70.260 141.490 ;
        RECT 70.415 141.630 70.705 141.675 ;
        RECT 98.460 141.630 98.780 141.690 ;
        RECT 70.415 141.490 98.780 141.630 ;
        RECT 70.415 141.445 70.705 141.490 ;
        RECT 98.460 141.430 98.780 141.490 ;
        RECT 104.900 141.630 105.220 141.690 ;
        RECT 105.835 141.630 106.125 141.675 ;
        RECT 104.900 141.490 106.125 141.630 ;
        RECT 104.900 141.430 105.220 141.490 ;
        RECT 105.835 141.445 106.125 141.490 ;
        RECT 113.180 141.630 113.500 141.690 ;
        RECT 122.840 141.630 123.160 141.690 ;
        RECT 126.060 141.630 126.380 141.690 ;
        RECT 113.180 141.490 126.380 141.630 ;
        RECT 38.200 141.290 38.520 141.350 ;
        RECT 41.895 141.290 42.185 141.335 ;
        RECT 38.200 141.150 42.185 141.290 ;
        RECT 38.200 141.090 38.520 141.150 ;
        RECT 41.895 141.105 42.185 141.150 ;
        RECT 55.695 141.105 55.985 141.335 ;
        RECT 57.100 141.290 57.390 141.335 ;
        RECT 59.200 141.290 59.490 141.335 ;
        RECT 60.770 141.290 61.060 141.335 ;
        RECT 57.100 141.150 61.060 141.290 ;
        RECT 70.030 141.290 70.170 141.430 ;
        RECT 71.780 141.290 72.100 141.350 ;
        RECT 70.030 141.150 72.100 141.290 ;
        RECT 57.100 141.105 57.390 141.150 ;
        RECT 59.200 141.105 59.490 141.150 ;
        RECT 60.770 141.105 61.060 141.150 ;
        RECT 27.620 140.810 31.605 140.950 ;
        RECT 27.620 140.750 27.940 140.810 ;
        RECT 19.800 140.610 20.120 140.670 ;
        RECT 20.735 140.610 21.025 140.655 ;
        RECT 27.160 140.610 27.480 140.670 ;
        RECT 29.090 140.655 29.230 140.810 ;
        RECT 31.315 140.765 31.605 140.810 ;
        RECT 33.690 140.810 34.750 140.950 ;
        RECT 35.070 140.810 36.590 140.950 ;
        RECT 19.800 140.470 27.480 140.610 ;
        RECT 19.800 140.410 20.120 140.470 ;
        RECT 20.735 140.425 21.025 140.470 ;
        RECT 27.160 140.410 27.480 140.470 ;
        RECT 29.015 140.425 29.305 140.655 ;
        RECT 29.920 140.410 30.240 140.670 ;
        RECT 30.380 140.610 30.700 140.670 ;
        RECT 30.855 140.610 31.145 140.655 ;
        RECT 30.380 140.470 31.145 140.610 ;
        RECT 30.380 140.410 30.700 140.470 ;
        RECT 30.855 140.425 31.145 140.470 ;
        RECT 31.760 140.410 32.080 140.670 ;
        RECT 32.220 140.410 32.540 140.670 ;
        RECT 22.070 140.270 22.360 140.315 ;
        RECT 22.560 140.270 22.880 140.330 ;
        RECT 22.070 140.130 22.880 140.270 ;
        RECT 30.010 140.270 30.150 140.410 ;
        RECT 33.690 140.270 33.830 140.810 ;
        RECT 34.075 140.425 34.365 140.655 ;
        RECT 30.010 140.130 33.830 140.270 ;
        RECT 22.070 140.085 22.360 140.130 ;
        RECT 22.560 140.070 22.880 140.130 ;
        RECT 34.150 139.930 34.290 140.425 ;
        RECT 34.610 140.270 34.750 140.810 ;
        RECT 35.440 140.410 35.760 140.670 ;
        RECT 35.900 140.610 36.220 140.670 ;
        RECT 36.450 140.655 36.590 140.810 ;
        RECT 37.370 140.810 37.970 140.950 ;
        RECT 38.660 140.950 38.980 141.010 ;
        RECT 42.340 140.950 42.660 141.010 ;
        RECT 38.660 140.810 42.660 140.950 ;
        RECT 36.375 140.610 36.665 140.655 ;
        RECT 35.900 140.470 36.665 140.610 ;
        RECT 35.900 140.410 36.220 140.470 ;
        RECT 36.375 140.425 36.665 140.470 ;
        RECT 36.820 140.410 37.140 140.670 ;
        RECT 37.370 140.655 37.510 140.810 ;
        RECT 38.660 140.750 38.980 140.810 ;
        RECT 42.340 140.750 42.660 140.810 ;
        RECT 37.295 140.425 37.585 140.655 ;
        RECT 39.580 140.610 39.900 140.670 ;
        RECT 37.830 140.470 39.900 140.610 ;
        RECT 37.370 140.270 37.510 140.425 ;
        RECT 34.610 140.130 37.510 140.270 ;
        RECT 37.830 139.930 37.970 140.470 ;
        RECT 39.580 140.410 39.900 140.470 ;
        RECT 42.800 140.610 43.120 140.670 ;
        RECT 43.275 140.610 43.565 140.655 ;
        RECT 42.800 140.470 43.565 140.610 ;
        RECT 42.800 140.410 43.120 140.470 ;
        RECT 43.275 140.425 43.565 140.470 ;
        RECT 43.735 140.610 44.025 140.655 ;
        RECT 44.640 140.610 44.960 140.670 ;
        RECT 43.735 140.470 44.960 140.610 ;
        RECT 43.735 140.425 44.025 140.470 ;
        RECT 44.640 140.410 44.960 140.470 ;
        RECT 45.100 140.610 45.420 140.670 ;
        RECT 47.415 140.610 47.705 140.655 ;
        RECT 45.100 140.470 47.705 140.610 ;
        RECT 45.100 140.410 45.420 140.470 ;
        RECT 47.415 140.425 47.705 140.470 ;
        RECT 48.795 140.610 49.085 140.655 ;
        RECT 52.000 140.610 52.320 140.670 ;
        RECT 48.795 140.470 52.320 140.610 ;
        RECT 48.795 140.425 49.085 140.470 ;
        RECT 52.000 140.410 52.320 140.470 ;
        RECT 54.760 140.410 55.080 140.670 ;
        RECT 55.770 140.610 55.910 141.105 ;
        RECT 71.780 141.090 72.100 141.150 ;
        RECT 86.040 141.290 86.330 141.335 ;
        RECT 87.610 141.290 87.900 141.335 ;
        RECT 89.710 141.290 90.000 141.335 ;
        RECT 86.040 141.150 90.000 141.290 ;
        RECT 86.040 141.105 86.330 141.150 ;
        RECT 87.610 141.105 87.900 141.150 ;
        RECT 89.710 141.105 90.000 141.150 ;
        RECT 91.140 141.290 91.430 141.335 ;
        RECT 93.240 141.290 93.530 141.335 ;
        RECT 94.810 141.290 95.100 141.335 ;
        RECT 91.140 141.150 95.100 141.290 ;
        RECT 91.140 141.105 91.430 141.150 ;
        RECT 93.240 141.105 93.530 141.150 ;
        RECT 94.810 141.105 95.100 141.150 ;
        RECT 97.540 141.090 97.860 141.350 ;
        RECT 99.420 141.290 99.710 141.335 ;
        RECT 101.520 141.290 101.810 141.335 ;
        RECT 103.090 141.290 103.380 141.335 ;
        RECT 99.420 141.150 103.380 141.290 ;
        RECT 99.420 141.105 99.710 141.150 ;
        RECT 101.520 141.105 101.810 141.150 ;
        RECT 103.090 141.105 103.380 141.150 ;
        RECT 57.495 140.950 57.785 140.995 ;
        RECT 58.685 140.950 58.975 140.995 ;
        RECT 61.205 140.950 61.495 140.995 ;
        RECT 57.495 140.810 61.495 140.950 ;
        RECT 57.495 140.765 57.785 140.810 ;
        RECT 58.685 140.765 58.975 140.810 ;
        RECT 61.205 140.765 61.495 140.810 ;
        RECT 68.560 140.950 68.880 141.010 ;
        RECT 72.700 140.950 73.020 141.010 ;
        RECT 68.560 140.810 75.690 140.950 ;
        RECT 68.560 140.750 68.880 140.810 ;
        RECT 72.700 140.750 73.020 140.810 ;
        RECT 56.615 140.610 56.905 140.655 ;
        RECT 60.740 140.610 61.060 140.670 ;
        RECT 55.770 140.470 56.370 140.610 ;
        RECT 38.675 140.270 38.965 140.315 ;
        RECT 40.960 140.270 41.280 140.330 ;
        RECT 38.675 140.130 41.280 140.270 ;
        RECT 38.675 140.085 38.965 140.130 ;
        RECT 40.960 140.070 41.280 140.130 ;
        RECT 49.715 140.270 50.005 140.315 ;
        RECT 53.855 140.270 54.145 140.315 ;
        RECT 54.850 140.270 54.990 140.410 ;
        RECT 49.715 140.130 54.990 140.270 ;
        RECT 56.230 140.270 56.370 140.470 ;
        RECT 56.615 140.470 61.060 140.610 ;
        RECT 56.615 140.425 56.905 140.470 ;
        RECT 60.740 140.410 61.060 140.470 ;
        RECT 70.860 140.610 71.180 140.670 ;
        RECT 71.335 140.610 71.625 140.655 ;
        RECT 70.860 140.470 71.625 140.610 ;
        RECT 70.860 140.410 71.180 140.470 ;
        RECT 71.335 140.425 71.625 140.470 ;
        RECT 71.780 140.610 72.100 140.670 ;
        RECT 75.550 140.655 75.690 140.810 ;
        RECT 76.840 140.750 77.160 141.010 ;
        RECT 81.440 140.750 81.760 141.010 ;
        RECT 85.605 140.950 85.895 140.995 ;
        RECT 88.125 140.950 88.415 140.995 ;
        RECT 89.315 140.950 89.605 140.995 ;
        RECT 85.605 140.810 89.605 140.950 ;
        RECT 85.605 140.765 85.895 140.810 ;
        RECT 88.125 140.765 88.415 140.810 ;
        RECT 89.315 140.765 89.605 140.810 ;
        RECT 91.535 140.950 91.825 140.995 ;
        RECT 92.725 140.950 93.015 140.995 ;
        RECT 95.245 140.950 95.535 140.995 ;
        RECT 91.535 140.810 95.535 140.950 ;
        RECT 91.535 140.765 91.825 140.810 ;
        RECT 92.725 140.765 93.015 140.810 ;
        RECT 95.245 140.765 95.535 140.810 ;
        RECT 99.815 140.950 100.105 140.995 ;
        RECT 101.005 140.950 101.295 140.995 ;
        RECT 103.525 140.950 103.815 140.995 ;
        RECT 99.815 140.810 103.815 140.950 ;
        RECT 105.910 140.950 106.050 141.445 ;
        RECT 113.180 141.430 113.500 141.490 ;
        RECT 122.840 141.430 123.160 141.490 ;
        RECT 126.060 141.430 126.380 141.490 ;
        RECT 115.940 141.290 116.260 141.350 ;
        RECT 134.380 141.290 134.670 141.335 ;
        RECT 136.480 141.290 136.770 141.335 ;
        RECT 138.050 141.290 138.340 141.335 ;
        RECT 115.940 141.150 120.310 141.290 ;
        RECT 115.940 141.090 116.260 141.150 ;
        RECT 110.895 140.950 111.185 140.995 ;
        RECT 119.175 140.950 119.465 140.995 ;
        RECT 105.910 140.810 111.185 140.950 ;
        RECT 99.815 140.765 100.105 140.810 ;
        RECT 101.005 140.765 101.295 140.810 ;
        RECT 103.525 140.765 103.815 140.810 ;
        RECT 110.895 140.765 111.185 140.810 ;
        RECT 116.490 140.810 119.465 140.950 ;
        RECT 74.555 140.610 74.845 140.655 ;
        RECT 71.780 140.470 74.845 140.610 ;
        RECT 71.780 140.410 72.100 140.470 ;
        RECT 74.555 140.425 74.845 140.470 ;
        RECT 75.475 140.425 75.765 140.655 ;
        RECT 88.860 140.425 89.150 140.655 ;
        RECT 90.180 140.610 90.500 140.670 ;
        RECT 90.655 140.610 90.945 140.655 ;
        RECT 96.620 140.610 96.940 140.670 ;
        RECT 98.935 140.610 99.225 140.655 ;
        RECT 90.180 140.470 99.225 140.610 ;
        RECT 57.840 140.270 58.130 140.315 ;
        RECT 56.230 140.130 58.130 140.270 ;
        RECT 49.715 140.085 50.005 140.130 ;
        RECT 53.855 140.085 54.145 140.130 ;
        RECT 57.840 140.085 58.130 140.130 ;
        RECT 68.575 140.270 68.865 140.315 ;
        RECT 70.950 140.270 71.090 140.410 ;
        RECT 68.575 140.130 71.090 140.270 ;
        RECT 75.000 140.270 75.320 140.330 ;
        RECT 87.880 140.270 88.200 140.330 ;
        RECT 75.000 140.130 88.200 140.270 ;
        RECT 68.575 140.085 68.865 140.130 ;
        RECT 75.000 140.070 75.320 140.130 ;
        RECT 87.880 140.070 88.200 140.130 ;
        RECT 88.935 139.990 89.075 140.425 ;
        RECT 90.180 140.410 90.500 140.470 ;
        RECT 90.655 140.425 90.945 140.470 ;
        RECT 96.620 140.410 96.940 140.470 ;
        RECT 98.935 140.425 99.225 140.470 ;
        RECT 104.440 140.610 104.760 140.670 ;
        RECT 116.490 140.655 116.630 140.810 ;
        RECT 119.175 140.765 119.465 140.810 ;
        RECT 114.575 140.610 114.865 140.655 ;
        RECT 104.440 140.470 114.865 140.610 ;
        RECT 104.440 140.410 104.760 140.470 ;
        RECT 114.575 140.425 114.865 140.470 ;
        RECT 115.495 140.425 115.785 140.655 ;
        RECT 116.415 140.425 116.705 140.655 ;
        RECT 116.875 140.425 117.165 140.655 ;
        RECT 91.990 140.270 92.280 140.315 ;
        RECT 95.240 140.270 95.560 140.330 ;
        RECT 91.990 140.130 95.560 140.270 ;
        RECT 91.990 140.085 92.280 140.130 ;
        RECT 95.240 140.070 95.560 140.130 ;
        RECT 100.270 140.270 100.560 140.315 ;
        RECT 104.900 140.270 105.220 140.330 ;
        RECT 100.270 140.130 105.220 140.270 ;
        RECT 100.270 140.085 100.560 140.130 ;
        RECT 104.900 140.070 105.220 140.130 ;
        RECT 114.100 140.270 114.420 140.330 ;
        RECT 115.570 140.270 115.710 140.425 ;
        RECT 114.100 140.130 115.710 140.270 ;
        RECT 114.100 140.070 114.420 140.130 ;
        RECT 34.150 139.790 37.970 139.930 ;
        RECT 39.120 139.730 39.440 139.990 ;
        RECT 40.040 139.730 40.360 139.990 ;
        RECT 43.735 139.930 44.025 139.975 ;
        RECT 44.180 139.930 44.500 139.990 ;
        RECT 43.735 139.790 44.500 139.930 ;
        RECT 43.735 139.745 44.025 139.790 ;
        RECT 44.180 139.730 44.500 139.790 ;
        RECT 47.875 139.930 48.165 139.975 ;
        RECT 49.240 139.930 49.560 139.990 ;
        RECT 47.875 139.790 49.560 139.930 ;
        RECT 47.875 139.745 48.165 139.790 ;
        RECT 49.240 139.730 49.560 139.790 ;
        RECT 54.905 139.930 55.195 139.975 ;
        RECT 58.440 139.930 58.760 139.990 ;
        RECT 54.905 139.790 58.760 139.930 ;
        RECT 54.905 139.745 55.195 139.790 ;
        RECT 58.440 139.730 58.760 139.790 ;
        RECT 59.820 139.930 60.140 139.990 ;
        RECT 63.515 139.930 63.805 139.975 ;
        RECT 59.820 139.790 63.805 139.930 ;
        RECT 59.820 139.730 60.140 139.790 ;
        RECT 63.515 139.745 63.805 139.790 ;
        RECT 69.625 139.930 69.915 139.975 ;
        RECT 73.620 139.930 73.940 139.990 ;
        RECT 69.625 139.790 73.940 139.930 ;
        RECT 69.625 139.745 69.915 139.790 ;
        RECT 73.620 139.730 73.940 139.790 ;
        RECT 78.235 139.930 78.525 139.975 ;
        RECT 79.600 139.930 79.920 139.990 ;
        RECT 78.235 139.790 79.920 139.930 ;
        RECT 78.235 139.745 78.525 139.790 ;
        RECT 79.600 139.730 79.920 139.790 ;
        RECT 83.295 139.930 83.585 139.975 ;
        RECT 88.340 139.930 88.660 139.990 ;
        RECT 83.295 139.790 88.660 139.930 ;
        RECT 83.295 139.745 83.585 139.790 ;
        RECT 88.340 139.730 88.660 139.790 ;
        RECT 88.800 139.730 89.120 139.990 ;
        RECT 106.740 139.930 107.060 139.990 ;
        RECT 108.135 139.930 108.425 139.975 ;
        RECT 106.740 139.790 108.425 139.930 ;
        RECT 106.740 139.730 107.060 139.790 ;
        RECT 108.135 139.745 108.425 139.790 ;
        RECT 110.880 139.930 111.200 139.990 ;
        RECT 111.815 139.930 112.105 139.975 ;
        RECT 110.880 139.790 112.105 139.930 ;
        RECT 110.880 139.730 111.200 139.790 ;
        RECT 111.815 139.745 112.105 139.790 ;
        RECT 115.480 139.930 115.800 139.990 ;
        RECT 116.950 139.930 117.090 140.425 ;
        RECT 117.320 140.410 117.640 140.670 ;
        RECT 120.170 140.655 120.310 141.150 ;
        RECT 134.380 141.150 138.340 141.290 ;
        RECT 134.380 141.105 134.670 141.150 ;
        RECT 136.480 141.105 136.770 141.150 ;
        RECT 138.050 141.105 138.340 141.150 ;
        RECT 134.775 140.950 135.065 140.995 ;
        RECT 135.965 140.950 136.255 140.995 ;
        RECT 138.485 140.950 138.775 140.995 ;
        RECT 134.775 140.810 138.775 140.950 ;
        RECT 134.775 140.765 135.065 140.810 ;
        RECT 135.965 140.765 136.255 140.810 ;
        RECT 138.485 140.765 138.775 140.810 ;
        RECT 120.095 140.610 120.385 140.655 ;
        RECT 128.820 140.610 129.140 140.670 ;
        RECT 120.095 140.470 129.140 140.610 ;
        RECT 120.095 140.425 120.385 140.470 ;
        RECT 128.820 140.410 129.140 140.470 ;
        RECT 133.880 140.410 134.200 140.670 ;
        RECT 117.410 140.270 117.550 140.410 ;
        RECT 117.410 140.130 120.770 140.270 ;
        RECT 115.480 139.790 117.090 139.930 ;
        RECT 115.480 139.730 115.800 139.790 ;
        RECT 118.700 139.730 119.020 139.990 ;
        RECT 120.630 139.930 120.770 140.130 ;
        RECT 121.000 140.070 121.320 140.330 ;
        RECT 133.420 140.270 133.740 140.330 ;
        RECT 135.120 140.270 135.410 140.315 ;
        RECT 133.420 140.130 135.410 140.270 ;
        RECT 133.420 140.070 133.740 140.130 ;
        RECT 135.120 140.085 135.410 140.130 ;
        RECT 127.900 139.930 128.220 139.990 ;
        RECT 132.040 139.930 132.360 139.990 ;
        RECT 120.630 139.790 132.360 139.930 ;
        RECT 127.900 139.730 128.220 139.790 ;
        RECT 132.040 139.730 132.360 139.790 ;
        RECT 140.320 139.930 140.640 139.990 ;
        RECT 140.795 139.930 141.085 139.975 ;
        RECT 140.320 139.790 141.085 139.930 ;
        RECT 140.320 139.730 140.640 139.790 ;
        RECT 140.795 139.745 141.085 139.790 ;
        RECT 17.430 139.110 143.010 139.590 ;
        RECT 12.440 138.910 12.760 138.970 ;
        RECT 12.440 138.770 78.450 138.910 ;
        RECT 12.440 138.710 12.760 138.770 ;
        RECT 27.635 138.570 27.925 138.615 ;
        RECT 38.200 138.570 38.520 138.630 ;
        RECT 40.515 138.570 40.805 138.615 ;
        RECT 43.260 138.570 43.580 138.630 ;
        RECT 43.735 138.570 44.025 138.615 ;
        RECT 27.635 138.430 28.770 138.570 ;
        RECT 27.635 138.385 27.925 138.430 ;
        RECT 19.800 138.030 20.120 138.290 ;
        RECT 21.180 138.275 21.500 138.290 ;
        RECT 21.150 138.230 21.500 138.275 ;
        RECT 20.985 138.090 21.500 138.230 ;
        RECT 21.150 138.045 21.500 138.090 ;
        RECT 21.180 138.030 21.500 138.045 ;
        RECT 26.700 138.230 27.020 138.290 ;
        RECT 27.175 138.230 27.465 138.275 ;
        RECT 26.700 138.090 27.465 138.230 ;
        RECT 26.700 138.030 27.020 138.090 ;
        RECT 27.175 138.045 27.465 138.090 ;
        RECT 28.080 138.030 28.400 138.290 ;
        RECT 28.630 138.275 28.770 138.430 ;
        RECT 38.200 138.430 39.350 138.570 ;
        RECT 38.200 138.370 38.520 138.430 ;
        RECT 28.555 138.045 28.845 138.275 ;
        RECT 29.475 138.230 29.765 138.275 ;
        RECT 30.840 138.230 31.160 138.290 ;
        RECT 29.475 138.090 31.160 138.230 ;
        RECT 29.475 138.045 29.765 138.090 ;
        RECT 20.695 137.890 20.985 137.935 ;
        RECT 21.885 137.890 22.175 137.935 ;
        RECT 24.405 137.890 24.695 137.935 ;
        RECT 20.695 137.750 24.695 137.890 ;
        RECT 20.695 137.705 20.985 137.750 ;
        RECT 21.885 137.705 22.175 137.750 ;
        RECT 24.405 137.705 24.695 137.750 ;
        RECT 26.240 137.890 26.560 137.950 ;
        RECT 27.620 137.890 27.940 137.950 ;
        RECT 29.550 137.890 29.690 138.045 ;
        RECT 30.840 138.030 31.160 138.090 ;
        RECT 35.900 138.230 36.220 138.290 ;
        RECT 36.375 138.230 36.665 138.275 ;
        RECT 35.900 138.090 36.665 138.230 ;
        RECT 35.900 138.030 36.220 138.090 ;
        RECT 36.375 138.045 36.665 138.090 ;
        RECT 37.755 138.045 38.045 138.275 ;
        RECT 26.240 137.750 26.930 137.890 ;
        RECT 26.240 137.690 26.560 137.750 ;
        RECT 26.790 137.595 26.930 137.750 ;
        RECT 27.620 137.750 29.690 137.890 ;
        RECT 27.620 137.690 27.940 137.750 ;
        RECT 20.300 137.550 20.590 137.595 ;
        RECT 22.400 137.550 22.690 137.595 ;
        RECT 23.970 137.550 24.260 137.595 ;
        RECT 20.300 137.410 24.260 137.550 ;
        RECT 20.300 137.365 20.590 137.410 ;
        RECT 22.400 137.365 22.690 137.410 ;
        RECT 23.970 137.365 24.260 137.410 ;
        RECT 26.715 137.365 27.005 137.595 ;
        RECT 28.540 137.010 28.860 137.270 ;
        RECT 36.820 137.010 37.140 137.270 ;
        RECT 37.830 137.210 37.970 138.045 ;
        RECT 38.660 138.030 38.980 138.290 ;
        RECT 39.210 138.275 39.350 138.430 ;
        RECT 40.515 138.430 44.025 138.570 ;
        RECT 40.515 138.385 40.805 138.430 ;
        RECT 43.260 138.370 43.580 138.430 ;
        RECT 43.735 138.385 44.025 138.430 ;
        RECT 44.180 138.570 44.500 138.630 ;
        RECT 44.735 138.570 45.025 138.615 ;
        RECT 44.180 138.430 45.025 138.570 ;
        RECT 44.180 138.370 44.500 138.430 ;
        RECT 44.735 138.385 45.025 138.430 ;
        RECT 45.190 138.430 50.850 138.570 ;
        RECT 39.135 138.045 39.425 138.275 ;
        RECT 39.580 138.030 39.900 138.290 ;
        RECT 40.960 138.030 41.280 138.290 ;
        RECT 41.435 138.045 41.725 138.275 ;
        RECT 41.880 138.230 42.200 138.290 ;
        RECT 45.190 138.230 45.330 138.430 ;
        RECT 50.710 138.290 50.850 138.430 ;
        RECT 52.000 138.370 52.320 138.630 ;
        RECT 53.380 138.370 53.700 138.630 ;
        RECT 55.680 138.570 56.000 138.630 ;
        RECT 54.850 138.430 56.000 138.570 ;
        RECT 47.415 138.230 47.705 138.275 ;
        RECT 41.880 138.090 45.330 138.230 ;
        RECT 45.650 138.090 47.705 138.230 ;
        RECT 38.215 137.890 38.505 137.935 ;
        RECT 41.510 137.890 41.650 138.045 ;
        RECT 41.880 138.030 42.200 138.090 ;
        RECT 45.100 137.890 45.420 137.950 ;
        RECT 38.215 137.750 41.650 137.890 ;
        RECT 42.430 137.750 45.420 137.890 ;
        RECT 38.215 137.705 38.505 137.750 ;
        RECT 38.660 137.550 38.980 137.610 ;
        RECT 40.040 137.550 40.360 137.610 ;
        RECT 41.880 137.550 42.200 137.610 ;
        RECT 42.430 137.595 42.570 137.750 ;
        RECT 45.100 137.690 45.420 137.750 ;
        RECT 45.650 137.595 45.790 138.090 ;
        RECT 47.415 138.045 47.705 138.090 ;
        RECT 48.795 138.230 49.085 138.275 ;
        RECT 49.240 138.230 49.560 138.290 ;
        RECT 48.795 138.090 49.560 138.230 ;
        RECT 48.795 138.045 49.085 138.090 ;
        RECT 49.240 138.030 49.560 138.090 ;
        RECT 50.160 138.030 50.480 138.290 ;
        RECT 50.620 138.230 50.940 138.290 ;
        RECT 50.620 138.090 53.150 138.230 ;
        RECT 53.390 138.155 53.680 138.370 ;
        RECT 54.850 138.275 54.990 138.430 ;
        RECT 55.680 138.370 56.000 138.430 ;
        RECT 58.900 138.370 59.220 138.630 ;
        RECT 59.360 138.570 59.680 138.630 ;
        RECT 59.915 138.570 60.205 138.615 ;
        RECT 61.675 138.570 61.965 138.615 ;
        RECT 59.360 138.430 60.205 138.570 ;
        RECT 59.360 138.370 59.680 138.430 ;
        RECT 59.915 138.385 60.205 138.430 ;
        RECT 60.370 138.430 61.965 138.570 ;
        RECT 50.620 138.030 50.940 138.090 ;
        RECT 52.000 137.690 52.320 137.950 ;
        RECT 38.660 137.410 40.360 137.550 ;
        RECT 38.660 137.350 38.980 137.410 ;
        RECT 40.040 137.350 40.360 137.410 ;
        RECT 40.590 137.410 42.200 137.550 ;
        RECT 40.590 137.210 40.730 137.410 ;
        RECT 41.880 137.350 42.200 137.410 ;
        RECT 42.355 137.365 42.645 137.595 ;
        RECT 45.575 137.365 45.865 137.595 ;
        RECT 48.320 137.550 48.640 137.610 ;
        RECT 52.460 137.550 52.780 137.610 ;
        RECT 48.320 137.410 52.780 137.550 ;
        RECT 53.010 137.550 53.150 138.090 ;
        RECT 53.855 138.035 54.145 138.265 ;
        RECT 54.775 138.045 55.065 138.275 ;
        RECT 55.265 138.045 55.555 138.275 ;
        RECT 53.930 137.890 54.070 138.035 ;
        RECT 54.300 137.890 54.620 137.950 ;
        RECT 53.930 137.750 54.620 137.890 ;
        RECT 54.300 137.690 54.620 137.750 ;
        RECT 54.850 137.550 54.990 138.045 ;
        RECT 55.340 137.890 55.480 138.045 ;
        RECT 56.140 138.030 56.460 138.290 ;
        RECT 56.615 138.230 56.905 138.275 ;
        RECT 56.615 138.045 56.910 138.230 ;
        RECT 57.075 138.220 57.365 138.275 ;
        RECT 57.520 138.220 57.840 138.290 ;
        RECT 57.075 138.080 57.840 138.220 ;
        RECT 57.075 138.045 57.365 138.080 ;
        RECT 55.340 137.750 55.495 137.890 ;
        RECT 53.010 137.410 54.990 137.550 ;
        RECT 48.320 137.350 48.640 137.410 ;
        RECT 52.460 137.350 52.780 137.410 ;
        RECT 37.830 137.070 40.730 137.210 ;
        RECT 40.960 137.210 41.280 137.270 ;
        RECT 44.655 137.210 44.945 137.255 ;
        RECT 40.960 137.070 44.945 137.210 ;
        RECT 40.960 137.010 41.280 137.070 ;
        RECT 44.655 137.025 44.945 137.070 ;
        RECT 51.080 137.210 51.400 137.270 ;
        RECT 52.935 137.210 53.225 137.255 ;
        RECT 51.080 137.070 53.225 137.210 ;
        RECT 51.080 137.010 51.400 137.070 ;
        RECT 52.935 137.025 53.225 137.070 ;
        RECT 53.380 137.210 53.700 137.270 ;
        RECT 54.315 137.210 54.605 137.255 ;
        RECT 53.380 137.070 54.605 137.210 ;
        RECT 55.355 137.210 55.495 137.750 ;
        RECT 56.770 137.850 56.910 138.045 ;
        RECT 57.520 138.030 57.840 138.080 ;
        RECT 58.440 138.230 58.760 138.290 ;
        RECT 60.370 138.230 60.510 138.430 ;
        RECT 61.675 138.385 61.965 138.430 ;
        RECT 72.700 138.370 73.020 138.630 ;
        RECT 78.310 138.615 78.450 138.770 ;
        RECT 85.580 138.710 85.900 138.970 ;
        RECT 91.100 138.910 91.420 138.970 ;
        RECT 92.940 138.910 93.260 138.970 ;
        RECT 94.335 138.910 94.625 138.955 ;
        RECT 91.100 138.770 94.625 138.910 ;
        RECT 91.100 138.710 91.420 138.770 ;
        RECT 92.940 138.710 93.260 138.770 ;
        RECT 94.335 138.725 94.625 138.770 ;
        RECT 104.440 138.710 104.760 138.970 ;
        RECT 104.900 138.710 105.220 138.970 ;
        RECT 106.740 138.710 107.060 138.970 ;
        RECT 109.055 138.725 109.345 138.955 ;
        RECT 88.800 138.615 89.120 138.630 ;
        RECT 74.095 138.385 74.385 138.615 ;
        RECT 75.175 138.570 75.465 138.615 ;
        RECT 76.855 138.570 77.145 138.615 ;
        RECT 75.175 138.430 77.145 138.570 ;
        RECT 75.175 138.385 75.465 138.430 ;
        RECT 76.855 138.385 77.145 138.430 ;
        RECT 78.235 138.385 78.525 138.615 ;
        RECT 88.660 138.385 89.120 138.615 ;
        RECT 98.890 138.570 99.180 138.615 ;
        RECT 109.130 138.570 109.270 138.725 ;
        RECT 110.880 138.710 111.200 138.970 ;
        RECT 112.260 138.910 112.580 138.970 ;
        RECT 117.320 138.910 117.640 138.970 ;
        RECT 112.260 138.770 117.640 138.910 ;
        RECT 112.260 138.710 112.580 138.770 ;
        RECT 117.320 138.710 117.640 138.770 ;
        RECT 118.700 138.910 119.020 138.970 ;
        RECT 127.915 138.910 128.205 138.955 ;
        RECT 128.820 138.910 129.140 138.970 ;
        RECT 118.700 138.770 122.380 138.910 ;
        RECT 118.700 138.710 119.020 138.770 ;
        RECT 122.240 138.615 122.380 138.770 ;
        RECT 127.915 138.770 129.140 138.910 ;
        RECT 127.915 138.725 128.205 138.770 ;
        RECT 128.820 138.710 129.140 138.770 ;
        RECT 133.420 138.710 133.740 138.970 ;
        RECT 138.940 138.710 139.260 138.970 ;
        RECT 140.780 138.710 141.100 138.970 ;
        RECT 98.890 138.430 109.270 138.570 ;
        RECT 113.270 138.430 116.630 138.570 ;
        RECT 98.890 138.385 99.180 138.430 ;
        RECT 58.440 138.090 60.510 138.230 ;
        RECT 58.440 138.030 58.760 138.090 ;
        RECT 61.215 138.045 61.505 138.275 ;
        RECT 61.290 137.890 61.430 138.045 ;
        RECT 62.120 138.030 62.440 138.290 ;
        RECT 70.860 138.030 71.180 138.290 ;
        RECT 74.170 138.230 74.310 138.385 ;
        RECT 88.800 138.370 89.120 138.385 ;
        RECT 75.920 138.230 76.240 138.290 ;
        RECT 74.170 138.090 76.240 138.230 ;
        RECT 75.920 138.030 76.240 138.090 ;
        RECT 77.300 138.030 77.620 138.290 ;
        RECT 87.420 138.030 87.740 138.290 ;
        RECT 96.160 138.230 96.480 138.290 ;
        RECT 87.970 138.090 96.480 138.230 ;
        RECT 75.000 137.890 75.320 137.950 ;
        RECT 80.060 137.890 80.380 137.950 ;
        RECT 87.970 137.890 88.110 138.090 ;
        RECT 96.160 138.030 96.480 138.090 ;
        RECT 96.620 138.230 96.940 138.290 ;
        RECT 97.555 138.230 97.845 138.275 ;
        RECT 96.620 138.090 97.845 138.230 ;
        RECT 96.620 138.030 96.940 138.090 ;
        RECT 97.555 138.045 97.845 138.090 ;
        RECT 107.215 138.230 107.505 138.275 ;
        RECT 109.500 138.230 109.820 138.290 ;
        RECT 107.215 138.090 109.820 138.230 ;
        RECT 107.215 138.045 107.505 138.090 ;
        RECT 109.500 138.030 109.820 138.090 ;
        RECT 111.355 138.230 111.645 138.275 ;
        RECT 112.720 138.230 113.040 138.290 ;
        RECT 113.270 138.275 113.410 138.430 ;
        RECT 116.490 138.290 116.630 138.430 ;
        RECT 122.240 138.385 122.530 138.615 ;
        RECT 130.660 138.570 130.980 138.630 ;
        RECT 134.340 138.570 134.660 138.630 ;
        RECT 130.660 138.430 131.810 138.570 ;
        RECT 130.660 138.370 130.980 138.430 ;
        RECT 111.355 138.090 113.040 138.230 ;
        RECT 111.355 138.045 111.645 138.090 ;
        RECT 112.720 138.030 113.040 138.090 ;
        RECT 113.195 138.045 113.485 138.275 ;
        RECT 113.640 138.230 113.960 138.290 ;
        RECT 114.475 138.230 114.765 138.275 ;
        RECT 113.640 138.090 114.765 138.230 ;
        RECT 113.640 138.030 113.960 138.090 ;
        RECT 114.475 138.045 114.765 138.090 ;
        RECT 116.400 138.230 116.720 138.290 ;
        RECT 120.080 138.230 120.400 138.290 ;
        RECT 121.015 138.230 121.305 138.275 ;
        RECT 116.400 138.090 121.305 138.230 ;
        RECT 116.400 138.030 116.720 138.090 ;
        RECT 120.080 138.030 120.400 138.090 ;
        RECT 121.015 138.045 121.305 138.090 ;
        RECT 121.460 138.030 121.780 138.290 ;
        RECT 131.670 138.275 131.810 138.430 ;
        RECT 132.130 138.430 134.660 138.570 ;
        RECT 132.130 138.290 132.270 138.430 ;
        RECT 134.340 138.370 134.660 138.430 ;
        RECT 134.815 138.570 135.105 138.615 ;
        RECT 140.320 138.570 140.640 138.630 ;
        RECT 134.815 138.430 140.640 138.570 ;
        RECT 134.815 138.385 135.105 138.430 ;
        RECT 140.320 138.370 140.640 138.430 ;
        RECT 130.215 138.045 130.505 138.275 ;
        RECT 131.135 138.045 131.425 138.275 ;
        RECT 131.595 138.045 131.885 138.275 ;
        RECT 57.915 137.850 61.430 137.890 ;
        RECT 56.770 137.750 61.430 137.850 ;
        RECT 73.710 137.750 75.320 137.890 ;
        RECT 56.770 137.710 58.055 137.750 ;
        RECT 60.830 137.595 60.970 137.750 ;
        RECT 73.710 137.595 73.850 137.750 ;
        RECT 75.000 137.690 75.320 137.750 ;
        RECT 76.010 137.750 88.110 137.890 ;
        RECT 88.315 137.890 88.605 137.935 ;
        RECT 89.505 137.890 89.795 137.935 ;
        RECT 92.025 137.890 92.315 137.935 ;
        RECT 88.315 137.750 92.315 137.890 ;
        RECT 76.010 137.595 76.150 137.750 ;
        RECT 80.060 137.690 80.380 137.750 ;
        RECT 88.315 137.705 88.605 137.750 ;
        RECT 89.505 137.705 89.795 137.750 ;
        RECT 92.025 137.705 92.315 137.750 ;
        RECT 98.435 137.890 98.725 137.935 ;
        RECT 99.625 137.890 99.915 137.935 ;
        RECT 102.145 137.890 102.435 137.935 ;
        RECT 98.435 137.750 102.435 137.890 ;
        RECT 98.435 137.705 98.725 137.750 ;
        RECT 99.625 137.705 99.915 137.750 ;
        RECT 102.145 137.705 102.435 137.750 ;
        RECT 107.675 137.705 107.965 137.935 ;
        RECT 111.815 137.705 112.105 137.935 ;
        RECT 114.075 137.890 114.365 137.935 ;
        RECT 115.265 137.890 115.555 137.935 ;
        RECT 117.785 137.890 118.075 137.935 ;
        RECT 121.550 137.890 121.690 138.030 ;
        RECT 114.075 137.750 118.075 137.890 ;
        RECT 114.075 137.705 114.365 137.750 ;
        RECT 115.265 137.705 115.555 137.750 ;
        RECT 117.785 137.705 118.075 137.750 ;
        RECT 118.790 137.750 121.690 137.890 ;
        RECT 121.895 137.890 122.185 137.935 ;
        RECT 123.085 137.890 123.375 137.935 ;
        RECT 125.605 137.890 125.895 137.935 ;
        RECT 121.895 137.750 125.895 137.890 ;
        RECT 60.755 137.550 61.045 137.595 ;
        RECT 60.755 137.410 61.155 137.550 ;
        RECT 60.755 137.365 61.045 137.410 ;
        RECT 73.635 137.365 73.925 137.595 ;
        RECT 75.935 137.365 76.225 137.595 ;
        RECT 87.920 137.550 88.210 137.595 ;
        RECT 90.020 137.550 90.310 137.595 ;
        RECT 91.590 137.550 91.880 137.595 ;
        RECT 87.920 137.410 91.880 137.550 ;
        RECT 87.920 137.365 88.210 137.410 ;
        RECT 90.020 137.365 90.310 137.410 ;
        RECT 91.590 137.365 91.880 137.410 ;
        RECT 98.040 137.550 98.330 137.595 ;
        RECT 100.140 137.550 100.430 137.595 ;
        RECT 101.710 137.550 102.000 137.595 ;
        RECT 98.040 137.410 102.000 137.550 ;
        RECT 98.040 137.365 98.330 137.410 ;
        RECT 100.140 137.365 100.430 137.410 ;
        RECT 101.710 137.365 102.000 137.410 ;
        RECT 103.520 137.550 103.840 137.610 ;
        RECT 107.750 137.550 107.890 137.705 ;
        RECT 111.890 137.550 112.030 137.705 ;
        RECT 103.520 137.410 112.030 137.550 ;
        RECT 113.680 137.550 113.970 137.595 ;
        RECT 115.780 137.550 116.070 137.595 ;
        RECT 117.350 137.550 117.640 137.595 ;
        RECT 113.680 137.410 117.640 137.550 ;
        RECT 103.520 137.350 103.840 137.410 ;
        RECT 113.680 137.365 113.970 137.410 ;
        RECT 115.780 137.365 116.070 137.410 ;
        RECT 117.350 137.365 117.640 137.410 ;
        RECT 57.060 137.210 57.380 137.270 ;
        RECT 55.355 137.070 57.380 137.210 ;
        RECT 53.380 137.010 53.700 137.070 ;
        RECT 54.315 137.025 54.605 137.070 ;
        RECT 57.060 137.010 57.380 137.070 ;
        RECT 57.980 137.210 58.300 137.270 ;
        RECT 58.455 137.210 58.745 137.255 ;
        RECT 57.980 137.070 58.745 137.210 ;
        RECT 57.980 137.010 58.300 137.070 ;
        RECT 58.455 137.025 58.745 137.070 ;
        RECT 59.820 137.010 60.140 137.270 ;
        RECT 71.320 137.210 71.640 137.270 ;
        RECT 72.240 137.210 72.560 137.270 ;
        RECT 72.715 137.210 73.005 137.255 ;
        RECT 71.320 137.070 73.005 137.210 ;
        RECT 71.320 137.010 71.640 137.070 ;
        RECT 72.240 137.010 72.560 137.070 ;
        RECT 72.715 137.025 73.005 137.070 ;
        RECT 74.080 137.210 74.400 137.270 ;
        RECT 75.015 137.210 75.305 137.255 ;
        RECT 74.080 137.070 75.305 137.210 ;
        RECT 74.080 137.010 74.400 137.070 ;
        RECT 75.015 137.025 75.305 137.070 ;
        RECT 114.100 137.210 114.420 137.270 ;
        RECT 118.790 137.210 118.930 137.750 ;
        RECT 121.895 137.705 122.185 137.750 ;
        RECT 123.085 137.705 123.375 137.750 ;
        RECT 125.605 137.705 125.895 137.750 ;
        RECT 119.160 137.550 119.480 137.610 ;
        RECT 120.095 137.550 120.385 137.595 ;
        RECT 120.540 137.550 120.860 137.610 ;
        RECT 119.160 137.410 120.860 137.550 ;
        RECT 119.160 137.350 119.480 137.410 ;
        RECT 120.095 137.365 120.385 137.410 ;
        RECT 120.540 137.350 120.860 137.410 ;
        RECT 121.500 137.550 121.790 137.595 ;
        RECT 123.600 137.550 123.890 137.595 ;
        RECT 125.170 137.550 125.460 137.595 ;
        RECT 130.290 137.550 130.430 138.045 ;
        RECT 131.210 137.890 131.350 138.045 ;
        RECT 132.040 138.030 132.360 138.290 ;
        RECT 132.500 138.230 132.820 138.290 ;
        RECT 133.895 138.230 134.185 138.275 ;
        RECT 132.500 138.090 134.185 138.230 ;
        RECT 132.500 138.030 132.820 138.090 ;
        RECT 133.895 138.045 134.185 138.090 ;
        RECT 138.020 138.030 138.340 138.290 ;
        RECT 139.875 138.045 140.165 138.275 ;
        RECT 135.735 137.890 136.025 137.935 ;
        RECT 131.210 137.750 136.025 137.890 ;
        RECT 135.735 137.705 136.025 137.750 ;
        RECT 121.500 137.410 125.460 137.550 ;
        RECT 121.500 137.365 121.790 137.410 ;
        RECT 123.600 137.365 123.890 137.410 ;
        RECT 125.170 137.365 125.460 137.410 ;
        RECT 126.150 137.410 130.430 137.550 ;
        RECT 114.100 137.070 118.930 137.210 ;
        RECT 119.620 137.210 119.940 137.270 ;
        RECT 126.150 137.210 126.290 137.410 ;
        RECT 119.620 137.070 126.290 137.210 ;
        RECT 126.520 137.210 126.840 137.270 ;
        RECT 139.950 137.210 140.090 138.045 ;
        RECT 126.520 137.070 140.090 137.210 ;
        RECT 114.100 137.010 114.420 137.070 ;
        RECT 119.620 137.010 119.940 137.070 ;
        RECT 126.520 137.010 126.840 137.070 ;
        RECT 17.430 136.390 143.010 136.870 ;
        RECT 22.560 135.990 22.880 136.250 ;
        RECT 23.495 136.190 23.785 136.235 ;
        RECT 24.860 136.190 25.180 136.250 ;
        RECT 23.495 136.050 25.180 136.190 ;
        RECT 23.495 136.005 23.785 136.050 ;
        RECT 24.860 135.990 25.180 136.050 ;
        RECT 37.755 136.190 38.045 136.235 ;
        RECT 38.200 136.190 38.520 136.250 ;
        RECT 37.755 136.050 38.520 136.190 ;
        RECT 37.755 136.005 38.045 136.050 ;
        RECT 38.200 135.990 38.520 136.050 ;
        RECT 43.260 135.990 43.580 136.250 ;
        RECT 46.940 136.190 47.260 136.250 ;
        RECT 47.415 136.190 47.705 136.235 ;
        RECT 46.940 136.050 47.705 136.190 ;
        RECT 46.940 135.990 47.260 136.050 ;
        RECT 47.415 136.005 47.705 136.050 ;
        RECT 49.240 135.990 49.560 136.250 ;
        RECT 52.000 136.190 52.320 136.250 ;
        RECT 52.935 136.190 53.225 136.235 ;
        RECT 52.000 136.050 53.225 136.190 ;
        RECT 52.000 135.990 52.320 136.050 ;
        RECT 52.935 136.005 53.225 136.050 ;
        RECT 55.235 136.190 55.525 136.235 ;
        RECT 55.680 136.190 56.000 136.250 ;
        RECT 55.235 136.050 56.000 136.190 ;
        RECT 55.235 136.005 55.525 136.050 ;
        RECT 55.680 135.990 56.000 136.050 ;
        RECT 57.995 136.190 58.285 136.235 ;
        RECT 62.120 136.190 62.440 136.250 ;
        RECT 57.995 136.050 62.440 136.190 ;
        RECT 57.995 136.005 58.285 136.050 ;
        RECT 62.120 135.990 62.440 136.050 ;
        RECT 81.455 136.190 81.745 136.235 ;
        RECT 81.900 136.190 82.220 136.250 ;
        RECT 81.455 136.050 82.220 136.190 ;
        RECT 81.455 136.005 81.745 136.050 ;
        RECT 81.900 135.990 82.220 136.050 ;
        RECT 88.800 136.190 89.120 136.250 ;
        RECT 89.735 136.190 90.025 136.235 ;
        RECT 88.800 136.050 90.025 136.190 ;
        RECT 88.800 135.990 89.120 136.050 ;
        RECT 89.735 136.005 90.025 136.050 ;
        RECT 103.060 136.190 103.380 136.250 ;
        RECT 104.455 136.190 104.745 136.235 ;
        RECT 103.060 136.050 104.745 136.190 ;
        RECT 103.060 135.990 103.380 136.050 ;
        RECT 104.455 136.005 104.745 136.050 ;
        RECT 112.735 136.190 113.025 136.235 ;
        RECT 113.640 136.190 113.960 136.250 ;
        RECT 112.735 136.050 113.960 136.190 ;
        RECT 112.735 136.005 113.025 136.050 ;
        RECT 39.120 135.650 39.440 135.910 ;
        RECT 39.595 135.850 39.885 135.895 ;
        RECT 42.800 135.850 43.120 135.910 ;
        RECT 39.595 135.710 43.120 135.850 ;
        RECT 39.595 135.665 39.885 135.710 ;
        RECT 42.800 135.650 43.120 135.710 ;
        RECT 46.495 135.850 46.785 135.895 ;
        RECT 98.040 135.850 98.330 135.895 ;
        RECT 100.140 135.850 100.430 135.895 ;
        RECT 101.710 135.850 102.000 135.895 ;
        RECT 46.495 135.710 54.070 135.850 ;
        RECT 46.495 135.665 46.785 135.710 ;
        RECT 50.050 135.510 50.340 135.555 ;
        RECT 53.380 135.510 53.700 135.570 ;
        RECT 40.130 135.370 42.570 135.510 ;
        RECT 40.130 135.230 40.270 135.370 ;
        RECT 36.820 135.170 37.140 135.230 ;
        RECT 38.675 135.170 38.965 135.215 ;
        RECT 36.820 135.030 38.965 135.170 ;
        RECT 36.820 134.970 37.140 135.030 ;
        RECT 38.675 134.985 38.965 135.030 ;
        RECT 40.040 134.970 40.360 135.230 ;
        RECT 40.500 135.170 40.820 135.230 ;
        RECT 42.430 135.215 42.570 135.370 ;
        RECT 50.050 135.370 53.700 135.510 ;
        RECT 50.050 135.325 50.340 135.370 ;
        RECT 53.380 135.310 53.700 135.370 ;
        RECT 40.975 135.170 41.265 135.215 ;
        RECT 41.435 135.170 41.725 135.215 ;
        RECT 40.500 135.030 41.725 135.170 ;
        RECT 40.500 134.970 40.820 135.030 ;
        RECT 40.975 134.985 41.265 135.030 ;
        RECT 41.435 134.985 41.725 135.030 ;
        RECT 42.355 134.985 42.645 135.215 ;
        RECT 46.020 135.170 46.340 135.230 ;
        RECT 47.415 135.170 47.705 135.215 ;
        RECT 46.020 135.030 47.705 135.170 ;
        RECT 46.020 134.970 46.340 135.030 ;
        RECT 47.415 134.985 47.705 135.030 ;
        RECT 47.875 134.985 48.165 135.215 ;
        RECT 49.240 135.170 49.560 135.230 ;
        RECT 50.635 135.170 50.925 135.215 ;
        RECT 49.240 135.030 50.925 135.170 ;
        RECT 24.415 134.830 24.705 134.875 ;
        RECT 25.320 134.830 25.640 134.890 ;
        RECT 24.415 134.690 25.640 134.830 ;
        RECT 24.415 134.645 24.705 134.690 ;
        RECT 25.320 134.630 25.640 134.690 ;
        RECT 23.415 134.490 23.705 134.535 ;
        RECT 28.540 134.490 28.860 134.550 ;
        RECT 23.415 134.350 28.860 134.490 ;
        RECT 47.950 134.490 48.090 134.985 ;
        RECT 49.240 134.970 49.560 135.030 ;
        RECT 50.635 134.985 50.925 135.030 ;
        RECT 51.080 134.970 51.400 135.230 ;
        RECT 52.460 135.170 52.780 135.230 ;
        RECT 53.930 135.215 54.070 135.710 ;
        RECT 98.040 135.710 102.000 135.850 ;
        RECT 98.040 135.665 98.330 135.710 ;
        RECT 100.140 135.665 100.430 135.710 ;
        RECT 101.710 135.665 102.000 135.710 ;
        RECT 57.520 135.510 57.840 135.570 ;
        RECT 55.770 135.370 57.840 135.510 ;
        RECT 55.770 135.215 55.910 135.370 ;
        RECT 57.520 135.310 57.840 135.370 ;
        RECT 78.680 135.510 79.000 135.570 ;
        RECT 86.515 135.510 86.805 135.555 ;
        RECT 78.680 135.370 86.805 135.510 ;
        RECT 78.680 135.310 79.000 135.370 ;
        RECT 86.515 135.325 86.805 135.370 ;
        RECT 51.630 135.030 52.780 135.170 ;
        RECT 48.795 134.830 49.085 134.875 ;
        RECT 51.630 134.830 51.770 135.030 ;
        RECT 52.460 134.970 52.780 135.030 ;
        RECT 53.855 134.985 54.145 135.215 ;
        RECT 54.315 134.985 54.605 135.215 ;
        RECT 55.695 134.985 55.985 135.215 ;
        RECT 56.615 135.170 56.905 135.215 ;
        RECT 59.360 135.170 59.680 135.230 ;
        RECT 56.615 135.030 59.680 135.170 ;
        RECT 56.615 134.985 56.905 135.030 ;
        RECT 48.795 134.690 51.770 134.830 ;
        RECT 52.920 134.830 53.240 134.890 ;
        RECT 54.390 134.830 54.530 134.985 ;
        RECT 59.360 134.970 59.680 135.030 ;
        RECT 73.175 134.985 73.465 135.215 ;
        RECT 52.920 134.690 54.530 134.830 ;
        RECT 55.220 134.830 55.540 134.890 ;
        RECT 57.995 134.830 58.285 134.875 ;
        RECT 59.820 134.830 60.140 134.890 ;
        RECT 55.220 134.690 60.140 134.830 ;
        RECT 73.250 134.830 73.390 134.985 ;
        RECT 74.080 134.970 74.400 135.230 ;
        RECT 79.600 134.970 79.920 135.230 ;
        RECT 86.590 135.170 86.730 135.325 ;
        RECT 92.940 135.310 93.260 135.570 ;
        RECT 96.620 135.510 96.940 135.570 ;
        RECT 97.555 135.510 97.845 135.555 ;
        RECT 96.620 135.370 97.845 135.510 ;
        RECT 96.620 135.310 96.940 135.370 ;
        RECT 97.555 135.325 97.845 135.370 ;
        RECT 98.435 135.510 98.725 135.555 ;
        RECT 99.625 135.510 99.915 135.555 ;
        RECT 102.145 135.510 102.435 135.555 ;
        RECT 98.435 135.370 102.435 135.510 ;
        RECT 104.530 135.510 104.670 136.005 ;
        RECT 113.640 135.990 113.960 136.050 ;
        RECT 115.940 135.990 116.260 136.250 ;
        RECT 117.320 136.190 117.640 136.250 ;
        RECT 119.620 136.190 119.940 136.250 ;
        RECT 117.320 136.050 119.940 136.190 ;
        RECT 117.320 135.990 117.640 136.050 ;
        RECT 119.620 135.990 119.940 136.050 ;
        RECT 121.460 136.190 121.780 136.250 ;
        RECT 121.460 136.050 122.380 136.190 ;
        RECT 121.460 135.990 121.780 136.050 ;
        RECT 111.340 135.850 111.660 135.910 ;
        RECT 116.030 135.850 116.170 135.990 ;
        RECT 111.340 135.710 116.170 135.850 ;
        RECT 116.900 135.850 117.190 135.895 ;
        RECT 119.000 135.850 119.290 135.895 ;
        RECT 120.570 135.850 120.860 135.895 ;
        RECT 116.900 135.710 120.860 135.850 ;
        RECT 111.340 135.650 111.660 135.710 ;
        RECT 116.900 135.665 117.190 135.710 ;
        RECT 119.000 135.665 119.290 135.710 ;
        RECT 120.570 135.665 120.860 135.710 ;
        RECT 110.895 135.510 111.185 135.555 ;
        RECT 104.530 135.370 111.185 135.510 ;
        RECT 98.435 135.325 98.725 135.370 ;
        RECT 99.625 135.325 99.915 135.370 ;
        RECT 102.145 135.325 102.435 135.370 ;
        RECT 110.895 135.325 111.185 135.370 ;
        RECT 116.400 135.310 116.720 135.570 ;
        RECT 117.295 135.510 117.585 135.555 ;
        RECT 118.485 135.510 118.775 135.555 ;
        RECT 121.005 135.510 121.295 135.555 ;
        RECT 117.295 135.370 121.295 135.510 ;
        RECT 117.295 135.325 117.585 135.370 ;
        RECT 118.485 135.325 118.775 135.370 ;
        RECT 121.005 135.325 121.295 135.370 ;
        RECT 103.060 135.170 103.380 135.230 ;
        RECT 86.590 135.030 103.380 135.170 ;
        RECT 103.060 134.970 103.380 135.030 ;
        RECT 113.180 135.170 113.500 135.230 ;
        RECT 114.115 135.170 114.405 135.215 ;
        RECT 113.180 135.030 114.405 135.170 ;
        RECT 113.180 134.970 113.500 135.030 ;
        RECT 114.115 134.985 114.405 135.030 ;
        RECT 114.560 134.970 114.880 135.230 ;
        RECT 115.035 134.985 115.325 135.215 ;
        RECT 115.955 135.170 116.245 135.215 ;
        RECT 119.620 135.170 119.940 135.230 ;
        RECT 115.955 135.030 119.940 135.170 ;
        RECT 122.240 135.170 122.380 136.050 ;
        RECT 127.900 135.850 128.220 135.910 ;
        RECT 132.500 135.850 132.820 135.910 ;
        RECT 127.900 135.710 132.820 135.850 ;
        RECT 127.900 135.650 128.220 135.710 ;
        RECT 132.500 135.650 132.820 135.710 ;
        RECT 134.380 135.850 134.670 135.895 ;
        RECT 136.480 135.850 136.770 135.895 ;
        RECT 138.050 135.850 138.340 135.895 ;
        RECT 134.380 135.710 138.340 135.850 ;
        RECT 134.380 135.665 134.670 135.710 ;
        RECT 136.480 135.665 136.770 135.710 ;
        RECT 138.050 135.665 138.340 135.710 ;
        RECT 129.295 135.510 129.585 135.555 ;
        RECT 134.775 135.510 135.065 135.555 ;
        RECT 135.965 135.510 136.255 135.555 ;
        RECT 138.485 135.510 138.775 135.555 ;
        RECT 129.295 135.370 130.890 135.510 ;
        RECT 129.295 135.325 129.585 135.370 ;
        RECT 128.820 135.170 129.140 135.230 ;
        RECT 130.750 135.215 130.890 135.370 ;
        RECT 134.775 135.370 138.775 135.510 ;
        RECT 134.775 135.325 135.065 135.370 ;
        RECT 135.965 135.325 136.255 135.370 ;
        RECT 138.485 135.325 138.775 135.370 ;
        RECT 129.755 135.170 130.045 135.215 ;
        RECT 122.240 135.030 130.045 135.170 ;
        RECT 115.955 134.985 116.245 135.030 ;
        RECT 76.840 134.830 77.160 134.890 ;
        RECT 73.250 134.690 77.160 134.830 ;
        RECT 48.795 134.645 49.085 134.690 ;
        RECT 52.920 134.630 53.240 134.690 ;
        RECT 55.220 134.630 55.540 134.690 ;
        RECT 57.995 134.645 58.285 134.690 ;
        RECT 59.820 134.630 60.140 134.690 ;
        RECT 76.840 134.630 77.160 134.690 ;
        RECT 79.155 134.830 79.445 134.875 ;
        RECT 83.280 134.830 83.600 134.890 ;
        RECT 79.155 134.690 83.600 134.830 ;
        RECT 79.155 134.645 79.445 134.690 ;
        RECT 83.280 134.630 83.600 134.690 ;
        RECT 87.435 134.830 87.725 134.875 ;
        RECT 88.340 134.830 88.660 134.890 ;
        RECT 87.435 134.690 88.660 134.830 ;
        RECT 87.435 134.645 87.725 134.690 ;
        RECT 88.340 134.630 88.660 134.690 ;
        RECT 98.890 134.830 99.180 134.875 ;
        RECT 101.220 134.830 101.540 134.890 ;
        RECT 98.890 134.690 101.540 134.830 ;
        RECT 98.890 134.645 99.180 134.690 ;
        RECT 101.220 134.630 101.540 134.690 ;
        RECT 52.000 134.490 52.320 134.550 ;
        RECT 54.300 134.490 54.620 134.550 ;
        RECT 57.075 134.490 57.365 134.535 ;
        RECT 58.440 134.490 58.760 134.550 ;
        RECT 47.950 134.350 58.760 134.490 ;
        RECT 23.415 134.305 23.705 134.350 ;
        RECT 28.540 134.290 28.860 134.350 ;
        RECT 52.000 134.290 52.320 134.350 ;
        RECT 54.300 134.290 54.620 134.350 ;
        RECT 57.075 134.305 57.365 134.350 ;
        RECT 58.440 134.290 58.760 134.350 ;
        RECT 72.240 134.290 72.560 134.550 ;
        RECT 87.895 134.490 88.185 134.535 ;
        RECT 90.195 134.490 90.485 134.535 ;
        RECT 87.895 134.350 90.485 134.490 ;
        RECT 87.895 134.305 88.185 134.350 ;
        RECT 90.195 134.305 90.485 134.350 ;
        RECT 108.120 134.290 108.440 134.550 ;
        RECT 115.110 134.490 115.250 134.985 ;
        RECT 119.620 134.970 119.940 135.030 ;
        RECT 128.820 134.970 129.140 135.030 ;
        RECT 129.755 134.985 130.045 135.030 ;
        RECT 130.675 134.985 130.965 135.215 ;
        RECT 131.135 134.985 131.425 135.215 ;
        RECT 117.780 134.875 118.100 134.890 ;
        RECT 117.750 134.645 118.100 134.875 ;
        RECT 117.780 134.630 118.100 134.645 ;
        RECT 121.000 134.830 121.320 134.890 ;
        RECT 123.775 134.830 124.065 134.875 ;
        RECT 121.000 134.690 124.065 134.830 ;
        RECT 121.000 134.630 121.320 134.690 ;
        RECT 123.775 134.645 124.065 134.690 ;
        RECT 124.695 134.830 124.985 134.875 ;
        RECT 126.520 134.830 126.840 134.890 ;
        RECT 124.695 134.690 126.840 134.830 ;
        RECT 124.695 134.645 124.985 134.690 ;
        RECT 118.240 134.490 118.560 134.550 ;
        RECT 115.110 134.350 118.560 134.490 ;
        RECT 118.240 134.290 118.560 134.350 ;
        RECT 122.380 134.490 122.700 134.550 ;
        RECT 123.315 134.490 123.605 134.535 ;
        RECT 124.770 134.490 124.910 134.645 ;
        RECT 126.520 134.630 126.840 134.690 ;
        RECT 127.455 134.830 127.745 134.875 ;
        RECT 127.900 134.830 128.220 134.890 ;
        RECT 127.455 134.690 128.220 134.830 ;
        RECT 127.455 134.645 127.745 134.690 ;
        RECT 127.900 134.630 128.220 134.690 ;
        RECT 128.375 134.645 128.665 134.875 ;
        RECT 130.200 134.830 130.520 134.890 ;
        RECT 131.210 134.830 131.350 134.985 ;
        RECT 131.580 134.970 131.900 135.230 ;
        RECT 132.040 135.170 132.360 135.230 ;
        RECT 133.880 135.170 134.200 135.230 ;
        RECT 132.040 135.030 134.200 135.170 ;
        RECT 132.040 134.970 132.360 135.030 ;
        RECT 133.880 134.970 134.200 135.030 ;
        RECT 130.200 134.690 131.350 134.830 ;
        RECT 131.670 134.830 131.810 134.970 ;
        RECT 132.500 134.830 132.820 134.890 ;
        RECT 131.670 134.690 132.820 134.830 ;
        RECT 122.380 134.350 124.910 134.490 ;
        RECT 122.380 134.290 122.700 134.350 ;
        RECT 123.315 134.305 123.605 134.350 ;
        RECT 125.600 134.290 125.920 134.550 ;
        RECT 128.450 134.490 128.590 134.645 ;
        RECT 130.200 134.630 130.520 134.690 ;
        RECT 132.500 134.630 132.820 134.690 ;
        RECT 132.975 134.830 133.265 134.875 ;
        RECT 135.120 134.830 135.410 134.875 ;
        RECT 132.975 134.690 135.410 134.830 ;
        RECT 132.975 134.645 133.265 134.690 ;
        RECT 135.120 134.645 135.410 134.690 ;
        RECT 131.580 134.490 131.900 134.550 ;
        RECT 139.860 134.490 140.180 134.550 ;
        RECT 140.795 134.490 141.085 134.535 ;
        RECT 128.450 134.350 141.085 134.490 ;
        RECT 131.580 134.290 131.900 134.350 ;
        RECT 139.860 134.290 140.180 134.350 ;
        RECT 140.795 134.305 141.085 134.350 ;
        RECT 17.430 133.670 143.010 134.150 ;
        RECT 37.295 133.470 37.585 133.515 ;
        RECT 42.800 133.470 43.120 133.530 ;
        RECT 37.295 133.330 43.120 133.470 ;
        RECT 37.295 133.285 37.585 133.330 ;
        RECT 42.800 133.270 43.120 133.330 ;
        RECT 51.080 133.470 51.400 133.530 ;
        RECT 52.015 133.470 52.305 133.515 ;
        RECT 51.080 133.330 52.305 133.470 ;
        RECT 51.080 133.270 51.400 133.330 ;
        RECT 52.015 133.285 52.305 133.330 ;
        RECT 52.460 133.270 52.780 133.530 ;
        RECT 53.840 133.470 54.160 133.530 ;
        RECT 55.220 133.470 55.540 133.530 ;
        RECT 53.470 133.330 55.540 133.470 ;
        RECT 39.595 133.130 39.885 133.175 ;
        RECT 40.960 133.130 41.280 133.190 ;
        RECT 39.595 132.990 41.280 133.130 ;
        RECT 39.595 132.945 39.885 132.990 ;
        RECT 40.960 132.930 41.280 132.990 ;
        RECT 50.175 133.130 50.465 133.175 ;
        RECT 50.620 133.130 50.940 133.190 ;
        RECT 53.470 133.175 53.610 133.330 ;
        RECT 53.840 133.270 54.160 133.330 ;
        RECT 55.220 133.270 55.540 133.330 ;
        RECT 57.535 133.285 57.825 133.515 ;
        RECT 50.175 132.990 50.940 133.130 ;
        RECT 50.175 132.945 50.465 132.990 ;
        RECT 50.620 132.930 50.940 132.990 ;
        RECT 53.395 132.945 53.685 133.175 ;
        RECT 54.760 133.130 55.080 133.190 ;
        RECT 56.600 133.175 56.920 133.190 ;
        RECT 55.695 133.130 55.985 133.175 ;
        RECT 54.760 132.990 55.985 133.130 ;
        RECT 54.760 132.930 55.080 132.990 ;
        RECT 55.695 132.945 55.985 132.990 ;
        RECT 56.600 132.945 56.985 133.175 ;
        RECT 57.610 133.130 57.750 133.285 ;
        RECT 101.220 133.270 101.540 133.530 ;
        RECT 103.075 133.470 103.365 133.515 ;
        RECT 108.120 133.470 108.440 133.530 ;
        RECT 103.075 133.330 108.440 133.470 ;
        RECT 103.075 133.285 103.365 133.330 ;
        RECT 108.120 133.270 108.440 133.330 ;
        RECT 109.500 133.270 109.820 133.530 ;
        RECT 117.780 133.270 118.100 133.530 ;
        RECT 118.240 133.270 118.560 133.530 ;
        RECT 132.500 133.470 132.820 133.530 ;
        RECT 128.910 133.330 132.820 133.470 ;
        RECT 63.560 133.130 63.850 133.175 ;
        RECT 125.600 133.130 125.920 133.190 ;
        RECT 57.610 132.990 63.850 133.130 ;
        RECT 63.560 132.945 63.850 132.990 ;
        RECT 111.890 132.990 115.250 133.130 ;
        RECT 56.600 132.930 56.920 132.945 ;
        RECT 26.240 132.590 26.560 132.850 ;
        RECT 27.175 132.790 27.465 132.835 ;
        RECT 34.980 132.790 35.300 132.850 ;
        RECT 27.175 132.650 35.300 132.790 ;
        RECT 27.175 132.605 27.465 132.650 ;
        RECT 34.980 132.590 35.300 132.650 ;
        RECT 38.675 132.605 38.965 132.835 ;
        RECT 35.900 132.450 36.220 132.510 ;
        RECT 37.295 132.450 37.585 132.495 ;
        RECT 35.900 132.310 37.585 132.450 ;
        RECT 38.750 132.450 38.890 132.605 ;
        RECT 39.120 132.590 39.440 132.850 ;
        RECT 40.500 132.590 40.820 132.850 ;
        RECT 51.095 132.790 51.385 132.835 ;
        RECT 52.000 132.790 52.320 132.850 ;
        RECT 51.095 132.650 52.320 132.790 ;
        RECT 51.095 132.605 51.385 132.650 ;
        RECT 52.000 132.590 52.320 132.650 ;
        RECT 54.300 132.590 54.620 132.850 ;
        RECT 71.750 132.790 72.040 132.835 ;
        RECT 76.380 132.790 76.700 132.850 ;
        RECT 71.750 132.650 76.700 132.790 ;
        RECT 71.750 132.605 72.040 132.650 ;
        RECT 76.380 132.590 76.700 132.650 ;
        RECT 103.535 132.790 103.825 132.835 ;
        RECT 109.960 132.790 110.280 132.850 ;
        RECT 103.535 132.650 110.280 132.790 ;
        RECT 103.535 132.605 103.825 132.650 ;
        RECT 109.960 132.590 110.280 132.650 ;
        RECT 110.420 132.590 110.740 132.850 ;
        RECT 110.895 132.790 111.185 132.835 ;
        RECT 111.340 132.790 111.660 132.850 ;
        RECT 111.890 132.835 112.030 132.990 ;
        RECT 110.895 132.650 111.660 132.790 ;
        RECT 110.895 132.605 111.185 132.650 ;
        RECT 111.340 132.590 111.660 132.650 ;
        RECT 111.815 132.605 112.105 132.835 ;
        RECT 112.275 132.605 112.565 132.835 ;
        RECT 114.100 132.790 114.420 132.850 ;
        RECT 114.575 132.790 114.865 132.835 ;
        RECT 114.100 132.650 114.865 132.790 ;
        RECT 46.020 132.450 46.340 132.510 ;
        RECT 38.750 132.310 46.340 132.450 ;
        RECT 35.900 132.250 36.220 132.310 ;
        RECT 37.295 132.265 37.585 132.310 ;
        RECT 46.020 132.250 46.340 132.310 ;
        RECT 60.305 132.450 60.595 132.495 ;
        RECT 62.825 132.450 63.115 132.495 ;
        RECT 64.015 132.450 64.305 132.495 ;
        RECT 60.305 132.310 64.305 132.450 ;
        RECT 60.305 132.265 60.595 132.310 ;
        RECT 62.825 132.265 63.115 132.310 ;
        RECT 64.015 132.265 64.305 132.310 ;
        RECT 64.895 132.450 65.185 132.495 ;
        RECT 66.720 132.450 67.040 132.510 ;
        RECT 70.415 132.450 70.705 132.495 ;
        RECT 64.895 132.310 70.705 132.450 ;
        RECT 64.895 132.265 65.185 132.310 ;
        RECT 66.720 132.250 67.040 132.310 ;
        RECT 70.415 132.265 70.705 132.310 ;
        RECT 71.295 132.450 71.585 132.495 ;
        RECT 72.485 132.450 72.775 132.495 ;
        RECT 75.005 132.450 75.295 132.495 ;
        RECT 71.295 132.310 75.295 132.450 ;
        RECT 71.295 132.265 71.585 132.310 ;
        RECT 72.485 132.265 72.775 132.310 ;
        RECT 75.005 132.265 75.295 132.310 ;
        RECT 103.060 132.450 103.380 132.510 ;
        RECT 103.995 132.450 104.285 132.495 ;
        RECT 107.200 132.450 107.520 132.510 ;
        RECT 103.060 132.310 107.520 132.450 ;
        RECT 103.060 132.250 103.380 132.310 ;
        RECT 103.995 132.265 104.285 132.310 ;
        RECT 107.200 132.250 107.520 132.310 ;
        RECT 109.500 132.450 109.820 132.510 ;
        RECT 112.350 132.450 112.490 132.605 ;
        RECT 114.100 132.590 114.420 132.650 ;
        RECT 114.575 132.605 114.865 132.650 ;
        RECT 109.500 132.310 112.490 132.450 ;
        RECT 109.500 132.250 109.820 132.310 ;
        RECT 39.580 132.110 39.900 132.170 ;
        RECT 40.515 132.110 40.805 132.155 ;
        RECT 39.580 131.970 40.805 132.110 ;
        RECT 39.580 131.910 39.900 131.970 ;
        RECT 40.515 131.925 40.805 131.970 ;
        RECT 60.740 132.110 61.030 132.155 ;
        RECT 62.310 132.110 62.600 132.155 ;
        RECT 64.410 132.110 64.700 132.155 ;
        RECT 60.740 131.970 64.700 132.110 ;
        RECT 60.740 131.925 61.030 131.970 ;
        RECT 62.310 131.925 62.600 131.970 ;
        RECT 64.410 131.925 64.700 131.970 ;
        RECT 70.900 132.110 71.190 132.155 ;
        RECT 73.000 132.110 73.290 132.155 ;
        RECT 74.570 132.110 74.860 132.155 ;
        RECT 70.900 131.970 74.860 132.110 ;
        RECT 115.110 132.110 115.250 132.990 ;
        RECT 115.570 132.990 125.920 133.130 ;
        RECT 115.570 132.835 115.710 132.990 ;
        RECT 125.600 132.930 125.920 132.990 ;
        RECT 115.495 132.605 115.785 132.835 ;
        RECT 115.940 132.590 116.260 132.850 ;
        RECT 116.415 132.790 116.705 132.835 ;
        RECT 117.780 132.790 118.100 132.850 ;
        RECT 116.415 132.650 118.100 132.790 ;
        RECT 116.415 132.605 116.705 132.650 ;
        RECT 117.780 132.590 118.100 132.650 ;
        RECT 119.160 132.590 119.480 132.850 ;
        RECT 120.080 132.590 120.400 132.850 ;
        RECT 128.910 132.790 129.050 133.330 ;
        RECT 132.500 133.270 132.820 133.330 ;
        RECT 140.780 133.270 141.100 133.530 ;
        RECT 129.280 133.130 129.600 133.190 ;
        RECT 130.675 133.130 130.965 133.175 ;
        RECT 129.280 132.990 130.965 133.130 ;
        RECT 129.280 132.930 129.600 132.990 ;
        RECT 130.675 132.945 130.965 132.990 ;
        RECT 120.630 132.650 129.050 132.790 ;
        RECT 117.870 132.450 118.010 132.590 ;
        RECT 120.630 132.450 120.770 132.650 ;
        RECT 129.740 132.590 130.060 132.850 ;
        RECT 130.200 132.590 130.520 132.850 ;
        RECT 131.580 132.590 131.900 132.850 ;
        RECT 132.040 132.590 132.360 132.850 ;
        RECT 133.390 132.790 133.680 132.835 ;
        RECT 137.100 132.790 137.420 132.850 ;
        RECT 133.390 132.650 137.420 132.790 ;
        RECT 133.390 132.605 133.680 132.650 ;
        RECT 137.100 132.590 137.420 132.650 ;
        RECT 139.860 132.835 140.180 132.850 ;
        RECT 139.860 132.790 140.195 132.835 ;
        RECT 139.860 132.650 140.375 132.790 ;
        RECT 139.860 132.605 140.195 132.650 ;
        RECT 139.860 132.590 140.180 132.605 ;
        RECT 117.870 132.310 120.770 132.450 ;
        RECT 121.920 132.450 122.240 132.510 ;
        RECT 130.660 132.450 130.980 132.510 ;
        RECT 121.920 132.310 130.980 132.450 ;
        RECT 121.920 132.250 122.240 132.310 ;
        RECT 130.660 132.250 130.980 132.310 ;
        RECT 132.935 132.450 133.225 132.495 ;
        RECT 134.125 132.450 134.415 132.495 ;
        RECT 136.645 132.450 136.935 132.495 ;
        RECT 132.935 132.310 136.935 132.450 ;
        RECT 132.935 132.265 133.225 132.310 ;
        RECT 134.125 132.265 134.415 132.310 ;
        RECT 136.645 132.265 136.935 132.310 ;
        RECT 132.540 132.110 132.830 132.155 ;
        RECT 134.640 132.110 134.930 132.155 ;
        RECT 136.210 132.110 136.500 132.155 ;
        RECT 115.110 131.970 129.970 132.110 ;
        RECT 70.900 131.925 71.190 131.970 ;
        RECT 73.000 131.925 73.290 131.970 ;
        RECT 74.570 131.925 74.860 131.970 ;
        RECT 27.175 131.770 27.465 131.815 ;
        RECT 29.000 131.770 29.320 131.830 ;
        RECT 27.175 131.630 29.320 131.770 ;
        RECT 27.175 131.585 27.465 131.630 ;
        RECT 29.000 131.570 29.320 131.630 ;
        RECT 35.440 131.770 35.760 131.830 ;
        RECT 38.215 131.770 38.505 131.815 ;
        RECT 35.440 131.630 38.505 131.770 ;
        RECT 35.440 131.570 35.760 131.630 ;
        RECT 38.215 131.585 38.505 131.630 ;
        RECT 48.320 131.770 48.640 131.830 ;
        RECT 56.615 131.770 56.905 131.815 ;
        RECT 48.320 131.630 56.905 131.770 ;
        RECT 48.320 131.570 48.640 131.630 ;
        RECT 56.615 131.585 56.905 131.630 ;
        RECT 57.995 131.770 58.285 131.815 ;
        RECT 58.440 131.770 58.760 131.830 ;
        RECT 57.995 131.630 58.760 131.770 ;
        RECT 57.995 131.585 58.285 131.630 ;
        RECT 58.440 131.570 58.760 131.630 ;
        RECT 77.315 131.770 77.605 131.815 ;
        RECT 78.220 131.770 78.540 131.830 ;
        RECT 77.315 131.630 78.540 131.770 ;
        RECT 77.315 131.585 77.605 131.630 ;
        RECT 78.220 131.570 78.540 131.630 ;
        RECT 115.480 131.770 115.800 131.830 ;
        RECT 128.835 131.770 129.125 131.815 ;
        RECT 115.480 131.630 129.125 131.770 ;
        RECT 129.830 131.770 129.970 131.970 ;
        RECT 132.540 131.970 136.500 132.110 ;
        RECT 132.540 131.925 132.830 131.970 ;
        RECT 134.640 131.925 134.930 131.970 ;
        RECT 136.210 131.925 136.500 131.970 ;
        RECT 137.560 131.770 137.880 131.830 ;
        RECT 129.830 131.630 137.880 131.770 ;
        RECT 115.480 131.570 115.800 131.630 ;
        RECT 128.835 131.585 129.125 131.630 ;
        RECT 137.560 131.570 137.880 131.630 ;
        RECT 138.940 131.570 139.260 131.830 ;
        RECT 17.430 130.950 143.010 131.430 ;
        RECT 24.860 130.750 25.180 130.810 ;
        RECT 29.015 130.750 29.305 130.795 ;
        RECT 37.755 130.750 38.045 130.795 ;
        RECT 40.040 130.750 40.360 130.810 ;
        RECT 24.860 130.610 37.510 130.750 ;
        RECT 24.860 130.550 25.180 130.610 ;
        RECT 29.015 130.565 29.305 130.610 ;
        RECT 29.920 130.410 30.240 130.470 ;
        RECT 37.370 130.410 37.510 130.610 ;
        RECT 37.755 130.610 40.360 130.750 ;
        RECT 37.755 130.565 38.045 130.610 ;
        RECT 40.040 130.550 40.360 130.610 ;
        RECT 56.600 130.550 56.920 130.810 ;
        RECT 109.960 130.750 110.280 130.810 ;
        RECT 111.355 130.750 111.645 130.795 ;
        RECT 109.960 130.610 111.645 130.750 ;
        RECT 109.960 130.550 110.280 130.610 ;
        RECT 111.355 130.565 111.645 130.610 ;
        RECT 112.720 130.750 113.040 130.810 ;
        RECT 114.575 130.750 114.865 130.795 ;
        RECT 129.740 130.750 130.060 130.810 ;
        RECT 135.720 130.750 136.040 130.810 ;
        RECT 112.720 130.610 114.865 130.750 ;
        RECT 112.720 130.550 113.040 130.610 ;
        RECT 114.575 130.565 114.865 130.610 ;
        RECT 122.930 130.610 136.040 130.750 ;
        RECT 69.060 130.410 69.350 130.455 ;
        RECT 71.160 130.410 71.450 130.455 ;
        RECT 72.730 130.410 73.020 130.455 ;
        RECT 76.395 130.410 76.685 130.455 ;
        RECT 29.920 130.270 31.990 130.410 ;
        RECT 37.370 130.270 40.270 130.410 ;
        RECT 29.920 130.210 30.240 130.270 ;
        RECT 26.240 130.070 26.560 130.130 ;
        RECT 26.240 129.930 31.070 130.070 ;
        RECT 26.240 129.870 26.560 129.930 ;
        RECT 30.930 129.775 31.070 129.930 ;
        RECT 31.850 129.775 31.990 130.270 ;
        RECT 40.130 130.130 40.270 130.270 ;
        RECT 69.060 130.270 73.020 130.410 ;
        RECT 69.060 130.225 69.350 130.270 ;
        RECT 71.160 130.225 71.450 130.270 ;
        RECT 72.730 130.225 73.020 130.270 ;
        RECT 73.940 130.270 76.685 130.410 ;
        RECT 40.040 129.870 40.360 130.130 ;
        RECT 47.860 130.070 48.180 130.130 ;
        RECT 57.060 130.070 57.380 130.130 ;
        RECT 47.860 129.930 57.380 130.070 ;
        RECT 47.860 129.870 48.180 129.930 ;
        RECT 57.060 129.870 57.380 129.930 ;
        RECT 57.995 130.070 58.285 130.115 ;
        RECT 59.360 130.070 59.680 130.130 ;
        RECT 57.995 129.930 59.680 130.070 ;
        RECT 57.995 129.885 58.285 129.930 ;
        RECT 23.495 129.730 23.785 129.775 ;
        RECT 25.795 129.730 26.085 129.775 ;
        RECT 23.495 129.590 26.085 129.730 ;
        RECT 23.495 129.545 23.785 129.590 ;
        RECT 25.795 129.545 26.085 129.590 ;
        RECT 26.330 129.590 30.150 129.730 ;
        RECT 18.880 129.390 19.200 129.450 ;
        RECT 25.320 129.390 25.640 129.450 ;
        RECT 26.330 129.390 26.470 129.590 ;
        RECT 18.880 129.250 25.090 129.390 ;
        RECT 18.880 129.190 19.200 129.250 ;
        RECT 21.640 129.050 21.960 129.110 ;
        RECT 22.575 129.050 22.865 129.095 ;
        RECT 21.640 128.910 22.865 129.050 ;
        RECT 21.640 128.850 21.960 128.910 ;
        RECT 22.575 128.865 22.865 128.910 ;
        RECT 23.940 128.850 24.260 129.110 ;
        RECT 24.400 128.850 24.720 129.110 ;
        RECT 24.950 129.050 25.090 129.250 ;
        RECT 25.320 129.250 26.470 129.390 ;
        RECT 25.320 129.190 25.640 129.250 ;
        RECT 26.700 129.190 27.020 129.450 ;
        RECT 27.620 129.390 27.940 129.450 ;
        RECT 29.000 129.435 29.320 129.450 ;
        RECT 30.010 129.435 30.150 129.590 ;
        RECT 30.855 129.545 31.145 129.775 ;
        RECT 31.775 129.730 32.065 129.775 ;
        RECT 34.060 129.730 34.380 129.790 ;
        RECT 31.775 129.590 34.380 129.730 ;
        RECT 31.775 129.545 32.065 129.590 ;
        RECT 34.060 129.530 34.380 129.590 ;
        RECT 39.120 129.530 39.440 129.790 ;
        RECT 53.380 129.530 53.700 129.790 ;
        RECT 54.300 129.530 54.620 129.790 ;
        RECT 54.775 129.545 55.065 129.775 ;
        RECT 55.680 129.730 56.000 129.790 ;
        RECT 58.070 129.730 58.210 129.885 ;
        RECT 59.360 129.870 59.680 129.930 ;
        RECT 66.720 130.070 67.040 130.130 ;
        RECT 68.575 130.070 68.865 130.115 ;
        RECT 66.720 129.930 68.865 130.070 ;
        RECT 66.720 129.870 67.040 129.930 ;
        RECT 68.575 129.885 68.865 129.930 ;
        RECT 69.455 130.070 69.745 130.115 ;
        RECT 70.645 130.070 70.935 130.115 ;
        RECT 73.165 130.070 73.455 130.115 ;
        RECT 69.455 129.930 73.455 130.070 ;
        RECT 69.455 129.885 69.745 129.930 ;
        RECT 70.645 129.885 70.935 129.930 ;
        RECT 73.165 129.885 73.455 129.930 ;
        RECT 55.680 129.590 58.210 129.730 ;
        RECT 27.620 129.250 28.770 129.390 ;
        RECT 27.620 129.190 27.940 129.250 ;
        RECT 27.710 129.050 27.850 129.190 ;
        RECT 24.950 128.910 27.850 129.050 ;
        RECT 28.080 128.850 28.400 129.110 ;
        RECT 28.630 129.050 28.770 129.250 ;
        RECT 28.910 129.205 29.320 129.435 ;
        RECT 29.935 129.390 30.225 129.435 ;
        RECT 37.755 129.390 38.045 129.435 ;
        RECT 38.200 129.390 38.520 129.450 ;
        RECT 29.935 129.250 31.070 129.390 ;
        RECT 29.935 129.205 30.225 129.250 ;
        RECT 29.000 129.190 29.320 129.205 ;
        RECT 30.930 129.110 31.070 129.250 ;
        RECT 37.755 129.250 38.520 129.390 ;
        RECT 37.755 129.205 38.045 129.250 ;
        RECT 38.200 129.190 38.520 129.250 ;
        RECT 53.855 129.390 54.145 129.435 ;
        RECT 54.850 129.390 54.990 129.545 ;
        RECT 55.680 129.530 56.000 129.590 ;
        RECT 58.440 129.530 58.760 129.790 ;
        RECT 69.910 129.730 70.200 129.775 ;
        RECT 73.940 129.730 74.080 130.270 ;
        RECT 76.395 130.225 76.685 130.270 ;
        RECT 82.860 130.410 83.150 130.455 ;
        RECT 84.960 130.410 85.250 130.455 ;
        RECT 86.530 130.410 86.820 130.455 ;
        RECT 115.480 130.410 115.800 130.470 ;
        RECT 119.160 130.410 119.480 130.470 ;
        RECT 82.860 130.270 86.820 130.410 ;
        RECT 82.860 130.225 83.150 130.270 ;
        RECT 84.960 130.225 85.250 130.270 ;
        RECT 86.530 130.225 86.820 130.270 ;
        RECT 114.190 130.270 115.800 130.410 ;
        RECT 77.300 130.070 77.620 130.130 ;
        RECT 79.155 130.070 79.445 130.115 ;
        RECT 77.300 129.930 79.445 130.070 ;
        RECT 77.300 129.870 77.620 129.930 ;
        RECT 79.155 129.885 79.445 129.930 ;
        RECT 83.255 130.070 83.545 130.115 ;
        RECT 84.445 130.070 84.735 130.115 ;
        RECT 86.965 130.070 87.255 130.115 ;
        RECT 83.255 129.930 87.255 130.070 ;
        RECT 83.255 129.885 83.545 129.930 ;
        RECT 84.445 129.885 84.735 129.930 ;
        RECT 86.965 129.885 87.255 129.930 ;
        RECT 92.955 129.885 93.245 130.115 ;
        RECT 96.160 130.070 96.480 130.130 ;
        RECT 101.235 130.070 101.525 130.115 ;
        RECT 110.880 130.070 111.200 130.130 ;
        RECT 113.180 130.070 113.500 130.130 ;
        RECT 96.160 129.930 111.200 130.070 ;
        RECT 69.910 129.590 74.080 129.730 ;
        RECT 78.235 129.730 78.525 129.775 ;
        RECT 78.680 129.730 79.000 129.790 ;
        RECT 78.235 129.590 79.000 129.730 ;
        RECT 69.910 129.545 70.200 129.590 ;
        RECT 78.235 129.545 78.525 129.590 ;
        RECT 53.855 129.250 54.990 129.390 ;
        RECT 53.855 129.205 54.145 129.250 ;
        RECT 30.380 129.050 30.700 129.110 ;
        RECT 28.630 128.910 30.700 129.050 ;
        RECT 30.380 128.850 30.700 128.910 ;
        RECT 30.840 128.850 31.160 129.110 ;
        RECT 31.315 129.050 31.605 129.095 ;
        RECT 32.220 129.050 32.540 129.110 ;
        RECT 31.315 128.910 32.540 129.050 ;
        RECT 31.315 128.865 31.605 128.910 ;
        RECT 32.220 128.850 32.540 128.910 ;
        RECT 38.660 129.050 38.980 129.110 ;
        RECT 40.960 129.050 41.280 129.110 ;
        RECT 45.560 129.050 45.880 129.110 ;
        RECT 38.660 128.910 45.880 129.050 ;
        RECT 38.660 128.850 38.980 128.910 ;
        RECT 40.960 128.850 41.280 128.910 ;
        RECT 45.560 128.850 45.880 128.910 ;
        RECT 55.220 128.850 55.540 129.110 ;
        RECT 75.475 129.050 75.765 129.095 ;
        RECT 78.310 129.050 78.450 129.545 ;
        RECT 78.680 129.530 79.000 129.590 ;
        RECT 82.375 129.730 82.665 129.775 ;
        RECT 85.580 129.730 85.900 129.790 ;
        RECT 82.375 129.590 85.900 129.730 ;
        RECT 82.375 129.545 82.665 129.590 ;
        RECT 85.580 129.530 85.900 129.590 ;
        RECT 86.040 129.730 86.360 129.790 ;
        RECT 93.030 129.730 93.170 129.885 ;
        RECT 96.160 129.870 96.480 129.930 ;
        RECT 101.235 129.885 101.525 129.930 ;
        RECT 110.880 129.870 111.200 129.930 ;
        RECT 112.350 129.930 113.500 130.070 ;
        RECT 86.040 129.590 93.170 129.730 ;
        RECT 86.040 129.530 86.360 129.590 ;
        RECT 105.835 129.545 106.125 129.775 ;
        RECT 110.420 129.730 110.740 129.790 ;
        RECT 112.350 129.775 112.490 129.930 ;
        RECT 113.180 129.870 113.500 129.930 ;
        RECT 112.275 129.730 112.565 129.775 ;
        RECT 110.420 129.590 112.565 129.730 ;
        RECT 83.710 129.390 84.000 129.435 ;
        RECT 84.660 129.390 84.980 129.450 ;
        RECT 83.710 129.250 84.980 129.390 ;
        RECT 83.710 129.205 84.000 129.250 ;
        RECT 84.660 129.190 84.980 129.250 ;
        RECT 100.315 129.390 100.605 129.435 ;
        RECT 102.615 129.390 102.905 129.435 ;
        RECT 100.315 129.250 102.905 129.390 ;
        RECT 100.315 129.205 100.605 129.250 ;
        RECT 102.615 129.205 102.905 129.250 ;
        RECT 75.475 128.910 78.450 129.050 ;
        RECT 78.695 129.050 78.985 129.095 ;
        RECT 82.820 129.050 83.140 129.110 ;
        RECT 78.695 128.910 83.140 129.050 ;
        RECT 75.475 128.865 75.765 128.910 ;
        RECT 78.695 128.865 78.985 128.910 ;
        RECT 82.820 128.850 83.140 128.910 ;
        RECT 84.200 129.050 84.520 129.110 ;
        RECT 89.275 129.050 89.565 129.095 ;
        RECT 84.200 128.910 89.565 129.050 ;
        RECT 84.200 128.850 84.520 128.910 ;
        RECT 89.275 128.865 89.565 128.910 ;
        RECT 89.720 129.050 90.040 129.110 ;
        RECT 90.195 129.050 90.485 129.095 ;
        RECT 89.720 128.910 90.485 129.050 ;
        RECT 89.720 128.850 90.040 128.910 ;
        RECT 90.195 128.865 90.485 128.910 ;
        RECT 92.020 128.850 92.340 129.110 ;
        RECT 92.495 129.050 92.785 129.095 ;
        RECT 94.780 129.050 95.100 129.110 ;
        RECT 92.495 128.910 95.100 129.050 ;
        RECT 92.495 128.865 92.785 128.910 ;
        RECT 94.780 128.850 95.100 128.910 ;
        RECT 98.460 128.850 98.780 129.110 ;
        RECT 100.760 128.850 101.080 129.110 ;
        RECT 105.910 129.050 106.050 129.545 ;
        RECT 110.420 129.530 110.740 129.590 ;
        RECT 112.275 129.545 112.565 129.590 ;
        RECT 112.735 129.545 113.025 129.775 ;
        RECT 112.810 129.390 112.950 129.545 ;
        RECT 113.640 129.530 113.960 129.790 ;
        RECT 114.190 129.775 114.330 130.270 ;
        RECT 115.480 130.210 115.800 130.270 ;
        RECT 116.030 130.270 119.480 130.410 ;
        RECT 114.115 129.545 114.405 129.775 ;
        RECT 114.560 129.730 114.880 129.790 ;
        RECT 116.030 129.775 116.170 130.270 ;
        RECT 119.160 130.210 119.480 130.270 ;
        RECT 121.935 130.225 122.225 130.455 ;
        RECT 122.010 130.070 122.150 130.225 ;
        RECT 116.950 129.930 122.150 130.070 ;
        RECT 116.950 129.775 117.090 129.930 ;
        RECT 115.495 129.730 115.785 129.775 ;
        RECT 114.560 129.590 115.785 129.730 ;
        RECT 114.560 129.530 114.880 129.590 ;
        RECT 115.495 129.545 115.785 129.590 ;
        RECT 115.955 129.545 116.245 129.775 ;
        RECT 116.875 129.545 117.165 129.775 ;
        RECT 117.320 129.530 117.640 129.790 ;
        RECT 118.700 129.530 119.020 129.790 ;
        RECT 119.635 129.730 119.925 129.775 ;
        RECT 121.000 129.730 121.320 129.790 ;
        RECT 122.930 129.775 123.070 130.610 ;
        RECT 129.740 130.550 130.060 130.610 ;
        RECT 135.720 130.550 136.040 130.610 ;
        RECT 137.100 130.550 137.420 130.810 ;
        RECT 137.560 130.550 137.880 130.810 ;
        RECT 129.280 130.410 129.600 130.470 ;
        RECT 133.880 130.410 134.200 130.470 ;
        RECT 129.280 130.270 139.630 130.410 ;
        RECT 129.280 130.210 129.600 130.270 ;
        RECT 133.880 130.210 134.200 130.270 ;
        RECT 129.370 130.070 129.510 130.210 ;
        RECT 123.850 129.930 129.510 130.070 ;
        RECT 131.120 130.070 131.440 130.130 ;
        RECT 133.420 130.070 133.740 130.130 ;
        RECT 131.120 129.930 133.740 130.070 ;
        RECT 123.850 129.775 123.990 129.930 ;
        RECT 131.120 129.870 131.440 129.930 ;
        RECT 133.420 129.870 133.740 129.930 ;
        RECT 134.340 130.070 134.660 130.130 ;
        RECT 134.340 129.930 135.950 130.070 ;
        RECT 134.340 129.870 134.660 129.930 ;
        RECT 119.635 129.590 121.320 129.730 ;
        RECT 119.635 129.545 119.925 129.590 ;
        RECT 121.000 129.530 121.320 129.590 ;
        RECT 122.855 129.545 123.145 129.775 ;
        RECT 123.775 129.545 124.065 129.775 ;
        RECT 124.695 129.730 124.985 129.775 ;
        RECT 125.140 129.730 125.460 129.790 ;
        RECT 124.695 129.590 125.460 129.730 ;
        RECT 124.695 129.545 124.985 129.590 ;
        RECT 125.140 129.530 125.460 129.590 ;
        RECT 128.820 129.730 129.140 129.790 ;
        RECT 133.895 129.730 134.185 129.775 ;
        RECT 128.820 129.590 134.185 129.730 ;
        RECT 128.820 129.530 129.140 129.590 ;
        RECT 133.895 129.545 134.185 129.590 ;
        RECT 134.815 129.545 135.105 129.775 ;
        RECT 112.810 129.250 118.470 129.390 ;
        RECT 108.580 129.050 108.900 129.110 ;
        RECT 112.720 129.050 113.040 129.110 ;
        RECT 105.910 128.910 113.040 129.050 ;
        RECT 108.580 128.850 108.900 128.910 ;
        RECT 112.720 128.850 113.040 128.910 ;
        RECT 114.100 129.050 114.420 129.110 ;
        RECT 117.795 129.050 118.085 129.095 ;
        RECT 114.100 128.910 118.085 129.050 ;
        RECT 118.330 129.050 118.470 129.250 ;
        RECT 123.315 129.205 123.605 129.435 ;
        RECT 126.520 129.390 126.840 129.450 ;
        RECT 131.135 129.390 131.425 129.435 ;
        RECT 126.520 129.250 131.425 129.390 ;
        RECT 122.380 129.050 122.700 129.110 ;
        RECT 118.330 128.910 122.700 129.050 ;
        RECT 123.390 129.050 123.530 129.205 ;
        RECT 126.520 129.190 126.840 129.250 ;
        RECT 131.135 129.205 131.425 129.250 ;
        RECT 132.055 129.205 132.345 129.435 ;
        RECT 132.975 129.390 133.265 129.435 ;
        RECT 134.890 129.390 135.030 129.545 ;
        RECT 135.260 129.530 135.580 129.790 ;
        RECT 135.810 129.775 135.950 129.930 ;
        RECT 135.735 129.545 136.025 129.775 ;
        RECT 136.180 129.730 136.500 129.790 ;
        RECT 139.490 129.775 139.630 130.270 ;
        RECT 138.495 129.730 138.785 129.775 ;
        RECT 136.180 129.590 138.785 129.730 ;
        RECT 136.180 129.530 136.500 129.590 ;
        RECT 138.495 129.545 138.785 129.590 ;
        RECT 139.415 129.545 139.705 129.775 ;
        RECT 140.320 129.530 140.640 129.790 ;
        RECT 132.975 129.250 135.030 129.390 ;
        RECT 132.975 129.205 133.265 129.250 ;
        RECT 127.900 129.050 128.220 129.110 ;
        RECT 123.390 128.910 128.220 129.050 ;
        RECT 132.130 129.050 132.270 129.205 ;
        RECT 138.940 129.190 139.260 129.450 ;
        RECT 139.030 129.050 139.170 129.190 ;
        RECT 139.860 129.050 140.180 129.110 ;
        RECT 132.130 128.910 140.180 129.050 ;
        RECT 114.100 128.850 114.420 128.910 ;
        RECT 117.795 128.865 118.085 128.910 ;
        RECT 122.380 128.850 122.700 128.910 ;
        RECT 127.900 128.850 128.220 128.910 ;
        RECT 139.860 128.850 140.180 128.910 ;
        RECT 17.430 128.230 143.010 128.710 ;
        RECT 19.815 128.030 20.105 128.075 ;
        RECT 23.940 128.030 24.260 128.090 ;
        RECT 19.815 127.890 24.260 128.030 ;
        RECT 19.815 127.845 20.105 127.890 ;
        RECT 23.940 127.830 24.260 127.890 ;
        RECT 26.240 128.030 26.560 128.090 ;
        RECT 27.635 128.030 27.925 128.075 ;
        RECT 26.240 127.890 27.925 128.030 ;
        RECT 26.240 127.830 26.560 127.890 ;
        RECT 27.635 127.845 27.925 127.890 ;
        RECT 28.475 128.030 28.765 128.075 ;
        RECT 30.380 128.030 30.700 128.090 ;
        RECT 31.760 128.030 32.080 128.090 ;
        RECT 28.475 127.890 32.080 128.030 ;
        RECT 28.475 127.845 28.765 127.890 ;
        RECT 30.380 127.830 30.700 127.890 ;
        RECT 31.760 127.830 32.080 127.890 ;
        RECT 33.615 128.030 33.905 128.075 ;
        RECT 35.900 128.030 36.220 128.090 ;
        RECT 33.615 127.890 36.220 128.030 ;
        RECT 33.615 127.845 33.905 127.890 ;
        RECT 27.160 127.690 27.480 127.750 ;
        RECT 20.350 127.550 27.480 127.690 ;
        RECT 18.880 127.150 19.200 127.410 ;
        RECT 20.350 127.395 20.490 127.550 ;
        RECT 27.160 127.490 27.480 127.550 ;
        RECT 29.000 127.690 29.320 127.750 ;
        RECT 29.475 127.690 29.765 127.735 ;
        RECT 31.300 127.690 31.620 127.750 ;
        RECT 33.690 127.690 33.830 127.845 ;
        RECT 35.900 127.830 36.220 127.890 ;
        RECT 37.295 128.030 37.585 128.075 ;
        RECT 38.200 128.030 38.520 128.090 ;
        RECT 37.295 127.890 38.520 128.030 ;
        RECT 37.295 127.845 37.585 127.890 ;
        RECT 38.200 127.830 38.520 127.890 ;
        RECT 40.500 127.830 40.820 128.090 ;
        RECT 51.095 128.030 51.385 128.075 ;
        RECT 53.395 128.030 53.685 128.075 ;
        RECT 54.300 128.030 54.620 128.090 ;
        RECT 51.095 127.890 54.620 128.030 ;
        RECT 51.095 127.845 51.385 127.890 ;
        RECT 53.395 127.845 53.685 127.890 ;
        RECT 54.300 127.830 54.620 127.890 ;
        RECT 74.080 128.030 74.400 128.090 ;
        RECT 76.395 128.030 76.685 128.075 ;
        RECT 74.080 127.890 76.685 128.030 ;
        RECT 74.080 127.830 74.400 127.890 ;
        RECT 76.395 127.845 76.685 127.890 ;
        RECT 29.000 127.550 31.070 127.690 ;
        RECT 29.000 127.490 29.320 127.550 ;
        RECT 29.475 127.505 29.765 127.550 ;
        RECT 21.640 127.395 21.960 127.410 ;
        RECT 30.930 127.395 31.070 127.550 ;
        RECT 31.300 127.550 33.830 127.690 ;
        RECT 34.060 127.690 34.380 127.750 ;
        RECT 52.935 127.690 53.225 127.735 ;
        RECT 55.680 127.690 56.000 127.750 ;
        RECT 34.060 127.550 36.590 127.690 ;
        RECT 31.300 127.490 31.620 127.550 ;
        RECT 34.060 127.490 34.380 127.550 ;
        RECT 19.815 127.165 20.105 127.395 ;
        RECT 20.275 127.165 20.565 127.395 ;
        RECT 21.610 127.350 21.960 127.395 ;
        RECT 21.445 127.210 21.960 127.350 ;
        RECT 21.610 127.165 21.960 127.210 ;
        RECT 30.855 127.165 31.145 127.395 ;
        RECT 31.760 127.350 32.080 127.410 ;
        RECT 33.155 127.350 33.445 127.395 ;
        RECT 31.760 127.210 33.445 127.350 ;
        RECT 19.890 127.010 20.030 127.165 ;
        RECT 21.640 127.150 21.960 127.165 ;
        RECT 21.155 127.010 21.445 127.055 ;
        RECT 22.345 127.010 22.635 127.055 ;
        RECT 24.865 127.010 25.155 127.055 ;
        RECT 19.890 126.870 20.490 127.010 ;
        RECT 20.350 126.330 20.490 126.870 ;
        RECT 21.155 126.870 25.155 127.010 ;
        RECT 30.930 127.010 31.070 127.165 ;
        RECT 31.760 127.150 32.080 127.210 ;
        RECT 33.155 127.165 33.445 127.210 ;
        RECT 34.535 127.350 34.825 127.395 ;
        RECT 35.440 127.350 35.760 127.410 ;
        RECT 36.450 127.395 36.590 127.550 ;
        RECT 52.935 127.550 56.000 127.690 ;
        RECT 76.470 127.690 76.610 127.845 ;
        RECT 77.300 127.830 77.620 128.090 ;
        RECT 84.660 128.030 84.980 128.090 ;
        RECT 85.135 128.030 85.425 128.075 ;
        RECT 84.660 127.890 85.425 128.030 ;
        RECT 84.660 127.830 84.980 127.890 ;
        RECT 85.135 127.845 85.425 127.890 ;
        RECT 103.995 128.030 104.285 128.075 ;
        RECT 108.580 128.030 108.900 128.090 ;
        RECT 103.995 127.890 108.900 128.030 ;
        RECT 103.995 127.845 104.285 127.890 ;
        RECT 108.580 127.830 108.900 127.890 ;
        RECT 116.875 128.030 117.165 128.075 ;
        RECT 118.700 128.030 119.020 128.090 ;
        RECT 116.875 127.890 119.020 128.030 ;
        RECT 116.875 127.845 117.165 127.890 ;
        RECT 118.700 127.830 119.020 127.890 ;
        RECT 140.780 127.830 141.100 128.090 ;
        RECT 76.470 127.550 79.830 127.690 ;
        RECT 52.935 127.505 53.225 127.550 ;
        RECT 55.680 127.490 56.000 127.550 ;
        RECT 34.535 127.210 35.760 127.350 ;
        RECT 34.535 127.165 34.825 127.210 ;
        RECT 34.610 127.010 34.750 127.165 ;
        RECT 35.440 127.150 35.760 127.210 ;
        RECT 36.375 127.165 36.665 127.395 ;
        RECT 30.930 126.870 34.750 127.010 ;
        RECT 34.995 127.010 35.285 127.055 ;
        RECT 35.900 127.010 36.220 127.070 ;
        RECT 34.995 126.870 36.220 127.010 ;
        RECT 21.155 126.825 21.445 126.870 ;
        RECT 22.345 126.825 22.635 126.870 ;
        RECT 24.865 126.825 25.155 126.870 ;
        RECT 34.995 126.825 35.285 126.870 ;
        RECT 35.900 126.810 36.220 126.870 ;
        RECT 20.760 126.670 21.050 126.715 ;
        RECT 22.860 126.670 23.150 126.715 ;
        RECT 24.430 126.670 24.720 126.715 ;
        RECT 20.760 126.530 24.720 126.670 ;
        RECT 20.760 126.485 21.050 126.530 ;
        RECT 22.860 126.485 23.150 126.530 ;
        RECT 24.430 126.485 24.720 126.530 ;
        RECT 29.920 126.470 30.240 126.730 ;
        RECT 32.695 126.670 32.985 126.715 ;
        RECT 35.440 126.670 35.760 126.730 ;
        RECT 32.695 126.530 35.760 126.670 ;
        RECT 36.450 126.670 36.590 127.165 ;
        RECT 37.740 127.150 38.060 127.410 ;
        RECT 38.200 127.350 38.520 127.410 ;
        RECT 39.135 127.350 39.425 127.395 ;
        RECT 38.200 127.210 39.425 127.350 ;
        RECT 38.200 127.150 38.520 127.210 ;
        RECT 39.135 127.165 39.425 127.210 ;
        RECT 39.595 127.165 39.885 127.395 ;
        RECT 45.560 127.350 45.880 127.410 ;
        RECT 51.080 127.350 51.400 127.410 ;
        RECT 51.555 127.350 51.845 127.395 ;
        RECT 45.560 127.210 51.845 127.350 ;
        RECT 38.660 127.010 38.980 127.070 ;
        RECT 39.670 127.010 39.810 127.165 ;
        RECT 45.560 127.150 45.880 127.210 ;
        RECT 51.080 127.150 51.400 127.210 ;
        RECT 51.555 127.165 51.845 127.210 ;
        RECT 52.000 127.150 52.320 127.410 ;
        RECT 56.140 127.350 56.460 127.410 ;
        RECT 58.960 127.350 59.250 127.395 ;
        RECT 56.140 127.210 59.250 127.350 ;
        RECT 56.140 127.150 56.460 127.210 ;
        RECT 58.960 127.165 59.250 127.210 ;
        RECT 60.295 127.350 60.585 127.395 ;
        RECT 66.720 127.350 67.040 127.410 ;
        RECT 70.860 127.395 71.180 127.410 ;
        RECT 69.495 127.350 69.785 127.395 ;
        RECT 60.295 127.210 69.785 127.350 ;
        RECT 60.295 127.165 60.585 127.210 ;
        RECT 66.720 127.150 67.040 127.210 ;
        RECT 69.495 127.165 69.785 127.210 ;
        RECT 70.830 127.165 71.180 127.395 ;
        RECT 70.860 127.150 71.180 127.165 ;
        RECT 76.840 127.150 77.160 127.410 ;
        RECT 77.850 127.395 77.990 127.550 ;
        RECT 77.775 127.165 78.065 127.395 ;
        RECT 78.220 127.150 78.540 127.410 ;
        RECT 38.660 126.870 39.810 127.010 ;
        RECT 50.160 127.010 50.480 127.070 ;
        RECT 52.920 127.010 53.240 127.070 ;
        RECT 50.160 126.870 53.240 127.010 ;
        RECT 38.660 126.810 38.980 126.870 ;
        RECT 50.160 126.810 50.480 126.870 ;
        RECT 52.920 126.810 53.240 126.870 ;
        RECT 55.705 127.010 55.995 127.055 ;
        RECT 58.225 127.010 58.515 127.055 ;
        RECT 59.415 127.010 59.705 127.055 ;
        RECT 55.705 126.870 59.705 127.010 ;
        RECT 55.705 126.825 55.995 126.870 ;
        RECT 58.225 126.825 58.515 126.870 ;
        RECT 59.415 126.825 59.705 126.870 ;
        RECT 70.375 127.010 70.665 127.055 ;
        RECT 71.565 127.010 71.855 127.055 ;
        RECT 74.085 127.010 74.375 127.055 ;
        RECT 70.375 126.870 74.375 127.010 ;
        RECT 76.930 127.010 77.070 127.150 ;
        RECT 76.930 126.870 77.990 127.010 ;
        RECT 70.375 126.825 70.665 126.870 ;
        RECT 71.565 126.825 71.855 126.870 ;
        RECT 74.085 126.825 74.375 126.870 ;
        RECT 77.850 126.730 77.990 126.870 ;
        RECT 38.215 126.670 38.505 126.715 ;
        RECT 36.450 126.530 38.505 126.670 ;
        RECT 32.695 126.485 32.985 126.530 ;
        RECT 35.440 126.470 35.760 126.530 ;
        RECT 38.215 126.485 38.505 126.530 ;
        RECT 56.140 126.670 56.430 126.715 ;
        RECT 57.710 126.670 58.000 126.715 ;
        RECT 59.810 126.670 60.100 126.715 ;
        RECT 56.140 126.530 60.100 126.670 ;
        RECT 56.140 126.485 56.430 126.530 ;
        RECT 57.710 126.485 58.000 126.530 ;
        RECT 59.810 126.485 60.100 126.530 ;
        RECT 69.980 126.670 70.270 126.715 ;
        RECT 72.080 126.670 72.370 126.715 ;
        RECT 73.650 126.670 73.940 126.715 ;
        RECT 69.980 126.530 73.940 126.670 ;
        RECT 69.980 126.485 70.270 126.530 ;
        RECT 72.080 126.485 72.370 126.530 ;
        RECT 73.650 126.485 73.940 126.530 ;
        RECT 77.760 126.470 78.080 126.730 ;
        RECT 26.700 126.330 27.020 126.390 ;
        RECT 27.175 126.330 27.465 126.375 ;
        RECT 28.555 126.330 28.845 126.375 ;
        RECT 31.300 126.330 31.620 126.390 ;
        RECT 20.350 126.190 31.620 126.330 ;
        RECT 26.700 126.130 27.020 126.190 ;
        RECT 27.175 126.145 27.465 126.190 ;
        RECT 28.555 126.145 28.845 126.190 ;
        RECT 31.300 126.130 31.620 126.190 ;
        RECT 34.535 126.330 34.825 126.375 ;
        RECT 34.980 126.330 35.300 126.390 ;
        RECT 34.535 126.190 35.300 126.330 ;
        RECT 34.535 126.145 34.825 126.190 ;
        RECT 34.980 126.130 35.300 126.190 ;
        RECT 35.900 126.330 36.220 126.390 ;
        RECT 40.040 126.330 40.360 126.390 ;
        RECT 56.600 126.330 56.920 126.390 ;
        RECT 35.900 126.190 56.920 126.330 ;
        RECT 79.690 126.330 79.830 127.550 ;
        RECT 80.060 127.490 80.380 127.750 ;
        RECT 98.460 127.735 98.780 127.750 ;
        RECT 98.430 127.690 98.780 127.735 ;
        RECT 116.400 127.690 116.720 127.750 ;
        RECT 130.200 127.690 130.520 127.750 ;
        RECT 134.800 127.690 135.120 127.750 ;
        RECT 85.670 127.550 97.310 127.690 ;
        RECT 98.265 127.550 98.780 127.690 ;
        RECT 85.670 127.410 85.810 127.550 ;
        RECT 97.170 127.410 97.310 127.550 ;
        RECT 98.430 127.505 98.780 127.550 ;
        RECT 98.460 127.490 98.780 127.505 ;
        RECT 110.050 127.550 121.230 127.690 ;
        RECT 81.440 127.350 81.760 127.410 ;
        RECT 83.295 127.350 83.585 127.395 ;
        RECT 84.200 127.350 84.520 127.410 ;
        RECT 81.440 127.210 84.520 127.350 ;
        RECT 81.440 127.150 81.760 127.210 ;
        RECT 83.295 127.165 83.585 127.210 ;
        RECT 84.200 127.150 84.520 127.210 ;
        RECT 85.580 127.150 85.900 127.410 ;
        RECT 86.930 127.350 87.220 127.395 ;
        RECT 89.720 127.350 90.040 127.410 ;
        RECT 86.930 127.210 90.040 127.350 ;
        RECT 86.930 127.165 87.220 127.210 ;
        RECT 89.720 127.150 90.040 127.210 ;
        RECT 97.080 127.150 97.400 127.410 ;
        RECT 106.295 127.350 106.585 127.395 ;
        RECT 108.120 127.350 108.440 127.410 ;
        RECT 110.050 127.395 110.190 127.550 ;
        RECT 116.400 127.490 116.720 127.550 ;
        RECT 111.340 127.395 111.660 127.410 ;
        RECT 106.295 127.210 108.440 127.350 ;
        RECT 106.295 127.165 106.585 127.210 ;
        RECT 108.120 127.150 108.440 127.210 ;
        RECT 109.975 127.165 110.265 127.395 ;
        RECT 111.310 127.165 111.660 127.395 ;
        RECT 111.340 127.150 111.660 127.165 ;
        RECT 112.720 127.350 113.040 127.410 ;
        RECT 121.090 127.395 121.230 127.550 ;
        RECT 130.200 127.550 135.950 127.690 ;
        RECT 130.200 127.490 130.520 127.550 ;
        RECT 134.800 127.490 135.120 127.550 ;
        RECT 117.795 127.350 118.085 127.395 ;
        RECT 112.720 127.210 118.085 127.350 ;
        RECT 112.720 127.150 113.040 127.210 ;
        RECT 117.795 127.165 118.085 127.210 ;
        RECT 121.015 127.165 121.305 127.395 ;
        RECT 121.460 127.350 121.780 127.410 ;
        RECT 132.500 127.395 132.820 127.410 ;
        RECT 122.295 127.350 122.585 127.395 ;
        RECT 121.460 127.210 122.585 127.350 ;
        RECT 121.460 127.150 121.780 127.210 ;
        RECT 122.295 127.165 122.585 127.210 ;
        RECT 132.470 127.165 132.820 127.395 ;
        RECT 135.810 127.350 135.950 127.550 ;
        RECT 135.810 127.210 136.410 127.350 ;
        RECT 132.500 127.150 132.820 127.165 ;
        RECT 81.915 126.825 82.205 127.055 ;
        RECT 82.820 127.010 83.140 127.070 ;
        RECT 86.475 127.010 86.765 127.055 ;
        RECT 87.665 127.010 87.955 127.055 ;
        RECT 90.185 127.010 90.475 127.055 ;
        RECT 82.820 126.870 85.810 127.010 ;
        RECT 80.995 126.670 81.285 126.715 ;
        RECT 81.990 126.670 82.130 126.825 ;
        RECT 82.820 126.810 83.140 126.870 ;
        RECT 80.995 126.530 82.130 126.670 ;
        RECT 80.995 126.485 81.285 126.530 ;
        RECT 80.075 126.330 80.365 126.375 ;
        RECT 82.820 126.330 83.140 126.390 ;
        RECT 79.690 126.190 83.140 126.330 ;
        RECT 85.670 126.330 85.810 126.870 ;
        RECT 86.475 126.870 90.475 127.010 ;
        RECT 86.475 126.825 86.765 126.870 ;
        RECT 87.665 126.825 87.955 126.870 ;
        RECT 90.185 126.825 90.475 126.870 ;
        RECT 97.975 127.010 98.265 127.055 ;
        RECT 99.165 127.010 99.455 127.055 ;
        RECT 101.685 127.010 101.975 127.055 ;
        RECT 97.975 126.870 101.975 127.010 ;
        RECT 97.975 126.825 98.265 126.870 ;
        RECT 99.165 126.825 99.455 126.870 ;
        RECT 101.685 126.825 101.975 126.870 ;
        RECT 106.740 126.810 107.060 127.070 ;
        RECT 107.200 126.810 107.520 127.070 ;
        RECT 110.855 127.010 111.145 127.055 ;
        RECT 112.045 127.010 112.335 127.055 ;
        RECT 114.565 127.010 114.855 127.055 ;
        RECT 110.855 126.870 114.855 127.010 ;
        RECT 110.855 126.825 111.145 126.870 ;
        RECT 112.045 126.825 112.335 126.870 ;
        RECT 114.565 126.825 114.855 126.870 ;
        RECT 121.895 127.010 122.185 127.055 ;
        RECT 123.085 127.010 123.375 127.055 ;
        RECT 125.605 127.010 125.895 127.055 ;
        RECT 121.895 126.870 125.895 127.010 ;
        RECT 121.895 126.825 122.185 126.870 ;
        RECT 123.085 126.825 123.375 126.870 ;
        RECT 125.605 126.825 125.895 126.870 ;
        RECT 131.120 126.810 131.440 127.070 ;
        RECT 132.015 127.010 132.305 127.055 ;
        RECT 133.205 127.010 133.495 127.055 ;
        RECT 135.725 127.010 136.015 127.055 ;
        RECT 132.015 126.870 136.015 127.010 ;
        RECT 132.015 126.825 132.305 126.870 ;
        RECT 133.205 126.825 133.495 126.870 ;
        RECT 135.725 126.825 136.015 126.870 ;
        RECT 86.080 126.670 86.370 126.715 ;
        RECT 88.180 126.670 88.470 126.715 ;
        RECT 89.750 126.670 90.040 126.715 ;
        RECT 86.080 126.530 90.040 126.670 ;
        RECT 86.080 126.485 86.370 126.530 ;
        RECT 88.180 126.485 88.470 126.530 ;
        RECT 89.750 126.485 90.040 126.530 ;
        RECT 97.580 126.670 97.870 126.715 ;
        RECT 99.680 126.670 99.970 126.715 ;
        RECT 101.250 126.670 101.540 126.715 ;
        RECT 97.580 126.530 101.540 126.670 ;
        RECT 97.580 126.485 97.870 126.530 ;
        RECT 99.680 126.485 99.970 126.530 ;
        RECT 101.250 126.485 101.540 126.530 ;
        RECT 110.460 126.670 110.750 126.715 ;
        RECT 112.560 126.670 112.850 126.715 ;
        RECT 114.130 126.670 114.420 126.715 ;
        RECT 110.460 126.530 114.420 126.670 ;
        RECT 110.460 126.485 110.750 126.530 ;
        RECT 112.560 126.485 112.850 126.530 ;
        RECT 114.130 126.485 114.420 126.530 ;
        RECT 115.480 126.670 115.800 126.730 ;
        RECT 121.000 126.670 121.320 126.730 ;
        RECT 115.480 126.530 121.320 126.670 ;
        RECT 115.480 126.470 115.800 126.530 ;
        RECT 121.000 126.470 121.320 126.530 ;
        RECT 121.500 126.670 121.790 126.715 ;
        RECT 123.600 126.670 123.890 126.715 ;
        RECT 125.170 126.670 125.460 126.715 ;
        RECT 130.200 126.670 130.520 126.730 ;
        RECT 121.500 126.530 125.460 126.670 ;
        RECT 121.500 126.485 121.790 126.530 ;
        RECT 123.600 126.485 123.890 126.530 ;
        RECT 125.170 126.485 125.460 126.530 ;
        RECT 125.690 126.530 130.520 126.670 ;
        RECT 90.180 126.330 90.500 126.390 ;
        RECT 92.020 126.330 92.340 126.390 ;
        RECT 85.670 126.190 92.340 126.330 ;
        RECT 35.900 126.130 36.220 126.190 ;
        RECT 40.040 126.130 40.360 126.190 ;
        RECT 56.600 126.130 56.920 126.190 ;
        RECT 80.075 126.145 80.365 126.190 ;
        RECT 82.820 126.130 83.140 126.190 ;
        RECT 90.180 126.130 90.500 126.190 ;
        RECT 92.020 126.130 92.340 126.190 ;
        RECT 92.495 126.330 92.785 126.375 ;
        RECT 94.780 126.330 95.100 126.390 ;
        RECT 98.920 126.330 99.240 126.390 ;
        RECT 92.495 126.190 99.240 126.330 ;
        RECT 92.495 126.145 92.785 126.190 ;
        RECT 94.780 126.130 95.100 126.190 ;
        RECT 98.920 126.130 99.240 126.190 ;
        RECT 104.440 126.130 104.760 126.390 ;
        RECT 114.560 126.330 114.880 126.390 ;
        RECT 118.255 126.330 118.545 126.375 ;
        RECT 114.560 126.190 118.545 126.330 ;
        RECT 114.560 126.130 114.880 126.190 ;
        RECT 118.255 126.145 118.545 126.190 ;
        RECT 122.380 126.330 122.700 126.390 ;
        RECT 125.690 126.330 125.830 126.530 ;
        RECT 130.200 126.470 130.520 126.530 ;
        RECT 131.620 126.670 131.910 126.715 ;
        RECT 133.720 126.670 134.010 126.715 ;
        RECT 135.290 126.670 135.580 126.715 ;
        RECT 131.620 126.530 135.580 126.670 ;
        RECT 136.270 126.670 136.410 127.210 ;
        RECT 139.860 127.150 140.180 127.410 ;
        RECT 138.035 126.670 138.325 126.715 ;
        RECT 139.860 126.670 140.180 126.730 ;
        RECT 136.270 126.530 140.180 126.670 ;
        RECT 131.620 126.485 131.910 126.530 ;
        RECT 133.720 126.485 134.010 126.530 ;
        RECT 135.290 126.485 135.580 126.530 ;
        RECT 138.035 126.485 138.325 126.530 ;
        RECT 139.860 126.470 140.180 126.530 ;
        RECT 122.380 126.190 125.830 126.330 ;
        RECT 127.900 126.330 128.220 126.390 ;
        RECT 138.480 126.330 138.800 126.390 ;
        RECT 127.900 126.190 138.800 126.330 ;
        RECT 122.380 126.130 122.700 126.190 ;
        RECT 127.900 126.130 128.220 126.190 ;
        RECT 138.480 126.130 138.800 126.190 ;
        RECT 17.430 125.510 143.010 125.990 ;
        RECT 29.000 125.110 29.320 125.370 ;
        RECT 31.775 125.310 32.065 125.355 ;
        RECT 35.900 125.310 36.220 125.370 ;
        RECT 31.775 125.170 36.220 125.310 ;
        RECT 31.775 125.125 32.065 125.170 ;
        RECT 35.900 125.110 36.220 125.170 ;
        RECT 38.215 125.310 38.505 125.355 ;
        RECT 39.580 125.310 39.900 125.370 ;
        RECT 38.215 125.170 39.900 125.310 ;
        RECT 38.215 125.125 38.505 125.170 ;
        RECT 39.580 125.110 39.900 125.170 ;
        RECT 45.560 125.110 45.880 125.370 ;
        RECT 48.320 125.310 48.640 125.370 ;
        RECT 48.795 125.310 49.085 125.355 ;
        RECT 46.570 125.170 48.090 125.310 ;
        RECT 22.600 124.970 22.890 125.015 ;
        RECT 24.700 124.970 24.990 125.015 ;
        RECT 26.270 124.970 26.560 125.015 ;
        RECT 22.600 124.830 26.560 124.970 ;
        RECT 22.600 124.785 22.890 124.830 ;
        RECT 24.700 124.785 24.990 124.830 ;
        RECT 26.270 124.785 26.560 124.830 ;
        RECT 39.160 124.970 39.450 125.015 ;
        RECT 41.260 124.970 41.550 125.015 ;
        RECT 42.830 124.970 43.120 125.015 ;
        RECT 39.160 124.830 43.120 124.970 ;
        RECT 39.160 124.785 39.450 124.830 ;
        RECT 41.260 124.785 41.550 124.830 ;
        RECT 42.830 124.785 43.120 124.830 ;
        RECT 22.995 124.630 23.285 124.675 ;
        RECT 24.185 124.630 24.475 124.675 ;
        RECT 26.705 124.630 26.995 124.675 ;
        RECT 33.615 124.630 33.905 124.675 ;
        RECT 35.440 124.630 35.760 124.690 ;
        RECT 36.835 124.630 37.125 124.675 ;
        RECT 39.555 124.630 39.845 124.675 ;
        RECT 40.745 124.630 41.035 124.675 ;
        RECT 43.265 124.630 43.555 124.675 ;
        RECT 22.995 124.490 26.995 124.630 ;
        RECT 22.995 124.445 23.285 124.490 ;
        RECT 24.185 124.445 24.475 124.490 ;
        RECT 26.705 124.445 26.995 124.490 ;
        RECT 32.310 124.490 33.905 124.630 ;
        RECT 22.115 124.290 22.405 124.335 ;
        RECT 27.160 124.290 27.480 124.350 ;
        RECT 22.115 124.150 27.480 124.290 ;
        RECT 22.115 124.105 22.405 124.150 ;
        RECT 27.160 124.090 27.480 124.150 ;
        RECT 23.450 123.950 23.740 123.995 ;
        RECT 28.080 123.950 28.400 124.010 ;
        RECT 23.450 123.810 28.400 123.950 ;
        RECT 23.450 123.765 23.740 123.810 ;
        RECT 28.080 123.750 28.400 123.810 ;
        RECT 30.840 123.750 31.160 124.010 ;
        RECT 31.880 123.950 32.170 123.995 ;
        RECT 32.310 123.950 32.450 124.490 ;
        RECT 33.615 124.445 33.905 124.490 ;
        RECT 34.150 124.490 39.350 124.630 ;
        RECT 33.140 124.090 33.460 124.350 ;
        RECT 34.150 124.335 34.290 124.490 ;
        RECT 35.440 124.430 35.760 124.490 ;
        RECT 36.835 124.445 37.125 124.490 ;
        RECT 34.075 124.105 34.365 124.335 ;
        RECT 36.375 124.290 36.665 124.335 ;
        RECT 38.200 124.290 38.520 124.350 ;
        RECT 36.375 124.150 38.520 124.290 ;
        RECT 36.375 124.105 36.665 124.150 ;
        RECT 38.200 124.090 38.520 124.150 ;
        RECT 38.675 124.105 38.965 124.335 ;
        RECT 39.210 124.290 39.350 124.490 ;
        RECT 39.555 124.490 43.555 124.630 ;
        RECT 39.555 124.445 39.845 124.490 ;
        RECT 40.745 124.445 41.035 124.490 ;
        RECT 43.265 124.445 43.555 124.490 ;
        RECT 46.035 124.290 46.325 124.335 ;
        RECT 46.570 124.290 46.710 125.170 ;
        RECT 47.415 124.785 47.705 125.015 ;
        RECT 39.210 124.150 46.710 124.290 ;
        RECT 47.490 124.290 47.630 124.785 ;
        RECT 47.950 124.630 48.090 125.170 ;
        RECT 48.320 125.170 49.085 125.310 ;
        RECT 48.320 125.110 48.640 125.170 ;
        RECT 48.795 125.125 49.085 125.170 ;
        RECT 51.080 125.110 51.400 125.370 ;
        RECT 52.015 125.310 52.305 125.355 ;
        RECT 53.380 125.310 53.700 125.370 ;
        RECT 52.015 125.170 53.700 125.310 ;
        RECT 52.015 125.125 52.305 125.170 ;
        RECT 53.380 125.110 53.700 125.170 ;
        RECT 54.775 125.125 55.065 125.355 ;
        RECT 55.695 125.310 55.985 125.355 ;
        RECT 56.140 125.310 56.460 125.370 ;
        RECT 55.695 125.170 56.460 125.310 ;
        RECT 55.695 125.125 55.985 125.170 ;
        RECT 49.715 124.970 50.005 125.015 ;
        RECT 54.300 124.970 54.620 125.030 ;
        RECT 49.715 124.830 54.620 124.970 ;
        RECT 54.850 124.970 54.990 125.125 ;
        RECT 56.140 125.110 56.460 125.170 ;
        RECT 70.860 125.310 71.180 125.370 ;
        RECT 71.795 125.310 72.085 125.355 ;
        RECT 70.860 125.170 72.085 125.310 ;
        RECT 70.860 125.110 71.180 125.170 ;
        RECT 71.795 125.125 72.085 125.170 ;
        RECT 76.380 125.110 76.700 125.370 ;
        RECT 82.820 125.310 83.140 125.370 ;
        RECT 83.295 125.310 83.585 125.355 ;
        RECT 82.820 125.170 83.585 125.310 ;
        RECT 82.820 125.110 83.140 125.170 ;
        RECT 83.295 125.125 83.585 125.170 ;
        RECT 85.595 125.310 85.885 125.355 ;
        RECT 86.040 125.310 86.360 125.370 ;
        RECT 85.595 125.170 86.360 125.310 ;
        RECT 85.595 125.125 85.885 125.170 ;
        RECT 56.600 124.970 56.920 125.030 ;
        RECT 77.300 124.970 77.620 125.030 ;
        RECT 54.850 124.830 56.920 124.970 ;
        RECT 49.715 124.785 50.005 124.830 ;
        RECT 54.300 124.770 54.620 124.830 ;
        RECT 56.600 124.770 56.920 124.830 ;
        RECT 73.940 124.830 77.620 124.970 ;
        RECT 83.370 124.970 83.510 125.125 ;
        RECT 86.040 125.110 86.360 125.170 ;
        RECT 86.930 125.125 87.220 125.355 ;
        RECT 103.980 125.310 104.300 125.370 ;
        RECT 105.375 125.310 105.665 125.355 ;
        RECT 103.980 125.170 105.665 125.310 ;
        RECT 86.500 124.970 86.820 125.030 ;
        RECT 87.005 124.970 87.145 125.125 ;
        RECT 103.980 125.110 104.300 125.170 ;
        RECT 105.375 125.125 105.665 125.170 ;
        RECT 83.370 124.830 87.145 124.970 ;
        RECT 88.840 124.970 89.130 125.015 ;
        RECT 90.940 124.970 91.230 125.015 ;
        RECT 92.510 124.970 92.800 125.015 ;
        RECT 88.840 124.830 92.800 124.970 ;
        RECT 52.000 124.630 52.320 124.690 ;
        RECT 54.760 124.630 55.080 124.690 ;
        RECT 47.950 124.490 52.320 124.630 ;
        RECT 52.000 124.430 52.320 124.490 ;
        RECT 53.930 124.490 55.080 124.630 ;
        RECT 52.475 124.290 52.765 124.335 ;
        RECT 47.490 124.150 52.765 124.290 ;
        RECT 46.035 124.105 46.325 124.150 ;
        RECT 52.475 124.105 52.765 124.150 ;
        RECT 31.880 123.810 32.450 123.950 ;
        RECT 33.600 123.950 33.920 124.010 ;
        RECT 38.750 123.950 38.890 124.105 ;
        RECT 52.920 124.090 53.240 124.350 ;
        RECT 53.380 124.090 53.700 124.350 ;
        RECT 33.600 123.810 38.890 123.950 ;
        RECT 40.010 123.950 40.300 123.995 ;
        RECT 40.500 123.950 40.820 124.010 ;
        RECT 40.010 123.810 40.820 123.950 ;
        RECT 31.880 123.765 32.170 123.810 ;
        RECT 33.600 123.750 33.920 123.810 ;
        RECT 40.010 123.765 40.300 123.810 ;
        RECT 40.500 123.750 40.820 123.810 ;
        RECT 45.560 123.950 45.880 124.010 ;
        RECT 46.495 123.950 46.785 123.995 ;
        RECT 45.560 123.810 46.785 123.950 ;
        RECT 45.560 123.750 45.880 123.810 ;
        RECT 46.495 123.765 46.785 123.810 ;
        RECT 47.415 123.765 47.705 123.995 ;
        RECT 32.680 123.410 33.000 123.670 ;
        RECT 47.490 123.610 47.630 123.765 ;
        RECT 47.860 123.750 48.180 124.010 ;
        RECT 48.780 123.995 49.100 124.010 ;
        RECT 48.780 123.765 49.165 123.995 ;
        RECT 48.780 123.750 49.100 123.765 ;
        RECT 50.160 123.750 50.480 124.010 ;
        RECT 53.930 123.995 54.070 124.490 ;
        RECT 54.760 124.430 55.080 124.490 ;
        RECT 72.715 124.290 73.005 124.335 ;
        RECT 73.940 124.290 74.080 124.830 ;
        RECT 77.300 124.770 77.620 124.830 ;
        RECT 86.500 124.770 86.820 124.830 ;
        RECT 88.840 124.785 89.130 124.830 ;
        RECT 90.940 124.785 91.230 124.830 ;
        RECT 92.510 124.785 92.800 124.830 ;
        RECT 98.960 124.970 99.250 125.015 ;
        RECT 101.060 124.970 101.350 125.015 ;
        RECT 102.630 124.970 102.920 125.015 ;
        RECT 98.960 124.830 102.920 124.970 ;
        RECT 98.960 124.785 99.250 124.830 ;
        RECT 101.060 124.785 101.350 124.830 ;
        RECT 102.630 124.785 102.920 124.830 ;
        RECT 78.220 124.630 78.540 124.690 ;
        RECT 84.215 124.630 84.505 124.675 ;
        RECT 75.090 124.490 84.505 124.630 ;
        RECT 75.090 124.350 75.230 124.490 ;
        RECT 78.220 124.430 78.540 124.490 ;
        RECT 84.215 124.445 84.505 124.490 ;
        RECT 85.580 124.630 85.900 124.690 ;
        RECT 88.355 124.630 88.645 124.675 ;
        RECT 85.580 124.490 88.645 124.630 ;
        RECT 72.715 124.150 74.080 124.290 ;
        RECT 72.715 124.105 73.005 124.150 ;
        RECT 75.000 124.090 75.320 124.350 ;
        RECT 75.935 124.290 76.225 124.335 ;
        RECT 77.315 124.290 77.605 124.335 ;
        RECT 75.935 124.150 77.605 124.290 ;
        RECT 75.935 124.105 76.225 124.150 ;
        RECT 77.315 124.105 77.605 124.150 ;
        RECT 77.760 124.090 78.080 124.350 ;
        RECT 80.060 124.290 80.380 124.350 ;
        RECT 82.835 124.290 83.125 124.335 ;
        RECT 78.310 124.150 83.125 124.290 ;
        RECT 55.220 123.995 55.540 124.010 ;
        RECT 53.855 123.765 54.145 123.995 ;
        RECT 54.935 123.765 55.540 123.995 ;
        RECT 55.220 123.750 55.540 123.765 ;
        RECT 72.240 123.950 72.560 124.010 ;
        RECT 73.635 123.950 73.925 123.995 ;
        RECT 72.240 123.810 73.925 123.950 ;
        RECT 72.240 123.750 72.560 123.810 ;
        RECT 73.635 123.765 73.925 123.810 ;
        RECT 74.080 123.750 74.400 124.010 ;
        RECT 50.250 123.610 50.390 123.750 ;
        RECT 47.490 123.470 50.390 123.610 ;
        RECT 51.225 123.610 51.515 123.655 ;
        RECT 52.000 123.610 52.320 123.670 ;
        RECT 51.225 123.470 52.320 123.610 ;
        RECT 74.170 123.610 74.310 123.750 ;
        RECT 78.310 123.610 78.450 124.150 ;
        RECT 80.060 124.090 80.380 124.150 ;
        RECT 82.835 124.105 83.125 124.150 ;
        RECT 84.290 123.950 84.430 124.445 ;
        RECT 85.580 124.430 85.900 124.490 ;
        RECT 88.355 124.445 88.645 124.490 ;
        RECT 89.235 124.630 89.525 124.675 ;
        RECT 90.425 124.630 90.715 124.675 ;
        RECT 92.945 124.630 93.235 124.675 ;
        RECT 89.235 124.490 93.235 124.630 ;
        RECT 89.235 124.445 89.525 124.490 ;
        RECT 90.425 124.445 90.715 124.490 ;
        RECT 92.945 124.445 93.235 124.490 ;
        RECT 97.080 124.630 97.400 124.690 ;
        RECT 98.475 124.630 98.765 124.675 ;
        RECT 97.080 124.490 98.765 124.630 ;
        RECT 97.080 124.430 97.400 124.490 ;
        RECT 98.475 124.445 98.765 124.490 ;
        RECT 99.355 124.630 99.645 124.675 ;
        RECT 100.545 124.630 100.835 124.675 ;
        RECT 103.065 124.630 103.355 124.675 ;
        RECT 99.355 124.490 103.355 124.630 ;
        RECT 105.450 124.630 105.590 125.125 ;
        RECT 108.120 125.110 108.440 125.370 ;
        RECT 111.340 125.310 111.660 125.370 ;
        RECT 111.815 125.310 112.105 125.355 ;
        RECT 111.340 125.170 112.105 125.310 ;
        RECT 111.340 125.110 111.660 125.170 ;
        RECT 111.815 125.125 112.105 125.170 ;
        RECT 120.555 125.310 120.845 125.355 ;
        RECT 121.460 125.310 121.780 125.370 ;
        RECT 120.555 125.170 121.780 125.310 ;
        RECT 120.555 125.125 120.845 125.170 ;
        RECT 121.460 125.110 121.780 125.170 ;
        RECT 126.520 125.310 126.840 125.370 ;
        RECT 126.520 125.170 136.870 125.310 ;
        RECT 126.520 125.110 126.840 125.170 ;
        RECT 106.740 124.970 107.060 125.030 ;
        RECT 115.495 124.970 115.785 125.015 ;
        RECT 122.840 124.970 123.160 125.030 ;
        RECT 106.740 124.830 112.030 124.970 ;
        RECT 106.740 124.770 107.060 124.830 ;
        RECT 110.895 124.630 111.185 124.675 ;
        RECT 105.450 124.490 111.185 124.630 ;
        RECT 111.890 124.630 112.030 124.830 ;
        RECT 113.730 124.830 115.785 124.970 ;
        RECT 113.730 124.630 113.870 124.830 ;
        RECT 115.495 124.785 115.785 124.830 ;
        RECT 122.240 124.830 123.160 124.970 ;
        RECT 111.890 124.490 113.870 124.630 ;
        RECT 114.560 124.630 114.880 124.690 ;
        RECT 118.700 124.630 119.020 124.690 ;
        RECT 122.240 124.630 122.380 124.830 ;
        RECT 122.840 124.770 123.160 124.830 ;
        RECT 129.740 124.970 130.060 125.030 ;
        RECT 136.195 124.970 136.485 125.015 ;
        RECT 129.740 124.830 136.485 124.970 ;
        RECT 129.740 124.770 130.060 124.830 ;
        RECT 136.195 124.785 136.485 124.830 ;
        RECT 124.235 124.630 124.525 124.675 ;
        RECT 127.900 124.630 128.220 124.690 ;
        RECT 114.560 124.490 116.630 124.630 ;
        RECT 99.355 124.445 99.645 124.490 ;
        RECT 100.545 124.445 100.835 124.490 ;
        RECT 103.065 124.445 103.355 124.490 ;
        RECT 110.895 124.445 111.185 124.490 ;
        RECT 114.560 124.430 114.880 124.490 ;
        RECT 99.810 124.290 100.100 124.335 ;
        RECT 104.440 124.290 104.760 124.350 ;
        RECT 99.810 124.150 104.760 124.290 ;
        RECT 99.810 124.105 100.100 124.150 ;
        RECT 104.440 124.090 104.760 124.150 ;
        RECT 113.180 124.090 113.500 124.350 ;
        RECT 113.655 124.105 113.945 124.335 ;
        RECT 84.660 123.950 84.980 124.010 ;
        RECT 86.055 123.950 86.345 123.995 ;
        RECT 84.290 123.810 86.345 123.950 ;
        RECT 84.660 123.750 84.980 123.810 ;
        RECT 86.055 123.765 86.345 123.810 ;
        RECT 88.800 123.950 89.120 124.010 ;
        RECT 89.580 123.950 89.870 123.995 ;
        RECT 88.800 123.810 89.870 123.950 ;
        RECT 88.800 123.750 89.120 123.810 ;
        RECT 89.580 123.765 89.870 123.810 ;
        RECT 98.920 123.950 99.240 124.010 ;
        RECT 113.730 123.950 113.870 124.105 ;
        RECT 114.100 124.090 114.420 124.350 ;
        RECT 116.490 124.335 116.630 124.490 ;
        RECT 116.950 124.490 119.020 124.630 ;
        RECT 116.950 124.335 117.090 124.490 ;
        RECT 118.700 124.430 119.020 124.490 ;
        RECT 122.010 124.490 122.380 124.630 ;
        RECT 122.930 124.490 124.525 124.630 ;
        RECT 115.035 124.105 115.325 124.335 ;
        RECT 116.415 124.105 116.705 124.335 ;
        RECT 116.875 124.105 117.165 124.335 ;
        RECT 115.110 123.950 115.250 124.105 ;
        RECT 117.780 124.090 118.100 124.350 ;
        RECT 118.255 124.290 118.545 124.335 ;
        RECT 119.160 124.290 119.480 124.350 ;
        RECT 118.255 124.150 119.480 124.290 ;
        RECT 118.255 124.105 118.545 124.150 ;
        RECT 119.160 124.090 119.480 124.150 ;
        RECT 119.620 124.290 119.940 124.350 ;
        RECT 122.010 124.335 122.150 124.490 ;
        RECT 121.935 124.290 122.225 124.335 ;
        RECT 119.620 124.150 122.225 124.290 ;
        RECT 119.620 124.090 119.940 124.150 ;
        RECT 121.935 124.105 122.225 124.150 ;
        RECT 122.380 124.090 122.700 124.350 ;
        RECT 122.930 124.335 123.070 124.490 ;
        RECT 124.235 124.445 124.525 124.490 ;
        RECT 125.230 124.490 128.220 124.630 ;
        RECT 122.855 124.105 123.145 124.335 ;
        RECT 123.760 124.090 124.080 124.350 ;
        RECT 125.230 124.335 125.370 124.490 ;
        RECT 127.900 124.430 128.220 124.490 ;
        RECT 128.820 124.630 129.140 124.690 ;
        RECT 130.200 124.630 130.520 124.690 ;
        RECT 128.820 124.490 129.970 124.630 ;
        RECT 128.820 124.430 129.140 124.490 ;
        RECT 129.830 124.335 129.970 124.490 ;
        RECT 130.200 124.490 131.350 124.630 ;
        RECT 130.200 124.430 130.520 124.490 ;
        RECT 131.210 124.335 131.350 124.490 ;
        RECT 132.975 124.445 133.265 124.675 ;
        RECT 136.730 124.630 136.870 125.170 ;
        RECT 140.780 125.110 141.100 125.370 ;
        RECT 135.810 124.490 138.250 124.630 ;
        RECT 125.155 124.105 125.445 124.335 ;
        RECT 129.755 124.105 130.045 124.335 ;
        RECT 130.675 124.105 130.965 124.335 ;
        RECT 131.135 124.105 131.425 124.335 ;
        RECT 121.000 123.950 121.320 124.010 ;
        RECT 98.920 123.810 114.790 123.950 ;
        RECT 115.110 123.810 121.320 123.950 ;
        RECT 98.920 123.750 99.240 123.810 ;
        RECT 74.170 123.470 78.450 123.610 ;
        RECT 86.500 123.610 86.820 123.670 ;
        RECT 87.055 123.610 87.345 123.655 ;
        RECT 86.500 123.470 87.345 123.610 ;
        RECT 51.225 123.425 51.515 123.470 ;
        RECT 52.000 123.410 52.320 123.470 ;
        RECT 86.500 123.410 86.820 123.470 ;
        RECT 87.055 123.425 87.345 123.470 ;
        RECT 87.895 123.610 88.185 123.655 ;
        RECT 91.560 123.610 91.880 123.670 ;
        RECT 87.895 123.470 91.880 123.610 ;
        RECT 87.895 123.425 88.185 123.470 ;
        RECT 91.560 123.410 91.880 123.470 ;
        RECT 95.255 123.610 95.545 123.655 ;
        RECT 97.540 123.610 97.860 123.670 ;
        RECT 95.255 123.470 97.860 123.610 ;
        RECT 114.650 123.610 114.790 123.810 ;
        RECT 116.950 123.670 117.090 123.810 ;
        RECT 121.000 123.750 121.320 123.810 ;
        RECT 126.075 123.950 126.365 123.995 ;
        RECT 126.520 123.950 126.840 124.010 ;
        RECT 126.075 123.810 126.840 123.950 ;
        RECT 130.750 123.950 130.890 124.105 ;
        RECT 131.580 124.090 131.900 124.350 ;
        RECT 132.500 124.290 132.820 124.350 ;
        RECT 133.050 124.290 133.190 124.445 ;
        RECT 135.810 124.335 135.950 124.490 ;
        RECT 132.500 124.150 133.190 124.290 ;
        RECT 132.500 124.090 132.820 124.150 ;
        RECT 135.735 124.105 136.025 124.335 ;
        RECT 133.895 123.950 134.185 123.995 ;
        RECT 130.750 123.810 134.185 123.950 ;
        RECT 126.075 123.765 126.365 123.810 ;
        RECT 126.520 123.750 126.840 123.810 ;
        RECT 133.895 123.765 134.185 123.810 ;
        RECT 134.800 123.750 135.120 124.010 ;
        RECT 136.180 123.950 136.500 124.010 ;
        RECT 138.110 123.995 138.250 124.490 ;
        RECT 138.480 124.290 138.800 124.350 ;
        RECT 139.875 124.290 140.165 124.335 ;
        RECT 138.480 124.150 140.165 124.290 ;
        RECT 138.480 124.090 138.800 124.150 ;
        RECT 139.875 124.105 140.165 124.150 ;
        RECT 137.115 123.950 137.405 123.995 ;
        RECT 136.180 123.810 137.405 123.950 ;
        RECT 136.180 123.750 136.500 123.810 ;
        RECT 137.115 123.765 137.405 123.810 ;
        RECT 138.035 123.765 138.325 123.995 ;
        RECT 115.020 123.610 115.340 123.670 ;
        RECT 114.650 123.470 115.340 123.610 ;
        RECT 95.255 123.425 95.545 123.470 ;
        RECT 97.540 123.410 97.860 123.470 ;
        RECT 115.020 123.410 115.340 123.470 ;
        RECT 116.860 123.410 117.180 123.670 ;
        RECT 17.430 122.790 143.010 123.270 ;
        RECT 26.255 122.590 26.545 122.635 ;
        RECT 29.920 122.590 30.240 122.650 ;
        RECT 26.255 122.450 30.240 122.590 ;
        RECT 26.255 122.405 26.545 122.450 ;
        RECT 29.920 122.390 30.240 122.450 ;
        RECT 30.840 122.590 31.160 122.650 ;
        RECT 39.135 122.590 39.425 122.635 ;
        RECT 40.500 122.590 40.820 122.650 ;
        RECT 30.840 122.450 34.585 122.590 ;
        RECT 30.840 122.390 31.160 122.450 ;
        RECT 27.160 122.250 27.480 122.310 ;
        RECT 33.600 122.250 33.920 122.310 ;
        RECT 27.160 122.110 33.920 122.250 ;
        RECT 27.160 122.050 27.480 122.110 ;
        RECT 31.875 121.910 32.165 121.955 ;
        RECT 32.680 121.910 33.000 121.970 ;
        RECT 33.230 121.955 33.370 122.110 ;
        RECT 33.600 122.050 33.920 122.110 ;
        RECT 31.875 121.770 33.000 121.910 ;
        RECT 31.875 121.725 32.165 121.770 ;
        RECT 32.680 121.710 33.000 121.770 ;
        RECT 33.155 121.725 33.445 121.955 ;
        RECT 34.445 121.910 34.585 122.450 ;
        RECT 39.135 122.450 40.820 122.590 ;
        RECT 39.135 122.405 39.425 122.450 ;
        RECT 40.500 122.390 40.820 122.450 ;
        RECT 47.875 122.590 48.165 122.635 ;
        RECT 49.240 122.590 49.560 122.650 ;
        RECT 47.875 122.450 49.560 122.590 ;
        RECT 47.875 122.405 48.165 122.450 ;
        RECT 49.240 122.390 49.560 122.450 ;
        RECT 49.715 122.590 50.005 122.635 ;
        RECT 50.160 122.590 50.480 122.650 ;
        RECT 49.715 122.450 50.480 122.590 ;
        RECT 49.715 122.405 50.005 122.450 ;
        RECT 39.580 122.295 39.900 122.310 ;
        RECT 39.580 122.065 40.185 122.295 ;
        RECT 40.975 122.250 41.265 122.295 ;
        RECT 47.400 122.250 47.720 122.310 ;
        RECT 40.975 122.110 47.720 122.250 ;
        RECT 40.975 122.065 41.265 122.110 ;
        RECT 39.580 122.050 39.900 122.065 ;
        RECT 41.050 121.910 41.190 122.065 ;
        RECT 47.400 122.050 47.720 122.110 ;
        RECT 34.445 121.770 41.190 121.910 ;
        RECT 46.035 121.910 46.325 121.955 ;
        RECT 49.790 121.910 49.930 122.405 ;
        RECT 50.160 122.390 50.480 122.450 ;
        RECT 69.955 122.590 70.245 122.635 ;
        RECT 73.620 122.590 73.940 122.650 ;
        RECT 69.955 122.450 73.940 122.590 ;
        RECT 69.955 122.405 70.245 122.450 ;
        RECT 73.620 122.390 73.940 122.450 ;
        RECT 75.015 122.590 75.305 122.635 ;
        RECT 77.760 122.590 78.080 122.650 ;
        RECT 75.015 122.450 78.080 122.590 ;
        RECT 75.015 122.405 75.305 122.450 ;
        RECT 77.760 122.390 78.080 122.450 ;
        RECT 83.755 122.590 84.045 122.635 ;
        RECT 86.500 122.590 86.820 122.650 ;
        RECT 83.755 122.450 86.820 122.590 ;
        RECT 83.755 122.405 84.045 122.450 ;
        RECT 86.500 122.390 86.820 122.450 ;
        RECT 88.800 122.390 89.120 122.650 ;
        RECT 94.320 122.590 94.640 122.650 ;
        RECT 112.260 122.590 112.580 122.650 ;
        RECT 119.620 122.590 119.940 122.650 ;
        RECT 123.300 122.590 123.620 122.650 ;
        RECT 125.140 122.590 125.460 122.650 ;
        RECT 94.320 122.450 112.580 122.590 ;
        RECT 94.320 122.390 94.640 122.450 ;
        RECT 112.260 122.390 112.580 122.450 ;
        RECT 118.790 122.450 119.940 122.590 ;
        RECT 54.300 122.250 54.620 122.310 ;
        RECT 55.280 122.250 55.570 122.295 ;
        RECT 66.720 122.250 67.040 122.310 ;
        RECT 85.120 122.250 85.440 122.310 ;
        RECT 95.240 122.250 95.560 122.310 ;
        RECT 118.790 122.250 118.930 122.450 ;
        RECT 119.620 122.390 119.940 122.450 ;
        RECT 122.010 122.450 125.460 122.590 ;
        RECT 122.010 122.295 122.150 122.450 ;
        RECT 123.300 122.390 123.620 122.450 ;
        RECT 125.140 122.390 125.460 122.450 ;
        RECT 130.200 122.590 130.520 122.650 ;
        RECT 135.260 122.590 135.580 122.650 ;
        RECT 130.200 122.450 135.580 122.590 ;
        RECT 130.200 122.390 130.520 122.450 ;
        RECT 135.260 122.390 135.580 122.450 ;
        RECT 140.780 122.390 141.100 122.650 ;
        RECT 121.015 122.250 121.305 122.295 ;
        RECT 54.300 122.110 55.570 122.250 ;
        RECT 54.300 122.050 54.620 122.110 ;
        RECT 55.280 122.065 55.570 122.110 ;
        RECT 56.690 122.110 67.040 122.250 ;
        RECT 56.690 121.955 56.830 122.110 ;
        RECT 66.720 122.050 67.040 122.110 ;
        RECT 67.270 122.110 95.560 122.250 ;
        RECT 46.035 121.770 49.930 121.910 ;
        RECT 46.035 121.725 46.325 121.770 ;
        RECT 56.615 121.725 56.905 121.955 ;
        RECT 60.280 121.910 60.600 121.970 ;
        RECT 63.055 121.910 63.345 121.955 ;
        RECT 67.270 121.910 67.410 122.110 ;
        RECT 85.120 122.050 85.440 122.110 ;
        RECT 95.240 122.050 95.560 122.110 ;
        RECT 97.630 122.110 118.930 122.250 ;
        RECT 119.250 122.110 121.305 122.250 ;
        RECT 97.630 121.970 97.770 122.110 ;
        RECT 60.280 121.770 67.410 121.910 ;
        RECT 68.100 121.910 68.420 121.970 ;
        RECT 69.495 121.910 69.785 121.955 ;
        RECT 68.100 121.770 69.785 121.910 ;
        RECT 60.280 121.710 60.600 121.770 ;
        RECT 63.055 121.725 63.345 121.770 ;
        RECT 68.100 121.710 68.420 121.770 ;
        RECT 69.495 121.725 69.785 121.770 ;
        RECT 70.415 121.725 70.705 121.955 ;
        RECT 72.255 121.725 72.545 121.955 ;
        RECT 28.565 121.570 28.855 121.615 ;
        RECT 31.085 121.570 31.375 121.615 ;
        RECT 32.275 121.570 32.565 121.615 ;
        RECT 28.565 121.430 32.565 121.570 ;
        RECT 28.565 121.385 28.855 121.430 ;
        RECT 31.085 121.385 31.375 121.430 ;
        RECT 32.275 121.385 32.565 121.430 ;
        RECT 45.560 121.370 45.880 121.630 ;
        RECT 52.025 121.570 52.315 121.615 ;
        RECT 54.545 121.570 54.835 121.615 ;
        RECT 55.735 121.570 56.025 121.615 ;
        RECT 52.025 121.430 56.025 121.570 ;
        RECT 52.025 121.385 52.315 121.430 ;
        RECT 54.545 121.385 54.835 121.430 ;
        RECT 55.735 121.385 56.025 121.430 ;
        RECT 29.000 121.230 29.290 121.275 ;
        RECT 30.570 121.230 30.860 121.275 ;
        RECT 32.670 121.230 32.960 121.275 ;
        RECT 29.000 121.090 32.960 121.230 ;
        RECT 29.000 121.045 29.290 121.090 ;
        RECT 30.570 121.045 30.860 121.090 ;
        RECT 32.670 121.045 32.960 121.090 ;
        RECT 52.460 121.230 52.750 121.275 ;
        RECT 54.030 121.230 54.320 121.275 ;
        RECT 56.130 121.230 56.420 121.275 ;
        RECT 52.460 121.090 56.420 121.230 ;
        RECT 70.490 121.230 70.630 121.725 ;
        RECT 72.330 121.570 72.470 121.725 ;
        RECT 73.160 121.710 73.480 121.970 ;
        RECT 74.080 121.710 74.400 121.970 ;
        RECT 75.000 121.710 75.320 121.970 ;
        RECT 83.295 121.725 83.585 121.955 ;
        RECT 80.520 121.570 80.840 121.630 ;
        RECT 83.370 121.570 83.510 121.725 ;
        RECT 84.660 121.710 84.980 121.970 ;
        RECT 86.040 121.710 86.360 121.970 ;
        RECT 90.655 121.910 90.945 121.955 ;
        RECT 97.540 121.910 97.860 121.970 ;
        RECT 90.655 121.770 97.860 121.910 ;
        RECT 90.655 121.725 90.945 121.770 ;
        RECT 97.540 121.710 97.860 121.770 ;
        RECT 103.535 121.910 103.825 121.955 ;
        RECT 106.740 121.910 107.060 121.970 ;
        RECT 118.330 121.955 118.470 122.110 ;
        RECT 119.250 121.955 119.390 122.110 ;
        RECT 121.015 122.065 121.305 122.110 ;
        RECT 121.935 122.065 122.225 122.295 ;
        RECT 122.855 122.250 123.145 122.295 ;
        RECT 128.360 122.250 128.680 122.310 ;
        RECT 122.855 122.110 128.680 122.250 ;
        RECT 122.855 122.065 123.145 122.110 ;
        RECT 128.360 122.050 128.680 122.110 ;
        RECT 103.535 121.770 107.060 121.910 ;
        RECT 103.535 121.725 103.825 121.770 ;
        RECT 106.740 121.710 107.060 121.770 ;
        RECT 118.255 121.725 118.545 121.955 ;
        RECT 118.715 121.725 119.005 121.955 ;
        RECT 119.175 121.725 119.465 121.955 ;
        RECT 120.095 121.910 120.385 121.955 ;
        RECT 123.760 121.910 124.080 121.970 ;
        RECT 128.820 121.910 129.140 121.970 ;
        RECT 120.095 121.770 122.380 121.910 ;
        RECT 120.095 121.725 120.385 121.770 ;
        RECT 72.330 121.430 83.510 121.570 ;
        RECT 80.520 121.370 80.840 121.430 ;
        RECT 72.240 121.230 72.560 121.290 ;
        RECT 70.490 121.090 72.560 121.230 ;
        RECT 52.460 121.045 52.750 121.090 ;
        RECT 54.030 121.045 54.320 121.090 ;
        RECT 56.130 121.045 56.420 121.090 ;
        RECT 72.240 121.030 72.560 121.090 ;
        RECT 40.040 120.690 40.360 120.950 ;
        RECT 72.700 120.690 73.020 120.950 ;
        RECT 83.370 120.890 83.510 121.430 ;
        RECT 90.180 121.570 90.500 121.630 ;
        RECT 91.115 121.570 91.405 121.615 ;
        RECT 90.180 121.430 91.405 121.570 ;
        RECT 90.180 121.370 90.500 121.430 ;
        RECT 91.115 121.385 91.405 121.430 ;
        RECT 91.560 121.370 91.880 121.630 ;
        RECT 103.980 121.370 104.300 121.630 ;
        RECT 104.915 121.570 105.205 121.615 ;
        RECT 107.200 121.570 107.520 121.630 ;
        RECT 104.915 121.430 107.520 121.570 ;
        RECT 118.790 121.570 118.930 121.725 ;
        RECT 121.460 121.570 121.780 121.630 ;
        RECT 118.790 121.430 121.780 121.570 ;
        RECT 122.240 121.570 122.380 121.770 ;
        RECT 123.760 121.770 129.140 121.910 ;
        RECT 123.760 121.710 124.080 121.770 ;
        RECT 128.820 121.710 129.140 121.770 ;
        RECT 129.740 121.710 130.060 121.970 ;
        RECT 130.290 121.955 130.430 122.390 ;
        RECT 132.055 122.250 132.345 122.295 ;
        RECT 133.740 122.250 134.030 122.295 ;
        RECT 132.055 122.110 134.030 122.250 ;
        RECT 132.055 122.065 132.345 122.110 ;
        RECT 133.740 122.065 134.030 122.110 ;
        RECT 130.215 121.725 130.505 121.955 ;
        RECT 130.660 121.910 130.980 121.970 ;
        RECT 132.960 121.910 133.280 121.970 ;
        RECT 139.875 121.910 140.165 121.955 ;
        RECT 130.660 121.770 133.280 121.910 ;
        RECT 130.660 121.710 130.980 121.770 ;
        RECT 132.960 121.710 133.280 121.770 ;
        RECT 139.490 121.770 140.165 121.910 ;
        RECT 123.850 121.570 123.990 121.710 ;
        RECT 132.515 121.570 132.805 121.615 ;
        RECT 122.240 121.430 123.990 121.570 ;
        RECT 131.210 121.430 132.805 121.570 ;
        RECT 104.915 121.385 105.205 121.430 ;
        RECT 107.200 121.370 107.520 121.430 ;
        RECT 121.460 121.370 121.780 121.430 ;
        RECT 131.210 121.290 131.350 121.430 ;
        RECT 132.515 121.385 132.805 121.430 ;
        RECT 133.395 121.570 133.685 121.615 ;
        RECT 134.585 121.570 134.875 121.615 ;
        RECT 137.105 121.570 137.395 121.615 ;
        RECT 133.395 121.430 137.395 121.570 ;
        RECT 133.395 121.385 133.685 121.430 ;
        RECT 134.585 121.385 134.875 121.430 ;
        RECT 137.105 121.385 137.395 121.430 ;
        RECT 111.800 121.230 112.120 121.290 ;
        RECT 113.180 121.230 113.500 121.290 ;
        RECT 130.660 121.230 130.980 121.290 ;
        RECT 111.800 121.090 130.980 121.230 ;
        RECT 111.800 121.030 112.120 121.090 ;
        RECT 113.180 121.030 113.500 121.090 ;
        RECT 130.660 121.030 130.980 121.090 ;
        RECT 131.120 121.030 131.440 121.290 ;
        RECT 133.000 121.230 133.290 121.275 ;
        RECT 135.100 121.230 135.390 121.275 ;
        RECT 136.670 121.230 136.960 121.275 ;
        RECT 133.000 121.090 136.960 121.230 ;
        RECT 133.000 121.045 133.290 121.090 ;
        RECT 135.100 121.045 135.390 121.090 ;
        RECT 136.670 121.045 136.960 121.090 ;
        RECT 85.135 120.890 85.425 120.935 ;
        RECT 83.370 120.750 85.425 120.890 ;
        RECT 85.135 120.705 85.425 120.750 ;
        RECT 87.435 120.890 87.725 120.935 ;
        RECT 93.860 120.890 94.180 120.950 ;
        RECT 87.435 120.750 94.180 120.890 ;
        RECT 87.435 120.705 87.725 120.750 ;
        RECT 93.860 120.690 94.180 120.750 ;
        RECT 101.220 120.890 101.540 120.950 ;
        RECT 101.695 120.890 101.985 120.935 ;
        RECT 101.220 120.750 101.985 120.890 ;
        RECT 101.220 120.690 101.540 120.750 ;
        RECT 101.695 120.705 101.985 120.750 ;
        RECT 116.860 120.690 117.180 120.950 ;
        RECT 136.180 120.890 136.500 120.950 ;
        RECT 139.490 120.935 139.630 121.770 ;
        RECT 139.875 121.725 140.165 121.770 ;
        RECT 139.415 120.890 139.705 120.935 ;
        RECT 136.180 120.750 139.705 120.890 ;
        RECT 136.180 120.690 136.500 120.750 ;
        RECT 139.415 120.705 139.705 120.750 ;
        RECT 17.430 120.070 143.010 120.550 ;
        RECT 73.160 119.870 73.480 119.930 ;
        RECT 75.475 119.870 75.765 119.915 ;
        RECT 73.160 119.730 75.765 119.870 ;
        RECT 73.160 119.670 73.480 119.730 ;
        RECT 75.475 119.685 75.765 119.730 ;
        RECT 80.075 119.870 80.365 119.915 ;
        RECT 82.820 119.870 83.140 119.930 ;
        RECT 80.075 119.730 83.140 119.870 ;
        RECT 80.075 119.685 80.365 119.730 ;
        RECT 82.820 119.670 83.140 119.730 ;
        RECT 84.660 119.870 84.980 119.930 ;
        RECT 85.595 119.870 85.885 119.915 ;
        RECT 84.660 119.730 85.885 119.870 ;
        RECT 84.660 119.670 84.980 119.730 ;
        RECT 85.595 119.685 85.885 119.730 ;
        RECT 106.740 119.670 107.060 119.930 ;
        RECT 119.620 119.870 119.940 119.930 ;
        RECT 133.895 119.870 134.185 119.915 ;
        RECT 119.620 119.730 134.185 119.870 ;
        RECT 119.620 119.670 119.940 119.730 ;
        RECT 133.895 119.685 134.185 119.730 ;
        RECT 140.780 119.670 141.100 119.930 ;
        RECT 68.100 119.190 68.420 119.250 ;
        RECT 61.290 119.050 68.420 119.190 ;
        RECT 82.910 119.190 83.050 119.670 ;
        RECT 87.895 119.530 88.185 119.575 ;
        RECT 100.340 119.530 100.630 119.575 ;
        RECT 102.440 119.530 102.730 119.575 ;
        RECT 104.010 119.530 104.300 119.575 ;
        RECT 87.895 119.390 91.790 119.530 ;
        RECT 87.895 119.345 88.185 119.390 ;
        RECT 91.650 119.235 91.790 119.390 ;
        RECT 100.340 119.390 104.300 119.530 ;
        RECT 100.340 119.345 100.630 119.390 ;
        RECT 102.440 119.345 102.730 119.390 ;
        RECT 104.010 119.345 104.300 119.390 ;
        RECT 116.900 119.530 117.190 119.575 ;
        RECT 119.000 119.530 119.290 119.575 ;
        RECT 120.570 119.530 120.860 119.575 ;
        RECT 116.900 119.390 120.860 119.530 ;
        RECT 116.900 119.345 117.190 119.390 ;
        RECT 119.000 119.345 119.290 119.390 ;
        RECT 120.570 119.345 120.860 119.390 ;
        RECT 123.300 119.330 123.620 119.590 ;
        RECT 82.910 119.050 85.350 119.190 ;
        RECT 27.160 118.850 27.480 118.910 ;
        RECT 29.935 118.850 30.225 118.895 ;
        RECT 31.315 118.850 31.605 118.895 ;
        RECT 27.160 118.710 31.605 118.850 ;
        RECT 27.160 118.650 27.480 118.710 ;
        RECT 29.935 118.665 30.225 118.710 ;
        RECT 31.315 118.665 31.605 118.710 ;
        RECT 35.440 118.850 35.760 118.910 ;
        RECT 61.290 118.895 61.430 119.050 ;
        RECT 68.100 118.990 68.420 119.050 ;
        RECT 35.440 118.710 43.950 118.850 ;
        RECT 35.440 118.650 35.760 118.710 ;
        RECT 43.810 118.170 43.950 118.710 ;
        RECT 60.295 118.665 60.585 118.895 ;
        RECT 61.215 118.665 61.505 118.895 ;
        RECT 63.975 118.850 64.265 118.895 ;
        RECT 66.720 118.850 67.040 118.910 ;
        RECT 63.975 118.710 67.040 118.850 ;
        RECT 63.975 118.665 64.265 118.710 ;
        RECT 60.370 118.510 60.510 118.665 ;
        RECT 66.720 118.650 67.040 118.710 ;
        RECT 78.680 118.650 79.000 118.910 ;
        RECT 80.520 118.850 80.840 118.910 ;
        RECT 82.375 118.850 82.665 118.895 ;
        RECT 80.520 118.710 82.665 118.850 ;
        RECT 80.520 118.650 80.840 118.710 ;
        RECT 82.375 118.665 82.665 118.710 ;
        RECT 83.295 118.850 83.585 118.895 ;
        RECT 84.660 118.850 84.980 118.910 ;
        RECT 85.210 118.895 85.350 119.050 ;
        RECT 91.575 119.005 91.865 119.235 ;
        RECT 100.735 119.190 101.025 119.235 ;
        RECT 101.925 119.190 102.215 119.235 ;
        RECT 104.445 119.190 104.735 119.235 ;
        RECT 100.735 119.050 104.735 119.190 ;
        RECT 100.735 119.005 101.025 119.050 ;
        RECT 101.925 119.005 102.215 119.050 ;
        RECT 104.445 119.005 104.735 119.050 ;
        RECT 110.880 118.990 111.200 119.250 ;
        RECT 116.400 118.990 116.720 119.250 ;
        RECT 117.295 119.190 117.585 119.235 ;
        RECT 118.485 119.190 118.775 119.235 ;
        RECT 121.005 119.190 121.295 119.235 ;
        RECT 135.720 119.190 136.040 119.250 ;
        RECT 117.295 119.050 121.295 119.190 ;
        RECT 117.295 119.005 117.585 119.050 ;
        RECT 118.485 119.005 118.775 119.050 ;
        RECT 121.005 119.005 121.295 119.050 ;
        RECT 134.890 119.050 136.040 119.190 ;
        RECT 83.295 118.710 84.980 118.850 ;
        RECT 83.295 118.665 83.585 118.710 ;
        RECT 67.180 118.510 67.500 118.570 ;
        RECT 60.370 118.370 67.500 118.510 ;
        RECT 67.180 118.310 67.500 118.370 ;
        RECT 74.080 118.510 74.400 118.570 ;
        RECT 79.915 118.510 80.205 118.555 ;
        RECT 74.080 118.370 80.205 118.510 ;
        RECT 74.080 118.310 74.400 118.370 ;
        RECT 79.915 118.325 80.205 118.370 ;
        RECT 60.280 118.170 60.600 118.230 ;
        RECT 43.810 118.030 60.600 118.170 ;
        RECT 60.280 117.970 60.600 118.030 ;
        RECT 60.755 118.170 61.045 118.215 ;
        RECT 61.660 118.170 61.980 118.230 ;
        RECT 60.755 118.030 61.980 118.170 ;
        RECT 60.755 117.985 61.045 118.030 ;
        RECT 61.660 117.970 61.980 118.030 ;
        RECT 79.140 117.970 79.460 118.230 ;
        RECT 80.610 118.170 80.750 118.650 ;
        RECT 80.995 118.510 81.285 118.555 ;
        RECT 83.370 118.510 83.510 118.665 ;
        RECT 84.660 118.650 84.980 118.710 ;
        RECT 85.135 118.665 85.425 118.895 ;
        RECT 86.515 118.665 86.805 118.895 ;
        RECT 86.590 118.510 86.730 118.665 ;
        RECT 99.840 118.650 100.160 118.910 ;
        RECT 101.220 118.895 101.540 118.910 ;
        RECT 101.190 118.850 101.540 118.895 ;
        RECT 101.025 118.710 101.540 118.850 ;
        RECT 101.190 118.665 101.540 118.710 ;
        RECT 101.220 118.650 101.540 118.665 ;
        RECT 103.980 118.850 104.300 118.910 ;
        RECT 105.820 118.850 106.140 118.910 ;
        RECT 103.980 118.710 112.950 118.850 ;
        RECT 103.980 118.650 104.300 118.710 ;
        RECT 105.820 118.650 106.140 118.710 ;
        RECT 80.995 118.370 83.510 118.510 ;
        RECT 83.830 118.370 86.730 118.510 ;
        RECT 87.880 118.510 88.200 118.570 ;
        RECT 90.180 118.510 90.500 118.570 ;
        RECT 90.655 118.510 90.945 118.555 ;
        RECT 87.880 118.370 90.945 118.510 ;
        RECT 80.995 118.325 81.285 118.370 ;
        RECT 83.830 118.170 83.970 118.370 ;
        RECT 87.880 118.310 88.200 118.370 ;
        RECT 90.180 118.310 90.500 118.370 ;
        RECT 90.655 118.325 90.945 118.370 ;
        RECT 99.380 118.510 99.700 118.570 ;
        RECT 109.975 118.510 110.265 118.555 ;
        RECT 112.275 118.510 112.565 118.555 ;
        RECT 99.380 118.370 108.810 118.510 ;
        RECT 99.380 118.310 99.700 118.370 ;
        RECT 80.610 118.030 83.970 118.170 ;
        RECT 84.215 118.170 84.505 118.215 ;
        RECT 85.120 118.170 85.440 118.230 ;
        RECT 84.215 118.030 85.440 118.170 ;
        RECT 84.215 117.985 84.505 118.030 ;
        RECT 85.120 117.970 85.440 118.030 ;
        RECT 88.800 117.970 89.120 118.230 ;
        RECT 91.115 118.170 91.405 118.215 ;
        RECT 94.320 118.170 94.640 118.230 ;
        RECT 91.115 118.030 94.640 118.170 ;
        RECT 91.115 117.985 91.405 118.030 ;
        RECT 94.320 117.970 94.640 118.030 ;
        RECT 108.120 117.970 108.440 118.230 ;
        RECT 108.670 118.170 108.810 118.370 ;
        RECT 109.975 118.370 112.565 118.510 ;
        RECT 112.810 118.510 112.950 118.710 ;
        RECT 115.020 118.650 115.340 118.910 ;
        RECT 116.860 118.850 117.180 118.910 ;
        RECT 117.695 118.850 117.985 118.895 ;
        RECT 116.860 118.710 117.985 118.850 ;
        RECT 116.860 118.650 117.180 118.710 ;
        RECT 117.695 118.665 117.985 118.710 ;
        RECT 132.040 118.850 132.360 118.910 ;
        RECT 134.890 118.895 135.030 119.050 ;
        RECT 135.720 118.990 136.040 119.050 ;
        RECT 134.815 118.850 135.105 118.895 ;
        RECT 132.040 118.710 135.105 118.850 ;
        RECT 132.040 118.650 132.360 118.710 ;
        RECT 134.815 118.665 135.105 118.710 ;
        RECT 135.275 118.850 135.565 118.895 ;
        RECT 136.180 118.850 136.500 118.910 ;
        RECT 135.275 118.710 136.500 118.850 ;
        RECT 135.275 118.665 135.565 118.710 ;
        RECT 136.180 118.650 136.500 118.710 ;
        RECT 136.655 118.850 136.945 118.895 ;
        RECT 137.560 118.850 137.880 118.910 ;
        RECT 136.655 118.710 137.880 118.850 ;
        RECT 136.655 118.665 136.945 118.710 ;
        RECT 137.560 118.650 137.880 118.710 ;
        RECT 138.035 118.665 138.325 118.895 ;
        RECT 124.220 118.510 124.540 118.570 ;
        RECT 131.580 118.510 131.900 118.570 ;
        RECT 112.810 118.370 131.900 118.510 ;
        RECT 109.975 118.325 110.265 118.370 ;
        RECT 112.275 118.325 112.565 118.370 ;
        RECT 124.220 118.310 124.540 118.370 ;
        RECT 131.580 118.310 131.900 118.370 ;
        RECT 133.880 118.510 134.200 118.570 ;
        RECT 135.735 118.510 136.025 118.555 ;
        RECT 133.880 118.370 136.025 118.510 ;
        RECT 133.880 118.310 134.200 118.370 ;
        RECT 135.735 118.325 136.025 118.370 ;
        RECT 110.435 118.170 110.725 118.215 ;
        RECT 118.240 118.170 118.560 118.230 ;
        RECT 108.670 118.030 118.560 118.170 ;
        RECT 110.435 117.985 110.725 118.030 ;
        RECT 118.240 117.970 118.560 118.030 ;
        RECT 129.280 118.170 129.600 118.230 ;
        RECT 138.110 118.170 138.250 118.665 ;
        RECT 139.860 118.650 140.180 118.910 ;
        RECT 129.280 118.030 138.250 118.170 ;
        RECT 129.280 117.970 129.600 118.030 ;
        RECT 138.940 117.970 139.260 118.230 ;
        RECT 17.430 117.350 143.010 117.830 ;
        RECT 109.975 116.965 110.265 117.195 ;
        RECT 122.395 117.150 122.685 117.195 ;
        RECT 123.760 117.150 124.080 117.210 ;
        RECT 122.395 117.010 124.080 117.150 ;
        RECT 122.395 116.965 122.685 117.010 ;
        RECT 20.720 116.810 21.040 116.870 ;
        RECT 28.395 116.810 28.685 116.855 ;
        RECT 20.720 116.670 28.685 116.810 ;
        RECT 20.720 116.610 21.040 116.670 ;
        RECT 28.395 116.625 28.685 116.670 ;
        RECT 29.475 116.625 29.765 116.855 ;
        RECT 70.830 116.810 71.120 116.855 ;
        RECT 72.700 116.810 73.020 116.870 ;
        RECT 61.750 116.670 66.950 116.810 ;
        RECT 24.860 116.130 25.180 116.190 ;
        RECT 29.550 116.130 29.690 116.625 ;
        RECT 61.750 116.515 61.890 116.670 ;
        RECT 66.810 116.530 66.950 116.670 ;
        RECT 70.830 116.670 73.020 116.810 ;
        RECT 70.830 116.625 71.120 116.670 ;
        RECT 72.700 116.610 73.020 116.670 ;
        RECT 84.215 116.810 84.505 116.855 ;
        RECT 87.420 116.810 87.740 116.870 ;
        RECT 84.215 116.670 87.740 116.810 ;
        RECT 84.215 116.625 84.505 116.670 ;
        RECT 87.420 116.610 87.740 116.670 ;
        RECT 88.310 116.810 88.600 116.855 ;
        RECT 88.800 116.810 89.120 116.870 ;
        RECT 88.310 116.670 89.120 116.810 ;
        RECT 88.310 116.625 88.600 116.670 ;
        RECT 88.800 116.610 89.120 116.670 ;
        RECT 93.860 116.810 94.180 116.870 ;
        RECT 101.190 116.810 101.480 116.855 ;
        RECT 108.120 116.810 108.440 116.870 ;
        RECT 93.860 116.670 98.230 116.810 ;
        RECT 93.860 116.610 94.180 116.670 ;
        RECT 63.040 116.515 63.360 116.530 ;
        RECT 32.235 116.285 32.525 116.515 ;
        RECT 61.675 116.285 61.965 116.515 ;
        RECT 63.010 116.470 63.360 116.515 ;
        RECT 62.845 116.330 63.360 116.470 ;
        RECT 63.010 116.285 63.360 116.330 ;
        RECT 24.860 115.990 29.690 116.130 ;
        RECT 24.860 115.930 25.180 115.990 ;
        RECT 26.700 115.790 27.020 115.850 ;
        RECT 32.310 115.790 32.450 116.285 ;
        RECT 63.040 116.270 63.360 116.285 ;
        RECT 66.720 116.470 67.040 116.530 ;
        RECT 69.495 116.470 69.785 116.515 ;
        RECT 66.720 116.330 69.785 116.470 ;
        RECT 66.720 116.270 67.040 116.330 ;
        RECT 69.495 116.285 69.785 116.330 ;
        RECT 85.580 116.470 85.900 116.530 ;
        RECT 86.975 116.470 87.265 116.515 ;
        RECT 85.580 116.330 87.265 116.470 ;
        RECT 87.510 116.470 87.650 116.610 ;
        RECT 97.095 116.470 97.385 116.515 ;
        RECT 87.510 116.330 97.385 116.470 ;
        RECT 85.580 116.270 85.900 116.330 ;
        RECT 86.975 116.285 87.265 116.330 ;
        RECT 97.095 116.285 97.385 116.330 ;
        RECT 58.455 116.130 58.745 116.175 ;
        RECT 59.820 116.130 60.140 116.190 ;
        RECT 58.455 115.990 60.140 116.130 ;
        RECT 58.455 115.945 58.745 115.990 ;
        RECT 59.820 115.930 60.140 115.990 ;
        RECT 62.555 116.130 62.845 116.175 ;
        RECT 63.745 116.130 64.035 116.175 ;
        RECT 66.265 116.130 66.555 116.175 ;
        RECT 62.555 115.990 66.555 116.130 ;
        RECT 62.555 115.945 62.845 115.990 ;
        RECT 63.745 115.945 64.035 115.990 ;
        RECT 66.265 115.945 66.555 115.990 ;
        RECT 70.375 116.130 70.665 116.175 ;
        RECT 71.565 116.130 71.855 116.175 ;
        RECT 74.085 116.130 74.375 116.175 ;
        RECT 76.855 116.130 77.145 116.175 ;
        RECT 70.375 115.990 74.375 116.130 ;
        RECT 70.375 115.945 70.665 115.990 ;
        RECT 71.565 115.945 71.855 115.990 ;
        RECT 74.085 115.945 74.375 115.990 ;
        RECT 76.470 115.990 77.145 116.130 ;
        RECT 36.360 115.790 36.680 115.850 ;
        RECT 26.700 115.650 36.680 115.790 ;
        RECT 26.700 115.590 27.020 115.650 ;
        RECT 36.360 115.590 36.680 115.650 ;
        RECT 62.160 115.790 62.450 115.835 ;
        RECT 64.260 115.790 64.550 115.835 ;
        RECT 65.830 115.790 66.120 115.835 ;
        RECT 62.160 115.650 66.120 115.790 ;
        RECT 62.160 115.605 62.450 115.650 ;
        RECT 64.260 115.605 64.550 115.650 ;
        RECT 65.830 115.605 66.120 115.650 ;
        RECT 69.980 115.790 70.270 115.835 ;
        RECT 72.080 115.790 72.370 115.835 ;
        RECT 73.650 115.790 73.940 115.835 ;
        RECT 69.980 115.650 73.940 115.790 ;
        RECT 69.980 115.605 70.270 115.650 ;
        RECT 72.080 115.605 72.370 115.650 ;
        RECT 73.650 115.605 73.940 115.650 ;
        RECT 76.470 115.510 76.610 115.990 ;
        RECT 76.855 115.945 77.145 115.990 ;
        RECT 84.660 115.930 84.980 116.190 ;
        RECT 85.120 115.930 85.440 116.190 ;
        RECT 87.855 116.130 88.145 116.175 ;
        RECT 89.045 116.130 89.335 116.175 ;
        RECT 91.565 116.130 91.855 116.175 ;
        RECT 94.320 116.130 94.640 116.190 ;
        RECT 98.090 116.175 98.230 116.670 ;
        RECT 101.190 116.670 108.440 116.810 ;
        RECT 110.050 116.810 110.190 116.965 ;
        RECT 123.760 116.950 124.080 117.010 ;
        RECT 112.260 116.810 112.580 116.870 ;
        RECT 110.050 116.670 112.580 116.810 ;
        RECT 101.190 116.625 101.480 116.670 ;
        RECT 108.120 116.610 108.440 116.670 ;
        RECT 112.260 116.610 112.580 116.670 ;
        RECT 106.740 116.470 107.060 116.530 ;
        RECT 108.595 116.470 108.885 116.515 ;
        RECT 106.740 116.330 108.885 116.470 ;
        RECT 106.740 116.270 107.060 116.330 ;
        RECT 108.595 116.285 108.885 116.330 ;
        RECT 110.435 116.470 110.725 116.515 ;
        RECT 112.720 116.470 113.040 116.530 ;
        RECT 110.435 116.330 113.040 116.470 ;
        RECT 110.435 116.285 110.725 116.330 ;
        RECT 112.720 116.270 113.040 116.330 ;
        RECT 121.460 116.270 121.780 116.530 ;
        RECT 123.850 116.470 123.990 116.950 ;
        RECT 130.675 116.810 130.965 116.855 ;
        RECT 132.360 116.810 132.650 116.855 ;
        RECT 130.675 116.670 132.650 116.810 ;
        RECT 130.675 116.625 130.965 116.670 ;
        RECT 132.360 116.625 132.650 116.670 ;
        RECT 127.455 116.470 127.745 116.515 ;
        RECT 123.850 116.330 127.745 116.470 ;
        RECT 127.455 116.285 127.745 116.330 ;
        RECT 128.360 116.270 128.680 116.530 ;
        RECT 128.835 116.285 129.125 116.515 ;
        RECT 129.295 116.470 129.585 116.515 ;
        RECT 130.200 116.470 130.520 116.530 ;
        RECT 129.295 116.330 130.520 116.470 ;
        RECT 129.295 116.285 129.585 116.330 ;
        RECT 87.855 115.990 91.855 116.130 ;
        RECT 87.855 115.945 88.145 115.990 ;
        RECT 89.045 115.945 89.335 115.990 ;
        RECT 91.565 115.945 91.855 115.990 ;
        RECT 93.950 115.990 94.640 116.130 ;
        RECT 93.950 115.835 94.090 115.990 ;
        RECT 94.320 115.930 94.640 115.990 ;
        RECT 97.555 115.945 97.845 116.175 ;
        RECT 98.015 115.945 98.305 116.175 ;
        RECT 87.460 115.790 87.750 115.835 ;
        RECT 89.560 115.790 89.850 115.835 ;
        RECT 91.130 115.790 91.420 115.835 ;
        RECT 87.460 115.650 91.420 115.790 ;
        RECT 87.460 115.605 87.750 115.650 ;
        RECT 89.560 115.605 89.850 115.650 ;
        RECT 91.130 115.605 91.420 115.650 ;
        RECT 93.875 115.605 94.165 115.835 ;
        RECT 94.780 115.790 95.100 115.850 ;
        RECT 97.630 115.790 97.770 115.945 ;
        RECT 99.840 115.930 100.160 116.190 ;
        RECT 100.735 116.130 101.025 116.175 ;
        RECT 101.925 116.130 102.215 116.175 ;
        RECT 104.445 116.130 104.735 116.175 ;
        RECT 100.735 115.990 104.735 116.130 ;
        RECT 100.735 115.945 101.025 115.990 ;
        RECT 101.925 115.945 102.215 115.990 ;
        RECT 104.445 115.945 104.735 115.990 ;
        RECT 108.135 116.130 108.425 116.175 ;
        RECT 115.020 116.130 115.340 116.190 ;
        RECT 108.135 115.990 115.340 116.130 ;
        RECT 108.135 115.945 108.425 115.990 ;
        RECT 100.340 115.790 100.630 115.835 ;
        RECT 102.440 115.790 102.730 115.835 ;
        RECT 104.010 115.790 104.300 115.835 ;
        RECT 94.780 115.650 98.230 115.790 ;
        RECT 94.780 115.590 95.100 115.650 ;
        RECT 25.780 115.450 26.100 115.510 ;
        RECT 27.635 115.450 27.925 115.495 ;
        RECT 25.780 115.310 27.925 115.450 ;
        RECT 25.780 115.250 26.100 115.310 ;
        RECT 27.635 115.265 27.925 115.310 ;
        RECT 28.540 115.250 28.860 115.510 ;
        RECT 29.000 115.450 29.320 115.510 ;
        RECT 35.900 115.450 36.220 115.510 ;
        RECT 44.640 115.450 44.960 115.510 ;
        RECT 29.000 115.310 44.960 115.450 ;
        RECT 29.000 115.250 29.320 115.310 ;
        RECT 35.900 115.250 36.220 115.310 ;
        RECT 44.640 115.250 44.960 115.310 ;
        RECT 61.215 115.450 61.505 115.495 ;
        RECT 67.180 115.450 67.500 115.510 ;
        RECT 61.215 115.310 67.500 115.450 ;
        RECT 61.215 115.265 61.505 115.310 ;
        RECT 67.180 115.250 67.500 115.310 ;
        RECT 68.575 115.450 68.865 115.495 ;
        RECT 72.700 115.450 73.020 115.510 ;
        RECT 68.575 115.310 73.020 115.450 ;
        RECT 68.575 115.265 68.865 115.310 ;
        RECT 72.700 115.250 73.020 115.310 ;
        RECT 76.380 115.250 76.700 115.510 ;
        RECT 80.075 115.450 80.365 115.495 ;
        RECT 80.520 115.450 80.840 115.510 ;
        RECT 80.075 115.310 80.840 115.450 ;
        RECT 80.075 115.265 80.365 115.310 ;
        RECT 80.520 115.250 80.840 115.310 ;
        RECT 82.360 115.250 82.680 115.510 ;
        RECT 94.320 115.450 94.640 115.510 ;
        RECT 95.255 115.450 95.545 115.495 ;
        RECT 94.320 115.310 95.545 115.450 ;
        RECT 98.090 115.450 98.230 115.650 ;
        RECT 100.340 115.650 104.300 115.790 ;
        RECT 100.340 115.605 100.630 115.650 ;
        RECT 102.440 115.605 102.730 115.650 ;
        RECT 104.010 115.605 104.300 115.650 ;
        RECT 106.755 115.790 107.045 115.835 ;
        RECT 108.210 115.790 108.350 115.945 ;
        RECT 115.020 115.930 115.340 115.990 ;
        RECT 121.920 116.130 122.240 116.190 ;
        RECT 128.910 116.130 129.050 116.285 ;
        RECT 130.200 116.270 130.520 116.330 ;
        RECT 131.120 116.270 131.440 116.530 ;
        RECT 121.920 115.990 129.050 116.130 ;
        RECT 132.015 116.130 132.305 116.175 ;
        RECT 133.205 116.130 133.495 116.175 ;
        RECT 135.725 116.130 136.015 116.175 ;
        RECT 132.015 115.990 136.015 116.130 ;
        RECT 121.920 115.930 122.240 115.990 ;
        RECT 132.015 115.945 132.305 115.990 ;
        RECT 133.205 115.945 133.495 115.990 ;
        RECT 135.725 115.945 136.015 115.990 ;
        RECT 108.580 115.790 108.900 115.850 ;
        RECT 106.755 115.650 108.900 115.790 ;
        RECT 106.755 115.605 107.045 115.650 ;
        RECT 108.580 115.590 108.900 115.650 ;
        RECT 131.620 115.790 131.910 115.835 ;
        RECT 133.720 115.790 134.010 115.835 ;
        RECT 135.290 115.790 135.580 115.835 ;
        RECT 131.620 115.650 135.580 115.790 ;
        RECT 131.620 115.605 131.910 115.650 ;
        RECT 133.720 115.605 134.010 115.650 ;
        RECT 135.290 115.605 135.580 115.650 ;
        RECT 100.760 115.450 101.080 115.510 ;
        RECT 111.800 115.450 112.120 115.510 ;
        RECT 98.090 115.310 112.120 115.450 ;
        RECT 94.320 115.250 94.640 115.310 ;
        RECT 95.255 115.265 95.545 115.310 ;
        RECT 100.760 115.250 101.080 115.310 ;
        RECT 111.800 115.250 112.120 115.310 ;
        RECT 114.100 115.450 114.420 115.510 ;
        RECT 115.940 115.450 116.260 115.510 ;
        RECT 114.100 115.310 116.260 115.450 ;
        RECT 114.100 115.250 114.420 115.310 ;
        RECT 115.940 115.250 116.260 115.310 ;
        RECT 138.020 115.250 138.340 115.510 ;
        RECT 17.430 114.630 143.010 115.110 ;
        RECT 20.275 114.430 20.565 114.475 ;
        RECT 21.640 114.430 21.960 114.490 ;
        RECT 29.460 114.430 29.780 114.490 ;
        RECT 39.120 114.430 39.440 114.490 ;
        RECT 44.180 114.430 44.500 114.490 ;
        RECT 61.660 114.430 61.980 114.490 ;
        RECT 76.380 114.430 76.700 114.490 ;
        RECT 78.235 114.430 78.525 114.475 ;
        RECT 20.275 114.290 38.890 114.430 ;
        RECT 20.275 114.245 20.565 114.290 ;
        RECT 21.640 114.230 21.960 114.290 ;
        RECT 23.020 114.090 23.310 114.135 ;
        RECT 24.590 114.090 24.880 114.135 ;
        RECT 26.690 114.090 26.980 114.135 ;
        RECT 23.020 113.950 26.980 114.090 ;
        RECT 23.020 113.905 23.310 113.950 ;
        RECT 24.590 113.905 24.880 113.950 ;
        RECT 26.690 113.905 26.980 113.950 ;
        RECT 22.585 113.750 22.875 113.795 ;
        RECT 25.105 113.750 25.395 113.795 ;
        RECT 26.295 113.750 26.585 113.795 ;
        RECT 22.585 113.610 26.585 113.750 ;
        RECT 22.585 113.565 22.875 113.610 ;
        RECT 25.105 113.565 25.395 113.610 ;
        RECT 26.295 113.565 26.585 113.610 ;
        RECT 25.780 113.455 26.100 113.470 ;
        RECT 25.780 113.410 26.130 113.455 ;
        RECT 26.700 113.410 27.020 113.470 ;
        RECT 27.710 113.455 27.850 114.290 ;
        RECT 29.460 114.230 29.780 114.290 ;
        RECT 29.920 114.090 30.240 114.150 ;
        RECT 29.920 113.950 38.430 114.090 ;
        RECT 29.920 113.890 30.240 113.950 ;
        RECT 27.175 113.410 27.465 113.455 ;
        RECT 25.780 113.270 26.295 113.410 ;
        RECT 26.700 113.270 27.465 113.410 ;
        RECT 25.780 113.225 26.130 113.270 ;
        RECT 25.780 113.210 26.100 113.225 ;
        RECT 26.700 113.210 27.020 113.270 ;
        RECT 27.175 113.225 27.465 113.270 ;
        RECT 27.635 113.225 27.925 113.455 ;
        RECT 29.015 113.225 29.305 113.455 ;
        RECT 32.235 113.410 32.525 113.455 ;
        RECT 35.440 113.410 35.760 113.470 ;
        RECT 38.290 113.455 38.430 113.950 ;
        RECT 38.750 113.750 38.890 114.290 ;
        RECT 39.120 114.290 44.500 114.430 ;
        RECT 39.120 114.230 39.440 114.290 ;
        RECT 44.180 114.230 44.500 114.290 ;
        RECT 56.690 114.290 61.980 114.430 ;
        RECT 41.420 113.890 41.740 114.150 ;
        RECT 41.895 113.905 42.185 114.135 ;
        RECT 42.800 114.090 43.120 114.150 ;
        RECT 45.115 114.090 45.405 114.135 ;
        RECT 42.800 113.950 45.405 114.090 ;
        RECT 41.510 113.750 41.650 113.890 ;
        RECT 38.750 113.610 41.650 113.750 ;
        RECT 41.970 113.750 42.110 113.905 ;
        RECT 42.800 113.890 43.120 113.950 ;
        RECT 45.115 113.905 45.405 113.950 ;
        RECT 47.860 114.090 48.180 114.150 ;
        RECT 51.540 114.090 51.860 114.150 ;
        RECT 47.860 113.950 51.860 114.090 ;
        RECT 47.860 113.890 48.180 113.950 ;
        RECT 51.540 113.890 51.860 113.950 ;
        RECT 44.640 113.750 44.960 113.810 ;
        RECT 45.575 113.750 45.865 113.795 ;
        RECT 41.970 113.610 46.715 113.750 ;
        RECT 38.750 113.455 38.890 113.610 ;
        RECT 44.640 113.550 44.960 113.610 ;
        RECT 45.575 113.565 45.865 113.610 ;
        RECT 32.235 113.270 35.760 113.410 ;
        RECT 32.235 113.225 32.525 113.270 ;
        RECT 29.090 113.070 29.230 113.225 ;
        RECT 35.440 113.210 35.760 113.270 ;
        RECT 38.215 113.225 38.505 113.455 ;
        RECT 38.675 113.225 38.965 113.455 ;
        RECT 39.120 113.210 39.440 113.470 ;
        RECT 40.500 113.410 40.820 113.470 ;
        RECT 40.500 113.270 43.950 113.410 ;
        RECT 40.500 113.210 40.820 113.270 ;
        RECT 34.980 113.070 35.300 113.130 ;
        RECT 29.090 112.930 35.300 113.070 ;
        RECT 34.980 112.870 35.300 112.930 ;
        RECT 36.360 112.870 36.680 113.130 ;
        RECT 37.295 113.070 37.585 113.115 ;
        RECT 39.580 113.070 39.900 113.130 ;
        RECT 37.295 112.930 39.900 113.070 ;
        RECT 37.295 112.885 37.585 112.930 ;
        RECT 39.580 112.870 39.900 112.930 ;
        RECT 40.040 112.870 40.360 113.130 ;
        RECT 41.420 113.070 41.740 113.130 ;
        RECT 43.275 113.070 43.565 113.115 ;
        RECT 41.420 112.930 43.565 113.070 ;
        RECT 43.810 113.070 43.950 113.270 ;
        RECT 44.180 113.210 44.500 113.470 ;
        RECT 46.020 113.410 46.340 113.470 ;
        RECT 46.575 113.455 46.715 113.610 ;
        RECT 56.690 113.455 56.830 114.290 ;
        RECT 61.660 114.230 61.980 114.290 ;
        RECT 73.940 114.290 78.525 114.430 ;
        RECT 57.995 113.905 58.285 114.135 ;
        RECT 58.940 114.090 59.230 114.135 ;
        RECT 61.040 114.090 61.330 114.135 ;
        RECT 62.610 114.090 62.900 114.135 ;
        RECT 58.940 113.950 62.900 114.090 ;
        RECT 58.940 113.905 59.230 113.950 ;
        RECT 61.040 113.905 61.330 113.950 ;
        RECT 62.610 113.905 62.900 113.950 ;
        RECT 58.070 113.750 58.210 113.905 ;
        RECT 59.335 113.750 59.625 113.795 ;
        RECT 60.525 113.750 60.815 113.795 ;
        RECT 63.045 113.750 63.335 113.795 ;
        RECT 58.070 113.610 59.130 113.750 ;
        RECT 44.730 113.270 46.340 113.410 ;
        RECT 44.730 113.070 44.870 113.270 ;
        RECT 46.020 113.210 46.340 113.270 ;
        RECT 46.500 113.225 46.790 113.455 ;
        RECT 56.615 113.225 56.905 113.455 ;
        RECT 58.440 113.210 58.760 113.470 ;
        RECT 43.810 112.930 44.870 113.070 ;
        RECT 57.995 113.070 58.285 113.115 ;
        RECT 58.990 113.070 59.130 113.610 ;
        RECT 59.335 113.610 63.335 113.750 ;
        RECT 59.335 113.565 59.625 113.610 ;
        RECT 60.525 113.565 60.815 113.610 ;
        RECT 63.045 113.565 63.335 113.610 ;
        RECT 72.700 113.550 73.020 113.810 ;
        RECT 73.300 113.750 73.590 113.795 ;
        RECT 73.940 113.750 74.080 114.290 ;
        RECT 76.380 114.230 76.700 114.290 ;
        RECT 78.235 114.245 78.525 114.290 ;
        RECT 80.060 114.230 80.380 114.490 ;
        RECT 94.780 114.230 95.100 114.490 ;
        RECT 106.740 114.430 107.060 114.490 ;
        RECT 109.055 114.430 109.345 114.475 ;
        RECT 124.695 114.430 124.985 114.475 ;
        RECT 106.740 114.290 109.345 114.430 ;
        RECT 106.740 114.230 107.060 114.290 ;
        RECT 109.055 114.245 109.345 114.290 ;
        RECT 116.030 114.290 124.985 114.430 ;
        RECT 88.380 114.090 88.670 114.135 ;
        RECT 90.480 114.090 90.770 114.135 ;
        RECT 92.050 114.090 92.340 114.135 ;
        RECT 88.380 113.950 92.340 114.090 ;
        RECT 88.380 113.905 88.670 113.950 ;
        RECT 90.480 113.905 90.770 113.950 ;
        RECT 92.050 113.905 92.340 113.950 ;
        RECT 73.300 113.610 74.080 113.750 ;
        RECT 77.775 113.750 78.065 113.795 ;
        RECT 85.580 113.750 85.900 113.810 ;
        RECT 87.895 113.750 88.185 113.795 ;
        RECT 77.775 113.610 83.510 113.750 ;
        RECT 73.300 113.565 73.590 113.610 ;
        RECT 77.775 113.565 78.065 113.610 ;
        RECT 69.480 113.410 69.800 113.470 ;
        RECT 70.875 113.410 71.165 113.455 ;
        RECT 69.480 113.270 71.165 113.410 ;
        RECT 72.790 113.410 72.930 113.550 ;
        RECT 77.850 113.410 77.990 113.565 ;
        RECT 72.790 113.270 77.990 113.410 ;
        RECT 69.480 113.210 69.800 113.270 ;
        RECT 70.875 113.225 71.165 113.270 ;
        RECT 78.235 113.225 78.525 113.455 ;
        RECT 79.155 113.410 79.445 113.455 ;
        RECT 80.060 113.410 80.380 113.470 ;
        RECT 79.155 113.270 80.380 113.410 ;
        RECT 79.155 113.225 79.445 113.270 ;
        RECT 59.680 113.070 59.970 113.115 ;
        RECT 57.995 112.930 58.670 113.070 ;
        RECT 58.990 112.930 59.970 113.070 ;
        RECT 41.420 112.870 41.740 112.930 ;
        RECT 43.275 112.885 43.565 112.930 ;
        RECT 57.995 112.885 58.285 112.930 ;
        RECT 28.095 112.730 28.385 112.775 ;
        RECT 29.000 112.730 29.320 112.790 ;
        RECT 28.095 112.590 29.320 112.730 ;
        RECT 28.095 112.545 28.385 112.590 ;
        RECT 29.000 112.530 29.320 112.590 ;
        RECT 29.935 112.730 30.225 112.775 ;
        RECT 35.440 112.730 35.760 112.790 ;
        RECT 29.935 112.590 35.760 112.730 ;
        RECT 29.935 112.545 30.225 112.590 ;
        RECT 35.440 112.530 35.760 112.590 ;
        RECT 40.500 112.730 40.820 112.790 ;
        RECT 42.815 112.730 43.105 112.775 ;
        RECT 45.560 112.730 45.880 112.790 ;
        RECT 40.500 112.590 45.880 112.730 ;
        RECT 40.500 112.530 40.820 112.590 ;
        RECT 42.815 112.545 43.105 112.590 ;
        RECT 45.560 112.530 45.880 112.590 ;
        RECT 57.060 112.530 57.380 112.790 ;
        RECT 58.530 112.730 58.670 112.930 ;
        RECT 59.680 112.885 59.970 112.930 ;
        RECT 64.420 113.070 64.740 113.130 ;
        RECT 65.815 113.070 66.105 113.115 ;
        RECT 64.420 112.930 66.105 113.070 ;
        RECT 64.420 112.870 64.740 112.930 ;
        RECT 65.815 112.885 66.105 112.930 ;
        RECT 72.255 113.070 72.545 113.115 ;
        RECT 78.310 113.070 78.450 113.225 ;
        RECT 80.060 113.210 80.380 113.270 ;
        RECT 80.980 113.410 81.300 113.470 ;
        RECT 83.370 113.455 83.510 113.610 ;
        RECT 85.580 113.610 88.185 113.750 ;
        RECT 85.580 113.550 85.900 113.610 ;
        RECT 87.895 113.565 88.185 113.610 ;
        RECT 88.775 113.750 89.065 113.795 ;
        RECT 89.965 113.750 90.255 113.795 ;
        RECT 92.485 113.750 92.775 113.795 ;
        RECT 88.775 113.610 92.775 113.750 ;
        RECT 88.775 113.565 89.065 113.610 ;
        RECT 89.965 113.565 90.255 113.610 ;
        RECT 92.485 113.565 92.775 113.610 ;
        RECT 100.300 113.750 100.620 113.810 ;
        RECT 109.960 113.750 110.280 113.810 ;
        RECT 114.560 113.750 114.880 113.810 ;
        RECT 100.300 113.610 114.880 113.750 ;
        RECT 100.300 113.550 100.620 113.610 ;
        RECT 109.960 113.550 110.280 113.610 ;
        RECT 114.560 113.550 114.880 113.610 ;
        RECT 82.375 113.410 82.665 113.455 ;
        RECT 80.980 113.270 82.665 113.410 ;
        RECT 80.980 113.210 81.300 113.270 ;
        RECT 82.375 113.225 82.665 113.270 ;
        RECT 83.295 113.225 83.585 113.455 ;
        RECT 89.230 113.410 89.520 113.455 ;
        RECT 94.320 113.410 94.640 113.470 ;
        RECT 89.230 113.270 94.640 113.410 ;
        RECT 89.230 113.225 89.520 113.270 ;
        RECT 94.320 113.210 94.640 113.270 ;
        RECT 106.755 113.410 107.045 113.455 ;
        RECT 108.580 113.410 108.900 113.470 ;
        RECT 114.100 113.410 114.420 113.470 ;
        RECT 115.035 113.410 115.325 113.455 ;
        RECT 106.755 113.270 109.270 113.410 ;
        RECT 106.755 113.225 107.045 113.270 ;
        RECT 108.580 113.210 108.900 113.270 ;
        RECT 79.600 113.070 79.920 113.130 ;
        RECT 82.835 113.070 83.125 113.115 ;
        RECT 72.255 112.930 76.610 113.070 ;
        RECT 78.310 112.930 83.125 113.070 ;
        RECT 72.255 112.885 72.545 112.930 ;
        RECT 63.040 112.730 63.360 112.790 ;
        RECT 58.530 112.590 63.360 112.730 ;
        RECT 63.040 112.530 63.360 112.590 ;
        RECT 65.355 112.730 65.645 112.775 ;
        RECT 68.100 112.730 68.420 112.790 ;
        RECT 65.355 112.590 68.420 112.730 ;
        RECT 65.355 112.545 65.645 112.590 ;
        RECT 68.100 112.530 68.420 112.590 ;
        RECT 68.560 112.730 68.880 112.790 ;
        RECT 73.620 112.730 73.940 112.790 ;
        RECT 68.560 112.590 73.940 112.730 ;
        RECT 68.560 112.530 68.880 112.590 ;
        RECT 73.620 112.530 73.940 112.590 ;
        RECT 74.080 112.530 74.400 112.790 ;
        RECT 74.540 112.530 74.860 112.790 ;
        RECT 76.470 112.730 76.610 112.930 ;
        RECT 79.600 112.870 79.920 112.930 ;
        RECT 82.835 112.885 83.125 112.930 ;
        RECT 105.360 113.070 105.680 113.130 ;
        RECT 109.130 113.115 109.270 113.270 ;
        RECT 114.100 113.270 115.325 113.410 ;
        RECT 114.100 113.210 114.420 113.270 ;
        RECT 115.035 113.225 115.325 113.270 ;
        RECT 115.480 113.210 115.800 113.470 ;
        RECT 116.030 113.455 116.170 114.290 ;
        RECT 124.695 114.245 124.985 114.290 ;
        RECT 128.360 114.430 128.680 114.490 ;
        RECT 135.735 114.430 136.025 114.475 ;
        RECT 128.360 114.290 136.025 114.430 ;
        RECT 128.360 114.230 128.680 114.290 ;
        RECT 135.735 114.245 136.025 114.290 ;
        RECT 117.820 114.090 118.110 114.135 ;
        RECT 119.920 114.090 120.210 114.135 ;
        RECT 121.490 114.090 121.780 114.135 ;
        RECT 117.820 113.950 121.780 114.090 ;
        RECT 117.820 113.905 118.110 113.950 ;
        RECT 119.920 113.905 120.210 113.950 ;
        RECT 121.490 113.905 121.780 113.950 ;
        RECT 122.380 114.090 122.700 114.150 ;
        RECT 124.235 114.090 124.525 114.135 ;
        RECT 126.060 114.090 126.380 114.150 ;
        RECT 133.880 114.090 134.200 114.150 ;
        RECT 122.380 113.950 125.830 114.090 ;
        RECT 122.380 113.890 122.700 113.950 ;
        RECT 124.235 113.905 124.525 113.950 ;
        RECT 116.400 113.750 116.720 113.810 ;
        RECT 117.335 113.750 117.625 113.795 ;
        RECT 116.400 113.610 117.625 113.750 ;
        RECT 116.400 113.550 116.720 113.610 ;
        RECT 117.335 113.565 117.625 113.610 ;
        RECT 118.215 113.750 118.505 113.795 ;
        RECT 119.405 113.750 119.695 113.795 ;
        RECT 121.925 113.750 122.215 113.795 ;
        RECT 118.215 113.610 122.215 113.750 ;
        RECT 118.215 113.565 118.505 113.610 ;
        RECT 119.405 113.565 119.695 113.610 ;
        RECT 121.925 113.565 122.215 113.610 ;
        RECT 115.955 113.225 116.245 113.455 ;
        RECT 116.875 113.410 117.165 113.455 ;
        RECT 123.760 113.410 124.080 113.470 ;
        RECT 125.690 113.455 125.830 113.950 ;
        RECT 126.060 113.950 134.200 114.090 ;
        RECT 126.060 113.890 126.380 113.950 ;
        RECT 133.880 113.890 134.200 113.950 ;
        RECT 128.820 113.750 129.140 113.810 ;
        RECT 138.020 113.750 138.340 113.810 ;
        RECT 128.820 113.610 133.605 113.750 ;
        RECT 128.820 113.550 129.140 113.610 ;
        RECT 116.875 113.270 124.080 113.410 ;
        RECT 116.875 113.225 117.165 113.270 ;
        RECT 123.760 113.210 124.080 113.270 ;
        RECT 125.615 113.410 125.905 113.455 ;
        RECT 129.280 113.410 129.600 113.470 ;
        RECT 125.615 113.270 129.600 113.410 ;
        RECT 133.465 113.410 133.605 113.610 ;
        RECT 134.890 113.610 138.340 113.750 ;
        RECT 134.890 113.455 135.030 113.610 ;
        RECT 138.020 113.550 138.340 113.610 ;
        RECT 133.895 113.410 134.185 113.455 ;
        RECT 133.465 113.270 134.185 113.410 ;
        RECT 125.615 113.225 125.905 113.270 ;
        RECT 129.280 113.210 129.600 113.270 ;
        RECT 133.895 113.225 134.185 113.270 ;
        RECT 134.815 113.225 135.105 113.455 ;
        RECT 135.350 113.270 138.250 113.410 ;
        RECT 108.135 113.070 108.425 113.115 ;
        RECT 105.360 112.930 108.425 113.070 ;
        RECT 105.360 112.870 105.680 112.930 ;
        RECT 108.135 112.885 108.425 112.930 ;
        RECT 109.055 112.885 109.345 113.115 ;
        RECT 113.655 113.070 113.945 113.115 ;
        RECT 118.560 113.070 118.850 113.115 ;
        RECT 113.655 112.930 118.850 113.070 ;
        RECT 113.655 112.885 113.945 112.930 ;
        RECT 118.560 112.885 118.850 112.930 ;
        RECT 126.520 112.870 126.840 113.130 ;
        RECT 135.350 113.070 135.490 113.270 ;
        RECT 130.290 112.930 135.490 113.070 ;
        RECT 78.220 112.730 78.540 112.790 ;
        RECT 76.470 112.590 78.540 112.730 ;
        RECT 78.220 112.530 78.540 112.590 ;
        RECT 106.295 112.730 106.585 112.775 ;
        RECT 107.200 112.730 107.520 112.790 ;
        RECT 106.295 112.590 107.520 112.730 ;
        RECT 106.295 112.545 106.585 112.590 ;
        RECT 107.200 112.530 107.520 112.590 ;
        RECT 109.975 112.730 110.265 112.775 ;
        RECT 119.620 112.730 119.940 112.790 ;
        RECT 109.975 112.590 119.940 112.730 ;
        RECT 126.610 112.730 126.750 112.870 ;
        RECT 130.290 112.730 130.430 112.930 ;
        RECT 137.100 112.870 137.420 113.130 ;
        RECT 138.110 113.115 138.250 113.270 ;
        RECT 139.860 113.210 140.180 113.470 ;
        RECT 138.035 113.070 138.325 113.115 ;
        RECT 138.480 113.070 138.800 113.130 ;
        RECT 138.035 112.930 138.800 113.070 ;
        RECT 138.035 112.885 138.325 112.930 ;
        RECT 138.480 112.870 138.800 112.930 ;
        RECT 126.610 112.590 130.430 112.730 ;
        RECT 134.340 112.730 134.660 112.790 ;
        RECT 136.195 112.730 136.485 112.775 ;
        RECT 134.340 112.590 136.485 112.730 ;
        RECT 109.975 112.545 110.265 112.590 ;
        RECT 119.620 112.530 119.940 112.590 ;
        RECT 134.340 112.530 134.660 112.590 ;
        RECT 136.195 112.545 136.485 112.590 ;
        RECT 140.780 112.530 141.100 112.790 ;
        RECT 17.430 111.910 143.010 112.390 ;
        RECT 20.720 111.510 21.040 111.770 ;
        RECT 24.860 111.510 25.180 111.770 ;
        RECT 25.795 111.710 26.085 111.755 ;
        RECT 35.455 111.710 35.745 111.755 ;
        RECT 40.960 111.710 41.280 111.770 ;
        RECT 25.795 111.570 27.850 111.710 ;
        RECT 25.795 111.525 26.085 111.570 ;
        RECT 21.640 111.170 21.960 111.430 ;
        RECT 22.575 111.370 22.865 111.415 ;
        RECT 27.160 111.370 27.480 111.430 ;
        RECT 22.575 111.230 27.480 111.370 ;
        RECT 22.575 111.185 22.865 111.230 ;
        RECT 27.160 111.170 27.480 111.230 ;
        RECT 26.700 111.030 27.020 111.090 ;
        RECT 27.710 111.075 27.850 111.570 ;
        RECT 35.455 111.570 41.280 111.710 ;
        RECT 35.455 111.525 35.745 111.570 ;
        RECT 40.960 111.510 41.280 111.570 ;
        RECT 42.800 111.510 43.120 111.770 ;
        RECT 55.680 111.710 56.000 111.770 ;
        RECT 52.550 111.570 56.000 111.710 ;
        RECT 28.080 111.370 28.400 111.430 ;
        RECT 29.920 111.370 30.240 111.430 ;
        RECT 28.080 111.230 30.240 111.370 ;
        RECT 28.080 111.170 28.400 111.230 ;
        RECT 29.920 111.170 30.240 111.230 ;
        RECT 34.520 111.170 34.840 111.430 ;
        RECT 38.200 111.370 38.520 111.430 ;
        RECT 38.200 111.230 42.570 111.370 ;
        RECT 38.200 111.170 38.520 111.230 ;
        RECT 26.330 110.890 27.020 111.030 ;
        RECT 23.035 110.690 23.325 110.735 ;
        RECT 25.780 110.690 26.100 110.750 ;
        RECT 26.330 110.735 26.470 110.890 ;
        RECT 26.700 110.830 27.020 110.890 ;
        RECT 27.590 110.845 27.880 111.075 ;
        RECT 33.615 111.030 33.905 111.075 ;
        RECT 31.390 110.890 33.905 111.030 ;
        RECT 23.035 110.550 26.100 110.690 ;
        RECT 23.035 110.505 23.325 110.550 ;
        RECT 25.780 110.490 26.100 110.550 ;
        RECT 26.255 110.505 26.545 110.735 ;
        RECT 27.135 110.690 27.425 110.735 ;
        RECT 28.325 110.690 28.615 110.735 ;
        RECT 30.845 110.690 31.135 110.735 ;
        RECT 27.135 110.550 31.135 110.690 ;
        RECT 27.135 110.505 27.425 110.550 ;
        RECT 28.325 110.505 28.615 110.550 ;
        RECT 30.845 110.505 31.135 110.550 ;
        RECT 26.330 110.350 26.470 110.505 ;
        RECT 24.490 110.210 26.470 110.350 ;
        RECT 26.740 110.350 27.030 110.395 ;
        RECT 28.840 110.350 29.130 110.395 ;
        RECT 30.410 110.350 30.700 110.395 ;
        RECT 26.740 110.210 30.700 110.350 ;
        RECT 21.640 110.010 21.960 110.070 ;
        RECT 24.490 110.010 24.630 110.210 ;
        RECT 26.740 110.165 27.030 110.210 ;
        RECT 28.840 110.165 29.130 110.210 ;
        RECT 30.410 110.165 30.700 110.210 ;
        RECT 21.640 109.870 24.630 110.010 ;
        RECT 24.875 110.010 25.165 110.055 ;
        RECT 27.620 110.010 27.940 110.070 ;
        RECT 24.875 109.870 27.940 110.010 ;
        RECT 21.640 109.810 21.960 109.870 ;
        RECT 24.875 109.825 25.165 109.870 ;
        RECT 27.620 109.810 27.940 109.870 ;
        RECT 28.080 110.010 28.400 110.070 ;
        RECT 30.840 110.010 31.160 110.070 ;
        RECT 31.390 110.010 31.530 110.890 ;
        RECT 33.615 110.845 33.905 110.890 ;
        RECT 35.900 110.830 36.220 111.090 ;
        RECT 37.250 111.030 37.540 111.075 ;
        RECT 40.040 111.030 40.360 111.090 ;
        RECT 37.250 110.890 40.360 111.030 ;
        RECT 37.250 110.845 37.540 110.890 ;
        RECT 40.040 110.830 40.360 110.890 ;
        RECT 36.795 110.690 37.085 110.735 ;
        RECT 37.985 110.690 38.275 110.735 ;
        RECT 40.505 110.690 40.795 110.735 ;
        RECT 36.795 110.550 40.795 110.690 ;
        RECT 36.795 110.505 37.085 110.550 ;
        RECT 37.985 110.505 38.275 110.550 ;
        RECT 40.505 110.505 40.795 110.550 ;
        RECT 36.400 110.350 36.690 110.395 ;
        RECT 38.500 110.350 38.790 110.395 ;
        RECT 40.070 110.350 40.360 110.395 ;
        RECT 36.400 110.210 40.360 110.350 ;
        RECT 42.430 110.350 42.570 111.230 ;
        RECT 42.890 111.030 43.030 111.510 ;
        RECT 48.780 111.370 49.100 111.430 ;
        RECT 52.550 111.415 52.690 111.570 ;
        RECT 55.680 111.510 56.000 111.570 ;
        RECT 57.060 111.710 57.380 111.770 ;
        RECT 57.060 111.570 68.330 111.710 ;
        RECT 57.060 111.510 57.380 111.570 ;
        RECT 51.555 111.370 51.845 111.415 ;
        RECT 48.780 111.230 51.845 111.370 ;
        RECT 48.780 111.170 49.100 111.230 ;
        RECT 51.555 111.185 51.845 111.230 ;
        RECT 52.475 111.185 52.765 111.415 ;
        RECT 53.010 111.230 54.990 111.370 ;
        RECT 53.010 111.075 53.150 111.230 ;
        RECT 44.655 111.030 44.945 111.075 ;
        RECT 46.495 111.030 46.785 111.075 ;
        RECT 42.890 110.890 46.785 111.030 ;
        RECT 44.655 110.845 44.945 110.890 ;
        RECT 46.495 110.845 46.785 110.890 ;
        RECT 47.415 110.845 47.705 111.075 ;
        RECT 51.095 110.845 51.385 111.075 ;
        RECT 52.935 110.845 53.225 111.075 ;
        RECT 54.215 111.030 54.505 111.075 ;
        RECT 53.470 110.890 54.505 111.030 ;
        RECT 54.850 111.030 54.990 111.230 ;
        RECT 60.280 111.170 60.600 111.430 ;
        RECT 68.190 111.370 68.330 111.570 ;
        RECT 68.560 111.510 68.880 111.770 ;
        RECT 69.480 111.710 69.800 111.770 ;
        RECT 75.460 111.710 75.780 111.770 ;
        RECT 80.980 111.710 81.300 111.770 ;
        RECT 69.480 111.570 75.780 111.710 ;
        RECT 69.480 111.510 69.800 111.570 ;
        RECT 75.460 111.510 75.780 111.570 ;
        RECT 80.610 111.570 81.300 111.710 ;
        RECT 72.240 111.370 72.560 111.430 ;
        RECT 76.855 111.370 77.145 111.415 ;
        RECT 80.610 111.370 80.750 111.570 ;
        RECT 80.980 111.510 81.300 111.570 ;
        RECT 104.455 111.525 104.745 111.755 ;
        RECT 110.895 111.710 111.185 111.755 ;
        RECT 113.180 111.710 113.500 111.770 ;
        RECT 110.895 111.570 113.500 111.710 ;
        RECT 110.895 111.525 111.185 111.570 ;
        RECT 82.820 111.370 83.140 111.430 ;
        RECT 85.580 111.370 85.900 111.430 ;
        RECT 92.035 111.370 92.325 111.415 ;
        RECT 98.935 111.370 99.225 111.415 ;
        RECT 99.840 111.370 100.160 111.430 ;
        RECT 68.190 111.230 77.145 111.370 ;
        RECT 72.240 111.170 72.560 111.230 ;
        RECT 76.855 111.185 77.145 111.230 ;
        RECT 78.770 111.230 80.750 111.370 ;
        RECT 81.070 111.230 100.160 111.370 ;
        RECT 58.440 111.030 58.760 111.090 ;
        RECT 69.495 111.030 69.785 111.075 ;
        RECT 54.850 110.890 69.785 111.030 ;
        RECT 46.020 110.490 46.340 110.750 ;
        RECT 47.490 110.350 47.630 110.845 ;
        RECT 51.170 110.690 51.310 110.845 ;
        RECT 52.000 110.690 52.320 110.750 ;
        RECT 53.470 110.690 53.610 110.890 ;
        RECT 54.215 110.845 54.505 110.890 ;
        RECT 58.440 110.830 58.760 110.890 ;
        RECT 64.510 110.750 64.650 110.890 ;
        RECT 69.495 110.845 69.785 110.890 ;
        RECT 69.940 111.030 70.260 111.090 ;
        RECT 70.775 111.030 71.065 111.075 ;
        RECT 77.775 111.030 78.065 111.075 ;
        RECT 69.940 110.890 71.065 111.030 ;
        RECT 69.940 110.830 70.260 110.890 ;
        RECT 70.775 110.845 71.065 110.890 ;
        RECT 76.470 110.890 78.065 111.030 ;
        RECT 51.170 110.550 52.320 110.690 ;
        RECT 52.000 110.490 52.320 110.550 ;
        RECT 52.550 110.550 53.610 110.690 ;
        RECT 53.815 110.690 54.105 110.735 ;
        RECT 55.005 110.690 55.295 110.735 ;
        RECT 57.525 110.690 57.815 110.735 ;
        RECT 53.815 110.550 57.815 110.690 ;
        RECT 52.550 110.395 52.690 110.550 ;
        RECT 53.815 110.505 54.105 110.550 ;
        RECT 55.005 110.505 55.295 110.550 ;
        RECT 57.525 110.505 57.815 110.550 ;
        RECT 64.420 110.490 64.740 110.750 ;
        RECT 65.815 110.690 66.105 110.735 ;
        RECT 68.100 110.690 68.420 110.750 ;
        RECT 65.815 110.550 68.420 110.690 ;
        RECT 65.815 110.505 66.105 110.550 ;
        RECT 68.100 110.490 68.420 110.550 ;
        RECT 70.375 110.690 70.665 110.735 ;
        RECT 71.565 110.690 71.855 110.735 ;
        RECT 74.085 110.690 74.375 110.735 ;
        RECT 70.375 110.550 74.375 110.690 ;
        RECT 70.375 110.505 70.665 110.550 ;
        RECT 71.565 110.505 71.855 110.550 ;
        RECT 74.085 110.505 74.375 110.550 ;
        RECT 42.430 110.210 47.630 110.350 ;
        RECT 36.400 110.165 36.690 110.210 ;
        RECT 38.500 110.165 38.790 110.210 ;
        RECT 40.070 110.165 40.360 110.210 ;
        RECT 52.475 110.165 52.765 110.395 ;
        RECT 53.420 110.350 53.710 110.395 ;
        RECT 55.520 110.350 55.810 110.395 ;
        RECT 57.090 110.350 57.380 110.395 ;
        RECT 53.420 110.210 57.380 110.350 ;
        RECT 53.420 110.165 53.710 110.210 ;
        RECT 55.520 110.165 55.810 110.210 ;
        RECT 57.090 110.165 57.380 110.210 ;
        RECT 59.820 110.150 60.140 110.410 ;
        RECT 63.040 110.350 63.360 110.410 ;
        RECT 69.980 110.350 70.270 110.395 ;
        RECT 72.080 110.350 72.370 110.395 ;
        RECT 73.650 110.350 73.940 110.395 ;
        RECT 63.040 110.210 69.250 110.350 ;
        RECT 63.040 110.150 63.360 110.210 ;
        RECT 28.080 109.870 31.530 110.010 ;
        RECT 33.155 110.010 33.445 110.055 ;
        RECT 34.980 110.010 35.300 110.070 ;
        RECT 39.120 110.010 39.440 110.070 ;
        RECT 33.155 109.870 39.440 110.010 ;
        RECT 28.080 109.810 28.400 109.870 ;
        RECT 30.840 109.810 31.160 109.870 ;
        RECT 33.155 109.825 33.445 109.870 ;
        RECT 34.980 109.810 35.300 109.870 ;
        RECT 39.120 109.810 39.440 109.870 ;
        RECT 43.720 109.810 44.040 110.070 ;
        RECT 44.180 110.010 44.500 110.070 ;
        RECT 45.575 110.010 45.865 110.055 ;
        RECT 46.020 110.010 46.340 110.070 ;
        RECT 44.180 109.870 46.340 110.010 ;
        RECT 44.180 109.810 44.500 109.870 ;
        RECT 45.575 109.825 45.865 109.870 ;
        RECT 46.020 109.810 46.340 109.870 ;
        RECT 48.320 109.810 48.640 110.070 ;
        RECT 69.110 110.010 69.250 110.210 ;
        RECT 69.980 110.210 73.940 110.350 ;
        RECT 69.980 110.165 70.270 110.210 ;
        RECT 72.080 110.165 72.370 110.210 ;
        RECT 73.650 110.165 73.940 110.210 ;
        RECT 70.860 110.010 71.180 110.070 ;
        RECT 69.110 109.870 71.180 110.010 ;
        RECT 70.860 109.810 71.180 109.870 ;
        RECT 72.700 110.010 73.020 110.070 ;
        RECT 74.080 110.010 74.400 110.070 ;
        RECT 72.700 109.870 74.400 110.010 ;
        RECT 72.700 109.810 73.020 109.870 ;
        RECT 74.080 109.810 74.400 109.870 ;
        RECT 75.460 110.010 75.780 110.070 ;
        RECT 76.470 110.055 76.610 110.890 ;
        RECT 77.775 110.845 78.065 110.890 ;
        RECT 78.220 111.030 78.540 111.090 ;
        RECT 78.770 111.075 78.910 111.230 ;
        RECT 78.695 111.030 78.985 111.075 ;
        RECT 78.220 110.890 78.985 111.030 ;
        RECT 77.850 110.690 77.990 110.845 ;
        RECT 78.220 110.830 78.540 110.890 ;
        RECT 78.695 110.845 78.985 110.890 ;
        RECT 79.155 110.845 79.445 111.075 ;
        RECT 79.230 110.690 79.370 110.845 ;
        RECT 79.600 110.830 79.920 111.090 ;
        RECT 81.070 111.075 81.210 111.230 ;
        RECT 82.820 111.170 83.140 111.230 ;
        RECT 85.580 111.170 85.900 111.230 ;
        RECT 92.035 111.185 92.325 111.230 ;
        RECT 98.935 111.185 99.225 111.230 ;
        RECT 99.840 111.170 100.160 111.230 ;
        RECT 100.775 111.370 101.065 111.415 ;
        RECT 101.220 111.370 101.540 111.430 ;
        RECT 103.980 111.370 104.300 111.430 ;
        RECT 100.775 111.230 104.300 111.370 ;
        RECT 100.775 111.185 101.065 111.230 ;
        RECT 101.220 111.170 101.540 111.230 ;
        RECT 103.980 111.170 104.300 111.230 ;
        RECT 82.360 111.075 82.680 111.090 ;
        RECT 80.995 110.845 81.285 111.075 ;
        RECT 82.330 111.030 82.680 111.075 ;
        RECT 82.165 110.890 82.680 111.030 ;
        RECT 82.330 110.845 82.680 110.890 ;
        RECT 82.360 110.830 82.680 110.845 ;
        RECT 84.660 111.030 84.980 111.090 ;
        RECT 84.660 110.890 88.110 111.030 ;
        RECT 84.660 110.830 84.980 110.890 ;
        RECT 80.060 110.690 80.380 110.750 ;
        RECT 77.850 110.550 80.380 110.690 ;
        RECT 80.060 110.490 80.380 110.550 ;
        RECT 80.520 110.490 80.840 110.750 ;
        RECT 81.875 110.690 82.165 110.735 ;
        RECT 83.065 110.690 83.355 110.735 ;
        RECT 85.585 110.690 85.875 110.735 ;
        RECT 81.875 110.550 85.875 110.690 ;
        RECT 81.875 110.505 82.165 110.550 ;
        RECT 83.065 110.505 83.355 110.550 ;
        RECT 85.585 110.505 85.875 110.550 ;
        RECT 87.970 110.690 88.110 110.890 ;
        RECT 95.240 110.830 95.560 111.090 ;
        RECT 96.160 111.030 96.480 111.090 ;
        RECT 100.300 111.030 100.620 111.090 ;
        RECT 96.160 110.890 100.620 111.030 ;
        RECT 104.530 111.030 104.670 111.525 ;
        RECT 113.180 111.510 113.500 111.570 ;
        RECT 115.480 111.710 115.800 111.770 ;
        RECT 116.860 111.710 117.180 111.770 ;
        RECT 115.480 111.570 117.180 111.710 ;
        RECT 115.480 111.510 115.800 111.570 ;
        RECT 116.860 111.510 117.180 111.570 ;
        RECT 122.840 111.710 123.160 111.770 ;
        RECT 126.980 111.710 127.300 111.770 ;
        RECT 128.820 111.710 129.140 111.770 ;
        RECT 122.840 111.570 129.140 111.710 ;
        RECT 122.840 111.510 123.160 111.570 ;
        RECT 126.980 111.510 127.300 111.570 ;
        RECT 128.820 111.510 129.140 111.570 ;
        RECT 130.675 111.710 130.965 111.755 ;
        RECT 130.675 111.570 131.810 111.710 ;
        RECT 130.675 111.525 130.965 111.570 ;
        RECT 105.360 111.170 105.680 111.430 ;
        RECT 116.400 111.370 116.720 111.430 ;
        RECT 124.695 111.370 124.985 111.415 ;
        RECT 131.670 111.370 131.810 111.570 ;
        RECT 132.360 111.370 132.650 111.415 ;
        RECT 140.335 111.370 140.625 111.415 ;
        RECT 116.400 111.230 131.350 111.370 ;
        RECT 131.670 111.230 132.650 111.370 ;
        RECT 116.400 111.170 116.720 111.230 ;
        RECT 124.695 111.185 124.985 111.230 ;
        RECT 131.210 111.090 131.350 111.230 ;
        RECT 132.360 111.185 132.650 111.230 ;
        RECT 134.430 111.230 140.625 111.370 ;
        RECT 107.200 111.030 107.520 111.090 ;
        RECT 104.530 110.890 107.520 111.030 ;
        RECT 96.160 110.830 96.480 110.890 ;
        RECT 100.300 110.830 100.620 110.890 ;
        RECT 107.200 110.830 107.520 110.890 ;
        RECT 109.960 110.830 110.280 111.090 ;
        RECT 112.260 110.830 112.580 111.090 ;
        RECT 113.195 111.030 113.485 111.075 ;
        RECT 113.195 110.890 118.470 111.030 ;
        RECT 113.195 110.845 113.485 110.890 ;
        RECT 103.980 110.690 104.300 110.750 ;
        RECT 106.740 110.690 107.060 110.750 ;
        RECT 87.970 110.550 104.300 110.690 ;
        RECT 78.680 110.350 79.000 110.410 ;
        RECT 87.970 110.395 88.110 110.550 ;
        RECT 103.980 110.490 104.300 110.550 ;
        RECT 104.530 110.550 107.060 110.690 ;
        RECT 118.330 110.690 118.470 110.890 ;
        RECT 118.700 110.830 119.020 111.090 ;
        RECT 119.620 111.030 119.940 111.090 ;
        RECT 121.935 111.030 122.225 111.075 ;
        RECT 119.620 110.890 122.225 111.030 ;
        RECT 119.620 110.830 119.940 110.890 ;
        RECT 121.935 110.845 122.225 110.890 ;
        RECT 122.380 110.830 122.700 111.090 ;
        RECT 122.855 110.845 123.145 111.075 ;
        RECT 122.930 110.690 123.070 110.845 ;
        RECT 123.760 110.830 124.080 111.090 ;
        RECT 127.440 110.830 127.760 111.090 ;
        RECT 128.375 110.845 128.665 111.075 ;
        RECT 126.060 110.690 126.380 110.750 ;
        RECT 118.330 110.550 126.380 110.690 ;
        RECT 128.450 110.690 128.590 110.845 ;
        RECT 128.820 110.830 129.140 111.090 ;
        RECT 129.295 111.030 129.585 111.075 ;
        RECT 130.660 111.030 130.980 111.090 ;
        RECT 129.295 110.890 130.980 111.030 ;
        RECT 129.295 110.845 129.585 110.890 ;
        RECT 130.660 110.830 130.980 110.890 ;
        RECT 131.120 110.830 131.440 111.090 ;
        RECT 134.430 111.030 134.570 111.230 ;
        RECT 140.335 111.185 140.625 111.230 ;
        RECT 131.670 110.890 134.570 111.030 ;
        RECT 131.670 110.690 131.810 110.890 ;
        RECT 138.480 110.830 138.800 111.090 ;
        RECT 139.415 111.030 139.705 111.075 ;
        RECT 139.860 111.030 140.180 111.090 ;
        RECT 139.415 110.890 140.180 111.030 ;
        RECT 139.415 110.845 139.705 110.890 ;
        RECT 128.450 110.550 131.810 110.690 ;
        RECT 132.015 110.690 132.305 110.735 ;
        RECT 133.205 110.690 133.495 110.735 ;
        RECT 135.725 110.690 136.015 110.735 ;
        RECT 139.490 110.690 139.630 110.845 ;
        RECT 139.860 110.830 140.180 110.890 ;
        RECT 132.015 110.550 136.015 110.690 ;
        RECT 81.480 110.350 81.770 110.395 ;
        RECT 83.580 110.350 83.870 110.395 ;
        RECT 85.150 110.350 85.440 110.395 ;
        RECT 78.680 110.210 80.290 110.350 ;
        RECT 78.680 110.150 79.000 110.210 ;
        RECT 80.150 110.055 80.290 110.210 ;
        RECT 81.480 110.210 85.440 110.350 ;
        RECT 81.480 110.165 81.770 110.210 ;
        RECT 83.580 110.165 83.870 110.210 ;
        RECT 85.150 110.165 85.440 110.210 ;
        RECT 87.895 110.165 88.185 110.395 ;
        RECT 100.760 110.350 101.080 110.410 ;
        RECT 103.535 110.350 103.825 110.395 ;
        RECT 100.760 110.210 103.825 110.350 ;
        RECT 100.760 110.150 101.080 110.210 ;
        RECT 103.535 110.165 103.825 110.210 ;
        RECT 104.530 110.055 104.670 110.550 ;
        RECT 106.740 110.490 107.060 110.550 ;
        RECT 126.060 110.490 126.380 110.550 ;
        RECT 132.015 110.505 132.305 110.550 ;
        RECT 133.205 110.505 133.495 110.550 ;
        RECT 135.725 110.505 136.015 110.550 ;
        RECT 138.110 110.550 139.630 110.690 ;
        RECT 116.860 110.350 117.180 110.410 ;
        RECT 119.635 110.350 119.925 110.395 ;
        RECT 129.280 110.350 129.600 110.410 ;
        RECT 116.860 110.210 129.600 110.350 ;
        RECT 116.860 110.150 117.180 110.210 ;
        RECT 119.635 110.165 119.925 110.210 ;
        RECT 129.280 110.150 129.600 110.210 ;
        RECT 131.620 110.350 131.910 110.395 ;
        RECT 133.720 110.350 134.010 110.395 ;
        RECT 135.290 110.350 135.580 110.395 ;
        RECT 131.620 110.210 135.580 110.350 ;
        RECT 131.620 110.165 131.910 110.210 ;
        RECT 133.720 110.165 134.010 110.210 ;
        RECT 135.290 110.165 135.580 110.210 ;
        RECT 136.180 110.350 136.500 110.410 ;
        RECT 138.110 110.395 138.250 110.550 ;
        RECT 138.035 110.350 138.325 110.395 ;
        RECT 136.180 110.210 138.325 110.350 ;
        RECT 136.180 110.150 136.500 110.210 ;
        RECT 138.035 110.165 138.325 110.210 ;
        RECT 76.395 110.010 76.685 110.055 ;
        RECT 75.460 109.870 76.685 110.010 ;
        RECT 75.460 109.810 75.780 109.870 ;
        RECT 76.395 109.825 76.685 109.870 ;
        RECT 80.075 109.825 80.365 110.055 ;
        RECT 104.455 109.825 104.745 110.055 ;
        RECT 106.290 110.010 106.585 110.085 ;
        RECT 109.050 110.010 109.345 110.085 ;
        RECT 106.290 109.870 109.345 110.010 ;
        RECT 106.290 109.815 106.585 109.870 ;
        RECT 109.050 109.815 109.345 109.870 ;
        RECT 115.480 110.010 115.800 110.070 ;
        RECT 121.015 110.010 121.305 110.055 ;
        RECT 115.480 109.870 121.305 110.010 ;
        RECT 115.480 109.810 115.800 109.870 ;
        RECT 121.015 109.825 121.305 109.870 ;
        RECT 17.430 109.190 143.010 109.670 ;
        RECT 23.955 108.990 24.245 109.035 ;
        RECT 25.780 108.990 26.100 109.050 ;
        RECT 23.955 108.850 26.100 108.990 ;
        RECT 23.955 108.805 24.245 108.850 ;
        RECT 25.780 108.790 26.100 108.850 ;
        RECT 27.620 108.790 27.940 109.050 ;
        RECT 40.040 108.790 40.360 109.050 ;
        RECT 40.960 108.790 41.280 109.050 ;
        RECT 48.780 108.990 49.100 109.050 ;
        RECT 50.175 108.990 50.465 109.035 ;
        RECT 48.780 108.850 50.465 108.990 ;
        RECT 48.780 108.790 49.100 108.850 ;
        RECT 50.175 108.805 50.465 108.850 ;
        RECT 69.480 108.990 69.800 109.050 ;
        RECT 70.415 108.990 70.705 109.035 ;
        RECT 69.480 108.850 70.705 108.990 ;
        RECT 69.480 108.790 69.800 108.850 ;
        RECT 70.415 108.805 70.705 108.850 ;
        RECT 70.860 108.990 71.180 109.050 ;
        RECT 71.795 108.990 72.085 109.035 ;
        RECT 70.860 108.850 72.085 108.990 ;
        RECT 70.860 108.790 71.180 108.850 ;
        RECT 71.795 108.805 72.085 108.850 ;
        RECT 72.715 108.805 73.005 109.035 ;
        RECT 87.880 108.990 88.200 109.050 ;
        RECT 81.070 108.850 88.200 108.990 ;
        RECT 26.715 108.650 27.005 108.695 ;
        RECT 28.540 108.650 28.860 108.710 ;
        RECT 39.580 108.650 39.900 108.710 ;
        RECT 42.340 108.650 42.660 108.710 ;
        RECT 42.815 108.650 43.105 108.695 ;
        RECT 26.715 108.510 28.860 108.650 ;
        RECT 26.715 108.465 27.005 108.510 ;
        RECT 28.540 108.450 28.860 108.510 ;
        RECT 32.770 108.510 39.350 108.650 ;
        RECT 26.330 108.170 30.150 108.310 ;
        RECT 26.330 108.015 26.470 108.170 ;
        RECT 30.010 108.030 30.150 108.170 ;
        RECT 25.795 107.970 26.085 108.015 ;
        RECT 26.255 107.970 26.545 108.015 ;
        RECT 25.795 107.830 26.545 107.970 ;
        RECT 25.795 107.785 26.085 107.830 ;
        RECT 26.255 107.785 26.545 107.830 ;
        RECT 27.175 107.785 27.465 108.015 ;
        RECT 28.555 107.785 28.845 108.015 ;
        RECT 23.955 107.630 24.245 107.675 ;
        RECT 24.860 107.630 25.180 107.690 ;
        RECT 23.955 107.490 25.180 107.630 ;
        RECT 23.955 107.445 24.245 107.490 ;
        RECT 24.860 107.430 25.180 107.490 ;
        RECT 23.035 107.290 23.325 107.335 ;
        RECT 23.480 107.290 23.800 107.350 ;
        RECT 23.035 107.150 23.800 107.290 ;
        RECT 27.250 107.290 27.390 107.785 ;
        RECT 28.630 107.630 28.770 107.785 ;
        RECT 29.460 107.770 29.780 108.030 ;
        RECT 29.920 107.770 30.240 108.030 ;
        RECT 31.300 107.770 31.620 108.030 ;
        RECT 31.775 107.785 32.065 108.015 ;
        RECT 31.850 107.630 31.990 107.785 ;
        RECT 32.220 107.770 32.540 108.030 ;
        RECT 32.770 108.015 32.910 108.510 ;
        RECT 33.615 108.310 33.905 108.355 ;
        RECT 37.755 108.310 38.045 108.355 ;
        RECT 33.615 108.170 38.045 108.310 ;
        RECT 39.210 108.310 39.350 108.510 ;
        RECT 39.580 108.510 43.105 108.650 ;
        RECT 39.580 108.450 39.900 108.510 ;
        RECT 42.340 108.450 42.660 108.510 ;
        RECT 42.815 108.465 43.105 108.510 ;
        RECT 49.255 108.465 49.545 108.695 ;
        RECT 56.615 108.650 56.905 108.695 ;
        RECT 53.010 108.510 56.905 108.650 ;
        RECT 40.500 108.310 40.820 108.370 ;
        RECT 39.210 108.170 40.820 108.310 ;
        RECT 33.615 108.125 33.905 108.170 ;
        RECT 37.755 108.125 38.045 108.170 ;
        RECT 40.500 108.110 40.820 108.170 ;
        RECT 40.960 108.310 41.280 108.370 ;
        RECT 49.330 108.310 49.470 108.465 ;
        RECT 53.010 108.355 53.150 108.510 ;
        RECT 56.615 108.465 56.905 108.510 ;
        RECT 59.360 108.650 59.650 108.695 ;
        RECT 60.930 108.650 61.220 108.695 ;
        RECT 63.030 108.650 63.320 108.695 ;
        RECT 59.360 108.510 63.320 108.650 ;
        RECT 59.360 108.465 59.650 108.510 ;
        RECT 60.930 108.465 61.220 108.510 ;
        RECT 63.030 108.465 63.320 108.510 ;
        RECT 67.180 108.650 67.500 108.710 ;
        RECT 72.790 108.650 72.930 108.805 ;
        RECT 67.180 108.510 72.930 108.650 ;
        RECT 67.180 108.450 67.500 108.510 ;
        RECT 40.960 108.170 49.470 108.310 ;
        RECT 52.015 108.310 52.305 108.355 ;
        RECT 52.935 108.310 53.225 108.355 ;
        RECT 52.015 108.170 53.225 108.310 ;
        RECT 40.960 108.110 41.280 108.170 ;
        RECT 52.015 108.125 52.305 108.170 ;
        RECT 52.935 108.125 53.225 108.170 ;
        RECT 58.925 108.310 59.215 108.355 ;
        RECT 61.445 108.310 61.735 108.355 ;
        RECT 62.635 108.310 62.925 108.355 ;
        RECT 58.925 108.170 62.925 108.310 ;
        RECT 58.925 108.125 59.215 108.170 ;
        RECT 61.445 108.125 61.735 108.170 ;
        RECT 62.635 108.125 62.925 108.170 ;
        RECT 63.960 108.310 64.280 108.370 ;
        RECT 66.720 108.310 67.040 108.370 ;
        RECT 67.655 108.310 67.945 108.355 ;
        RECT 63.960 108.170 67.945 108.310 ;
        RECT 63.960 108.110 64.280 108.170 ;
        RECT 66.720 108.110 67.040 108.170 ;
        RECT 67.655 108.125 67.945 108.170 ;
        RECT 70.400 108.310 70.720 108.370 ;
        RECT 74.540 108.310 74.860 108.370 ;
        RECT 70.400 108.170 74.860 108.310 ;
        RECT 70.400 108.110 70.720 108.170 ;
        RECT 74.540 108.110 74.860 108.170 ;
        RECT 77.315 108.310 77.605 108.355 ;
        RECT 78.220 108.310 78.540 108.370 ;
        RECT 77.315 108.170 78.540 108.310 ;
        RECT 77.315 108.125 77.605 108.170 ;
        RECT 32.695 107.785 32.985 108.015 ;
        RECT 35.440 107.970 35.760 108.030 ;
        RECT 35.915 107.970 36.205 108.015 ;
        RECT 35.440 107.830 36.205 107.970 ;
        RECT 35.440 107.770 35.760 107.830 ;
        RECT 35.915 107.785 36.205 107.830 ;
        RECT 36.835 107.785 37.125 108.015 ;
        RECT 37.295 107.970 37.585 108.015 ;
        RECT 38.200 107.970 38.520 108.030 ;
        RECT 37.295 107.830 38.520 107.970 ;
        RECT 37.295 107.785 37.585 107.830 ;
        RECT 33.600 107.630 33.920 107.690 ;
        RECT 28.630 107.490 30.150 107.630 ;
        RECT 31.850 107.490 33.920 107.630 ;
        RECT 36.910 107.630 37.050 107.785 ;
        RECT 38.200 107.770 38.520 107.830 ;
        RECT 38.675 107.970 38.965 108.015 ;
        RECT 41.420 107.970 41.740 108.030 ;
        RECT 38.675 107.830 41.740 107.970 ;
        RECT 38.675 107.785 38.965 107.830 ;
        RECT 41.420 107.770 41.740 107.830 ;
        RECT 44.640 107.770 44.960 108.030 ;
        RECT 45.100 107.970 45.420 108.030 ;
        RECT 45.100 107.830 45.615 107.970 ;
        RECT 45.100 107.770 45.420 107.830 ;
        RECT 46.480 107.770 46.800 108.030 ;
        RECT 47.185 107.970 47.475 108.015 ;
        RECT 47.860 107.970 48.180 108.030 ;
        RECT 47.185 107.830 48.180 107.970 ;
        RECT 47.185 107.785 47.475 107.830 ;
        RECT 47.860 107.770 48.180 107.830 ;
        RECT 63.515 107.970 63.805 108.015 ;
        RECT 64.420 107.970 64.740 108.030 ;
        RECT 63.515 107.830 64.740 107.970 ;
        RECT 63.515 107.785 63.805 107.830 ;
        RECT 64.420 107.770 64.740 107.830 ;
        RECT 66.275 107.785 66.565 108.015 ;
        RECT 67.195 107.785 67.485 108.015 ;
        RECT 68.100 107.970 68.420 108.030 ;
        RECT 70.875 107.970 71.165 108.015 ;
        RECT 68.100 107.830 71.165 107.970 ;
        RECT 43.720 107.630 44.040 107.690 ;
        RECT 36.910 107.490 44.040 107.630 ;
        RECT 29.460 107.290 29.780 107.350 ;
        RECT 27.250 107.150 29.780 107.290 ;
        RECT 30.010 107.290 30.150 107.490 ;
        RECT 33.600 107.430 33.920 107.490 ;
        RECT 43.720 107.430 44.040 107.490 ;
        RECT 46.035 107.445 46.325 107.675 ;
        RECT 57.520 107.630 57.840 107.690 ;
        RECT 47.030 107.490 57.840 107.630 ;
        RECT 34.980 107.290 35.300 107.350 ;
        RECT 30.010 107.150 35.300 107.290 ;
        RECT 23.035 107.105 23.325 107.150 ;
        RECT 23.480 107.090 23.800 107.150 ;
        RECT 29.460 107.090 29.780 107.150 ;
        RECT 34.980 107.090 35.300 107.150 ;
        RECT 39.580 107.090 39.900 107.350 ;
        RECT 40.960 107.090 41.280 107.350 ;
        RECT 46.110 107.290 46.250 107.445 ;
        RECT 47.030 107.290 47.170 107.490 ;
        RECT 57.520 107.430 57.840 107.490 ;
        RECT 62.290 107.630 62.580 107.675 ;
        RECT 65.355 107.630 65.645 107.675 ;
        RECT 62.290 107.490 65.645 107.630 ;
        RECT 62.290 107.445 62.580 107.490 ;
        RECT 65.355 107.445 65.645 107.490 ;
        RECT 46.110 107.150 47.170 107.290 ;
        RECT 47.400 107.290 47.720 107.350 ;
        RECT 47.875 107.290 48.165 107.335 ;
        RECT 47.400 107.150 48.165 107.290 ;
        RECT 47.400 107.090 47.720 107.150 ;
        RECT 47.875 107.105 48.165 107.150 ;
        RECT 50.175 107.290 50.465 107.335 ;
        RECT 52.000 107.290 52.320 107.350 ;
        RECT 50.175 107.150 52.320 107.290 ;
        RECT 50.175 107.105 50.465 107.150 ;
        RECT 52.000 107.090 52.320 107.150 ;
        RECT 55.680 107.290 56.000 107.350 ;
        RECT 66.350 107.290 66.490 107.785 ;
        RECT 66.720 107.630 67.040 107.690 ;
        RECT 67.270 107.630 67.410 107.785 ;
        RECT 68.100 107.770 68.420 107.830 ;
        RECT 70.875 107.785 71.165 107.830 ;
        RECT 71.335 107.970 71.625 108.015 ;
        RECT 75.000 107.970 75.320 108.030 ;
        RECT 77.390 107.970 77.530 108.125 ;
        RECT 78.220 108.110 78.540 108.170 ;
        RECT 78.695 108.310 78.985 108.355 ;
        RECT 79.140 108.310 79.460 108.370 ;
        RECT 78.695 108.170 79.460 108.310 ;
        RECT 78.695 108.125 78.985 108.170 ;
        RECT 79.140 108.110 79.460 108.170 ;
        RECT 81.070 107.970 81.210 108.850 ;
        RECT 87.880 108.790 88.200 108.850 ;
        RECT 98.920 108.790 99.240 109.050 ;
        RECT 108.120 108.990 108.440 109.050 ;
        RECT 108.595 108.990 108.885 109.035 ;
        RECT 116.400 108.990 116.720 109.050 ;
        RECT 108.120 108.850 116.720 108.990 ;
        RECT 108.120 108.790 108.440 108.850 ;
        RECT 108.595 108.805 108.885 108.850 ;
        RECT 116.400 108.790 116.720 108.850 ;
        RECT 81.455 108.465 81.745 108.695 ;
        RECT 82.860 108.650 83.150 108.695 ;
        RECT 84.960 108.650 85.250 108.695 ;
        RECT 86.530 108.650 86.820 108.695 ;
        RECT 82.860 108.510 86.820 108.650 ;
        RECT 82.860 108.465 83.150 108.510 ;
        RECT 84.960 108.465 85.250 108.510 ;
        RECT 86.530 108.465 86.820 108.510 ;
        RECT 102.140 108.650 102.460 108.710 ;
        RECT 115.020 108.650 115.340 108.710 ;
        RECT 102.140 108.510 115.340 108.650 ;
        RECT 71.335 107.830 77.530 107.970 ;
        RECT 79.230 107.830 81.210 107.970 ;
        RECT 71.335 107.785 71.625 107.830 ;
        RECT 75.000 107.770 75.320 107.830 ;
        RECT 72.240 107.675 72.560 107.690 ;
        RECT 72.240 107.630 72.845 107.675 ;
        RECT 66.720 107.490 72.995 107.630 ;
        RECT 66.720 107.430 67.040 107.490 ;
        RECT 72.240 107.445 72.845 107.490 ;
        RECT 72.240 107.430 72.560 107.445 ;
        RECT 73.620 107.430 73.940 107.690 ;
        RECT 74.540 107.630 74.860 107.690 ;
        RECT 79.230 107.675 79.370 107.830 ;
        RECT 79.155 107.630 79.445 107.675 ;
        RECT 74.540 107.490 79.445 107.630 ;
        RECT 81.530 107.630 81.670 108.465 ;
        RECT 102.140 108.450 102.460 108.510 ;
        RECT 115.020 108.450 115.340 108.510 ;
        RECT 115.980 108.650 116.270 108.695 ;
        RECT 118.080 108.650 118.370 108.695 ;
        RECT 119.650 108.650 119.940 108.695 ;
        RECT 115.980 108.510 119.940 108.650 ;
        RECT 115.980 108.465 116.270 108.510 ;
        RECT 118.080 108.465 118.370 108.510 ;
        RECT 119.650 108.465 119.940 108.510 ;
        RECT 134.380 108.650 134.670 108.695 ;
        RECT 136.480 108.650 136.770 108.695 ;
        RECT 138.050 108.650 138.340 108.695 ;
        RECT 134.380 108.510 138.340 108.650 ;
        RECT 134.380 108.465 134.670 108.510 ;
        RECT 136.480 108.465 136.770 108.510 ;
        RECT 138.050 108.465 138.340 108.510 ;
        RECT 83.255 108.310 83.545 108.355 ;
        RECT 84.445 108.310 84.735 108.355 ;
        RECT 86.965 108.310 87.255 108.355 ;
        RECT 83.255 108.170 87.255 108.310 ;
        RECT 83.255 108.125 83.545 108.170 ;
        RECT 84.445 108.125 84.735 108.170 ;
        RECT 86.965 108.125 87.255 108.170 ;
        RECT 97.080 108.310 97.400 108.370 ;
        RECT 112.260 108.310 112.580 108.370 ;
        RECT 97.080 108.170 106.510 108.310 ;
        RECT 97.080 108.110 97.400 108.170 ;
        RECT 82.375 107.970 82.665 108.015 ;
        RECT 82.820 107.970 83.140 108.030 ;
        RECT 82.375 107.830 83.140 107.970 ;
        RECT 82.375 107.785 82.665 107.830 ;
        RECT 82.820 107.770 83.140 107.830 ;
        RECT 99.395 107.970 99.685 108.015 ;
        RECT 101.220 107.970 101.540 108.030 ;
        RECT 106.370 108.015 106.510 108.170 ;
        RECT 108.210 108.170 112.580 108.310 ;
        RECT 108.210 108.015 108.350 108.170 ;
        RECT 112.260 108.110 112.580 108.170 ;
        RECT 116.375 108.310 116.665 108.355 ;
        RECT 117.565 108.310 117.855 108.355 ;
        RECT 120.085 108.310 120.375 108.355 ;
        RECT 131.580 108.310 131.900 108.370 ;
        RECT 133.895 108.310 134.185 108.355 ;
        RECT 116.375 108.170 120.375 108.310 ;
        RECT 116.375 108.125 116.665 108.170 ;
        RECT 117.565 108.125 117.855 108.170 ;
        RECT 120.085 108.125 120.375 108.170 ;
        RECT 126.610 108.170 134.185 108.310 ;
        RECT 99.395 107.830 101.540 107.970 ;
        RECT 99.395 107.785 99.685 107.830 ;
        RECT 101.220 107.770 101.540 107.830 ;
        RECT 101.695 107.970 101.985 108.015 ;
        RECT 103.075 107.970 103.365 108.015 ;
        RECT 101.695 107.830 103.365 107.970 ;
        RECT 101.695 107.785 101.985 107.830 ;
        RECT 103.075 107.785 103.365 107.830 ;
        RECT 105.835 107.785 106.125 108.015 ;
        RECT 106.295 107.970 106.585 108.015 ;
        RECT 108.135 107.970 108.425 108.015 ;
        RECT 106.295 107.830 108.425 107.970 ;
        RECT 106.295 107.785 106.585 107.830 ;
        RECT 108.135 107.785 108.425 107.830 ;
        RECT 109.515 107.785 109.805 108.015 ;
        RECT 115.495 107.970 115.785 108.015 ;
        RECT 115.940 107.970 116.260 108.030 ;
        RECT 126.610 108.015 126.750 108.170 ;
        RECT 131.580 108.110 131.900 108.170 ;
        RECT 133.895 108.125 134.185 108.170 ;
        RECT 134.775 108.310 135.065 108.355 ;
        RECT 135.965 108.310 136.255 108.355 ;
        RECT 138.485 108.310 138.775 108.355 ;
        RECT 134.775 108.170 138.775 108.310 ;
        RECT 134.775 108.125 135.065 108.170 ;
        RECT 135.965 108.125 136.255 108.170 ;
        RECT 138.485 108.125 138.775 108.170 ;
        RECT 126.535 107.970 126.825 108.015 ;
        RECT 115.495 107.830 126.825 107.970 ;
        RECT 115.495 107.785 115.785 107.830 ;
        RECT 83.600 107.630 83.890 107.675 ;
        RECT 81.530 107.490 83.890 107.630 ;
        RECT 74.540 107.430 74.860 107.490 ;
        RECT 79.155 107.445 79.445 107.490 ;
        RECT 83.600 107.445 83.890 107.490 ;
        RECT 89.720 107.630 90.040 107.690 ;
        RECT 92.495 107.630 92.785 107.675 ;
        RECT 89.720 107.490 92.785 107.630 ;
        RECT 89.720 107.430 90.040 107.490 ;
        RECT 92.495 107.445 92.785 107.490 ;
        RECT 100.315 107.630 100.605 107.675 ;
        RECT 101.770 107.630 101.910 107.785 ;
        RECT 100.315 107.490 101.910 107.630 ;
        RECT 103.535 107.630 103.825 107.675 ;
        RECT 105.910 107.630 106.050 107.785 ;
        RECT 109.590 107.630 109.730 107.785 ;
        RECT 115.940 107.770 116.260 107.830 ;
        RECT 126.535 107.785 126.825 107.830 ;
        RECT 127.440 107.970 127.760 108.030 ;
        RECT 127.915 107.970 128.205 108.015 ;
        RECT 127.440 107.830 128.205 107.970 ;
        RECT 127.440 107.770 127.760 107.830 ;
        RECT 127.915 107.785 128.205 107.830 ;
        RECT 128.835 107.785 129.125 108.015 ;
        RECT 116.860 107.675 117.180 107.690 ;
        RECT 103.535 107.490 109.730 107.630 ;
        RECT 100.315 107.445 100.605 107.490 ;
        RECT 103.535 107.445 103.825 107.490 ;
        RECT 55.680 107.150 66.490 107.290 ;
        RECT 69.020 107.290 69.340 107.350 ;
        RECT 69.495 107.290 69.785 107.335 ;
        RECT 69.020 107.150 69.785 107.290 ;
        RECT 55.680 107.090 56.000 107.150 ;
        RECT 69.020 107.090 69.340 107.150 ;
        RECT 69.495 107.105 69.785 107.150 ;
        RECT 74.080 107.090 74.400 107.350 ;
        RECT 79.615 107.290 79.905 107.335 ;
        RECT 89.275 107.290 89.565 107.335 ;
        RECT 91.100 107.290 91.420 107.350 ;
        RECT 79.615 107.150 91.420 107.290 ;
        RECT 79.615 107.105 79.905 107.150 ;
        RECT 89.275 107.105 89.565 107.150 ;
        RECT 91.100 107.090 91.420 107.150 ;
        RECT 94.780 107.290 95.100 107.350 ;
        RECT 100.390 107.290 100.530 107.445 ;
        RECT 94.780 107.150 100.530 107.290 ;
        RECT 94.780 107.090 95.100 107.150 ;
        RECT 107.200 107.090 107.520 107.350 ;
        RECT 109.590 107.290 109.730 107.490 ;
        RECT 116.830 107.445 117.180 107.675 ;
        RECT 116.860 107.430 117.180 107.445 ;
        RECT 121.000 107.630 121.320 107.690 ;
        RECT 122.855 107.630 123.145 107.675 ;
        RECT 121.000 107.490 123.145 107.630 ;
        RECT 128.910 107.630 129.050 107.785 ;
        RECT 129.280 107.770 129.600 108.030 ;
        RECT 129.755 107.970 130.045 108.015 ;
        RECT 130.660 107.970 130.980 108.030 ;
        RECT 134.340 107.970 134.660 108.030 ;
        RECT 129.755 107.830 130.980 107.970 ;
        RECT 129.755 107.785 130.045 107.830 ;
        RECT 130.660 107.770 130.980 107.830 ;
        RECT 131.210 107.830 134.660 107.970 ;
        RECT 131.210 107.630 131.350 107.830 ;
        RECT 134.340 107.770 134.660 107.830 ;
        RECT 128.910 107.490 131.350 107.630 ;
        RECT 132.040 107.630 132.360 107.690 ;
        RECT 135.120 107.630 135.410 107.675 ;
        RECT 132.040 107.490 135.410 107.630 ;
        RECT 121.000 107.430 121.320 107.490 ;
        RECT 122.855 107.445 123.145 107.490 ;
        RECT 132.040 107.430 132.360 107.490 ;
        RECT 135.120 107.445 135.410 107.490 ;
        RECT 118.240 107.290 118.560 107.350 ;
        RECT 109.590 107.150 118.560 107.290 ;
        RECT 118.240 107.090 118.560 107.150 ;
        RECT 122.380 107.290 122.700 107.350 ;
        RECT 123.760 107.290 124.080 107.350 ;
        RECT 122.380 107.150 124.080 107.290 ;
        RECT 122.380 107.090 122.700 107.150 ;
        RECT 123.760 107.090 124.080 107.150 ;
        RECT 131.120 107.090 131.440 107.350 ;
        RECT 140.320 107.290 140.640 107.350 ;
        RECT 140.795 107.290 141.085 107.335 ;
        RECT 140.320 107.150 141.085 107.290 ;
        RECT 140.320 107.090 140.640 107.150 ;
        RECT 140.795 107.105 141.085 107.150 ;
        RECT 17.430 106.470 143.010 106.950 ;
        RECT 30.840 106.270 31.160 106.330 ;
        RECT 31.315 106.270 31.605 106.315 ;
        RECT 30.840 106.130 31.605 106.270 ;
        RECT 30.840 106.070 31.160 106.130 ;
        RECT 31.315 106.085 31.605 106.130 ;
        RECT 33.600 106.070 33.920 106.330 ;
        RECT 34.980 106.070 35.300 106.330 ;
        RECT 45.100 106.270 45.420 106.330 ;
        RECT 45.100 106.130 48.550 106.270 ;
        RECT 45.100 106.070 45.420 106.130 ;
        RECT 29.920 105.930 30.240 105.990 ;
        RECT 32.075 105.930 32.365 105.975 ;
        RECT 29.920 105.790 32.365 105.930 ;
        RECT 29.920 105.730 30.240 105.790 ;
        RECT 32.075 105.745 32.365 105.790 ;
        RECT 33.155 105.930 33.445 105.975 ;
        RECT 35.070 105.930 35.210 106.070 ;
        RECT 33.155 105.790 35.210 105.930 ;
        RECT 39.580 105.930 39.900 105.990 ;
        RECT 48.410 105.930 48.550 106.130 ;
        RECT 48.780 106.070 49.100 106.330 ;
        RECT 52.000 106.070 52.320 106.330 ;
        RECT 57.520 106.070 57.840 106.330 ;
        RECT 65.355 106.270 65.645 106.315 ;
        RECT 69.940 106.270 70.260 106.330 ;
        RECT 65.355 106.130 70.260 106.270 ;
        RECT 65.355 106.085 65.645 106.130 ;
        RECT 69.940 106.070 70.260 106.130 ;
        RECT 72.715 106.270 73.005 106.315 ;
        RECT 94.780 106.270 95.100 106.330 ;
        RECT 72.715 106.130 95.100 106.270 ;
        RECT 72.715 106.085 73.005 106.130 ;
        RECT 94.780 106.070 95.100 106.130 ;
        RECT 95.255 106.270 95.545 106.315 ;
        RECT 95.700 106.270 96.020 106.330 ;
        RECT 95.255 106.130 96.020 106.270 ;
        RECT 95.255 106.085 95.545 106.130 ;
        RECT 95.700 106.070 96.020 106.130 ;
        RECT 107.200 106.270 107.520 106.330 ;
        RECT 115.955 106.270 116.245 106.315 ;
        RECT 116.860 106.270 117.180 106.330 ;
        RECT 121.920 106.270 122.240 106.330 ;
        RECT 133.420 106.270 133.740 106.330 ;
        RECT 107.200 106.130 112.030 106.270 ;
        RECT 107.200 106.070 107.520 106.130 ;
        RECT 56.615 105.930 56.905 105.975 ;
        RECT 74.080 105.930 74.400 105.990 ;
        RECT 89.720 105.930 90.040 105.990 ;
        RECT 39.580 105.790 46.710 105.930 ;
        RECT 48.410 105.790 50.390 105.930 ;
        RECT 33.155 105.745 33.445 105.790 ;
        RECT 39.580 105.730 39.900 105.790 ;
        RECT 23.480 105.635 23.800 105.650 ;
        RECT 23.450 105.590 23.800 105.635 ;
        RECT 23.285 105.450 23.800 105.590 ;
        RECT 23.450 105.405 23.800 105.450 ;
        RECT 34.535 105.590 34.825 105.635 ;
        RECT 34.980 105.590 35.300 105.650 ;
        RECT 34.535 105.450 35.300 105.590 ;
        RECT 34.535 105.405 34.825 105.450 ;
        RECT 23.480 105.390 23.800 105.405 ;
        RECT 34.980 105.390 35.300 105.450 ;
        RECT 46.035 105.405 46.325 105.635 ;
        RECT 46.570 105.590 46.710 105.790 ;
        RECT 46.860 105.590 47.150 105.635 ;
        RECT 46.570 105.450 47.150 105.590 ;
        RECT 46.860 105.405 47.150 105.450 ;
        RECT 21.640 105.250 21.960 105.310 ;
        RECT 22.115 105.250 22.405 105.295 ;
        RECT 21.640 105.110 22.405 105.250 ;
        RECT 21.640 105.050 21.960 105.110 ;
        RECT 22.115 105.065 22.405 105.110 ;
        RECT 22.995 105.250 23.285 105.295 ;
        RECT 24.185 105.250 24.475 105.295 ;
        RECT 26.705 105.250 26.995 105.295 ;
        RECT 22.995 105.110 26.995 105.250 ;
        RECT 22.995 105.065 23.285 105.110 ;
        RECT 24.185 105.065 24.475 105.110 ;
        RECT 26.705 105.065 26.995 105.110 ;
        RECT 29.000 105.250 29.320 105.310 ;
        RECT 35.455 105.250 35.745 105.295 ;
        RECT 29.000 105.110 35.745 105.250 ;
        RECT 29.000 105.050 29.320 105.110 ;
        RECT 35.455 105.065 35.745 105.110 ;
        RECT 22.600 104.910 22.890 104.955 ;
        RECT 24.700 104.910 24.990 104.955 ;
        RECT 26.270 104.910 26.560 104.955 ;
        RECT 22.600 104.770 26.560 104.910 ;
        RECT 22.600 104.725 22.890 104.770 ;
        RECT 24.700 104.725 24.990 104.770 ;
        RECT 26.270 104.725 26.560 104.770 ;
        RECT 28.080 104.570 28.400 104.630 ;
        RECT 29.015 104.570 29.305 104.615 ;
        RECT 28.080 104.430 29.305 104.570 ;
        RECT 28.080 104.370 28.400 104.430 ;
        RECT 29.015 104.385 29.305 104.430 ;
        RECT 29.460 104.570 29.780 104.630 ;
        RECT 32.235 104.570 32.525 104.615 ;
        RECT 29.460 104.430 32.525 104.570 ;
        RECT 46.110 104.570 46.250 105.405 ;
        RECT 47.400 105.390 47.720 105.650 ;
        RECT 47.875 105.590 48.165 105.635 ;
        RECT 48.320 105.590 48.640 105.650 ;
        RECT 50.250 105.635 50.390 105.790 ;
        RECT 51.170 105.790 56.905 105.930 ;
        RECT 51.170 105.650 51.310 105.790 ;
        RECT 56.615 105.745 56.905 105.790 ;
        RECT 66.810 105.790 74.400 105.930 ;
        RECT 47.875 105.450 48.640 105.590 ;
        RECT 47.875 105.405 48.165 105.450 ;
        RECT 48.320 105.390 48.640 105.450 ;
        RECT 48.795 105.590 49.085 105.635 ;
        RECT 49.255 105.590 49.545 105.635 ;
        RECT 48.795 105.450 49.545 105.590 ;
        RECT 48.795 105.405 49.085 105.450 ;
        RECT 49.255 105.405 49.545 105.450 ;
        RECT 50.175 105.405 50.465 105.635 ;
        RECT 50.250 105.250 50.390 105.405 ;
        RECT 51.080 105.390 51.400 105.650 ;
        RECT 51.540 105.390 51.860 105.650 ;
        RECT 52.460 105.590 52.780 105.650 ;
        RECT 52.935 105.590 53.225 105.635 ;
        RECT 52.460 105.450 53.225 105.590 ;
        RECT 52.460 105.390 52.780 105.450 ;
        RECT 52.935 105.405 53.225 105.450 ;
        RECT 54.300 105.590 54.620 105.650 ;
        RECT 55.235 105.590 55.525 105.635 ;
        RECT 54.300 105.450 55.525 105.590 ;
        RECT 54.300 105.390 54.620 105.450 ;
        RECT 55.235 105.405 55.525 105.450 ;
        RECT 55.695 105.405 55.985 105.635 ;
        RECT 53.395 105.250 53.685 105.295 ;
        RECT 50.250 105.110 53.685 105.250 ;
        RECT 53.395 105.065 53.685 105.110 ;
        RECT 51.540 104.910 51.860 104.970 ;
        RECT 55.770 104.910 55.910 105.405 ;
        RECT 63.960 105.390 64.280 105.650 ;
        RECT 64.435 105.590 64.725 105.635 ;
        RECT 66.260 105.590 66.580 105.650 ;
        RECT 66.810 105.635 66.950 105.790 ;
        RECT 74.080 105.730 74.400 105.790 ;
        RECT 87.510 105.790 90.040 105.930 ;
        RECT 64.435 105.450 66.580 105.590 ;
        RECT 64.435 105.405 64.725 105.450 ;
        RECT 66.260 105.390 66.580 105.450 ;
        RECT 66.735 105.405 67.025 105.635 ;
        RECT 69.480 105.390 69.800 105.650 ;
        RECT 70.400 105.390 70.720 105.650 ;
        RECT 75.460 105.390 75.780 105.650 ;
        RECT 87.510 105.635 87.650 105.790 ;
        RECT 89.720 105.730 90.040 105.790 ;
        RECT 105.360 105.930 105.680 105.990 ;
        RECT 109.975 105.930 110.265 105.975 ;
        RECT 105.360 105.790 108.350 105.930 ;
        RECT 105.360 105.730 105.680 105.790 ;
        RECT 108.210 105.650 108.350 105.790 ;
        RECT 108.670 105.790 110.265 105.930 ;
        RECT 88.800 105.635 89.120 105.650 ;
        RECT 87.435 105.405 87.725 105.635 ;
        RECT 88.770 105.405 89.120 105.635 ;
        RECT 88.800 105.390 89.120 105.405 ;
        RECT 96.160 105.390 96.480 105.650 ;
        RECT 96.620 105.390 96.940 105.650 ;
        RECT 97.555 105.405 97.845 105.635 ;
        RECT 98.015 105.405 98.305 105.635 ;
        RECT 65.355 105.065 65.645 105.295 ;
        RECT 67.195 105.250 67.485 105.295 ;
        RECT 71.320 105.250 71.640 105.310 ;
        RECT 71.795 105.250 72.085 105.295 ;
        RECT 67.195 105.110 70.170 105.250 ;
        RECT 67.195 105.065 67.485 105.110 ;
        RECT 51.540 104.770 55.910 104.910 ;
        RECT 51.540 104.710 51.860 104.770 ;
        RECT 54.300 104.570 54.620 104.630 ;
        RECT 46.110 104.430 54.620 104.570 ;
        RECT 29.460 104.370 29.780 104.430 ;
        RECT 32.235 104.385 32.525 104.430 ;
        RECT 54.300 104.370 54.620 104.430 ;
        RECT 54.775 104.570 55.065 104.615 ;
        RECT 55.770 104.570 55.910 104.770 ;
        RECT 54.775 104.430 55.910 104.570 ;
        RECT 65.430 104.570 65.570 105.065 ;
        RECT 70.030 104.970 70.170 105.110 ;
        RECT 71.320 105.110 72.085 105.250 ;
        RECT 71.320 105.050 71.640 105.110 ;
        RECT 71.795 105.065 72.085 105.110 ;
        RECT 72.240 105.250 72.560 105.310 ;
        RECT 73.635 105.250 73.925 105.295 ;
        RECT 72.240 105.110 73.925 105.250 ;
        RECT 72.240 105.050 72.560 105.110 ;
        RECT 73.635 105.065 73.925 105.110 ;
        RECT 74.080 105.050 74.400 105.310 ;
        RECT 75.015 105.250 75.305 105.295 ;
        RECT 79.140 105.250 79.460 105.310 ;
        RECT 75.015 105.110 79.460 105.250 ;
        RECT 75.015 105.065 75.305 105.110 ;
        RECT 79.140 105.050 79.460 105.110 ;
        RECT 88.315 105.250 88.605 105.295 ;
        RECT 89.505 105.250 89.795 105.295 ;
        RECT 92.025 105.250 92.315 105.295 ;
        RECT 88.315 105.110 92.315 105.250 ;
        RECT 88.315 105.065 88.605 105.110 ;
        RECT 89.505 105.065 89.795 105.110 ;
        RECT 92.025 105.065 92.315 105.110 ;
        RECT 68.560 104.710 68.880 104.970 ;
        RECT 69.940 104.710 70.260 104.970 ;
        RECT 74.555 104.910 74.845 104.955 ;
        RECT 71.410 104.770 74.845 104.910 ;
        RECT 71.410 104.570 71.550 104.770 ;
        RECT 74.555 104.725 74.845 104.770 ;
        RECT 87.920 104.910 88.210 104.955 ;
        RECT 90.020 104.910 90.310 104.955 ;
        RECT 91.590 104.910 91.880 104.955 ;
        RECT 87.920 104.770 91.880 104.910 ;
        RECT 97.630 104.910 97.770 105.405 ;
        RECT 98.090 105.250 98.230 105.405 ;
        RECT 107.660 105.390 107.980 105.650 ;
        RECT 108.120 105.390 108.440 105.650 ;
        RECT 108.670 105.635 108.810 105.790 ;
        RECT 109.975 105.745 110.265 105.790 ;
        RECT 108.595 105.405 108.885 105.635 ;
        RECT 109.040 105.590 109.360 105.650 ;
        RECT 109.515 105.590 109.805 105.635 ;
        RECT 109.040 105.450 109.805 105.590 ;
        RECT 109.040 105.390 109.360 105.450 ;
        RECT 109.515 105.405 109.805 105.450 ;
        RECT 110.880 105.390 111.200 105.650 ;
        RECT 111.890 105.635 112.030 106.130 ;
        RECT 115.955 106.130 117.180 106.270 ;
        RECT 115.955 106.085 116.245 106.130 ;
        RECT 116.860 106.070 117.180 106.130 ;
        RECT 117.870 106.130 122.240 106.270 ;
        RECT 114.100 105.930 114.420 105.990 ;
        RECT 114.100 105.790 117.550 105.930 ;
        RECT 114.100 105.730 114.420 105.790 ;
        RECT 116.030 105.650 116.170 105.790 ;
        RECT 111.815 105.590 112.105 105.635 ;
        RECT 113.655 105.590 113.945 105.635 ;
        RECT 111.815 105.450 113.945 105.590 ;
        RECT 111.815 105.405 112.105 105.450 ;
        RECT 113.655 105.405 113.945 105.450 ;
        RECT 98.090 105.110 112.490 105.250 ;
        RECT 111.800 104.910 112.120 104.970 ;
        RECT 97.630 104.770 112.120 104.910 ;
        RECT 87.920 104.725 88.210 104.770 ;
        RECT 90.020 104.725 90.310 104.770 ;
        RECT 91.590 104.725 91.880 104.770 ;
        RECT 111.800 104.710 112.120 104.770 ;
        RECT 65.430 104.430 71.550 104.570 ;
        RECT 54.775 104.385 55.065 104.430 ;
        RECT 71.780 104.370 72.100 104.630 ;
        RECT 94.335 104.570 94.625 104.615 ;
        RECT 96.620 104.570 96.940 104.630 ;
        RECT 94.335 104.430 96.940 104.570 ;
        RECT 94.335 104.385 94.625 104.430 ;
        RECT 96.620 104.370 96.940 104.430 ;
        RECT 106.295 104.570 106.585 104.615 ;
        RECT 108.580 104.570 108.900 104.630 ;
        RECT 106.295 104.430 108.900 104.570 ;
        RECT 112.350 104.570 112.490 105.110 ;
        RECT 113.730 104.910 113.870 105.405 ;
        RECT 114.560 105.390 114.880 105.650 ;
        RECT 115.940 105.390 116.260 105.650 ;
        RECT 117.410 105.635 117.550 105.790 ;
        RECT 117.870 105.635 118.010 106.130 ;
        RECT 121.920 106.070 122.240 106.130 ;
        RECT 129.830 106.130 133.740 106.270 ;
        RECT 121.000 105.730 121.320 105.990 ;
        RECT 128.360 105.930 128.680 105.990 ;
        RECT 129.830 105.930 129.970 106.130 ;
        RECT 133.420 106.070 133.740 106.130 ;
        RECT 137.100 106.270 137.420 106.330 ;
        RECT 138.495 106.270 138.785 106.315 ;
        RECT 139.860 106.270 140.180 106.330 ;
        RECT 137.100 106.130 140.180 106.270 ;
        RECT 137.100 106.070 137.420 106.130 ;
        RECT 138.495 106.085 138.785 106.130 ;
        RECT 139.860 106.070 140.180 106.130 ;
        RECT 140.795 106.270 141.085 106.315 ;
        RECT 142.620 106.270 142.940 106.330 ;
        RECT 140.795 106.130 142.940 106.270 ;
        RECT 140.795 106.085 141.085 106.130 ;
        RECT 142.620 106.070 142.940 106.130 ;
        RECT 128.360 105.790 129.970 105.930 ;
        RECT 128.360 105.730 128.680 105.790 ;
        RECT 117.335 105.405 117.625 105.635 ;
        RECT 117.795 105.405 118.085 105.635 ;
        RECT 118.255 105.405 118.545 105.635 ;
        RECT 119.160 105.590 119.480 105.650 ;
        RECT 127.915 105.590 128.205 105.635 ;
        RECT 119.160 105.450 128.205 105.590 ;
        RECT 116.860 105.250 117.180 105.310 ;
        RECT 117.870 105.250 118.010 105.405 ;
        RECT 116.860 105.110 118.010 105.250 ;
        RECT 118.330 105.250 118.470 105.405 ;
        RECT 119.160 105.390 119.480 105.450 ;
        RECT 127.915 105.405 128.205 105.450 ;
        RECT 128.835 105.405 129.125 105.635 ;
        RECT 124.220 105.250 124.540 105.310 ;
        RECT 118.330 105.110 124.540 105.250 ;
        RECT 116.860 105.050 117.180 105.110 ;
        RECT 124.220 105.050 124.540 105.110 ;
        RECT 125.140 105.050 125.460 105.310 ;
        RECT 122.840 104.910 123.160 104.970 ;
        RECT 113.730 104.770 123.160 104.910 ;
        RECT 128.910 104.910 129.050 105.405 ;
        RECT 129.280 105.390 129.600 105.650 ;
        RECT 129.830 105.635 129.970 105.790 ;
        RECT 131.120 105.930 131.440 105.990 ;
        RECT 132.820 105.930 133.110 105.975 ;
        RECT 131.120 105.790 133.110 105.930 ;
        RECT 131.120 105.730 131.440 105.790 ;
        RECT 132.820 105.745 133.110 105.790 ;
        RECT 129.755 105.405 130.045 105.635 ;
        RECT 131.580 105.390 131.900 105.650 ;
        RECT 132.040 105.390 132.360 105.650 ;
        RECT 135.260 105.590 135.580 105.650 ;
        RECT 139.875 105.590 140.165 105.635 ;
        RECT 140.320 105.590 140.640 105.650 ;
        RECT 135.260 105.450 140.640 105.590 ;
        RECT 135.260 105.390 135.580 105.450 ;
        RECT 139.875 105.405 140.165 105.450 ;
        RECT 140.320 105.390 140.640 105.450 ;
        RECT 131.135 105.250 131.425 105.295 ;
        RECT 132.130 105.250 132.270 105.390 ;
        RECT 131.135 105.110 132.270 105.250 ;
        RECT 132.475 105.250 132.765 105.295 ;
        RECT 133.665 105.250 133.955 105.295 ;
        RECT 136.185 105.250 136.475 105.295 ;
        RECT 132.475 105.110 136.475 105.250 ;
        RECT 131.135 105.065 131.425 105.110 ;
        RECT 132.475 105.065 132.765 105.110 ;
        RECT 133.665 105.065 133.955 105.110 ;
        RECT 136.185 105.065 136.475 105.110 ;
        RECT 129.280 104.910 129.600 104.970 ;
        RECT 128.910 104.770 129.600 104.910 ;
        RECT 122.840 104.710 123.160 104.770 ;
        RECT 129.280 104.710 129.600 104.770 ;
        RECT 132.080 104.910 132.370 104.955 ;
        RECT 134.180 104.910 134.470 104.955 ;
        RECT 135.750 104.910 136.040 104.955 ;
        RECT 132.080 104.770 136.040 104.910 ;
        RECT 132.080 104.725 132.370 104.770 ;
        RECT 134.180 104.725 134.470 104.770 ;
        RECT 135.750 104.725 136.040 104.770 ;
        RECT 115.020 104.570 115.340 104.630 ;
        RECT 112.350 104.430 115.340 104.570 ;
        RECT 106.295 104.385 106.585 104.430 ;
        RECT 108.580 104.370 108.900 104.430 ;
        RECT 115.020 104.370 115.340 104.430 ;
        RECT 115.495 104.570 115.785 104.615 ;
        RECT 116.400 104.570 116.720 104.630 ;
        RECT 115.495 104.430 116.720 104.570 ;
        RECT 115.495 104.385 115.785 104.430 ;
        RECT 116.400 104.370 116.720 104.430 ;
        RECT 17.430 103.750 143.010 104.230 ;
        RECT 48.795 103.550 49.085 103.595 ;
        RECT 51.080 103.550 51.400 103.610 ;
        RECT 65.815 103.550 66.105 103.595 ;
        RECT 69.020 103.550 69.340 103.610 ;
        RECT 71.780 103.550 72.100 103.610 ;
        RECT 48.795 103.410 55.910 103.550 ;
        RECT 48.795 103.365 49.085 103.410 ;
        RECT 51.080 103.350 51.400 103.410 ;
        RECT 22.140 103.210 22.430 103.255 ;
        RECT 24.240 103.210 24.530 103.255 ;
        RECT 25.810 103.210 26.100 103.255 ;
        RECT 22.140 103.070 26.100 103.210 ;
        RECT 22.140 103.025 22.430 103.070 ;
        RECT 24.240 103.025 24.530 103.070 ;
        RECT 25.810 103.025 26.100 103.070 ;
        RECT 51.540 103.210 51.830 103.255 ;
        RECT 53.110 103.210 53.400 103.255 ;
        RECT 55.210 103.210 55.500 103.255 ;
        RECT 51.540 103.070 55.500 103.210 ;
        RECT 51.540 103.025 51.830 103.070 ;
        RECT 53.110 103.025 53.400 103.070 ;
        RECT 55.210 103.025 55.500 103.070 ;
        RECT 21.640 102.670 21.960 102.930 ;
        RECT 22.535 102.870 22.825 102.915 ;
        RECT 23.725 102.870 24.015 102.915 ;
        RECT 26.245 102.870 26.535 102.915 ;
        RECT 22.535 102.730 26.535 102.870 ;
        RECT 22.535 102.685 22.825 102.730 ;
        RECT 23.725 102.685 24.015 102.730 ;
        RECT 26.245 102.685 26.535 102.730 ;
        RECT 29.920 102.870 30.240 102.930 ;
        RECT 33.615 102.870 33.905 102.915 ;
        RECT 29.920 102.730 33.905 102.870 ;
        RECT 29.920 102.670 30.240 102.730 ;
        RECT 33.615 102.685 33.905 102.730 ;
        RECT 51.105 102.870 51.395 102.915 ;
        RECT 53.625 102.870 53.915 102.915 ;
        RECT 54.815 102.870 55.105 102.915 ;
        RECT 51.105 102.730 55.105 102.870 ;
        RECT 55.770 102.870 55.910 103.410 ;
        RECT 65.815 103.410 72.100 103.550 ;
        RECT 65.815 103.365 66.105 103.410 ;
        RECT 69.020 103.350 69.340 103.410 ;
        RECT 71.780 103.350 72.100 103.410 ;
        RECT 74.095 103.550 74.385 103.595 ;
        RECT 75.000 103.550 75.320 103.610 ;
        RECT 74.095 103.410 75.320 103.550 ;
        RECT 74.095 103.365 74.385 103.410 ;
        RECT 75.000 103.350 75.320 103.410 ;
        RECT 83.280 103.550 83.600 103.610 ;
        RECT 86.515 103.550 86.805 103.595 ;
        RECT 83.280 103.410 86.805 103.550 ;
        RECT 83.280 103.350 83.600 103.410 ;
        RECT 86.515 103.365 86.805 103.410 ;
        RECT 92.480 103.550 92.800 103.610 ;
        RECT 107.660 103.550 107.980 103.610 ;
        RECT 109.040 103.550 109.360 103.610 ;
        RECT 92.480 103.410 107.980 103.550 ;
        RECT 92.480 103.350 92.800 103.410 ;
        RECT 107.660 103.350 107.980 103.410 ;
        RECT 108.210 103.410 115.710 103.550 ;
        RECT 67.180 103.210 67.500 103.270 ;
        RECT 66.350 103.070 67.500 103.210 ;
        RECT 56.615 102.870 56.905 102.915 ;
        RECT 55.770 102.730 56.905 102.870 ;
        RECT 51.105 102.685 51.395 102.730 ;
        RECT 53.625 102.685 53.915 102.730 ;
        RECT 54.815 102.685 55.105 102.730 ;
        RECT 56.615 102.685 56.905 102.730 ;
        RECT 28.080 102.530 28.400 102.590 ;
        RECT 31.300 102.530 31.620 102.590 ;
        RECT 31.775 102.530 32.065 102.575 ;
        RECT 28.080 102.390 32.065 102.530 ;
        RECT 28.080 102.330 28.400 102.390 ;
        RECT 31.300 102.330 31.620 102.390 ;
        RECT 31.775 102.345 32.065 102.390 ;
        RECT 32.680 102.530 33.000 102.590 ;
        RECT 34.980 102.530 35.300 102.590 ;
        RECT 32.680 102.390 35.300 102.530 ;
        RECT 32.680 102.330 33.000 102.390 ;
        RECT 34.980 102.330 35.300 102.390 ;
        RECT 40.960 102.530 41.280 102.590 ;
        RECT 47.415 102.530 47.705 102.575 ;
        RECT 40.960 102.390 47.705 102.530 ;
        RECT 40.960 102.330 41.280 102.390 ;
        RECT 47.415 102.345 47.705 102.390 ;
        RECT 55.680 102.330 56.000 102.590 ;
        RECT 59.835 102.530 60.125 102.575 ;
        RECT 60.295 102.530 60.585 102.575 ;
        RECT 59.835 102.390 60.585 102.530 ;
        RECT 59.835 102.345 60.125 102.390 ;
        RECT 60.295 102.345 60.585 102.390 ;
        RECT 65.355 102.530 65.645 102.575 ;
        RECT 66.350 102.530 66.490 103.070 ;
        RECT 67.180 103.010 67.500 103.070 ;
        RECT 67.680 103.210 67.970 103.255 ;
        RECT 69.780 103.210 70.070 103.255 ;
        RECT 71.350 103.210 71.640 103.255 ;
        RECT 101.695 103.210 101.985 103.255 ;
        RECT 104.900 103.210 105.220 103.270 ;
        RECT 67.680 103.070 71.640 103.210 ;
        RECT 67.680 103.025 67.970 103.070 ;
        RECT 69.780 103.025 70.070 103.070 ;
        RECT 71.350 103.025 71.640 103.070 ;
        RECT 87.050 103.070 96.850 103.210 ;
        RECT 66.720 102.670 67.040 102.930 ;
        RECT 67.270 102.870 67.410 103.010 ;
        RECT 68.075 102.870 68.365 102.915 ;
        RECT 69.265 102.870 69.555 102.915 ;
        RECT 71.785 102.870 72.075 102.915 ;
        RECT 67.270 102.730 67.870 102.870 ;
        RECT 65.355 102.390 66.490 102.530 ;
        RECT 65.355 102.345 65.645 102.390 ;
        RECT 67.195 102.345 67.485 102.575 ;
        RECT 22.990 102.190 23.280 102.235 ;
        RECT 23.480 102.190 23.800 102.250 ;
        RECT 22.990 102.050 23.800 102.190 ;
        RECT 22.990 102.005 23.280 102.050 ;
        RECT 23.480 101.990 23.800 102.050 ;
        RECT 27.620 102.190 27.940 102.250 ;
        RECT 30.855 102.190 31.145 102.235 ;
        RECT 32.235 102.190 32.525 102.235 ;
        RECT 27.620 102.050 31.145 102.190 ;
        RECT 27.620 101.990 27.940 102.050 ;
        RECT 30.855 102.005 31.145 102.050 ;
        RECT 31.390 102.050 32.525 102.190 ;
        RECT 22.560 101.850 22.880 101.910 ;
        RECT 28.555 101.850 28.845 101.895 ;
        RECT 30.380 101.850 30.700 101.910 ;
        RECT 31.390 101.850 31.530 102.050 ;
        RECT 32.235 102.005 32.525 102.050 ;
        RECT 54.470 102.190 54.760 102.235 ;
        RECT 56.140 102.190 56.460 102.250 ;
        RECT 54.470 102.050 56.460 102.190 ;
        RECT 54.470 102.005 54.760 102.050 ;
        RECT 56.140 101.990 56.460 102.050 ;
        RECT 64.420 102.190 64.740 102.250 ;
        RECT 67.270 102.190 67.410 102.345 ;
        RECT 64.420 102.050 67.410 102.190 ;
        RECT 67.730 102.190 67.870 102.730 ;
        RECT 68.075 102.730 72.075 102.870 ;
        RECT 68.075 102.685 68.365 102.730 ;
        RECT 69.265 102.685 69.555 102.730 ;
        RECT 71.785 102.685 72.075 102.730 ;
        RECT 68.560 102.575 68.880 102.590 ;
        RECT 68.530 102.530 68.880 102.575 ;
        RECT 68.365 102.390 68.880 102.530 ;
        RECT 68.530 102.345 68.880 102.390 ;
        RECT 68.560 102.330 68.880 102.345 ;
        RECT 80.980 102.530 81.300 102.590 ;
        RECT 82.375 102.530 82.665 102.575 ;
        RECT 85.120 102.530 85.440 102.590 ;
        RECT 87.050 102.530 87.190 103.070 ;
        RECT 96.160 102.870 96.480 102.930 ;
        RECT 87.510 102.730 96.480 102.870 ;
        RECT 96.710 102.870 96.850 103.070 ;
        RECT 101.695 103.070 105.220 103.210 ;
        RECT 101.695 103.025 101.985 103.070 ;
        RECT 104.900 103.010 105.220 103.070 ;
        RECT 106.280 102.870 106.600 102.930 ;
        RECT 108.210 102.870 108.350 103.410 ;
        RECT 109.040 103.350 109.360 103.410 ;
        RECT 108.620 103.210 108.910 103.255 ;
        RECT 110.720 103.210 111.010 103.255 ;
        RECT 112.290 103.210 112.580 103.255 ;
        RECT 108.620 103.070 112.580 103.210 ;
        RECT 108.620 103.025 108.910 103.070 ;
        RECT 110.720 103.025 111.010 103.070 ;
        RECT 112.290 103.025 112.580 103.070 ;
        RECT 96.710 102.730 97.770 102.870 ;
        RECT 87.510 102.590 87.650 102.730 ;
        RECT 96.160 102.670 96.480 102.730 ;
        RECT 80.980 102.390 87.190 102.530 ;
        RECT 80.980 102.330 81.300 102.390 ;
        RECT 82.375 102.345 82.665 102.390 ;
        RECT 85.120 102.330 85.440 102.390 ;
        RECT 87.420 102.330 87.740 102.590 ;
        RECT 87.895 102.345 88.185 102.575 ;
        RECT 88.815 102.345 89.105 102.575 ;
        RECT 71.320 102.190 71.640 102.250 ;
        RECT 67.730 102.050 71.640 102.190 ;
        RECT 64.420 101.990 64.740 102.050 ;
        RECT 71.320 101.990 71.640 102.050 ;
        RECT 83.280 102.190 83.600 102.250 ;
        RECT 87.970 102.190 88.110 102.345 ;
        RECT 83.280 102.050 88.110 102.190 ;
        RECT 83.280 101.990 83.600 102.050 ;
        RECT 22.560 101.710 31.530 101.850 ;
        RECT 34.980 101.850 35.300 101.910 ;
        RECT 47.875 101.850 48.165 101.895 ;
        RECT 50.620 101.850 50.940 101.910 ;
        RECT 34.980 101.710 50.940 101.850 ;
        RECT 22.560 101.650 22.880 101.710 ;
        RECT 28.555 101.665 28.845 101.710 ;
        RECT 30.380 101.650 30.700 101.710 ;
        RECT 34.980 101.650 35.300 101.710 ;
        RECT 47.875 101.665 48.165 101.710 ;
        RECT 50.620 101.650 50.940 101.710 ;
        RECT 52.460 101.850 52.780 101.910 ;
        RECT 60.755 101.850 61.045 101.895 ;
        RECT 52.460 101.710 61.045 101.850 ;
        RECT 52.460 101.650 52.780 101.710 ;
        RECT 60.755 101.665 61.045 101.710 ;
        RECT 66.735 101.850 67.025 101.895 ;
        RECT 68.560 101.850 68.880 101.910 ;
        RECT 66.735 101.710 68.880 101.850 ;
        RECT 66.735 101.665 67.025 101.710 ;
        RECT 68.560 101.650 68.880 101.710 ;
        RECT 84.215 101.850 84.505 101.895 ;
        RECT 84.660 101.850 84.980 101.910 ;
        RECT 84.215 101.710 84.980 101.850 ;
        RECT 88.890 101.850 89.030 102.345 ;
        RECT 89.260 102.330 89.580 102.590 ;
        RECT 95.240 102.330 95.560 102.590 ;
        RECT 97.630 102.575 97.770 102.730 ;
        RECT 104.025 102.730 108.350 102.870 ;
        RECT 109.015 102.870 109.305 102.915 ;
        RECT 110.205 102.870 110.495 102.915 ;
        RECT 112.725 102.870 113.015 102.915 ;
        RECT 109.015 102.730 113.015 102.870 ;
        RECT 97.555 102.530 97.845 102.575 ;
        RECT 102.140 102.530 102.460 102.590 ;
        RECT 104.025 102.575 104.165 102.730 ;
        RECT 106.280 102.670 106.600 102.730 ;
        RECT 109.015 102.685 109.305 102.730 ;
        RECT 110.205 102.685 110.495 102.730 ;
        RECT 112.725 102.685 113.015 102.730 ;
        RECT 115.570 102.870 115.710 103.410 ;
        RECT 119.620 103.350 119.940 103.610 ;
        RECT 132.960 103.550 133.280 103.610 ;
        RECT 134.800 103.550 135.120 103.610 ;
        RECT 123.850 103.410 135.120 103.550 ;
        RECT 119.160 102.870 119.480 102.930 ;
        RECT 115.570 102.730 119.480 102.870 ;
        RECT 119.710 102.870 119.850 103.350 ;
        RECT 123.850 102.870 123.990 103.410 ;
        RECT 132.960 103.350 133.280 103.410 ;
        RECT 134.800 103.350 135.120 103.410 ;
        RECT 135.260 103.210 135.580 103.270 ;
        RECT 130.290 103.070 135.580 103.210 ;
        RECT 119.710 102.730 123.990 102.870 ;
        RECT 97.555 102.390 102.460 102.530 ;
        RECT 97.555 102.345 97.845 102.390 ;
        RECT 102.140 102.330 102.460 102.390 ;
        RECT 103.935 102.345 104.225 102.575 ;
        RECT 104.900 102.330 105.220 102.590 ;
        RECT 105.360 102.330 105.680 102.590 ;
        RECT 105.820 102.330 106.140 102.590 ;
        RECT 107.660 102.530 107.980 102.590 ;
        RECT 115.570 102.575 115.710 102.730 ;
        RECT 119.160 102.670 119.480 102.730 ;
        RECT 108.135 102.530 108.425 102.575 ;
        RECT 107.660 102.390 108.425 102.530 ;
        RECT 107.660 102.330 107.980 102.390 ;
        RECT 108.135 102.345 108.425 102.390 ;
        RECT 115.495 102.345 115.785 102.575 ;
        RECT 116.400 102.330 116.720 102.590 ;
        RECT 116.860 102.330 117.180 102.590 ;
        RECT 117.335 102.345 117.625 102.575 ;
        RECT 118.240 102.530 118.560 102.590 ;
        RECT 123.850 102.575 123.990 102.730 ;
        RECT 124.220 102.870 124.540 102.930 ;
        RECT 125.155 102.870 125.445 102.915 ;
        RECT 124.220 102.730 125.445 102.870 ;
        RECT 124.220 102.670 124.540 102.730 ;
        RECT 125.155 102.685 125.445 102.730 ;
        RECT 129.280 102.670 129.600 102.930 ;
        RECT 122.855 102.530 123.145 102.575 ;
        RECT 118.240 102.390 123.145 102.530 ;
        RECT 89.720 102.190 90.040 102.250 ;
        RECT 91.115 102.190 91.405 102.235 ;
        RECT 89.720 102.050 91.405 102.190 ;
        RECT 89.720 101.990 90.040 102.050 ;
        RECT 91.115 102.005 91.405 102.050 ;
        RECT 96.160 102.190 96.480 102.250 ;
        RECT 96.635 102.190 96.925 102.235 ;
        RECT 96.160 102.050 96.925 102.190 ;
        RECT 96.160 101.990 96.480 102.050 ;
        RECT 96.635 102.005 96.925 102.050 ;
        RECT 102.615 102.005 102.905 102.235 ;
        RECT 103.535 102.190 103.825 102.235 ;
        RECT 106.740 102.190 107.060 102.250 ;
        RECT 103.535 102.050 107.060 102.190 ;
        RECT 103.535 102.005 103.825 102.050 ;
        RECT 91.560 101.850 91.880 101.910 ;
        RECT 88.890 101.710 91.880 101.850 ;
        RECT 84.215 101.665 84.505 101.710 ;
        RECT 84.660 101.650 84.980 101.710 ;
        RECT 91.560 101.650 91.880 101.710 ;
        RECT 92.020 101.850 92.340 101.910 ;
        RECT 95.715 101.850 96.005 101.895 ;
        RECT 92.020 101.710 96.005 101.850 ;
        RECT 92.020 101.650 92.340 101.710 ;
        RECT 95.715 101.665 96.005 101.710 ;
        RECT 101.680 101.850 102.000 101.910 ;
        RECT 102.690 101.850 102.830 102.005 ;
        RECT 106.740 101.990 107.060 102.050 ;
        RECT 107.215 102.190 107.505 102.235 ;
        RECT 109.360 102.190 109.650 102.235 ;
        RECT 107.215 102.050 109.650 102.190 ;
        RECT 117.410 102.190 117.550 102.345 ;
        RECT 118.240 102.330 118.560 102.390 ;
        RECT 122.855 102.345 123.145 102.390 ;
        RECT 123.775 102.345 124.065 102.575 ;
        RECT 124.695 102.530 124.985 102.575 ;
        RECT 126.520 102.530 126.840 102.590 ;
        RECT 130.290 102.575 130.430 103.070 ;
        RECT 135.260 103.010 135.580 103.070 ;
        RECT 124.695 102.390 129.970 102.530 ;
        RECT 124.695 102.345 124.985 102.390 ;
        RECT 126.520 102.330 126.840 102.390 ;
        RECT 120.540 102.190 120.860 102.250 ;
        RECT 117.410 102.050 120.860 102.190 ;
        RECT 107.215 102.005 107.505 102.050 ;
        RECT 109.360 102.005 109.650 102.050 ;
        RECT 120.540 101.990 120.860 102.050 ;
        RECT 122.380 102.190 122.700 102.250 ;
        RECT 126.075 102.190 126.365 102.235 ;
        RECT 122.380 102.050 126.365 102.190 ;
        RECT 122.380 101.990 122.700 102.050 ;
        RECT 126.075 102.005 126.365 102.050 ;
        RECT 115.035 101.850 115.325 101.895 ;
        RECT 115.480 101.850 115.800 101.910 ;
        RECT 101.680 101.710 115.800 101.850 ;
        RECT 101.680 101.650 102.000 101.710 ;
        RECT 115.035 101.665 115.325 101.710 ;
        RECT 115.480 101.650 115.800 101.710 ;
        RECT 118.700 101.650 119.020 101.910 ;
        RECT 126.150 101.850 126.290 102.005 ;
        RECT 126.980 101.990 127.300 102.250 ;
        RECT 129.830 102.190 129.970 102.390 ;
        RECT 130.215 102.345 130.505 102.575 ;
        RECT 134.800 102.330 135.120 102.590 ;
        RECT 135.260 102.330 135.580 102.590 ;
        RECT 136.640 102.330 136.960 102.590 ;
        RECT 138.035 102.345 138.325 102.575 ;
        RECT 131.135 102.190 131.425 102.235 ;
        RECT 129.830 102.050 131.425 102.190 ;
        RECT 131.135 102.005 131.425 102.050 ;
        RECT 131.670 102.050 134.570 102.190 ;
        RECT 131.670 101.850 131.810 102.050 ;
        RECT 126.150 101.710 131.810 101.850 ;
        RECT 133.880 101.650 134.200 101.910 ;
        RECT 134.430 101.850 134.570 102.050 ;
        RECT 135.720 101.990 136.040 102.250 ;
        RECT 138.110 101.850 138.250 102.345 ;
        RECT 139.860 102.330 140.180 102.590 ;
        RECT 134.430 101.710 138.250 101.850 ;
        RECT 138.940 101.650 139.260 101.910 ;
        RECT 140.780 101.650 141.100 101.910 ;
        RECT 17.430 101.030 143.010 101.510 ;
        RECT 23.035 100.645 23.325 100.875 ;
        RECT 22.560 100.290 22.880 100.550 ;
        RECT 23.110 100.490 23.250 100.645 ;
        RECT 23.480 100.630 23.800 100.890 ;
        RECT 25.780 100.630 26.100 100.890 ;
        RECT 31.315 100.830 31.605 100.875 ;
        RECT 32.220 100.830 32.540 100.890 ;
        RECT 26.790 100.690 32.540 100.830 ;
        RECT 24.255 100.490 24.545 100.535 ;
        RECT 23.110 100.350 24.545 100.490 ;
        RECT 24.255 100.305 24.545 100.350 ;
        RECT 25.335 100.490 25.625 100.535 ;
        RECT 26.790 100.490 26.930 100.690 ;
        RECT 31.315 100.645 31.605 100.690 ;
        RECT 32.220 100.630 32.540 100.690 ;
        RECT 41.895 100.830 42.185 100.875 ;
        RECT 44.180 100.830 44.500 100.890 ;
        RECT 41.895 100.690 44.500 100.830 ;
        RECT 41.895 100.645 42.185 100.690 ;
        RECT 44.180 100.630 44.500 100.690 ;
        RECT 44.640 100.630 44.960 100.890 ;
        RECT 52.460 100.630 52.780 100.890 ;
        RECT 56.140 100.830 56.460 100.890 ;
        RECT 56.615 100.830 56.905 100.875 ;
        RECT 66.720 100.830 67.040 100.890 ;
        RECT 82.820 100.830 83.140 100.890 ;
        RECT 56.140 100.690 56.905 100.830 ;
        RECT 56.140 100.630 56.460 100.690 ;
        RECT 56.615 100.645 56.905 100.690 ;
        RECT 66.350 100.690 83.140 100.830 ;
        RECT 34.980 100.490 35.300 100.550 ;
        RECT 37.755 100.490 38.045 100.535 ;
        RECT 25.335 100.350 26.930 100.490 ;
        RECT 27.250 100.350 30.610 100.490 ;
        RECT 25.335 100.305 25.625 100.350 ;
        RECT 21.655 99.965 21.945 100.195 ;
        RECT 23.035 100.150 23.325 100.195 ;
        RECT 24.860 100.150 25.180 100.210 ;
        RECT 27.250 100.195 27.390 100.350 ;
        RECT 30.470 100.210 30.610 100.350 ;
        RECT 34.980 100.350 38.045 100.490 ;
        RECT 34.980 100.290 35.300 100.350 ;
        RECT 37.755 100.305 38.045 100.350 ;
        RECT 38.200 100.490 38.520 100.550 ;
        RECT 38.755 100.490 39.045 100.535 ;
        RECT 44.730 100.490 44.870 100.630 ;
        RECT 51.540 100.490 51.860 100.550 ;
        RECT 38.200 100.350 39.045 100.490 ;
        RECT 38.200 100.290 38.520 100.350 ;
        RECT 38.755 100.305 39.045 100.350 ;
        RECT 41.050 100.350 44.870 100.490 ;
        RECT 48.870 100.350 51.860 100.490 ;
        RECT 23.035 100.010 25.180 100.150 ;
        RECT 23.035 99.965 23.325 100.010 ;
        RECT 21.730 99.810 21.870 99.965 ;
        RECT 24.860 99.950 25.180 100.010 ;
        RECT 27.175 99.965 27.465 100.195 ;
        RECT 27.620 99.950 27.940 100.210 ;
        RECT 28.080 99.950 28.400 100.210 ;
        RECT 29.000 99.950 29.320 100.210 ;
        RECT 29.475 99.965 29.765 100.195 ;
        RECT 26.715 99.810 27.005 99.855 ;
        RECT 21.730 99.670 27.005 99.810 ;
        RECT 27.710 99.810 27.850 99.950 ;
        RECT 29.550 99.810 29.690 99.965 ;
        RECT 30.380 99.950 30.700 100.210 ;
        RECT 41.050 100.195 41.190 100.350 ;
        RECT 40.975 99.965 41.265 100.195 ;
        RECT 42.340 99.950 42.660 100.210 ;
        RECT 43.735 100.150 44.025 100.195 ;
        RECT 44.180 100.150 44.500 100.210 ;
        RECT 48.870 100.195 49.010 100.350 ;
        RECT 51.540 100.290 51.860 100.350 ;
        RECT 53.380 100.490 53.700 100.550 ;
        RECT 57.075 100.490 57.365 100.535 ;
        RECT 53.380 100.350 57.365 100.490 ;
        RECT 53.380 100.290 53.700 100.350 ;
        RECT 57.075 100.305 57.365 100.350 ;
        RECT 58.915 100.490 59.205 100.535 ;
        RECT 60.135 100.490 60.425 100.535 ;
        RECT 58.915 100.350 60.425 100.490 ;
        RECT 58.915 100.305 59.205 100.350 ;
        RECT 60.135 100.305 60.425 100.350 ;
        RECT 61.215 100.305 61.505 100.535 ;
        RECT 43.735 100.010 44.500 100.150 ;
        RECT 43.735 99.965 44.025 100.010 ;
        RECT 44.180 99.950 44.500 100.010 ;
        RECT 44.655 99.965 44.945 100.195 ;
        RECT 48.795 99.965 49.085 100.195 ;
        RECT 27.710 99.670 29.690 99.810 ;
        RECT 42.430 99.810 42.570 99.950 ;
        RECT 44.730 99.810 44.870 99.965 ;
        RECT 49.240 99.950 49.560 100.210 ;
        RECT 50.620 99.950 50.940 100.210 ;
        RECT 52.935 100.150 53.225 100.195 ;
        RECT 53.840 100.150 54.160 100.210 ;
        RECT 52.935 100.010 54.160 100.150 ;
        RECT 52.935 99.965 53.225 100.010 ;
        RECT 53.840 99.950 54.160 100.010 ;
        RECT 54.300 100.150 54.620 100.210 ;
        RECT 56.600 100.150 56.920 100.210 ;
        RECT 57.995 100.150 58.285 100.195 ;
        RECT 54.300 100.010 58.285 100.150 ;
        RECT 54.300 99.950 54.620 100.010 ;
        RECT 56.600 99.950 56.920 100.010 ;
        RECT 57.995 99.965 58.285 100.010 ;
        RECT 58.440 100.150 58.760 100.210 ;
        RECT 61.290 100.150 61.430 100.305 ;
        RECT 66.350 100.195 66.490 100.690 ;
        RECT 66.720 100.630 67.040 100.690 ;
        RECT 82.820 100.630 83.140 100.690 ;
        RECT 88.800 100.830 89.120 100.890 ;
        RECT 89.735 100.830 90.025 100.875 ;
        RECT 88.800 100.690 90.025 100.830 ;
        RECT 88.800 100.630 89.120 100.690 ;
        RECT 89.735 100.645 90.025 100.690 ;
        RECT 91.560 100.830 91.880 100.890 ;
        RECT 95.255 100.830 95.545 100.875 ;
        RECT 133.880 100.830 134.200 100.890 ;
        RECT 91.560 100.690 95.545 100.830 ;
        RECT 91.560 100.630 91.880 100.690 ;
        RECT 95.255 100.645 95.545 100.690 ;
        RECT 105.910 100.690 134.200 100.830 ;
        RECT 67.195 100.490 67.485 100.535 ;
        RECT 72.240 100.490 72.560 100.550 ;
        RECT 89.260 100.490 89.580 100.550 ;
        RECT 105.910 100.490 106.050 100.690 ;
        RECT 133.880 100.630 134.200 100.690 ;
        RECT 108.580 100.535 108.900 100.550 ;
        RECT 108.550 100.490 108.900 100.535 ;
        RECT 129.755 100.490 130.045 100.535 ;
        RECT 131.440 100.490 131.730 100.535 ;
        RECT 67.195 100.350 72.560 100.490 ;
        RECT 67.195 100.305 67.485 100.350 ;
        RECT 72.240 100.290 72.560 100.350 ;
        RECT 78.310 100.350 83.050 100.490 ;
        RECT 58.440 100.010 61.430 100.150 ;
        RECT 58.440 99.950 58.760 100.010 ;
        RECT 66.275 99.965 66.565 100.195 ;
        RECT 66.720 99.950 67.040 100.210 ;
        RECT 78.310 100.195 78.450 100.350 ;
        RECT 67.885 100.150 68.175 100.195 ;
        RECT 70.875 100.150 71.165 100.195 ;
        RECT 67.885 100.010 71.165 100.150 ;
        RECT 67.885 99.965 68.175 100.010 ;
        RECT 70.875 99.965 71.165 100.010 ;
        RECT 78.235 99.965 78.525 100.195 ;
        RECT 79.570 100.150 79.860 100.195 ;
        RECT 82.360 100.150 82.680 100.210 ;
        RECT 79.570 100.010 82.680 100.150 ;
        RECT 82.910 100.150 83.050 100.350 ;
        RECT 89.260 100.350 106.050 100.490 ;
        RECT 108.385 100.350 108.900 100.490 ;
        RECT 89.260 100.290 89.580 100.350 ;
        RECT 108.550 100.305 108.900 100.350 ;
        RECT 108.580 100.290 108.900 100.305 ;
        RECT 122.240 100.350 129.050 100.490 ;
        RECT 89.720 100.150 90.040 100.210 ;
        RECT 82.910 100.010 90.040 100.150 ;
        RECT 79.570 99.965 79.860 100.010 ;
        RECT 82.360 99.950 82.680 100.010 ;
        RECT 89.720 99.950 90.040 100.010 ;
        RECT 91.100 99.950 91.420 100.210 ;
        RECT 91.560 99.950 91.880 100.210 ;
        RECT 92.020 99.950 92.340 100.210 ;
        RECT 92.955 99.965 93.245 100.195 ;
        RECT 95.700 100.150 96.020 100.210 ;
        RECT 96.175 100.150 96.465 100.195 ;
        RECT 95.700 100.010 96.465 100.150 ;
        RECT 42.430 99.670 44.870 99.810 ;
        RECT 51.555 99.810 51.845 99.855 ;
        RECT 53.395 99.810 53.685 99.855 ;
        RECT 51.555 99.670 53.685 99.810 ;
        RECT 24.950 99.190 25.090 99.670 ;
        RECT 26.715 99.625 27.005 99.670 ;
        RECT 51.555 99.625 51.845 99.670 ;
        RECT 53.395 99.625 53.685 99.670 ;
        RECT 26.790 99.470 26.930 99.625 ;
        RECT 68.560 99.610 68.880 99.870 ;
        RECT 71.780 99.810 72.100 99.870 ;
        RECT 73.635 99.810 73.925 99.855 ;
        RECT 71.780 99.670 73.925 99.810 ;
        RECT 71.780 99.610 72.100 99.670 ;
        RECT 73.635 99.625 73.925 99.670 ;
        RECT 79.115 99.810 79.405 99.855 ;
        RECT 80.305 99.810 80.595 99.855 ;
        RECT 82.825 99.810 83.115 99.855 ;
        RECT 79.115 99.670 83.115 99.810 ;
        RECT 79.115 99.625 79.405 99.670 ;
        RECT 80.305 99.625 80.595 99.670 ;
        RECT 82.825 99.625 83.115 99.670 ;
        RECT 85.580 99.810 85.900 99.870 ;
        RECT 93.030 99.810 93.170 99.965 ;
        RECT 95.700 99.950 96.020 100.010 ;
        RECT 96.175 99.965 96.465 100.010 ;
        RECT 96.620 99.950 96.940 100.210 ;
        RECT 97.080 99.950 97.400 100.210 ;
        RECT 98.015 100.150 98.305 100.195 ;
        RECT 110.880 100.150 111.200 100.210 ;
        RECT 98.015 100.010 111.200 100.150 ;
        RECT 98.015 99.965 98.305 100.010 ;
        RECT 110.880 99.950 111.200 100.010 ;
        RECT 118.240 99.950 118.560 100.210 ;
        RECT 118.715 99.965 119.005 100.195 ;
        RECT 119.160 100.150 119.480 100.210 ;
        RECT 120.540 100.150 120.860 100.210 ;
        RECT 122.240 100.150 122.380 100.350 ;
        RECT 119.160 100.010 122.380 100.150 ;
        RECT 126.535 100.150 126.825 100.195 ;
        RECT 126.980 100.150 127.300 100.210 ;
        RECT 126.535 100.010 127.300 100.150 ;
        RECT 93.860 99.810 94.180 99.870 ;
        RECT 97.170 99.810 97.310 99.950 ;
        RECT 85.580 99.670 94.180 99.810 ;
        RECT 85.580 99.610 85.900 99.670 ;
        RECT 93.860 99.610 94.180 99.670 ;
        RECT 96.710 99.670 97.310 99.810 ;
        RECT 29.000 99.470 29.320 99.530 ;
        RECT 32.680 99.470 33.000 99.530 ;
        RECT 44.195 99.470 44.485 99.515 ;
        RECT 26.790 99.330 33.000 99.470 ;
        RECT 29.000 99.270 29.320 99.330 ;
        RECT 32.680 99.270 33.000 99.330 ;
        RECT 38.750 99.330 44.485 99.470 ;
        RECT 24.400 98.930 24.720 99.190 ;
        RECT 24.860 98.930 25.180 99.190 ;
        RECT 38.750 99.175 38.890 99.330 ;
        RECT 44.195 99.285 44.485 99.330 ;
        RECT 53.840 99.470 54.160 99.530 ;
        RECT 78.720 99.470 79.010 99.515 ;
        RECT 80.820 99.470 81.110 99.515 ;
        RECT 82.390 99.470 82.680 99.515 ;
        RECT 53.840 99.330 60.510 99.470 ;
        RECT 53.840 99.270 54.160 99.330 ;
        RECT 38.675 98.945 38.965 99.175 ;
        RECT 39.580 98.930 39.900 99.190 ;
        RECT 40.055 99.130 40.345 99.175 ;
        RECT 40.500 99.130 40.820 99.190 ;
        RECT 40.055 98.990 40.820 99.130 ;
        RECT 40.055 98.945 40.345 98.990 ;
        RECT 40.500 98.930 40.820 98.990 ;
        RECT 50.175 99.130 50.465 99.175 ;
        RECT 53.380 99.130 53.700 99.190 ;
        RECT 50.175 98.990 53.700 99.130 ;
        RECT 50.175 98.945 50.465 98.990 ;
        RECT 53.380 98.930 53.700 98.990 ;
        RECT 59.360 98.930 59.680 99.190 ;
        RECT 60.370 99.175 60.510 99.330 ;
        RECT 78.720 99.330 82.680 99.470 ;
        RECT 78.720 99.285 79.010 99.330 ;
        RECT 80.820 99.285 81.110 99.330 ;
        RECT 82.390 99.285 82.680 99.330 ;
        RECT 84.200 99.470 84.520 99.530 ;
        RECT 92.940 99.470 93.260 99.530 ;
        RECT 96.710 99.470 96.850 99.670 ;
        RECT 107.200 99.610 107.520 99.870 ;
        RECT 108.095 99.810 108.385 99.855 ;
        RECT 109.285 99.810 109.575 99.855 ;
        RECT 111.805 99.810 112.095 99.855 ;
        RECT 108.095 99.670 112.095 99.810 ;
        RECT 108.095 99.625 108.385 99.670 ;
        RECT 109.285 99.625 109.575 99.670 ;
        RECT 111.805 99.625 112.095 99.670 ;
        RECT 113.180 99.810 113.500 99.870 ;
        RECT 118.790 99.810 118.930 99.965 ;
        RECT 119.160 99.950 119.480 100.010 ;
        RECT 120.540 99.950 120.860 100.010 ;
        RECT 126.535 99.965 126.825 100.010 ;
        RECT 126.980 99.950 127.300 100.010 ;
        RECT 127.440 99.950 127.760 100.210 ;
        RECT 127.900 99.950 128.220 100.210 ;
        RECT 128.360 99.950 128.680 100.210 ;
        RECT 128.910 100.150 129.050 100.350 ;
        RECT 129.755 100.350 131.730 100.490 ;
        RECT 129.755 100.305 130.045 100.350 ;
        RECT 131.440 100.305 131.730 100.350 ;
        RECT 138.955 100.490 139.245 100.535 ;
        RECT 139.860 100.490 140.180 100.550 ;
        RECT 138.955 100.350 140.180 100.490 ;
        RECT 138.955 100.305 139.245 100.350 ;
        RECT 139.860 100.290 140.180 100.350 ;
        RECT 130.660 100.150 130.980 100.210 ;
        RECT 128.910 100.010 130.980 100.150 ;
        RECT 130.660 99.950 130.980 100.010 ;
        RECT 135.260 100.150 135.580 100.210 ;
        RECT 138.495 100.150 138.785 100.195 ;
        RECT 135.260 100.010 138.785 100.150 ;
        RECT 135.260 99.950 135.580 100.010 ;
        RECT 138.495 99.965 138.785 100.010 ;
        RECT 139.415 99.965 139.705 100.195 ;
        RECT 140.335 99.965 140.625 100.195 ;
        RECT 124.680 99.810 125.000 99.870 ;
        RECT 113.180 99.670 125.000 99.810 ;
        RECT 113.180 99.610 113.500 99.670 ;
        RECT 124.680 99.610 125.000 99.670 ;
        RECT 125.140 99.810 125.460 99.870 ;
        RECT 130.215 99.810 130.505 99.855 ;
        RECT 125.140 99.670 130.505 99.810 ;
        RECT 125.140 99.610 125.460 99.670 ;
        RECT 130.215 99.625 130.505 99.670 ;
        RECT 131.095 99.810 131.385 99.855 ;
        RECT 132.285 99.810 132.575 99.855 ;
        RECT 134.805 99.810 135.095 99.855 ;
        RECT 131.095 99.670 135.095 99.810 ;
        RECT 131.095 99.625 131.385 99.670 ;
        RECT 132.285 99.625 132.575 99.670 ;
        RECT 134.805 99.625 135.095 99.670 ;
        RECT 135.720 99.810 136.040 99.870 ;
        RECT 139.490 99.810 139.630 99.965 ;
        RECT 135.720 99.670 139.630 99.810 ;
        RECT 135.720 99.610 136.040 99.670 ;
        RECT 84.200 99.330 91.790 99.470 ;
        RECT 84.200 99.270 84.520 99.330 ;
        RECT 91.650 99.190 91.790 99.330 ;
        RECT 92.940 99.330 96.850 99.470 ;
        RECT 107.700 99.470 107.990 99.515 ;
        RECT 109.800 99.470 110.090 99.515 ;
        RECT 111.370 99.470 111.660 99.515 ;
        RECT 107.700 99.330 111.660 99.470 ;
        RECT 92.940 99.270 93.260 99.330 ;
        RECT 107.700 99.285 107.990 99.330 ;
        RECT 109.800 99.285 110.090 99.330 ;
        RECT 111.370 99.285 111.660 99.330 ;
        RECT 114.560 99.470 114.880 99.530 ;
        RECT 120.540 99.470 120.860 99.530 ;
        RECT 114.560 99.330 120.860 99.470 ;
        RECT 114.560 99.270 114.880 99.330 ;
        RECT 120.540 99.270 120.860 99.330 ;
        RECT 130.700 99.470 130.990 99.515 ;
        RECT 132.800 99.470 133.090 99.515 ;
        RECT 134.370 99.470 134.660 99.515 ;
        RECT 130.700 99.330 134.660 99.470 ;
        RECT 130.700 99.285 130.990 99.330 ;
        RECT 132.800 99.285 133.090 99.330 ;
        RECT 134.370 99.285 134.660 99.330 ;
        RECT 136.640 99.470 136.960 99.530 ;
        RECT 138.480 99.470 138.800 99.530 ;
        RECT 140.410 99.470 140.550 99.965 ;
        RECT 136.640 99.330 138.250 99.470 ;
        RECT 136.640 99.270 136.960 99.330 ;
        RECT 60.295 98.945 60.585 99.175 ;
        RECT 65.355 99.130 65.645 99.175 ;
        RECT 65.800 99.130 66.120 99.190 ;
        RECT 65.355 98.990 66.120 99.130 ;
        RECT 65.355 98.945 65.645 98.990 ;
        RECT 65.800 98.930 66.120 98.990 ;
        RECT 81.440 99.130 81.760 99.190 ;
        RECT 83.280 99.130 83.600 99.190 ;
        RECT 85.135 99.130 85.425 99.175 ;
        RECT 81.440 98.990 85.425 99.130 ;
        RECT 81.440 98.930 81.760 98.990 ;
        RECT 83.280 98.930 83.600 98.990 ;
        RECT 85.135 98.945 85.425 98.990 ;
        RECT 91.560 99.130 91.880 99.190 ;
        RECT 98.920 99.130 99.240 99.190 ;
        RECT 91.560 98.990 99.240 99.130 ;
        RECT 91.560 98.930 91.880 98.990 ;
        RECT 98.920 98.930 99.240 98.990 ;
        RECT 110.880 99.130 111.200 99.190 ;
        RECT 114.115 99.130 114.405 99.175 ;
        RECT 116.400 99.130 116.720 99.190 ;
        RECT 110.880 98.990 116.720 99.130 ;
        RECT 110.880 98.930 111.200 98.990 ;
        RECT 114.115 98.945 114.405 98.990 ;
        RECT 116.400 98.930 116.720 98.990 ;
        RECT 119.620 98.930 119.940 99.190 ;
        RECT 132.040 99.130 132.360 99.190 ;
        RECT 137.190 99.175 137.330 99.330 ;
        RECT 137.115 99.130 137.405 99.175 ;
        RECT 132.040 98.990 137.405 99.130 ;
        RECT 132.040 98.930 132.360 98.990 ;
        RECT 137.115 98.945 137.405 98.990 ;
        RECT 137.560 98.930 137.880 99.190 ;
        RECT 138.110 99.130 138.250 99.330 ;
        RECT 138.480 99.330 140.550 99.470 ;
        RECT 138.480 99.270 138.800 99.330 ;
        RECT 139.860 99.130 140.180 99.190 ;
        RECT 138.110 98.990 140.180 99.130 ;
        RECT 139.860 98.930 140.180 98.990 ;
        RECT 17.430 98.310 143.010 98.790 ;
        RECT 24.400 98.110 24.720 98.170 ;
        RECT 34.060 98.110 34.380 98.170 ;
        RECT 24.400 97.970 34.380 98.110 ;
        RECT 24.400 97.910 24.720 97.970 ;
        RECT 34.060 97.910 34.380 97.970 ;
        RECT 35.915 98.110 36.205 98.155 ;
        RECT 38.200 98.110 38.520 98.170 ;
        RECT 35.915 97.970 38.520 98.110 ;
        RECT 35.915 97.925 36.205 97.970 ;
        RECT 38.200 97.910 38.520 97.970 ;
        RECT 39.580 98.110 39.900 98.170 ;
        RECT 39.580 97.970 45.790 98.110 ;
        RECT 39.580 97.910 39.900 97.970 ;
        RECT 38.700 97.770 38.990 97.815 ;
        RECT 40.800 97.770 41.090 97.815 ;
        RECT 42.370 97.770 42.660 97.815 ;
        RECT 38.700 97.630 42.660 97.770 ;
        RECT 38.700 97.585 38.990 97.630 ;
        RECT 40.800 97.585 41.090 97.630 ;
        RECT 42.370 97.585 42.660 97.630 ;
        RECT 44.640 97.770 44.960 97.830 ;
        RECT 45.115 97.770 45.405 97.815 ;
        RECT 44.640 97.630 45.405 97.770 ;
        RECT 44.640 97.570 44.960 97.630 ;
        RECT 45.115 97.585 45.405 97.630 ;
        RECT 39.095 97.430 39.385 97.475 ;
        RECT 40.285 97.430 40.575 97.475 ;
        RECT 42.805 97.430 43.095 97.475 ;
        RECT 39.095 97.290 43.095 97.430 ;
        RECT 39.095 97.245 39.385 97.290 ;
        RECT 40.285 97.245 40.575 97.290 ;
        RECT 42.805 97.245 43.095 97.290 ;
        RECT 25.320 97.090 25.640 97.150 ;
        RECT 27.175 97.090 27.465 97.135 ;
        RECT 27.620 97.090 27.940 97.150 ;
        RECT 25.320 96.950 27.940 97.090 ;
        RECT 25.320 96.890 25.640 96.950 ;
        RECT 27.175 96.905 27.465 96.950 ;
        RECT 27.620 96.890 27.940 96.950 ;
        RECT 38.200 96.890 38.520 97.150 ;
        RECT 42.340 97.090 42.660 97.150 ;
        RECT 39.210 96.950 42.660 97.090 ;
        RECT 45.650 97.090 45.790 97.970 ;
        RECT 54.760 97.910 55.080 98.170 ;
        RECT 56.600 97.910 56.920 98.170 ;
        RECT 82.360 97.910 82.680 98.170 ;
        RECT 86.515 98.110 86.805 98.155 ;
        RECT 88.340 98.110 88.660 98.170 ;
        RECT 86.515 97.970 88.660 98.110 ;
        RECT 86.515 97.925 86.805 97.970 ;
        RECT 88.340 97.910 88.660 97.970 ;
        RECT 91.100 98.110 91.420 98.170 ;
        RECT 103.520 98.110 103.840 98.170 ;
        RECT 91.100 97.970 103.840 98.110 ;
        RECT 91.100 97.910 91.420 97.970 ;
        RECT 103.520 97.910 103.840 97.970 ;
        RECT 120.540 98.110 120.860 98.170 ;
        RECT 122.380 98.110 122.700 98.170 ;
        RECT 120.540 97.970 122.700 98.110 ;
        RECT 120.540 97.910 120.860 97.970 ;
        RECT 122.380 97.910 122.700 97.970 ;
        RECT 127.440 98.110 127.760 98.170 ;
        RECT 131.135 98.110 131.425 98.155 ;
        RECT 127.440 97.970 131.425 98.110 ;
        RECT 127.440 97.910 127.760 97.970 ;
        RECT 131.135 97.925 131.425 97.970 ;
        RECT 131.580 98.110 131.900 98.170 ;
        RECT 138.480 98.110 138.800 98.170 ;
        RECT 131.580 97.970 138.800 98.110 ;
        RECT 131.580 97.910 131.900 97.970 ;
        RECT 138.480 97.910 138.800 97.970 ;
        RECT 140.780 97.910 141.100 98.170 ;
        RECT 48.320 97.770 48.610 97.815 ;
        RECT 49.890 97.770 50.180 97.815 ;
        RECT 51.990 97.770 52.280 97.815 ;
        RECT 48.320 97.630 52.280 97.770 ;
        RECT 48.320 97.585 48.610 97.630 ;
        RECT 49.890 97.585 50.180 97.630 ;
        RECT 51.990 97.585 52.280 97.630 ;
        RECT 52.935 97.770 53.225 97.815 ;
        RECT 53.380 97.770 53.700 97.830 ;
        RECT 52.935 97.630 53.700 97.770 ;
        RECT 52.935 97.585 53.225 97.630 ;
        RECT 53.380 97.570 53.700 97.630 ;
        RECT 59.360 97.770 59.650 97.815 ;
        RECT 60.930 97.770 61.220 97.815 ;
        RECT 63.030 97.770 63.320 97.815 ;
        RECT 59.360 97.630 63.320 97.770 ;
        RECT 59.360 97.585 59.650 97.630 ;
        RECT 60.930 97.585 61.220 97.630 ;
        RECT 63.030 97.585 63.320 97.630 ;
        RECT 64.920 97.770 65.210 97.815 ;
        RECT 67.020 97.770 67.310 97.815 ;
        RECT 68.590 97.770 68.880 97.815 ;
        RECT 64.920 97.630 68.880 97.770 ;
        RECT 64.920 97.585 65.210 97.630 ;
        RECT 67.020 97.585 67.310 97.630 ;
        RECT 68.590 97.585 68.880 97.630 ;
        RECT 80.980 97.570 81.300 97.830 ;
        RECT 82.820 97.770 83.140 97.830 ;
        RECT 85.580 97.770 85.900 97.830 ;
        RECT 82.820 97.630 85.900 97.770 ;
        RECT 82.820 97.570 83.140 97.630 ;
        RECT 85.580 97.570 85.900 97.630 ;
        RECT 90.220 97.770 90.510 97.815 ;
        RECT 92.320 97.770 92.610 97.815 ;
        RECT 93.890 97.770 94.180 97.815 ;
        RECT 90.220 97.630 94.180 97.770 ;
        RECT 90.220 97.585 90.510 97.630 ;
        RECT 92.320 97.585 92.610 97.630 ;
        RECT 93.890 97.585 94.180 97.630 ;
        RECT 96.620 97.770 96.940 97.830 ;
        RECT 98.000 97.770 98.320 97.830 ;
        RECT 96.620 97.630 98.320 97.770 ;
        RECT 96.620 97.570 96.940 97.630 ;
        RECT 98.000 97.570 98.320 97.630 ;
        RECT 100.300 97.570 100.620 97.830 ;
        RECT 108.580 97.770 108.900 97.830 ;
        RECT 114.560 97.770 114.880 97.830 ;
        RECT 108.580 97.630 114.880 97.770 ;
        RECT 108.580 97.570 108.900 97.630 ;
        RECT 114.560 97.570 114.880 97.630 ;
        RECT 115.980 97.770 116.270 97.815 ;
        RECT 118.080 97.770 118.370 97.815 ;
        RECT 119.650 97.770 119.940 97.815 ;
        RECT 115.980 97.630 119.940 97.770 ;
        RECT 115.980 97.585 116.270 97.630 ;
        RECT 118.080 97.585 118.370 97.630 ;
        RECT 119.650 97.585 119.940 97.630 ;
        RECT 130.660 97.770 130.980 97.830 ;
        RECT 138.955 97.770 139.245 97.815 ;
        RECT 130.660 97.630 139.245 97.770 ;
        RECT 130.660 97.570 130.980 97.630 ;
        RECT 138.955 97.585 139.245 97.630 ;
        RECT 47.885 97.430 48.175 97.475 ;
        RECT 50.405 97.430 50.695 97.475 ;
        RECT 51.595 97.430 51.885 97.475 ;
        RECT 47.885 97.290 51.885 97.430 ;
        RECT 47.885 97.245 48.175 97.290 ;
        RECT 50.405 97.245 50.695 97.290 ;
        RECT 51.595 97.245 51.885 97.290 ;
        RECT 52.475 97.430 52.765 97.475 ;
        RECT 55.680 97.430 56.000 97.490 ;
        RECT 52.475 97.290 56.000 97.430 ;
        RECT 52.475 97.245 52.765 97.290 ;
        RECT 55.680 97.230 56.000 97.290 ;
        RECT 58.925 97.430 59.215 97.475 ;
        RECT 61.445 97.430 61.735 97.475 ;
        RECT 62.635 97.430 62.925 97.475 ;
        RECT 58.925 97.290 62.925 97.430 ;
        RECT 58.925 97.245 59.215 97.290 ;
        RECT 61.445 97.245 61.735 97.290 ;
        RECT 62.635 97.245 62.925 97.290 ;
        RECT 65.315 97.430 65.605 97.475 ;
        RECT 66.505 97.430 66.795 97.475 ;
        RECT 69.025 97.430 69.315 97.475 ;
        RECT 65.315 97.290 69.315 97.430 ;
        RECT 65.315 97.245 65.605 97.290 ;
        RECT 66.505 97.245 66.795 97.290 ;
        RECT 69.025 97.245 69.315 97.290 ;
        RECT 51.140 97.090 51.430 97.135 ;
        RECT 45.650 96.950 51.430 97.090 ;
        RECT 55.770 97.090 55.910 97.230 ;
        RECT 63.515 97.090 63.805 97.135 ;
        RECT 64.420 97.090 64.740 97.150 ;
        RECT 65.800 97.135 66.120 97.150 ;
        RECT 65.770 97.090 66.120 97.135 ;
        RECT 55.770 96.950 64.740 97.090 ;
        RECT 65.605 96.950 66.120 97.090 ;
        RECT 81.070 97.090 81.210 97.570 ;
        RECT 81.900 97.430 82.220 97.490 ;
        RECT 81.900 97.290 88.570 97.430 ;
        RECT 81.900 97.230 82.220 97.290 ;
        RECT 83.830 97.135 83.970 97.290 ;
        RECT 81.455 97.090 81.745 97.135 ;
        RECT 81.070 96.950 81.745 97.090 ;
        RECT 24.860 96.750 25.180 96.810 ;
        RECT 26.255 96.750 26.545 96.795 ;
        RECT 24.860 96.610 26.545 96.750 ;
        RECT 24.860 96.550 25.180 96.610 ;
        RECT 26.255 96.565 26.545 96.610 ;
        RECT 36.835 96.565 37.125 96.795 ;
        RECT 37.755 96.750 38.045 96.795 ;
        RECT 39.210 96.750 39.350 96.950 ;
        RECT 42.340 96.890 42.660 96.950 ;
        RECT 51.140 96.905 51.430 96.950 ;
        RECT 63.515 96.905 63.805 96.950 ;
        RECT 64.420 96.890 64.740 96.950 ;
        RECT 65.770 96.905 66.120 96.950 ;
        RECT 81.455 96.905 81.745 96.950 ;
        RECT 83.755 96.905 84.045 97.135 ;
        RECT 65.800 96.890 66.120 96.905 ;
        RECT 84.200 96.890 84.520 97.150 ;
        RECT 84.660 96.890 84.980 97.150 ;
        RECT 85.580 96.890 85.900 97.150 ;
        RECT 87.420 96.890 87.740 97.150 ;
        RECT 87.895 96.905 88.185 97.135 ;
        RECT 39.580 96.795 39.900 96.810 ;
        RECT 37.755 96.610 39.350 96.750 ;
        RECT 37.755 96.565 38.045 96.610 ;
        RECT 39.550 96.565 39.900 96.795 ;
        RECT 28.080 96.210 28.400 96.470 ;
        RECT 36.910 96.410 37.050 96.565 ;
        RECT 39.580 96.550 39.900 96.565 ;
        RECT 50.620 96.750 50.940 96.810 ;
        RECT 54.775 96.750 55.065 96.795 ;
        RECT 58.440 96.750 58.760 96.810 ;
        RECT 50.620 96.610 58.760 96.750 ;
        RECT 50.620 96.550 50.940 96.610 ;
        RECT 54.775 96.565 55.065 96.610 ;
        RECT 58.440 96.550 58.760 96.610 ;
        RECT 59.360 96.750 59.680 96.810 ;
        RECT 62.180 96.750 62.470 96.795 ;
        RECT 59.360 96.610 62.470 96.750 ;
        RECT 59.360 96.550 59.680 96.610 ;
        RECT 62.180 96.565 62.470 96.610 ;
        RECT 80.535 96.750 80.825 96.795 ;
        RECT 80.980 96.750 81.300 96.810 ;
        RECT 80.535 96.610 81.300 96.750 ;
        RECT 80.535 96.565 80.825 96.610 ;
        RECT 80.980 96.550 81.300 96.610 ;
        RECT 82.360 96.750 82.680 96.810 ;
        RECT 87.970 96.750 88.110 96.905 ;
        RECT 82.360 96.610 88.110 96.750 ;
        RECT 82.360 96.550 82.680 96.610 ;
        RECT 44.180 96.410 44.500 96.470 ;
        RECT 45.100 96.410 45.420 96.470 ;
        RECT 45.575 96.410 45.865 96.455 ;
        RECT 36.910 96.270 45.865 96.410 ;
        RECT 44.180 96.210 44.500 96.270 ;
        RECT 45.100 96.210 45.420 96.270 ;
        RECT 45.575 96.225 45.865 96.270 ;
        RECT 55.220 96.410 55.540 96.470 ;
        RECT 55.695 96.410 55.985 96.455 ;
        RECT 55.220 96.270 55.985 96.410 ;
        RECT 55.220 96.210 55.540 96.270 ;
        RECT 55.695 96.225 55.985 96.270 ;
        RECT 71.335 96.410 71.625 96.455 ;
        RECT 71.780 96.410 72.100 96.470 ;
        RECT 71.335 96.270 72.100 96.410 ;
        RECT 71.335 96.225 71.625 96.270 ;
        RECT 71.780 96.210 72.100 96.270 ;
        RECT 79.615 96.410 79.905 96.455 ;
        RECT 84.660 96.410 84.980 96.470 ;
        RECT 79.615 96.270 84.980 96.410 ;
        RECT 88.430 96.410 88.570 97.290 ;
        RECT 89.720 97.230 90.040 97.490 ;
        RECT 90.615 97.430 90.905 97.475 ;
        RECT 91.805 97.430 92.095 97.475 ;
        RECT 94.325 97.430 94.615 97.475 ;
        RECT 90.615 97.290 94.615 97.430 ;
        RECT 90.615 97.245 90.905 97.290 ;
        RECT 91.805 97.245 92.095 97.290 ;
        RECT 94.325 97.245 94.615 97.290 ;
        RECT 95.700 97.430 96.020 97.490 ;
        RECT 100.760 97.430 101.080 97.490 ;
        RECT 107.200 97.430 107.520 97.490 ;
        RECT 116.375 97.430 116.665 97.475 ;
        RECT 117.565 97.430 117.855 97.475 ;
        RECT 120.085 97.430 120.375 97.475 ;
        RECT 95.700 97.290 103.290 97.430 ;
        RECT 95.700 97.230 96.020 97.290 ;
        RECT 88.800 96.890 89.120 97.150 ;
        RECT 89.275 97.090 89.565 97.135 ;
        RECT 90.180 97.090 90.500 97.150 ;
        RECT 100.390 97.135 100.530 97.290 ;
        RECT 100.760 97.230 101.080 97.290 ;
        RECT 103.150 97.150 103.290 97.290 ;
        RECT 107.200 97.290 115.710 97.430 ;
        RECT 107.200 97.230 107.520 97.290 ;
        RECT 89.275 96.950 90.500 97.090 ;
        RECT 89.275 96.905 89.565 96.950 ;
        RECT 90.180 96.890 90.500 96.950 ;
        RECT 100.315 96.905 100.605 97.135 ;
        RECT 101.235 97.090 101.525 97.135 ;
        RECT 101.235 96.950 102.830 97.090 ;
        RECT 101.235 96.905 101.525 96.950 ;
        RECT 91.100 96.795 91.420 96.810 ;
        RECT 91.070 96.565 91.420 96.795 ;
        RECT 91.100 96.550 91.420 96.565 ;
        RECT 98.000 96.550 98.320 96.810 ;
        RECT 98.920 96.750 99.240 96.810 ;
        RECT 102.155 96.750 102.445 96.795 ;
        RECT 98.920 96.610 102.445 96.750 ;
        RECT 102.690 96.750 102.830 96.950 ;
        RECT 103.060 96.890 103.380 97.150 ;
        RECT 103.995 96.905 104.285 97.135 ;
        RECT 104.070 96.750 104.210 96.905 ;
        RECT 113.180 96.890 113.500 97.150 ;
        RECT 115.570 97.135 115.710 97.290 ;
        RECT 116.375 97.290 120.375 97.430 ;
        RECT 116.375 97.245 116.665 97.290 ;
        RECT 117.565 97.245 117.855 97.290 ;
        RECT 120.085 97.245 120.375 97.290 ;
        RECT 133.970 97.290 137.330 97.430 ;
        RECT 114.575 96.905 114.865 97.135 ;
        RECT 115.495 97.090 115.785 97.135 ;
        RECT 122.840 97.090 123.160 97.150 ;
        RECT 125.140 97.090 125.460 97.150 ;
        RECT 130.675 97.090 130.965 97.135 ;
        RECT 115.495 96.950 125.460 97.090 ;
        RECT 115.495 96.905 115.785 96.950 ;
        RECT 114.650 96.750 114.790 96.905 ;
        RECT 122.840 96.890 123.160 96.950 ;
        RECT 125.140 96.890 125.460 96.950 ;
        RECT 129.370 96.950 132.730 97.090 ;
        RECT 102.690 96.610 114.790 96.750 ;
        RECT 98.920 96.550 99.240 96.610 ;
        RECT 102.155 96.565 102.445 96.610 ;
        RECT 92.480 96.410 92.800 96.470 ;
        RECT 88.430 96.270 92.800 96.410 ;
        RECT 79.615 96.225 79.905 96.270 ;
        RECT 84.660 96.210 84.980 96.270 ;
        RECT 92.480 96.210 92.800 96.270 ;
        RECT 97.080 96.210 97.400 96.470 ;
        RECT 114.650 96.410 114.790 96.610 ;
        RECT 115.035 96.750 115.325 96.795 ;
        RECT 115.940 96.750 116.260 96.810 ;
        RECT 115.035 96.610 116.260 96.750 ;
        RECT 115.035 96.565 115.325 96.610 ;
        RECT 115.940 96.550 116.260 96.610 ;
        RECT 116.830 96.750 117.120 96.795 ;
        RECT 118.700 96.750 119.020 96.810 ;
        RECT 116.830 96.610 119.020 96.750 ;
        RECT 116.830 96.565 117.120 96.610 ;
        RECT 118.700 96.550 119.020 96.610 ;
        RECT 119.620 96.750 119.940 96.810 ;
        RECT 129.370 96.750 129.510 96.950 ;
        RECT 130.675 96.905 130.965 96.950 ;
        RECT 119.620 96.610 129.510 96.750 ;
        RECT 129.755 96.750 130.045 96.795 ;
        RECT 131.580 96.750 131.900 96.810 ;
        RECT 129.755 96.610 131.900 96.750 ;
        RECT 119.620 96.550 119.940 96.610 ;
        RECT 129.755 96.565 130.045 96.610 ;
        RECT 131.580 96.550 131.900 96.610 ;
        RECT 132.040 96.550 132.360 96.810 ;
        RECT 132.590 96.750 132.730 96.950 ;
        RECT 132.975 96.750 133.265 96.795 ;
        RECT 133.970 96.750 134.110 97.290 ;
        RECT 134.800 96.890 135.120 97.150 ;
        RECT 135.275 97.090 135.565 97.135 ;
        RECT 136.180 97.090 136.500 97.150 ;
        RECT 137.190 97.135 137.330 97.290 ;
        RECT 135.275 96.950 136.500 97.090 ;
        RECT 135.275 96.905 135.565 96.950 ;
        RECT 136.180 96.890 136.500 96.950 ;
        RECT 136.655 96.905 136.945 97.135 ;
        RECT 137.115 96.905 137.405 97.135 ;
        RECT 132.590 96.610 134.110 96.750 ;
        RECT 132.975 96.565 133.265 96.610 ;
        RECT 135.720 96.550 136.040 96.810 ;
        RECT 136.730 96.750 136.870 96.905 ;
        RECT 139.860 96.890 140.180 97.150 ;
        RECT 138.035 96.750 138.325 96.795 ;
        RECT 139.400 96.750 139.720 96.810 ;
        RECT 136.730 96.610 139.720 96.750 ;
        RECT 138.035 96.565 138.325 96.610 ;
        RECT 139.400 96.550 139.720 96.610 ;
        RECT 118.240 96.410 118.560 96.470 ;
        RECT 114.650 96.270 118.560 96.410 ;
        RECT 118.240 96.210 118.560 96.270 ;
        RECT 122.380 96.410 122.700 96.470 ;
        RECT 128.360 96.410 128.680 96.470 ;
        RECT 122.380 96.270 128.680 96.410 ;
        RECT 122.380 96.210 122.700 96.270 ;
        RECT 128.360 96.210 128.680 96.270 ;
        RECT 128.835 96.410 129.125 96.455 ;
        RECT 129.280 96.410 129.600 96.470 ;
        RECT 128.835 96.270 129.600 96.410 ;
        RECT 128.835 96.225 129.125 96.270 ;
        RECT 129.280 96.210 129.600 96.270 ;
        RECT 130.200 96.410 130.520 96.470 ;
        RECT 133.895 96.410 134.185 96.455 ;
        RECT 130.200 96.270 134.185 96.410 ;
        RECT 130.200 96.210 130.520 96.270 ;
        RECT 133.895 96.225 134.185 96.270 ;
        RECT 17.430 95.590 143.010 96.070 ;
        RECT 21.640 95.190 21.960 95.450 ;
        RECT 28.080 95.390 28.400 95.450 ;
        RECT 33.945 95.390 34.235 95.435 ;
        RECT 28.080 95.250 34.235 95.390 ;
        RECT 28.080 95.190 28.400 95.250 ;
        RECT 33.945 95.205 34.235 95.250 ;
        RECT 39.580 95.190 39.900 95.450 ;
        RECT 40.515 95.390 40.805 95.435 ;
        RECT 40.960 95.390 41.280 95.450 ;
        RECT 40.515 95.250 41.280 95.390 ;
        RECT 40.515 95.205 40.805 95.250 ;
        RECT 40.960 95.190 41.280 95.250 ;
        RECT 42.340 95.390 42.660 95.450 ;
        RECT 44.735 95.390 45.025 95.435 ;
        RECT 42.340 95.250 45.025 95.390 ;
        RECT 42.340 95.190 42.660 95.250 ;
        RECT 44.735 95.205 45.025 95.250 ;
        RECT 45.575 95.205 45.865 95.435 ;
        RECT 51.095 95.390 51.385 95.435 ;
        RECT 54.760 95.390 55.080 95.450 ;
        RECT 84.200 95.390 84.520 95.450 ;
        RECT 51.095 95.250 55.080 95.390 ;
        RECT 51.095 95.205 51.385 95.250 ;
        RECT 21.730 95.050 21.870 95.190 ;
        RECT 21.730 94.910 32.910 95.050 ;
        RECT 21.655 94.525 21.945 94.755 ;
        RECT 22.575 94.710 22.865 94.755 ;
        RECT 25.320 94.710 25.640 94.770 ;
        RECT 32.770 94.755 32.910 94.910 ;
        RECT 34.980 94.850 35.300 95.110 ;
        RECT 43.735 95.050 44.025 95.095 ;
        RECT 44.180 95.050 44.500 95.110 ;
        RECT 43.735 94.910 44.500 95.050 ;
        RECT 43.735 94.865 44.025 94.910 ;
        RECT 44.180 94.850 44.500 94.910 ;
        RECT 45.650 95.050 45.790 95.205 ;
        RECT 54.760 95.190 55.080 95.250 ;
        RECT 80.150 95.250 84.520 95.390 ;
        RECT 49.240 95.050 49.560 95.110 ;
        RECT 45.650 94.910 49.560 95.050 ;
        RECT 22.575 94.570 25.640 94.710 ;
        RECT 22.575 94.525 22.865 94.570 ;
        RECT 21.730 94.370 21.870 94.525 ;
        RECT 25.320 94.510 25.640 94.570 ;
        RECT 31.415 94.710 31.705 94.755 ;
        RECT 32.695 94.710 32.985 94.755 ;
        RECT 38.200 94.710 38.520 94.770 ;
        RECT 31.415 94.570 32.450 94.710 ;
        RECT 31.415 94.525 31.705 94.570 ;
        RECT 28.105 94.370 28.395 94.415 ;
        RECT 30.625 94.370 30.915 94.415 ;
        RECT 31.815 94.370 32.105 94.415 ;
        RECT 21.730 94.230 25.090 94.370 ;
        RECT 24.950 94.090 25.090 94.230 ;
        RECT 28.105 94.230 32.105 94.370 ;
        RECT 32.310 94.370 32.450 94.570 ;
        RECT 32.695 94.570 38.520 94.710 ;
        RECT 32.695 94.525 32.985 94.570 ;
        RECT 38.200 94.510 38.520 94.570 ;
        RECT 42.355 94.710 42.645 94.755 ;
        RECT 45.650 94.710 45.790 94.910 ;
        RECT 49.240 94.850 49.560 94.910 ;
        RECT 50.175 95.050 50.465 95.095 ;
        RECT 51.540 95.050 51.860 95.110 ;
        RECT 50.175 94.910 51.860 95.050 ;
        RECT 50.175 94.865 50.465 94.910 ;
        RECT 51.540 94.850 51.860 94.910 ;
        RECT 55.680 95.050 56.000 95.110 ;
        RECT 55.680 94.910 58.670 95.050 ;
        RECT 55.680 94.850 56.000 94.910 ;
        RECT 42.355 94.570 45.790 94.710 ;
        RECT 55.220 94.710 55.540 94.770 ;
        RECT 58.530 94.755 58.670 94.910 ;
        RECT 57.120 94.710 57.410 94.755 ;
        RECT 55.220 94.570 57.410 94.710 ;
        RECT 42.355 94.525 42.645 94.570 ;
        RECT 55.220 94.510 55.540 94.570 ;
        RECT 57.120 94.525 57.410 94.570 ;
        RECT 58.455 94.525 58.745 94.755 ;
        RECT 77.760 94.710 78.080 94.770 ;
        RECT 80.150 94.755 80.290 95.250 ;
        RECT 84.200 95.190 84.520 95.250 ;
        RECT 90.655 95.390 90.945 95.435 ;
        RECT 91.100 95.390 91.420 95.450 ;
        RECT 90.655 95.250 91.420 95.390 ;
        RECT 90.655 95.205 90.945 95.250 ;
        RECT 91.100 95.190 91.420 95.250 ;
        RECT 109.040 95.390 109.360 95.450 ;
        RECT 109.515 95.390 109.805 95.435 ;
        RECT 116.860 95.390 117.180 95.450 ;
        RECT 118.240 95.390 118.560 95.450 ;
        RECT 122.380 95.390 122.700 95.450 ;
        RECT 109.040 95.250 114.330 95.390 ;
        RECT 109.040 95.190 109.360 95.250 ;
        RECT 109.515 95.205 109.805 95.250 ;
        RECT 81.915 95.050 82.205 95.095 ;
        RECT 80.610 94.910 82.205 95.050 ;
        RECT 80.610 94.755 80.750 94.910 ;
        RECT 81.915 94.865 82.205 94.910 ;
        RECT 83.755 95.050 84.045 95.095 ;
        RECT 85.120 95.050 85.440 95.110 ;
        RECT 83.755 94.910 85.440 95.050 ;
        RECT 83.755 94.865 84.045 94.910 ;
        RECT 85.120 94.850 85.440 94.910 ;
        RECT 86.975 95.050 87.265 95.095 ;
        RECT 97.080 95.050 97.400 95.110 ;
        RECT 86.975 94.910 90.870 95.050 ;
        RECT 86.975 94.865 87.265 94.910 ;
        RECT 90.730 94.770 90.870 94.910 ;
        RECT 93.030 94.910 97.400 95.050 ;
        RECT 79.615 94.710 79.905 94.755 ;
        RECT 77.760 94.570 79.905 94.710 ;
        RECT 77.760 94.510 78.080 94.570 ;
        RECT 79.615 94.525 79.905 94.570 ;
        RECT 80.075 94.525 80.365 94.755 ;
        RECT 80.535 94.525 80.825 94.755 ;
        RECT 81.455 94.525 81.745 94.755 ;
        RECT 82.360 94.710 82.680 94.770 ;
        RECT 82.835 94.710 83.125 94.755 ;
        RECT 82.360 94.570 83.125 94.710 ;
        RECT 53.865 94.370 54.155 94.415 ;
        RECT 56.385 94.370 56.675 94.415 ;
        RECT 57.575 94.370 57.865 94.415 ;
        RECT 32.310 94.230 33.370 94.370 ;
        RECT 28.105 94.185 28.395 94.230 ;
        RECT 30.625 94.185 30.915 94.230 ;
        RECT 31.815 94.185 32.105 94.230 ;
        RECT 22.115 94.030 22.405 94.075 ;
        RECT 23.955 94.030 24.245 94.075 ;
        RECT 24.400 94.030 24.720 94.090 ;
        RECT 22.115 93.890 23.710 94.030 ;
        RECT 22.115 93.845 22.405 93.890 ;
        RECT 23.020 93.490 23.340 93.750 ;
        RECT 23.570 93.690 23.710 93.890 ;
        RECT 23.955 93.890 24.720 94.030 ;
        RECT 23.955 93.845 24.245 93.890 ;
        RECT 24.400 93.830 24.720 93.890 ;
        RECT 24.860 94.030 25.180 94.090 ;
        RECT 33.230 94.075 33.370 94.230 ;
        RECT 53.865 94.230 57.865 94.370 ;
        RECT 79.690 94.370 79.830 94.525 ;
        RECT 79.690 94.230 80.290 94.370 ;
        RECT 53.865 94.185 54.155 94.230 ;
        RECT 56.385 94.185 56.675 94.230 ;
        RECT 57.575 94.185 57.865 94.230 ;
        RECT 25.795 94.030 26.085 94.075 ;
        RECT 24.860 93.890 26.085 94.030 ;
        RECT 24.860 93.830 25.180 93.890 ;
        RECT 25.795 93.845 26.085 93.890 ;
        RECT 28.540 94.030 28.830 94.075 ;
        RECT 30.110 94.030 30.400 94.075 ;
        RECT 32.210 94.030 32.500 94.075 ;
        RECT 28.540 93.890 32.500 94.030 ;
        RECT 28.540 93.845 28.830 93.890 ;
        RECT 30.110 93.845 30.400 93.890 ;
        RECT 32.210 93.845 32.500 93.890 ;
        RECT 33.155 93.845 33.445 94.075 ;
        RECT 34.980 94.030 35.300 94.090 ;
        RECT 33.690 93.890 35.300 94.030 ;
        RECT 33.690 93.690 33.830 93.890 ;
        RECT 34.980 93.830 35.300 93.890 ;
        RECT 51.540 93.830 51.860 94.090 ;
        RECT 54.300 94.030 54.590 94.075 ;
        RECT 55.870 94.030 56.160 94.075 ;
        RECT 57.970 94.030 58.260 94.075 ;
        RECT 54.300 93.890 58.260 94.030 ;
        RECT 54.300 93.845 54.590 93.890 ;
        RECT 55.870 93.845 56.160 93.890 ;
        RECT 57.970 93.845 58.260 93.890 ;
        RECT 23.570 93.550 33.830 93.690 ;
        RECT 34.060 93.490 34.380 93.750 ;
        RECT 40.500 93.490 40.820 93.750 ;
        RECT 44.655 93.690 44.945 93.735 ;
        RECT 45.100 93.690 45.420 93.750 ;
        RECT 44.655 93.550 45.420 93.690 ;
        RECT 44.655 93.505 44.945 93.550 ;
        RECT 45.100 93.490 45.420 93.550 ;
        RECT 78.220 93.490 78.540 93.750 ;
        RECT 80.150 93.690 80.290 94.230 ;
        RECT 81.530 94.030 81.670 94.525 ;
        RECT 82.360 94.510 82.680 94.570 ;
        RECT 82.835 94.525 83.125 94.570 ;
        RECT 87.420 94.710 87.740 94.770 ;
        RECT 87.895 94.710 88.185 94.755 ;
        RECT 87.420 94.570 88.185 94.710 ;
        RECT 87.420 94.510 87.740 94.570 ;
        RECT 87.895 94.525 88.185 94.570 ;
        RECT 88.355 94.525 88.645 94.755 ;
        RECT 85.120 94.370 85.440 94.430 ;
        RECT 88.430 94.370 88.570 94.525 ;
        RECT 89.260 94.510 89.580 94.770 ;
        RECT 89.735 94.710 90.025 94.755 ;
        RECT 89.735 94.570 90.410 94.710 ;
        RECT 89.735 94.525 90.025 94.570 ;
        RECT 85.120 94.230 88.570 94.370 ;
        RECT 85.120 94.170 85.440 94.230 ;
        RECT 82.820 94.030 83.140 94.090 ;
        RECT 81.530 93.890 83.140 94.030 ;
        RECT 82.820 93.830 83.140 93.890 ;
        RECT 88.800 93.690 89.120 93.750 ;
        RECT 80.150 93.550 89.120 93.690 ;
        RECT 90.270 93.690 90.410 94.570 ;
        RECT 90.640 94.510 90.960 94.770 ;
        RECT 92.020 94.510 92.340 94.770 ;
        RECT 93.030 94.755 93.170 94.910 ;
        RECT 97.080 94.850 97.400 94.910 ;
        RECT 103.060 95.050 103.380 95.110 ;
        RECT 113.655 95.050 113.945 95.095 ;
        RECT 103.060 94.910 113.945 95.050 ;
        RECT 103.060 94.850 103.380 94.910 ;
        RECT 113.655 94.865 113.945 94.910 ;
        RECT 92.495 94.525 92.785 94.755 ;
        RECT 92.955 94.525 93.245 94.755 ;
        RECT 91.100 94.370 91.420 94.430 ;
        RECT 92.570 94.370 92.710 94.525 ;
        RECT 93.860 94.510 94.180 94.770 ;
        RECT 102.140 94.710 102.460 94.770 ;
        RECT 103.895 94.710 104.185 94.755 ;
        RECT 102.140 94.570 104.185 94.710 ;
        RECT 102.140 94.510 102.460 94.570 ;
        RECT 103.895 94.525 104.185 94.570 ;
        RECT 112.720 94.510 113.040 94.770 ;
        RECT 113.180 94.510 113.500 94.770 ;
        RECT 91.100 94.230 92.710 94.370 ;
        RECT 91.100 94.170 91.420 94.230 ;
        RECT 102.600 94.170 102.920 94.430 ;
        RECT 103.495 94.370 103.785 94.415 ;
        RECT 104.685 94.370 104.975 94.415 ;
        RECT 107.205 94.370 107.495 94.415 ;
        RECT 103.495 94.230 107.495 94.370 ;
        RECT 103.495 94.185 103.785 94.230 ;
        RECT 104.685 94.185 104.975 94.230 ;
        RECT 107.205 94.185 107.495 94.230 ;
        RECT 103.100 94.030 103.390 94.075 ;
        RECT 105.200 94.030 105.490 94.075 ;
        RECT 106.770 94.030 107.060 94.075 ;
        RECT 113.730 94.030 113.870 94.865 ;
        RECT 114.190 94.770 114.330 95.250 ;
        RECT 116.860 95.250 118.560 95.390 ;
        RECT 116.860 95.190 117.180 95.250 ;
        RECT 118.240 95.190 118.560 95.250 ;
        RECT 118.790 95.250 122.700 95.390 ;
        RECT 115.940 95.050 116.260 95.110 ;
        RECT 118.790 95.050 118.930 95.250 ;
        RECT 122.380 95.190 122.700 95.250 ;
        RECT 132.055 95.390 132.345 95.435 ;
        RECT 138.480 95.390 138.800 95.450 ;
        RECT 139.415 95.390 139.705 95.435 ;
        RECT 132.055 95.250 133.190 95.390 ;
        RECT 132.055 95.205 132.345 95.250 ;
        RECT 122.840 95.050 123.160 95.110 ;
        RECT 128.360 95.050 128.680 95.110 ;
        RECT 133.050 95.050 133.190 95.250 ;
        RECT 138.480 95.250 139.705 95.390 ;
        RECT 138.480 95.190 138.800 95.250 ;
        RECT 139.415 95.205 139.705 95.250 ;
        RECT 133.740 95.050 134.030 95.095 ;
        RECT 115.940 94.910 118.930 95.050 ;
        RECT 115.940 94.850 116.260 94.910 ;
        RECT 114.100 94.710 114.420 94.770 ;
        RECT 114.575 94.710 114.865 94.755 ;
        RECT 114.100 94.570 114.865 94.710 ;
        RECT 114.100 94.510 114.420 94.570 ;
        RECT 114.575 94.525 114.865 94.570 ;
        RECT 118.240 94.510 118.560 94.770 ;
        RECT 118.790 94.755 118.930 94.910 ;
        RECT 121.090 94.910 132.730 95.050 ;
        RECT 133.050 94.910 134.030 95.050 ;
        RECT 118.715 94.525 119.005 94.755 ;
        RECT 119.160 94.510 119.480 94.770 ;
        RECT 120.095 94.710 120.385 94.755 ;
        RECT 120.540 94.710 120.860 94.770 ;
        RECT 121.090 94.755 121.230 94.910 ;
        RECT 122.840 94.850 123.160 94.910 ;
        RECT 128.360 94.850 128.680 94.910 ;
        RECT 120.095 94.570 120.860 94.710 ;
        RECT 120.095 94.525 120.385 94.570 ;
        RECT 120.540 94.510 120.860 94.570 ;
        RECT 121.015 94.525 121.305 94.755 ;
        RECT 122.295 94.710 122.585 94.755 ;
        RECT 121.550 94.570 122.585 94.710 ;
        RECT 116.875 94.370 117.165 94.415 ;
        RECT 121.550 94.370 121.690 94.570 ;
        RECT 122.295 94.525 122.585 94.570 ;
        RECT 126.980 94.710 127.300 94.770 ;
        RECT 128.835 94.710 129.125 94.755 ;
        RECT 126.980 94.570 129.125 94.710 ;
        RECT 126.980 94.510 127.300 94.570 ;
        RECT 128.835 94.525 129.125 94.570 ;
        RECT 129.280 94.710 129.600 94.770 ;
        RECT 129.755 94.710 130.045 94.755 ;
        RECT 129.280 94.570 130.045 94.710 ;
        RECT 129.280 94.510 129.600 94.570 ;
        RECT 129.755 94.525 130.045 94.570 ;
        RECT 130.215 94.525 130.505 94.755 ;
        RECT 130.675 94.710 130.965 94.755 ;
        RECT 131.120 94.710 131.440 94.770 ;
        RECT 132.590 94.755 132.730 94.910 ;
        RECT 133.740 94.865 134.030 94.910 ;
        RECT 130.675 94.570 131.440 94.710 ;
        RECT 130.675 94.525 130.965 94.570 ;
        RECT 116.875 94.230 121.690 94.370 ;
        RECT 121.895 94.370 122.185 94.415 ;
        RECT 123.085 94.370 123.375 94.415 ;
        RECT 125.605 94.370 125.895 94.415 ;
        RECT 121.895 94.230 125.895 94.370 ;
        RECT 116.875 94.185 117.165 94.230 ;
        RECT 121.895 94.185 122.185 94.230 ;
        RECT 123.085 94.185 123.375 94.230 ;
        RECT 125.605 94.185 125.895 94.230 ;
        RECT 127.900 94.370 128.220 94.430 ;
        RECT 130.290 94.370 130.430 94.525 ;
        RECT 131.120 94.510 131.440 94.570 ;
        RECT 132.515 94.525 132.805 94.755 ;
        RECT 139.490 94.710 139.630 95.205 ;
        RECT 140.780 95.190 141.100 95.450 ;
        RECT 139.875 94.710 140.165 94.755 ;
        RECT 139.490 94.570 140.165 94.710 ;
        RECT 139.875 94.525 140.165 94.570 ;
        RECT 133.395 94.370 133.685 94.415 ;
        RECT 134.585 94.370 134.875 94.415 ;
        RECT 137.105 94.370 137.395 94.415 ;
        RECT 127.900 94.230 131.350 94.370 ;
        RECT 127.900 94.170 128.220 94.230 ;
        RECT 131.210 94.090 131.350 94.230 ;
        RECT 133.395 94.230 137.395 94.370 ;
        RECT 133.395 94.185 133.685 94.230 ;
        RECT 134.585 94.185 134.875 94.230 ;
        RECT 137.105 94.185 137.395 94.230 ;
        RECT 114.560 94.030 114.880 94.090 ;
        RECT 103.100 93.890 107.060 94.030 ;
        RECT 103.100 93.845 103.390 93.890 ;
        RECT 105.200 93.845 105.490 93.890 ;
        RECT 106.770 93.845 107.060 93.890 ;
        RECT 111.430 93.890 112.490 94.030 ;
        RECT 113.730 93.890 114.880 94.030 ;
        RECT 111.430 93.690 111.570 93.890 ;
        RECT 90.270 93.550 111.570 93.690 ;
        RECT 88.800 93.490 89.120 93.550 ;
        RECT 111.800 93.490 112.120 93.750 ;
        RECT 112.350 93.690 112.490 93.890 ;
        RECT 114.560 93.830 114.880 93.890 ;
        RECT 121.500 94.030 121.790 94.075 ;
        RECT 123.600 94.030 123.890 94.075 ;
        RECT 125.170 94.030 125.460 94.075 ;
        RECT 130.200 94.030 130.520 94.090 ;
        RECT 121.500 93.890 125.460 94.030 ;
        RECT 121.500 93.845 121.790 93.890 ;
        RECT 123.600 93.845 123.890 93.890 ;
        RECT 125.170 93.845 125.460 93.890 ;
        RECT 127.530 93.890 130.520 94.030 ;
        RECT 127.530 93.690 127.670 93.890 ;
        RECT 130.200 93.830 130.520 93.890 ;
        RECT 131.120 93.830 131.440 94.090 ;
        RECT 133.000 94.030 133.290 94.075 ;
        RECT 135.100 94.030 135.390 94.075 ;
        RECT 136.670 94.030 136.960 94.075 ;
        RECT 133.000 93.890 136.960 94.030 ;
        RECT 133.000 93.845 133.290 93.890 ;
        RECT 135.100 93.845 135.390 93.890 ;
        RECT 136.670 93.845 136.960 93.890 ;
        RECT 112.350 93.550 127.670 93.690 ;
        RECT 127.900 93.490 128.220 93.750 ;
        RECT 17.430 92.870 143.010 93.350 ;
        RECT 25.780 92.670 26.100 92.730 ;
        RECT 29.475 92.670 29.765 92.715 ;
        RECT 25.780 92.530 29.765 92.670 ;
        RECT 25.780 92.470 26.100 92.530 ;
        RECT 29.475 92.485 29.765 92.530 ;
        RECT 53.395 92.670 53.685 92.715 ;
        RECT 53.840 92.670 54.160 92.730 ;
        RECT 53.395 92.530 54.160 92.670 ;
        RECT 53.395 92.485 53.685 92.530 ;
        RECT 53.840 92.470 54.160 92.530 ;
        RECT 80.980 92.670 81.300 92.730 ;
        RECT 85.120 92.670 85.440 92.730 ;
        RECT 80.980 92.530 85.440 92.670 ;
        RECT 80.980 92.470 81.300 92.530 ;
        RECT 85.120 92.470 85.440 92.530 ;
        RECT 85.580 92.670 85.900 92.730 ;
        RECT 87.435 92.670 87.725 92.715 ;
        RECT 85.580 92.530 87.725 92.670 ;
        RECT 85.580 92.470 85.900 92.530 ;
        RECT 87.435 92.485 87.725 92.530 ;
        RECT 89.260 92.670 89.580 92.730 ;
        RECT 91.115 92.670 91.405 92.715 ;
        RECT 89.260 92.530 91.405 92.670 ;
        RECT 89.260 92.470 89.580 92.530 ;
        RECT 91.115 92.485 91.405 92.530 ;
        RECT 102.140 92.470 102.460 92.730 ;
        RECT 106.280 92.470 106.600 92.730 ;
        RECT 116.860 92.670 117.180 92.730 ;
        RECT 106.830 92.530 117.180 92.670 ;
        RECT 23.060 92.330 23.350 92.375 ;
        RECT 25.160 92.330 25.450 92.375 ;
        RECT 26.730 92.330 27.020 92.375 ;
        RECT 23.060 92.190 27.020 92.330 ;
        RECT 23.060 92.145 23.350 92.190 ;
        RECT 25.160 92.145 25.450 92.190 ;
        RECT 26.730 92.145 27.020 92.190 ;
        RECT 75.040 92.330 75.330 92.375 ;
        RECT 77.140 92.330 77.430 92.375 ;
        RECT 78.710 92.330 79.000 92.375 ;
        RECT 103.520 92.330 103.840 92.390 ;
        RECT 106.830 92.330 106.970 92.530 ;
        RECT 116.860 92.470 117.180 92.530 ;
        RECT 119.160 92.670 119.480 92.730 ;
        RECT 120.095 92.670 120.385 92.715 ;
        RECT 119.160 92.530 120.385 92.670 ;
        RECT 119.160 92.470 119.480 92.530 ;
        RECT 120.095 92.485 120.385 92.530 ;
        RECT 120.540 92.670 120.860 92.730 ;
        RECT 121.475 92.670 121.765 92.715 ;
        RECT 120.540 92.530 121.765 92.670 ;
        RECT 120.540 92.470 120.860 92.530 ;
        RECT 121.475 92.485 121.765 92.530 ;
        RECT 139.400 92.670 139.720 92.730 ;
        RECT 140.795 92.670 141.085 92.715 ;
        RECT 139.400 92.530 141.085 92.670 ;
        RECT 139.400 92.470 139.720 92.530 ;
        RECT 140.795 92.485 141.085 92.530 ;
        RECT 121.000 92.330 121.320 92.390 ;
        RECT 75.040 92.190 79.000 92.330 ;
        RECT 75.040 92.145 75.330 92.190 ;
        RECT 77.140 92.145 77.430 92.190 ;
        RECT 78.710 92.145 79.000 92.190 ;
        RECT 103.150 92.190 106.970 92.330 ;
        RECT 108.670 92.190 121.320 92.330 ;
        RECT 21.640 91.990 21.960 92.050 ;
        RECT 22.575 91.990 22.865 92.035 ;
        RECT 21.640 91.850 22.865 91.990 ;
        RECT 21.640 91.790 21.960 91.850 ;
        RECT 22.575 91.805 22.865 91.850 ;
        RECT 23.455 91.990 23.745 92.035 ;
        RECT 24.645 91.990 24.935 92.035 ;
        RECT 27.165 91.990 27.455 92.035 ;
        RECT 54.300 91.990 54.620 92.050 ;
        RECT 23.455 91.850 27.455 91.990 ;
        RECT 23.455 91.805 23.745 91.850 ;
        RECT 24.645 91.805 24.935 91.850 ;
        RECT 27.165 91.805 27.455 91.850 ;
        RECT 53.010 91.850 54.620 91.990 ;
        RECT 23.020 91.650 23.340 91.710 ;
        RECT 53.010 91.695 53.150 91.850 ;
        RECT 54.300 91.790 54.620 91.850 ;
        RECT 75.435 91.990 75.725 92.035 ;
        RECT 76.625 91.990 76.915 92.035 ;
        RECT 79.145 91.990 79.435 92.035 ;
        RECT 95.700 91.990 96.020 92.050 ;
        RECT 75.435 91.850 79.435 91.990 ;
        RECT 75.435 91.805 75.725 91.850 ;
        RECT 76.625 91.805 76.915 91.850 ;
        RECT 79.145 91.805 79.435 91.850 ;
        RECT 92.110 91.850 96.020 91.990 ;
        RECT 92.110 91.710 92.250 91.850 ;
        RECT 95.700 91.790 96.020 91.850 ;
        RECT 23.855 91.650 24.145 91.695 ;
        RECT 23.020 91.510 24.145 91.650 ;
        RECT 23.020 91.450 23.340 91.510 ;
        RECT 23.855 91.465 24.145 91.510 ;
        RECT 52.935 91.465 53.225 91.695 ;
        RECT 53.380 91.650 53.700 91.710 ;
        RECT 53.855 91.650 54.145 91.695 ;
        RECT 53.380 91.510 54.145 91.650 ;
        RECT 53.380 91.450 53.700 91.510 ;
        RECT 53.855 91.465 54.145 91.510 ;
        RECT 74.540 91.450 74.860 91.710 ;
        RECT 75.890 91.650 76.180 91.695 ;
        RECT 78.220 91.650 78.540 91.710 ;
        RECT 75.890 91.510 78.540 91.650 ;
        RECT 75.890 91.465 76.180 91.510 ;
        RECT 78.220 91.450 78.540 91.510 ;
        RECT 83.740 91.450 84.060 91.710 ;
        RECT 84.200 91.450 84.520 91.710 ;
        RECT 84.660 91.450 84.980 91.710 ;
        RECT 85.580 91.450 85.900 91.710 ;
        RECT 86.515 91.465 86.805 91.695 ;
        RECT 86.590 91.310 86.730 91.465 ;
        RECT 92.020 91.450 92.340 91.710 ;
        RECT 93.875 91.650 94.165 91.695 ;
        RECT 101.680 91.650 102.000 91.710 ;
        RECT 93.875 91.510 102.000 91.650 ;
        RECT 103.150 91.650 103.290 92.190 ;
        RECT 103.520 92.130 103.840 92.190 ;
        RECT 103.435 91.650 103.725 91.695 ;
        RECT 103.150 91.510 103.725 91.650 ;
        RECT 93.875 91.465 94.165 91.510 ;
        RECT 101.680 91.450 102.000 91.510 ;
        RECT 103.435 91.465 103.725 91.510 ;
        RECT 103.995 91.465 104.285 91.695 ;
        RECT 104.455 91.465 104.745 91.695 ;
        RECT 105.375 91.650 105.665 91.695 ;
        RECT 106.280 91.650 106.600 91.710 ;
        RECT 105.375 91.510 106.600 91.650 ;
        RECT 105.375 91.465 105.665 91.510 ;
        RECT 76.010 91.170 86.730 91.310 ;
        RECT 76.010 91.030 76.150 91.170 ;
        RECT 75.920 90.770 76.240 91.030 ;
        RECT 81.455 90.970 81.745 91.015 ;
        RECT 81.900 90.970 82.220 91.030 ;
        RECT 81.455 90.830 82.220 90.970 ;
        RECT 81.455 90.785 81.745 90.830 ;
        RECT 81.900 90.770 82.220 90.830 ;
        RECT 82.360 90.770 82.680 91.030 ;
        RECT 86.590 90.970 86.730 91.170 ;
        RECT 92.480 91.110 92.800 91.370 ;
        RECT 92.940 91.110 93.260 91.370 ;
        RECT 100.300 91.310 100.620 91.370 ;
        RECT 104.070 91.310 104.210 91.465 ;
        RECT 100.300 91.170 104.210 91.310 ;
        RECT 104.530 91.310 104.670 91.465 ;
        RECT 106.280 91.450 106.600 91.510 ;
        RECT 106.740 91.650 107.060 91.710 ;
        RECT 107.215 91.650 107.505 91.695 ;
        RECT 108.670 91.650 108.810 92.190 ;
        RECT 121.000 92.130 121.320 92.190 ;
        RECT 134.380 92.330 134.670 92.375 ;
        RECT 136.480 92.330 136.770 92.375 ;
        RECT 138.050 92.330 138.340 92.375 ;
        RECT 134.380 92.190 138.340 92.330 ;
        RECT 134.380 92.145 134.670 92.190 ;
        RECT 136.480 92.145 136.770 92.190 ;
        RECT 138.050 92.145 138.340 92.190 ;
        RECT 127.900 91.990 128.220 92.050 ;
        RECT 119.250 91.850 128.220 91.990 ;
        RECT 106.740 91.510 108.810 91.650 ;
        RECT 106.740 91.450 107.060 91.510 ;
        RECT 107.215 91.465 107.505 91.510 ;
        RECT 109.040 91.450 109.360 91.710 ;
        RECT 113.180 91.650 113.500 91.710 ;
        RECT 119.250 91.695 119.390 91.850 ;
        RECT 127.900 91.790 128.220 91.850 ;
        RECT 128.360 91.990 128.680 92.050 ;
        RECT 133.895 91.990 134.185 92.035 ;
        RECT 128.360 91.850 134.185 91.990 ;
        RECT 128.360 91.790 128.680 91.850 ;
        RECT 133.895 91.805 134.185 91.850 ;
        RECT 134.775 91.990 135.065 92.035 ;
        RECT 135.965 91.990 136.255 92.035 ;
        RECT 138.485 91.990 138.775 92.035 ;
        RECT 134.775 91.850 138.775 91.990 ;
        RECT 134.775 91.805 135.065 91.850 ;
        RECT 135.965 91.805 136.255 91.850 ;
        RECT 138.485 91.805 138.775 91.850 ;
        RECT 119.175 91.650 119.465 91.695 ;
        RECT 113.180 91.510 119.465 91.650 ;
        RECT 113.180 91.450 113.500 91.510 ;
        RECT 119.175 91.465 119.465 91.510 ;
        RECT 120.080 91.650 120.400 91.710 ;
        RECT 120.555 91.650 120.845 91.695 ;
        RECT 120.080 91.510 120.845 91.650 ;
        RECT 120.080 91.450 120.400 91.510 ;
        RECT 120.555 91.465 120.845 91.510 ;
        RECT 126.980 91.650 127.300 91.710 ;
        RECT 129.755 91.650 130.045 91.695 ;
        RECT 126.980 91.510 130.045 91.650 ;
        RECT 126.980 91.450 127.300 91.510 ;
        RECT 108.135 91.310 108.425 91.355 ;
        RECT 104.530 91.170 108.425 91.310 ;
        RECT 100.300 91.110 100.620 91.170 ;
        RECT 97.080 90.970 97.400 91.030 ;
        RECT 86.590 90.830 97.400 90.970 ;
        RECT 104.070 90.970 104.210 91.170 ;
        RECT 108.135 91.125 108.425 91.170 ;
        RECT 109.500 91.310 109.820 91.370 ;
        RECT 109.975 91.310 110.265 91.355 ;
        RECT 109.500 91.170 110.265 91.310 ;
        RECT 109.500 91.110 109.820 91.170 ;
        RECT 109.975 91.125 110.265 91.170 ;
        RECT 118.255 91.310 118.545 91.355 ;
        RECT 119.620 91.310 119.940 91.370 ;
        RECT 118.255 91.170 119.940 91.310 ;
        RECT 118.255 91.125 118.545 91.170 ;
        RECT 119.620 91.110 119.940 91.170 ;
        RECT 109.040 90.970 109.360 91.030 ;
        RECT 104.070 90.830 109.360 90.970 ;
        RECT 97.080 90.770 97.400 90.830 ;
        RECT 109.040 90.770 109.360 90.830 ;
        RECT 120.540 90.970 120.860 91.030 ;
        RECT 127.070 90.970 127.210 91.450 ;
        RECT 128.450 91.370 128.590 91.510 ;
        RECT 129.755 91.465 130.045 91.510 ;
        RECT 130.660 91.450 130.980 91.710 ;
        RECT 131.120 91.450 131.440 91.710 ;
        RECT 131.595 91.650 131.885 91.695 ;
        RECT 132.500 91.650 132.820 91.710 ;
        RECT 131.595 91.510 132.820 91.650 ;
        RECT 133.970 91.650 134.110 91.805 ;
        RECT 133.970 91.510 136.410 91.650 ;
        RECT 131.595 91.465 131.885 91.510 ;
        RECT 132.500 91.450 132.820 91.510 ;
        RECT 128.360 91.110 128.680 91.370 ;
        RECT 120.540 90.830 127.210 90.970 ;
        RECT 127.440 90.970 127.760 91.030 ;
        RECT 131.210 90.970 131.350 91.450 ;
        RECT 136.270 91.370 136.410 91.510 ;
        RECT 132.975 91.310 133.265 91.355 ;
        RECT 135.120 91.310 135.410 91.355 ;
        RECT 132.975 91.170 135.410 91.310 ;
        RECT 132.975 91.125 133.265 91.170 ;
        RECT 135.120 91.125 135.410 91.170 ;
        RECT 136.180 91.110 136.500 91.370 ;
        RECT 135.720 90.970 136.040 91.030 ;
        RECT 127.440 90.830 136.040 90.970 ;
        RECT 120.540 90.770 120.860 90.830 ;
        RECT 127.440 90.770 127.760 90.830 ;
        RECT 135.720 90.770 136.040 90.830 ;
        RECT 17.430 90.150 143.010 90.630 ;
        RECT 85.580 89.750 85.900 90.010 ;
        RECT 98.920 89.950 99.240 90.010 ;
        RECT 95.330 89.810 99.240 89.950 ;
        RECT 85.670 89.610 85.810 89.750 ;
        RECT 95.330 89.655 95.470 89.810 ;
        RECT 98.920 89.750 99.240 89.810 ;
        RECT 109.960 89.750 110.280 90.010 ;
        RECT 112.720 89.950 113.040 90.010 ;
        RECT 119.620 89.950 119.940 90.010 ;
        RECT 112.720 89.810 115.250 89.950 ;
        RECT 112.720 89.750 113.040 89.810 ;
        RECT 85.670 89.470 94.550 89.610 ;
        RECT 76.350 89.270 76.640 89.315 ;
        RECT 82.360 89.270 82.680 89.330 ;
        RECT 76.350 89.130 82.680 89.270 ;
        RECT 76.350 89.085 76.640 89.130 ;
        RECT 82.360 89.070 82.680 89.130 ;
        RECT 83.740 89.270 84.060 89.330 ;
        RECT 87.050 89.315 87.190 89.470 ;
        RECT 85.135 89.270 85.425 89.315 ;
        RECT 83.740 89.130 85.425 89.270 ;
        RECT 83.740 89.070 84.060 89.130 ;
        RECT 85.135 89.085 85.425 89.130 ;
        RECT 85.595 89.085 85.885 89.315 ;
        RECT 86.055 89.085 86.345 89.315 ;
        RECT 86.975 89.085 87.265 89.315 ;
        RECT 74.540 88.930 74.860 88.990 ;
        RECT 75.015 88.930 75.305 88.975 ;
        RECT 74.540 88.790 75.305 88.930 ;
        RECT 74.540 88.730 74.860 88.790 ;
        RECT 75.015 88.745 75.305 88.790 ;
        RECT 75.895 88.930 76.185 88.975 ;
        RECT 77.085 88.930 77.375 88.975 ;
        RECT 79.605 88.930 79.895 88.975 ;
        RECT 75.895 88.790 79.895 88.930 ;
        RECT 75.895 88.745 76.185 88.790 ;
        RECT 77.085 88.745 77.375 88.790 ;
        RECT 79.605 88.745 79.895 88.790 ;
        RECT 75.090 88.250 75.230 88.745 ;
        RECT 75.500 88.590 75.790 88.635 ;
        RECT 77.600 88.590 77.890 88.635 ;
        RECT 79.170 88.590 79.460 88.635 ;
        RECT 75.500 88.450 79.460 88.590 ;
        RECT 85.670 88.590 85.810 89.085 ;
        RECT 86.130 88.930 86.270 89.085 ;
        RECT 88.800 89.070 89.120 89.330 ;
        RECT 89.275 89.085 89.565 89.315 ;
        RECT 88.340 88.930 88.660 88.990 ;
        RECT 86.130 88.790 88.660 88.930 ;
        RECT 88.340 88.730 88.660 88.790 ;
        RECT 89.350 88.930 89.490 89.085 ;
        RECT 89.720 89.070 90.040 89.330 ;
        RECT 90.730 89.315 90.870 89.470 ;
        RECT 90.655 89.085 90.945 89.315 ;
        RECT 91.100 89.070 91.420 89.330 ;
        RECT 92.020 89.070 92.340 89.330 ;
        RECT 92.495 89.085 92.785 89.315 ;
        RECT 91.190 88.930 91.330 89.070 ;
        RECT 89.350 88.790 91.330 88.930 ;
        RECT 91.560 88.930 91.880 88.990 ;
        RECT 92.570 88.930 92.710 89.085 ;
        RECT 92.940 89.070 93.260 89.330 ;
        RECT 93.860 89.070 94.180 89.330 ;
        RECT 91.560 88.790 92.710 88.930 ;
        RECT 94.410 88.930 94.550 89.470 ;
        RECT 95.255 89.425 95.545 89.655 ;
        RECT 95.700 89.610 96.020 89.670 ;
        RECT 97.095 89.610 97.385 89.655 ;
        RECT 95.700 89.470 97.385 89.610 ;
        RECT 95.700 89.410 96.020 89.470 ;
        RECT 97.095 89.425 97.385 89.470 ;
        RECT 106.280 89.610 106.600 89.670 ;
        RECT 110.880 89.610 111.200 89.670 ;
        RECT 106.280 89.470 113.410 89.610 ;
        RECT 106.280 89.410 106.600 89.470 ;
        RECT 110.880 89.410 111.200 89.470 ;
        RECT 96.175 89.270 96.465 89.315 ;
        RECT 96.620 89.270 96.940 89.330 ;
        RECT 96.175 89.130 96.940 89.270 ;
        RECT 96.175 89.085 96.465 89.130 ;
        RECT 96.620 89.070 96.940 89.130 ;
        RECT 97.555 89.085 97.845 89.315 ;
        RECT 97.630 88.930 97.770 89.085 ;
        RECT 98.460 89.070 98.780 89.330 ;
        RECT 98.935 89.085 99.225 89.315 ;
        RECT 94.410 88.790 97.770 88.930 ;
        RECT 99.010 88.930 99.150 89.085 ;
        RECT 99.380 89.070 99.700 89.330 ;
        RECT 102.600 89.070 102.920 89.330 ;
        RECT 103.950 89.270 104.240 89.315 ;
        RECT 108.120 89.270 108.440 89.330 ;
        RECT 111.355 89.270 111.645 89.315 ;
        RECT 103.950 89.130 108.440 89.270 ;
        RECT 103.950 89.085 104.240 89.130 ;
        RECT 108.120 89.070 108.440 89.130 ;
        RECT 108.670 89.130 111.645 89.270 ;
        RECT 100.300 88.930 100.620 88.990 ;
        RECT 99.010 88.790 100.620 88.930 ;
        RECT 89.350 88.590 89.490 88.790 ;
        RECT 91.560 88.730 91.880 88.790 ;
        RECT 85.670 88.450 89.490 88.590 ;
        RECT 75.500 88.405 75.790 88.450 ;
        RECT 77.600 88.405 77.890 88.450 ;
        RECT 79.170 88.405 79.460 88.450 ;
        RECT 80.520 88.250 80.840 88.310 ;
        RECT 75.090 88.110 80.840 88.250 ;
        RECT 80.520 88.050 80.840 88.110 ;
        RECT 80.980 88.250 81.300 88.310 ;
        RECT 81.915 88.250 82.205 88.295 ;
        RECT 80.980 88.110 82.205 88.250 ;
        RECT 80.980 88.050 81.300 88.110 ;
        RECT 81.915 88.065 82.205 88.110 ;
        RECT 83.740 88.050 84.060 88.310 ;
        RECT 87.420 88.050 87.740 88.310 ;
        RECT 89.350 88.250 89.490 88.450 ;
        RECT 90.180 88.590 90.500 88.650 ;
        RECT 91.115 88.590 91.405 88.635 ;
        RECT 94.780 88.590 95.100 88.650 ;
        RECT 99.010 88.590 99.150 88.790 ;
        RECT 100.300 88.730 100.620 88.790 ;
        RECT 103.495 88.930 103.785 88.975 ;
        RECT 104.685 88.930 104.975 88.975 ;
        RECT 107.205 88.930 107.495 88.975 ;
        RECT 103.495 88.790 107.495 88.930 ;
        RECT 103.495 88.745 103.785 88.790 ;
        RECT 104.685 88.745 104.975 88.790 ;
        RECT 107.205 88.745 107.495 88.790 ;
        RECT 103.100 88.590 103.390 88.635 ;
        RECT 105.200 88.590 105.490 88.635 ;
        RECT 106.770 88.590 107.060 88.635 ;
        RECT 90.180 88.450 91.405 88.590 ;
        RECT 90.180 88.390 90.500 88.450 ;
        RECT 91.115 88.405 91.405 88.450 ;
        RECT 93.950 88.450 99.150 88.590 ;
        RECT 100.390 88.450 102.830 88.590 ;
        RECT 93.950 88.250 94.090 88.450 ;
        RECT 94.780 88.390 95.100 88.450 ;
        RECT 89.350 88.110 94.090 88.250 ;
        RECT 94.320 88.250 94.640 88.310 ;
        RECT 100.390 88.250 100.530 88.450 ;
        RECT 94.320 88.110 100.530 88.250 ;
        RECT 94.320 88.050 94.640 88.110 ;
        RECT 100.760 88.050 101.080 88.310 ;
        RECT 102.690 88.250 102.830 88.450 ;
        RECT 103.100 88.450 107.060 88.590 ;
        RECT 103.100 88.405 103.390 88.450 ;
        RECT 105.200 88.405 105.490 88.450 ;
        RECT 106.770 88.405 107.060 88.450 ;
        RECT 108.670 88.250 108.810 89.130 ;
        RECT 111.355 89.085 111.645 89.130 ;
        RECT 111.815 89.085 112.105 89.315 ;
        RECT 109.040 88.930 109.360 88.990 ;
        RECT 111.890 88.930 112.030 89.085 ;
        RECT 112.260 89.070 112.580 89.330 ;
        RECT 113.270 89.315 113.410 89.470 ;
        RECT 114.560 89.410 114.880 89.670 ;
        RECT 115.110 89.610 115.250 89.810 ;
        RECT 118.330 89.810 119.940 89.950 ;
        RECT 118.330 89.655 118.470 89.810 ;
        RECT 119.620 89.750 119.940 89.810 ;
        RECT 122.380 89.950 122.700 90.010 ;
        RECT 124.680 89.950 125.000 90.010 ;
        RECT 126.980 89.950 127.300 90.010 ;
        RECT 122.380 89.810 127.300 89.950 ;
        RECT 122.380 89.750 122.700 89.810 ;
        RECT 124.680 89.750 125.000 89.810 ;
        RECT 126.980 89.750 127.300 89.810 ;
        RECT 127.440 89.750 127.760 90.010 ;
        RECT 115.110 89.470 115.710 89.610 ;
        RECT 113.195 89.085 113.485 89.315 ;
        RECT 113.655 89.085 113.945 89.315 ;
        RECT 109.040 88.790 112.030 88.930 ;
        RECT 109.040 88.730 109.360 88.790 ;
        RECT 109.515 88.590 109.805 88.635 ;
        RECT 110.420 88.590 110.740 88.650 ;
        RECT 113.730 88.590 113.870 89.085 ;
        RECT 114.100 89.070 114.420 89.330 ;
        RECT 115.570 89.315 115.710 89.470 ;
        RECT 118.255 89.425 118.545 89.655 ;
        RECT 119.160 89.610 119.480 89.670 ;
        RECT 127.530 89.610 127.670 89.750 ;
        RECT 129.740 89.610 130.060 89.670 ;
        RECT 119.160 89.470 127.670 89.610 ;
        RECT 127.990 89.470 130.060 89.610 ;
        RECT 119.160 89.410 119.480 89.470 ;
        RECT 115.035 89.085 115.325 89.315 ;
        RECT 115.495 89.270 115.785 89.315 ;
        RECT 118.700 89.270 119.020 89.330 ;
        RECT 115.495 89.130 119.020 89.270 ;
        RECT 115.495 89.085 115.785 89.130 ;
        RECT 114.190 88.650 114.330 89.070 ;
        RECT 114.560 88.930 114.880 88.990 ;
        RECT 115.110 88.930 115.250 89.085 ;
        RECT 118.700 89.070 119.020 89.130 ;
        RECT 120.540 89.270 120.860 89.330 ;
        RECT 121.015 89.270 121.305 89.315 ;
        RECT 121.935 89.270 122.225 89.315 ;
        RECT 120.540 89.130 121.305 89.270 ;
        RECT 120.540 89.070 120.860 89.130 ;
        RECT 121.015 89.085 121.305 89.130 ;
        RECT 121.550 89.130 122.225 89.270 ;
        RECT 120.095 88.930 120.385 88.975 ;
        RECT 121.550 88.930 121.690 89.130 ;
        RECT 121.935 89.085 122.225 89.130 ;
        RECT 122.380 89.070 122.700 89.330 ;
        RECT 122.855 89.085 123.145 89.315 ;
        RECT 126.060 89.270 126.380 89.330 ;
        RECT 126.535 89.270 126.825 89.315 ;
        RECT 126.060 89.130 126.825 89.270 ;
        RECT 114.560 88.790 115.250 88.930 ;
        RECT 116.030 88.790 119.390 88.930 ;
        RECT 114.560 88.730 114.880 88.790 ;
        RECT 109.515 88.450 113.870 88.590 ;
        RECT 109.515 88.405 109.805 88.450 ;
        RECT 110.420 88.390 110.740 88.450 ;
        RECT 114.100 88.390 114.420 88.650 ;
        RECT 116.030 88.250 116.170 88.790 ;
        RECT 119.250 88.590 119.390 88.790 ;
        RECT 120.095 88.790 121.690 88.930 ;
        RECT 120.095 88.745 120.385 88.790 ;
        RECT 122.930 88.590 123.070 89.085 ;
        RECT 126.060 89.070 126.380 89.130 ;
        RECT 126.535 89.085 126.825 89.130 ;
        RECT 126.980 89.070 127.300 89.330 ;
        RECT 127.455 89.270 127.745 89.315 ;
        RECT 127.990 89.270 128.130 89.470 ;
        RECT 129.740 89.410 130.060 89.470 ;
        RECT 134.430 89.470 136.870 89.610 ;
        RECT 127.455 89.130 128.130 89.270 ;
        RECT 127.455 89.085 127.745 89.130 ;
        RECT 128.360 89.070 128.680 89.330 ;
        RECT 134.430 89.270 134.570 89.470 ;
        RECT 128.910 89.130 134.570 89.270 ;
        RECT 134.915 89.270 135.205 89.315 ;
        RECT 135.720 89.270 136.040 89.330 ;
        RECT 134.915 89.130 136.040 89.270 ;
        RECT 123.300 88.930 123.620 88.990 ;
        RECT 128.910 88.930 129.050 89.130 ;
        RECT 134.915 89.085 135.205 89.130 ;
        RECT 135.720 89.070 136.040 89.130 ;
        RECT 136.180 89.070 136.500 89.330 ;
        RECT 136.730 89.270 136.870 89.470 ;
        RECT 138.035 89.270 138.325 89.315 ;
        RECT 136.730 89.130 138.325 89.270 ;
        RECT 138.035 89.085 138.325 89.130 ;
        RECT 139.400 89.270 139.720 89.330 ;
        RECT 139.875 89.270 140.165 89.315 ;
        RECT 139.400 89.130 140.165 89.270 ;
        RECT 139.400 89.070 139.720 89.130 ;
        RECT 139.875 89.085 140.165 89.130 ;
        RECT 123.300 88.790 129.050 88.930 ;
        RECT 131.605 88.930 131.895 88.975 ;
        RECT 134.125 88.930 134.415 88.975 ;
        RECT 135.315 88.930 135.605 88.975 ;
        RECT 131.605 88.790 135.605 88.930 ;
        RECT 123.300 88.730 123.620 88.790 ;
        RECT 131.605 88.745 131.895 88.790 ;
        RECT 134.125 88.745 134.415 88.790 ;
        RECT 135.315 88.745 135.605 88.790 ;
        RECT 119.250 88.450 123.070 88.590 ;
        RECT 132.040 88.590 132.330 88.635 ;
        RECT 133.610 88.590 133.900 88.635 ;
        RECT 135.710 88.590 136.000 88.635 ;
        RECT 132.040 88.450 136.000 88.590 ;
        RECT 132.040 88.405 132.330 88.450 ;
        RECT 133.610 88.405 133.900 88.450 ;
        RECT 135.710 88.405 136.000 88.450 ;
        RECT 138.940 88.390 139.260 88.650 ;
        RECT 140.780 88.390 141.100 88.650 ;
        RECT 102.690 88.110 116.170 88.250 ;
        RECT 116.415 88.250 116.705 88.295 ;
        RECT 117.780 88.250 118.100 88.310 ;
        RECT 116.415 88.110 118.100 88.250 ;
        RECT 116.415 88.065 116.705 88.110 ;
        RECT 117.780 88.050 118.100 88.110 ;
        RECT 124.220 88.050 124.540 88.310 ;
        RECT 125.155 88.250 125.445 88.295 ;
        RECT 126.520 88.250 126.840 88.310 ;
        RECT 125.155 88.110 126.840 88.250 ;
        RECT 125.155 88.065 125.445 88.110 ;
        RECT 126.520 88.050 126.840 88.110 ;
        RECT 127.440 88.250 127.760 88.310 ;
        RECT 129.295 88.250 129.585 88.295 ;
        RECT 127.440 88.110 129.585 88.250 ;
        RECT 127.440 88.050 127.760 88.110 ;
        RECT 129.295 88.065 129.585 88.110 ;
        RECT 17.430 87.430 143.010 87.910 ;
        RECT 89.275 87.230 89.565 87.275 ;
        RECT 92.480 87.230 92.800 87.290 ;
        RECT 89.275 87.090 92.800 87.230 ;
        RECT 89.275 87.045 89.565 87.090 ;
        RECT 92.480 87.030 92.800 87.090 ;
        RECT 94.320 87.230 94.640 87.290 ;
        RECT 94.320 87.090 105.130 87.230 ;
        RECT 94.320 87.030 94.640 87.090 ;
        RECT 82.860 86.890 83.150 86.935 ;
        RECT 84.960 86.890 85.250 86.935 ;
        RECT 86.530 86.890 86.820 86.935 ;
        RECT 82.860 86.750 86.820 86.890 ;
        RECT 82.860 86.705 83.150 86.750 ;
        RECT 84.960 86.705 85.250 86.750 ;
        RECT 86.530 86.705 86.820 86.750 ;
        RECT 91.600 86.890 91.890 86.935 ;
        RECT 93.700 86.890 93.990 86.935 ;
        RECT 95.270 86.890 95.560 86.935 ;
        RECT 91.600 86.750 95.560 86.890 ;
        RECT 91.600 86.705 91.890 86.750 ;
        RECT 93.700 86.705 93.990 86.750 ;
        RECT 95.270 86.705 95.560 86.750 ;
        RECT 98.960 86.890 99.250 86.935 ;
        RECT 101.060 86.890 101.350 86.935 ;
        RECT 102.630 86.890 102.920 86.935 ;
        RECT 98.960 86.750 102.920 86.890 ;
        RECT 98.960 86.705 99.250 86.750 ;
        RECT 101.060 86.705 101.350 86.750 ;
        RECT 102.630 86.705 102.920 86.750 ;
        RECT 83.255 86.550 83.545 86.595 ;
        RECT 84.445 86.550 84.735 86.595 ;
        RECT 86.965 86.550 87.255 86.595 ;
        RECT 83.255 86.410 87.255 86.550 ;
        RECT 83.255 86.365 83.545 86.410 ;
        RECT 84.445 86.365 84.735 86.410 ;
        RECT 86.965 86.365 87.255 86.410 ;
        RECT 91.995 86.550 92.285 86.595 ;
        RECT 93.185 86.550 93.475 86.595 ;
        RECT 95.705 86.550 95.995 86.595 ;
        RECT 91.995 86.410 95.995 86.550 ;
        RECT 91.995 86.365 92.285 86.410 ;
        RECT 93.185 86.365 93.475 86.410 ;
        RECT 95.705 86.365 95.995 86.410 ;
        RECT 99.355 86.550 99.645 86.595 ;
        RECT 100.545 86.550 100.835 86.595 ;
        RECT 103.065 86.550 103.355 86.595 ;
        RECT 99.355 86.410 103.355 86.550 ;
        RECT 104.990 86.550 105.130 87.090 ;
        RECT 106.740 87.030 107.060 87.290 ;
        RECT 108.120 87.030 108.440 87.290 ;
        RECT 127.440 87.230 127.760 87.290 ;
        RECT 112.810 87.090 127.760 87.230 ;
        RECT 105.360 86.890 105.680 86.950 ;
        RECT 105.360 86.750 111.570 86.890 ;
        RECT 105.360 86.690 105.680 86.750 ;
        RECT 108.580 86.550 108.900 86.610 ;
        RECT 104.990 86.410 108.900 86.550 ;
        RECT 99.355 86.365 99.645 86.410 ;
        RECT 100.545 86.365 100.835 86.410 ;
        RECT 103.065 86.365 103.355 86.410 ;
        RECT 108.580 86.350 108.900 86.410 ;
        RECT 109.040 86.550 109.360 86.610 ;
        RECT 109.040 86.410 110.190 86.550 ;
        RECT 109.040 86.350 109.360 86.410 ;
        RECT 80.520 86.210 80.840 86.270 ;
        RECT 82.375 86.210 82.665 86.255 ;
        RECT 89.260 86.210 89.580 86.270 ;
        RECT 91.115 86.210 91.405 86.255 ;
        RECT 98.475 86.210 98.765 86.255 ;
        RECT 102.600 86.210 102.920 86.270 ;
        RECT 110.050 86.255 110.190 86.410 ;
        RECT 110.880 86.350 111.200 86.610 ;
        RECT 111.430 86.550 111.570 86.750 ;
        RECT 112.810 86.550 112.950 87.090 ;
        RECT 127.440 87.030 127.760 87.090 ;
        RECT 129.740 87.230 130.060 87.290 ;
        RECT 130.215 87.230 130.505 87.275 ;
        RECT 129.740 87.090 130.505 87.230 ;
        RECT 129.740 87.030 130.060 87.090 ;
        RECT 130.215 87.045 130.505 87.090 ;
        RECT 135.720 87.230 136.040 87.290 ;
        RECT 137.115 87.230 137.405 87.275 ;
        RECT 135.720 87.090 137.405 87.230 ;
        RECT 135.720 87.030 136.040 87.090 ;
        RECT 137.115 87.045 137.405 87.090 ;
        RECT 118.240 86.890 118.530 86.935 ;
        RECT 119.810 86.890 120.100 86.935 ;
        RECT 121.910 86.890 122.200 86.935 ;
        RECT 118.240 86.750 122.200 86.890 ;
        RECT 118.240 86.705 118.530 86.750 ;
        RECT 119.810 86.705 120.100 86.750 ;
        RECT 121.910 86.705 122.200 86.750 ;
        RECT 123.340 86.890 123.630 86.935 ;
        RECT 125.440 86.890 125.730 86.935 ;
        RECT 127.010 86.890 127.300 86.935 ;
        RECT 123.340 86.750 127.300 86.890 ;
        RECT 123.340 86.705 123.630 86.750 ;
        RECT 125.440 86.705 125.730 86.750 ;
        RECT 127.010 86.705 127.300 86.750 ;
        RECT 128.820 86.890 129.140 86.950 ;
        RECT 128.820 86.750 140.090 86.890 ;
        RECT 128.820 86.690 129.140 86.750 ;
        RECT 117.805 86.550 118.095 86.595 ;
        RECT 120.325 86.550 120.615 86.595 ;
        RECT 121.515 86.550 121.805 86.595 ;
        RECT 111.430 86.410 112.030 86.550 ;
        RECT 112.810 86.410 113.410 86.550 ;
        RECT 109.515 86.210 109.805 86.255 ;
        RECT 80.520 86.070 102.920 86.210 ;
        RECT 80.520 86.010 80.840 86.070 ;
        RECT 82.375 86.025 82.665 86.070 ;
        RECT 89.260 86.010 89.580 86.070 ;
        RECT 91.115 86.025 91.405 86.070 ;
        RECT 98.475 86.025 98.765 86.070 ;
        RECT 102.600 86.010 102.920 86.070 ;
        RECT 108.670 86.070 109.805 86.210 ;
        RECT 108.670 85.930 108.810 86.070 ;
        RECT 109.515 86.025 109.805 86.070 ;
        RECT 109.975 86.025 110.265 86.255 ;
        RECT 110.420 86.010 110.740 86.270 ;
        RECT 110.970 86.195 111.110 86.350 ;
        RECT 111.890 86.255 112.030 86.410 ;
        RECT 111.355 86.195 111.645 86.255 ;
        RECT 110.970 86.055 111.645 86.195 ;
        RECT 111.355 86.025 111.645 86.055 ;
        RECT 111.815 86.025 112.105 86.255 ;
        RECT 112.720 86.010 113.040 86.270 ;
        RECT 113.270 86.255 113.410 86.410 ;
        RECT 117.805 86.410 121.805 86.550 ;
        RECT 117.805 86.365 118.095 86.410 ;
        RECT 120.325 86.365 120.615 86.410 ;
        RECT 121.515 86.365 121.805 86.410 ;
        RECT 122.395 86.550 122.685 86.595 ;
        RECT 122.840 86.550 123.160 86.610 ;
        RECT 122.395 86.410 123.160 86.550 ;
        RECT 122.395 86.365 122.685 86.410 ;
        RECT 122.840 86.350 123.160 86.410 ;
        RECT 123.735 86.550 124.025 86.595 ;
        RECT 124.925 86.550 125.215 86.595 ;
        RECT 127.445 86.550 127.735 86.595 ;
        RECT 123.735 86.410 127.735 86.550 ;
        RECT 123.735 86.365 124.025 86.410 ;
        RECT 124.925 86.365 125.215 86.410 ;
        RECT 127.445 86.365 127.735 86.410 ;
        RECT 129.280 86.550 129.600 86.610 ;
        RECT 129.280 86.410 135.950 86.550 ;
        RECT 129.280 86.350 129.600 86.410 ;
        RECT 113.195 86.025 113.485 86.255 ;
        RECT 113.775 86.210 114.065 86.255 ;
        RECT 113.730 86.025 114.065 86.210 ;
        RECT 114.560 86.210 114.880 86.270 ;
        RECT 119.620 86.210 119.940 86.270 ;
        RECT 124.220 86.255 124.540 86.270 ;
        RECT 124.190 86.210 124.540 86.255 ;
        RECT 132.055 86.210 132.345 86.255 ;
        RECT 132.500 86.210 132.820 86.270 ;
        RECT 114.560 86.070 118.470 86.210 ;
        RECT 83.740 85.915 84.060 85.930 ;
        RECT 83.710 85.870 84.060 85.915 ;
        RECT 83.545 85.730 84.060 85.870 ;
        RECT 83.710 85.685 84.060 85.730 ;
        RECT 92.450 85.870 92.740 85.915 ;
        RECT 95.240 85.870 95.560 85.930 ;
        RECT 92.450 85.730 95.560 85.870 ;
        RECT 92.450 85.685 92.740 85.730 ;
        RECT 83.740 85.670 84.060 85.685 ;
        RECT 95.240 85.670 95.560 85.730 ;
        RECT 99.810 85.870 100.100 85.915 ;
        RECT 100.760 85.870 101.080 85.930 ;
        RECT 99.810 85.730 101.080 85.870 ;
        RECT 99.810 85.685 100.100 85.730 ;
        RECT 100.760 85.670 101.080 85.730 ;
        RECT 105.820 85.870 106.140 85.930 ;
        RECT 106.295 85.870 106.585 85.915 ;
        RECT 105.820 85.730 106.585 85.870 ;
        RECT 105.820 85.670 106.140 85.730 ;
        RECT 106.295 85.685 106.585 85.730 ;
        RECT 108.580 85.670 108.900 85.930 ;
        RECT 113.730 85.870 113.870 86.025 ;
        RECT 114.560 86.010 114.880 86.070 ;
        RECT 113.270 85.730 113.870 85.870 ;
        RECT 113.270 85.590 113.410 85.730 ;
        RECT 96.620 85.530 96.940 85.590 ;
        RECT 98.015 85.530 98.305 85.575 ;
        RECT 100.300 85.530 100.620 85.590 ;
        RECT 109.040 85.530 109.360 85.590 ;
        RECT 96.620 85.390 109.360 85.530 ;
        RECT 96.620 85.330 96.940 85.390 ;
        RECT 98.015 85.345 98.305 85.390 ;
        RECT 100.300 85.330 100.620 85.390 ;
        RECT 109.040 85.330 109.360 85.390 ;
        RECT 113.180 85.330 113.500 85.590 ;
        RECT 113.640 85.530 113.960 85.590 ;
        RECT 114.575 85.530 114.865 85.575 ;
        RECT 113.640 85.390 114.865 85.530 ;
        RECT 113.640 85.330 113.960 85.390 ;
        RECT 114.575 85.345 114.865 85.390 ;
        RECT 115.495 85.530 115.785 85.575 ;
        RECT 117.780 85.530 118.100 85.590 ;
        RECT 115.495 85.390 118.100 85.530 ;
        RECT 118.330 85.530 118.470 86.070 ;
        RECT 119.620 86.070 122.380 86.210 ;
        RECT 124.025 86.070 124.540 86.210 ;
        RECT 119.620 86.010 119.940 86.070 ;
        RECT 121.000 85.915 121.320 85.930 ;
        RECT 121.000 85.685 121.350 85.915 ;
        RECT 122.240 85.870 122.380 86.070 ;
        RECT 124.190 86.025 124.540 86.070 ;
        RECT 124.220 86.010 124.540 86.025 ;
        RECT 128.910 86.070 132.820 86.210 ;
        RECT 128.910 85.870 129.050 86.070 ;
        RECT 132.055 86.025 132.345 86.070 ;
        RECT 132.500 86.010 132.820 86.070 ;
        RECT 133.895 86.025 134.185 86.255 ;
        RECT 134.340 86.210 134.660 86.270 ;
        RECT 134.815 86.210 135.105 86.255 ;
        RECT 134.340 86.070 135.105 86.210 ;
        RECT 122.240 85.730 129.050 85.870 ;
        RECT 129.280 85.870 129.600 85.930 ;
        RECT 129.280 85.730 130.890 85.870 ;
        RECT 121.000 85.670 121.320 85.685 ;
        RECT 129.280 85.670 129.600 85.730 ;
        RECT 126.060 85.530 126.380 85.590 ;
        RECT 118.330 85.390 126.380 85.530 ;
        RECT 115.495 85.345 115.785 85.390 ;
        RECT 117.780 85.330 118.100 85.390 ;
        RECT 126.060 85.330 126.380 85.390 ;
        RECT 126.980 85.530 127.300 85.590 ;
        RECT 129.755 85.530 130.045 85.575 ;
        RECT 126.980 85.390 130.045 85.530 ;
        RECT 130.750 85.530 130.890 85.730 ;
        RECT 131.120 85.670 131.440 85.930 ;
        RECT 133.970 85.530 134.110 86.025 ;
        RECT 134.340 86.010 134.660 86.070 ;
        RECT 134.815 86.025 135.105 86.070 ;
        RECT 135.260 86.010 135.580 86.270 ;
        RECT 135.810 86.255 135.950 86.410 ;
        RECT 139.950 86.255 140.090 86.750 ;
        RECT 135.735 86.025 136.025 86.255 ;
        RECT 139.875 86.025 140.165 86.255 ;
        RECT 130.750 85.390 134.110 85.530 ;
        RECT 126.980 85.330 127.300 85.390 ;
        RECT 129.755 85.345 130.045 85.390 ;
        RECT 140.780 85.330 141.100 85.590 ;
        RECT 17.430 84.710 143.010 85.190 ;
        RECT 87.895 84.510 88.185 84.555 ;
        RECT 89.720 84.510 90.040 84.570 ;
        RECT 87.895 84.370 90.040 84.510 ;
        RECT 87.895 84.325 88.185 84.370 ;
        RECT 89.720 84.310 90.040 84.370 ;
        RECT 95.240 84.310 95.560 84.570 ;
        RECT 95.700 84.510 96.020 84.570 ;
        RECT 98.460 84.510 98.780 84.570 ;
        RECT 99.395 84.510 99.685 84.555 ;
        RECT 109.960 84.510 110.280 84.570 ;
        RECT 95.700 84.370 97.770 84.510 ;
        RECT 95.700 84.310 96.020 84.370 ;
        RECT 81.870 84.170 82.160 84.215 ;
        RECT 87.420 84.170 87.740 84.230 ;
        RECT 81.870 84.030 87.740 84.170 ;
        RECT 81.870 83.985 82.160 84.030 ;
        RECT 87.420 83.970 87.740 84.030 ;
        RECT 88.340 84.170 88.660 84.230 ;
        RECT 90.195 84.170 90.485 84.215 ;
        RECT 88.340 84.030 90.485 84.170 ;
        RECT 88.340 83.970 88.660 84.030 ;
        RECT 90.195 83.985 90.485 84.030 ;
        RECT 91.115 84.170 91.405 84.215 ;
        RECT 92.480 84.170 92.800 84.230 ;
        RECT 91.115 84.030 92.800 84.170 ;
        RECT 91.115 83.985 91.405 84.030 ;
        RECT 92.480 83.970 92.800 84.030 ;
        RECT 94.780 84.170 95.100 84.230 ;
        RECT 94.780 84.030 97.310 84.170 ;
        RECT 94.780 83.970 95.100 84.030 ;
        RECT 80.520 83.630 80.840 83.890 ;
        RECT 88.870 83.830 89.160 83.875 ;
        RECT 89.735 83.830 90.025 83.875 ;
        RECT 92.035 83.830 92.325 83.875 ;
        RECT 88.870 83.690 89.445 83.830 ;
        RECT 88.870 83.645 89.160 83.690 ;
        RECT 81.415 83.490 81.705 83.535 ;
        RECT 82.605 83.490 82.895 83.535 ;
        RECT 85.125 83.490 85.415 83.535 ;
        RECT 81.415 83.350 85.415 83.490 ;
        RECT 81.415 83.305 81.705 83.350 ;
        RECT 82.605 83.305 82.895 83.350 ;
        RECT 85.125 83.305 85.415 83.350 ;
        RECT 89.305 83.490 89.445 83.690 ;
        RECT 89.735 83.690 92.325 83.830 ;
        RECT 89.735 83.645 90.025 83.690 ;
        RECT 92.035 83.645 92.325 83.690 ;
        RECT 91.560 83.490 91.880 83.550 ;
        RECT 89.305 83.350 91.880 83.490 ;
        RECT 92.110 83.490 92.250 83.645 ;
        RECT 96.620 83.630 96.940 83.890 ;
        RECT 97.170 83.875 97.310 84.030 ;
        RECT 97.630 83.875 97.770 84.370 ;
        RECT 98.460 84.370 99.685 84.510 ;
        RECT 98.460 84.310 98.780 84.370 ;
        RECT 99.395 84.325 99.685 84.370 ;
        RECT 108.210 84.370 110.280 84.510 ;
        RECT 100.315 84.170 100.605 84.215 ;
        RECT 103.520 84.170 103.840 84.230 ;
        RECT 105.360 84.170 105.680 84.230 ;
        RECT 100.315 84.030 105.680 84.170 ;
        RECT 100.315 83.985 100.605 84.030 ;
        RECT 103.520 83.970 103.840 84.030 ;
        RECT 105.360 83.970 105.680 84.030 ;
        RECT 107.370 84.170 107.660 84.215 ;
        RECT 108.210 84.170 108.350 84.370 ;
        RECT 109.960 84.310 110.280 84.370 ;
        RECT 110.880 84.310 111.200 84.570 ;
        RECT 111.340 84.510 111.660 84.570 ;
        RECT 113.195 84.510 113.485 84.555 ;
        RECT 111.340 84.370 113.485 84.510 ;
        RECT 111.340 84.310 111.660 84.370 ;
        RECT 113.195 84.325 113.485 84.370 ;
        RECT 113.640 84.510 113.960 84.570 ;
        RECT 117.320 84.510 117.640 84.570 ;
        RECT 119.175 84.510 119.465 84.555 ;
        RECT 113.640 84.370 116.170 84.510 ;
        RECT 113.640 84.310 113.960 84.370 ;
        RECT 107.370 84.030 108.350 84.170 ;
        RECT 113.270 84.030 114.330 84.170 ;
        RECT 107.370 83.985 107.660 84.030 ;
        RECT 113.270 83.890 113.410 84.030 ;
        RECT 97.095 83.645 97.385 83.875 ;
        RECT 97.555 83.645 97.845 83.875 ;
        RECT 98.460 83.630 98.780 83.890 ;
        RECT 98.920 83.830 99.240 83.890 ;
        RECT 101.220 83.830 101.540 83.890 ;
        RECT 105.820 83.830 106.140 83.890 ;
        RECT 98.920 83.690 101.540 83.830 ;
        RECT 98.920 83.630 99.240 83.690 ;
        RECT 101.220 83.630 101.540 83.690 ;
        RECT 103.610 83.690 106.140 83.830 ;
        RECT 99.010 83.490 99.150 83.630 ;
        RECT 92.110 83.350 99.150 83.490 ;
        RECT 81.020 83.150 81.310 83.195 ;
        RECT 83.120 83.150 83.410 83.195 ;
        RECT 84.690 83.150 84.980 83.195 ;
        RECT 81.020 83.010 84.980 83.150 ;
        RECT 81.020 82.965 81.310 83.010 ;
        RECT 83.120 82.965 83.410 83.010 ;
        RECT 84.690 82.965 84.980 83.010 ;
        RECT 87.435 83.150 87.725 83.195 ;
        RECT 87.880 83.150 88.200 83.210 ;
        RECT 89.305 83.150 89.445 83.350 ;
        RECT 91.560 83.290 91.880 83.350 ;
        RECT 87.435 83.010 89.445 83.150 ;
        RECT 97.080 83.150 97.400 83.210 ;
        RECT 98.460 83.150 98.780 83.210 ;
        RECT 103.610 83.150 103.750 83.690 ;
        RECT 105.820 83.630 106.140 83.690 ;
        RECT 109.055 83.830 109.345 83.875 ;
        RECT 109.500 83.830 109.820 83.890 ;
        RECT 109.055 83.690 109.820 83.830 ;
        RECT 109.055 83.645 109.345 83.690 ;
        RECT 109.500 83.630 109.820 83.690 ;
        RECT 109.975 83.830 110.265 83.875 ;
        RECT 110.420 83.830 110.740 83.890 ;
        RECT 109.975 83.690 110.740 83.830 ;
        RECT 109.975 83.645 110.265 83.690 ;
        RECT 110.420 83.630 110.740 83.690 ;
        RECT 113.180 83.630 113.500 83.890 ;
        RECT 114.190 83.875 114.330 84.030 ;
        RECT 115.020 83.970 115.340 84.230 ;
        RECT 116.030 83.875 116.170 84.370 ;
        RECT 117.320 84.370 119.465 84.510 ;
        RECT 117.320 84.310 117.640 84.370 ;
        RECT 119.175 84.325 119.465 84.370 ;
        RECT 121.000 84.310 121.320 84.570 ;
        RECT 122.840 84.510 123.160 84.570 ;
        RECT 122.240 84.370 123.160 84.510 ;
        RECT 116.860 84.170 117.180 84.230 ;
        RECT 122.240 84.170 122.380 84.370 ;
        RECT 122.840 84.310 123.160 84.370 ;
        RECT 124.220 84.510 124.540 84.570 ;
        RECT 128.360 84.510 128.680 84.570 ;
        RECT 124.220 84.370 128.680 84.510 ;
        RECT 124.220 84.310 124.540 84.370 ;
        RECT 128.360 84.310 128.680 84.370 ;
        RECT 131.120 84.510 131.440 84.570 ;
        RECT 132.055 84.510 132.345 84.555 ;
        RECT 131.120 84.370 132.345 84.510 ;
        RECT 131.120 84.310 131.440 84.370 ;
        RECT 132.055 84.325 132.345 84.370 ;
        RECT 134.340 84.310 134.660 84.570 ;
        RECT 126.520 84.215 126.840 84.230 ;
        RECT 126.490 84.170 126.840 84.215 ;
        RECT 116.860 84.030 125.370 84.170 ;
        RECT 126.325 84.030 126.840 84.170 ;
        RECT 116.860 83.970 117.180 84.030 ;
        RECT 113.995 83.690 114.330 83.875 ;
        RECT 113.995 83.645 114.285 83.690 ;
        RECT 114.575 83.645 114.865 83.875 ;
        RECT 115.955 83.645 116.245 83.875 ;
        RECT 104.005 83.490 104.295 83.535 ;
        RECT 106.525 83.490 106.815 83.535 ;
        RECT 107.715 83.490 108.005 83.535 ;
        RECT 104.005 83.350 108.005 83.490 ;
        RECT 104.005 83.305 104.295 83.350 ;
        RECT 106.525 83.305 106.815 83.350 ;
        RECT 107.715 83.305 108.005 83.350 ;
        RECT 108.595 83.305 108.885 83.535 ;
        RECT 112.720 83.490 113.040 83.550 ;
        RECT 114.650 83.490 114.790 83.645 ;
        RECT 116.400 83.630 116.720 83.890 ;
        RECT 117.320 83.630 117.640 83.890 ;
        RECT 117.780 83.630 118.100 83.890 ;
        RECT 118.255 83.830 118.545 83.875 ;
        RECT 118.700 83.830 119.020 83.890 ;
        RECT 118.255 83.690 119.020 83.830 ;
        RECT 118.255 83.645 118.545 83.690 ;
        RECT 118.700 83.630 119.020 83.690 ;
        RECT 122.380 83.630 122.700 83.890 ;
        RECT 122.855 83.645 123.145 83.875 ;
        RECT 112.720 83.350 114.790 83.490 ;
        RECT 122.930 83.490 123.070 83.645 ;
        RECT 123.300 83.630 123.620 83.890 ;
        RECT 124.220 83.630 124.540 83.890 ;
        RECT 125.230 83.875 125.370 84.030 ;
        RECT 126.490 83.985 126.840 84.030 ;
        RECT 126.520 83.970 126.840 83.985 ;
        RECT 127.440 83.970 127.760 84.230 ;
        RECT 132.500 83.970 132.820 84.230 ;
        RECT 125.155 83.645 125.445 83.875 ;
        RECT 127.530 83.830 127.670 83.970 ;
        RECT 133.435 83.830 133.725 83.875 ;
        RECT 136.180 83.830 136.500 83.890 ;
        RECT 127.530 83.690 136.500 83.830 ;
        RECT 133.435 83.645 133.725 83.690 ;
        RECT 136.180 83.630 136.500 83.690 ;
        RECT 138.020 83.830 138.340 83.890 ;
        RECT 139.875 83.830 140.165 83.875 ;
        RECT 138.020 83.690 140.165 83.830 ;
        RECT 138.020 83.630 138.340 83.690 ;
        RECT 139.875 83.645 140.165 83.690 ;
        RECT 124.680 83.490 125.000 83.550 ;
        RECT 122.930 83.350 125.000 83.490 ;
        RECT 97.080 83.010 103.750 83.150 ;
        RECT 104.440 83.150 104.730 83.195 ;
        RECT 106.010 83.150 106.300 83.195 ;
        RECT 108.110 83.150 108.400 83.195 ;
        RECT 104.440 83.010 108.400 83.150 ;
        RECT 108.670 83.150 108.810 83.305 ;
        RECT 112.720 83.290 113.040 83.350 ;
        RECT 124.680 83.290 125.000 83.350 ;
        RECT 126.035 83.490 126.325 83.535 ;
        RECT 127.225 83.490 127.515 83.535 ;
        RECT 129.745 83.490 130.035 83.535 ;
        RECT 126.035 83.350 130.035 83.490 ;
        RECT 126.035 83.305 126.325 83.350 ;
        RECT 127.225 83.305 127.515 83.350 ;
        RECT 129.745 83.305 130.035 83.350 ;
        RECT 125.640 83.150 125.930 83.195 ;
        RECT 127.740 83.150 128.030 83.195 ;
        RECT 129.310 83.150 129.600 83.195 ;
        RECT 108.670 83.010 115.710 83.150 ;
        RECT 87.435 82.965 87.725 83.010 ;
        RECT 87.880 82.950 88.200 83.010 ;
        RECT 97.080 82.950 97.400 83.010 ;
        RECT 98.460 82.950 98.780 83.010 ;
        RECT 104.440 82.965 104.730 83.010 ;
        RECT 106.010 82.965 106.300 83.010 ;
        RECT 108.110 82.965 108.400 83.010 ;
        RECT 101.695 82.810 101.985 82.855 ;
        RECT 104.900 82.810 105.220 82.870 ;
        RECT 101.695 82.670 105.220 82.810 ;
        RECT 101.695 82.625 101.985 82.670 ;
        RECT 104.900 82.610 105.220 82.670 ;
        RECT 108.580 82.810 108.900 82.870 ;
        RECT 111.340 82.810 111.660 82.870 ;
        RECT 114.560 82.810 114.880 82.870 ;
        RECT 108.580 82.670 114.880 82.810 ;
        RECT 115.570 82.810 115.710 83.010 ;
        RECT 125.640 83.010 129.600 83.150 ;
        RECT 125.640 82.965 125.930 83.010 ;
        RECT 127.740 82.965 128.030 83.010 ;
        RECT 129.310 82.965 129.600 83.010 ;
        RECT 116.860 82.810 117.180 82.870 ;
        RECT 115.570 82.670 117.180 82.810 ;
        RECT 108.580 82.610 108.900 82.670 ;
        RECT 111.340 82.610 111.660 82.670 ;
        RECT 114.560 82.610 114.880 82.670 ;
        RECT 116.860 82.610 117.180 82.670 ;
        RECT 117.320 82.810 117.640 82.870 ;
        RECT 119.620 82.810 119.940 82.870 ;
        RECT 117.320 82.670 119.940 82.810 ;
        RECT 117.320 82.610 117.640 82.670 ;
        RECT 119.620 82.610 119.940 82.670 ;
        RECT 140.780 82.610 141.100 82.870 ;
        RECT 17.430 81.990 143.010 82.470 ;
        RECT 63.960 81.790 64.280 81.850 ;
        RECT 64.895 81.790 65.185 81.835 ;
        RECT 63.960 81.650 65.185 81.790 ;
        RECT 63.960 81.590 64.280 81.650 ;
        RECT 64.895 81.605 65.185 81.650 ;
        RECT 104.900 81.790 105.220 81.850 ;
        RECT 118.240 81.790 118.560 81.850 ;
        RECT 121.935 81.790 122.225 81.835 ;
        RECT 104.900 81.650 109.730 81.790 ;
        RECT 104.900 81.590 105.220 81.650 ;
        RECT 105.360 81.450 105.680 81.510 ;
        RECT 108.595 81.450 108.885 81.495 ;
        RECT 105.360 81.310 108.885 81.450 ;
        RECT 105.360 81.250 105.680 81.310 ;
        RECT 108.595 81.265 108.885 81.310 ;
        RECT 75.000 80.910 75.320 81.170 ;
        RECT 101.680 81.110 102.000 81.170 ;
        RECT 109.040 81.110 109.360 81.170 ;
        RECT 101.680 80.970 109.360 81.110 ;
        RECT 101.680 80.910 102.000 80.970 ;
        RECT 63.500 80.770 63.820 80.830 ;
        RECT 63.975 80.770 64.265 80.815 ;
        RECT 63.500 80.630 64.265 80.770 ;
        RECT 63.500 80.570 63.820 80.630 ;
        RECT 63.975 80.585 64.265 80.630 ;
        RECT 71.780 80.570 72.100 80.830 ;
        RECT 73.160 80.770 73.480 80.830 ;
        RECT 73.635 80.770 73.925 80.815 ;
        RECT 73.160 80.630 73.925 80.770 ;
        RECT 73.160 80.570 73.480 80.630 ;
        RECT 73.635 80.585 73.925 80.630 ;
        RECT 79.615 80.770 79.905 80.815 ;
        RECT 80.980 80.770 81.300 80.830 ;
        RECT 79.615 80.630 81.300 80.770 ;
        RECT 79.615 80.585 79.905 80.630 ;
        RECT 80.980 80.570 81.300 80.630 ;
        RECT 81.440 80.570 81.760 80.830 ;
        RECT 81.900 80.770 82.220 80.830 ;
        RECT 84.675 80.770 84.965 80.815 ;
        RECT 81.900 80.630 84.965 80.770 ;
        RECT 81.900 80.570 82.220 80.630 ;
        RECT 84.675 80.585 84.965 80.630 ;
        RECT 87.880 80.570 88.200 80.830 ;
        RECT 91.115 80.770 91.405 80.815 ;
        RECT 92.480 80.770 92.800 80.830 ;
        RECT 91.115 80.630 92.800 80.770 ;
        RECT 91.115 80.585 91.405 80.630 ;
        RECT 92.480 80.570 92.800 80.630 ;
        RECT 94.335 80.770 94.625 80.815 ;
        RECT 96.160 80.770 96.480 80.830 ;
        RECT 94.335 80.630 96.480 80.770 ;
        RECT 94.335 80.585 94.625 80.630 ;
        RECT 96.160 80.570 96.480 80.630 ;
        RECT 97.555 80.770 97.845 80.815 ;
        RECT 98.000 80.770 98.320 80.830 ;
        RECT 97.555 80.630 98.320 80.770 ;
        RECT 97.555 80.585 97.845 80.630 ;
        RECT 98.000 80.570 98.320 80.630 ;
        RECT 100.760 80.570 101.080 80.830 ;
        RECT 103.520 80.570 103.840 80.830 ;
        RECT 104.070 80.815 104.210 80.970 ;
        RECT 109.040 80.910 109.360 80.970 ;
        RECT 109.590 81.110 109.730 81.650 ;
        RECT 118.240 81.650 122.225 81.790 ;
        RECT 118.240 81.590 118.560 81.650 ;
        RECT 121.935 81.605 122.225 81.650 ;
        RECT 113.640 81.250 113.960 81.510 ;
        RECT 119.635 81.450 119.925 81.495 ;
        RECT 123.300 81.450 123.620 81.510 ;
        RECT 119.635 81.310 123.620 81.450 ;
        RECT 119.635 81.265 119.925 81.310 ;
        RECT 123.300 81.250 123.620 81.310 ;
        RECT 123.775 81.265 124.065 81.495 ;
        RECT 113.730 81.110 113.870 81.250 ;
        RECT 109.590 80.970 113.870 81.110 ;
        RECT 116.400 81.110 116.720 81.170 ;
        RECT 123.850 81.110 123.990 81.265 ;
        RECT 116.400 80.970 121.230 81.110 ;
        RECT 103.995 80.770 104.285 80.815 ;
        RECT 103.995 80.630 104.395 80.770 ;
        RECT 103.995 80.585 104.285 80.630 ;
        RECT 104.900 80.570 105.220 80.830 ;
        RECT 109.590 80.815 109.730 80.970 ;
        RECT 116.400 80.910 116.720 80.970 ;
        RECT 109.515 80.585 109.805 80.815 ;
        RECT 110.420 80.770 110.740 80.830 ;
        RECT 111.355 80.770 111.645 80.815 ;
        RECT 110.420 80.630 111.645 80.770 ;
        RECT 110.420 80.570 110.740 80.630 ;
        RECT 111.355 80.585 111.645 80.630 ;
        RECT 113.655 80.770 113.945 80.815 ;
        RECT 114.100 80.770 114.420 80.830 ;
        RECT 113.655 80.630 114.420 80.770 ;
        RECT 113.655 80.585 113.945 80.630 ;
        RECT 114.100 80.570 114.420 80.630 ;
        RECT 115.480 80.570 115.800 80.830 ;
        RECT 117.320 80.770 117.640 80.830 ;
        RECT 121.090 80.815 121.230 80.970 ;
        RECT 122.240 80.970 123.990 81.110 ;
        RECT 117.795 80.770 118.085 80.815 ;
        RECT 117.320 80.630 118.085 80.770 ;
        RECT 117.320 80.570 117.640 80.630 ;
        RECT 117.795 80.585 118.085 80.630 ;
        RECT 121.015 80.585 121.305 80.815 ;
        RECT 121.460 80.770 121.780 80.830 ;
        RECT 122.240 80.770 122.380 80.970 ;
        RECT 121.460 80.630 122.380 80.770 ;
        RECT 121.460 80.570 121.780 80.630 ;
        RECT 122.855 80.585 123.145 80.815 ;
        RECT 126.535 80.770 126.825 80.815 ;
        RECT 126.980 80.770 127.300 80.830 ;
        RECT 126.535 80.630 127.300 80.770 ;
        RECT 126.535 80.585 126.825 80.630 ;
        RECT 105.835 80.430 106.125 80.475 ;
        RECT 112.260 80.430 112.580 80.490 ;
        RECT 118.715 80.430 119.005 80.475 ;
        RECT 122.930 80.430 123.070 80.585 ;
        RECT 126.980 80.570 127.300 80.630 ;
        RECT 127.900 80.770 128.220 80.830 ;
        RECT 128.375 80.770 128.665 80.815 ;
        RECT 127.900 80.630 128.665 80.770 ;
        RECT 127.900 80.570 128.220 80.630 ;
        RECT 128.375 80.585 128.665 80.630 ;
        RECT 131.120 80.770 131.440 80.830 ;
        RECT 131.595 80.770 131.885 80.815 ;
        RECT 131.120 80.630 131.885 80.770 ;
        RECT 131.120 80.570 131.440 80.630 ;
        RECT 131.595 80.585 131.885 80.630 ;
        RECT 136.180 80.570 136.500 80.830 ;
        RECT 105.835 80.290 112.580 80.430 ;
        RECT 105.835 80.245 106.125 80.290 ;
        RECT 112.260 80.230 112.580 80.290 ;
        RECT 117.870 80.290 123.070 80.430 ;
        RECT 117.870 80.150 118.010 80.290 ;
        RECT 118.715 80.245 119.005 80.290 ;
        RECT 69.940 80.090 70.260 80.150 ;
        RECT 70.875 80.090 71.165 80.135 ;
        RECT 69.940 79.950 71.165 80.090 ;
        RECT 69.940 79.890 70.260 79.950 ;
        RECT 70.875 79.905 71.165 79.950 ;
        RECT 76.380 80.090 76.700 80.150 ;
        RECT 78.695 80.090 78.985 80.135 ;
        RECT 76.380 79.950 78.985 80.090 ;
        RECT 76.380 79.890 76.700 79.950 ;
        RECT 78.695 79.905 78.985 79.950 ;
        RECT 79.600 80.090 79.920 80.150 ;
        RECT 80.535 80.090 80.825 80.135 ;
        RECT 79.600 79.950 80.825 80.090 ;
        RECT 79.600 79.890 79.920 79.950 ;
        RECT 80.535 79.905 80.825 79.950 ;
        RECT 82.820 80.090 83.140 80.150 ;
        RECT 83.755 80.090 84.045 80.135 ;
        RECT 82.820 79.950 84.045 80.090 ;
        RECT 82.820 79.890 83.140 79.950 ;
        RECT 83.755 79.905 84.045 79.950 ;
        RECT 86.040 80.090 86.360 80.150 ;
        RECT 86.975 80.090 87.265 80.135 ;
        RECT 86.040 79.950 87.265 80.090 ;
        RECT 86.040 79.890 86.360 79.950 ;
        RECT 86.975 79.905 87.265 79.950 ;
        RECT 89.260 80.090 89.580 80.150 ;
        RECT 90.195 80.090 90.485 80.135 ;
        RECT 89.260 79.950 90.485 80.090 ;
        RECT 89.260 79.890 89.580 79.950 ;
        RECT 90.195 79.905 90.485 79.950 ;
        RECT 92.480 80.090 92.800 80.150 ;
        RECT 93.415 80.090 93.705 80.135 ;
        RECT 92.480 79.950 93.705 80.090 ;
        RECT 92.480 79.890 92.800 79.950 ;
        RECT 93.415 79.905 93.705 79.950 ;
        RECT 95.700 80.090 96.020 80.150 ;
        RECT 96.635 80.090 96.925 80.135 ;
        RECT 95.700 79.950 96.925 80.090 ;
        RECT 95.700 79.890 96.020 79.950 ;
        RECT 96.635 79.905 96.925 79.950 ;
        RECT 98.920 80.090 99.240 80.150 ;
        RECT 99.855 80.090 100.145 80.135 ;
        RECT 98.920 79.950 100.145 80.090 ;
        RECT 98.920 79.890 99.240 79.950 ;
        RECT 99.855 79.905 100.145 79.950 ;
        RECT 102.140 80.090 102.460 80.150 ;
        RECT 102.615 80.090 102.905 80.135 ;
        RECT 102.140 79.950 102.905 80.090 ;
        RECT 102.140 79.890 102.460 79.950 ;
        RECT 102.615 79.905 102.905 79.950 ;
        RECT 109.040 80.090 109.360 80.150 ;
        RECT 110.435 80.090 110.725 80.135 ;
        RECT 109.040 79.950 110.725 80.090 ;
        RECT 109.040 79.890 109.360 79.950 ;
        RECT 110.435 79.905 110.725 79.950 ;
        RECT 111.800 80.090 112.120 80.150 ;
        RECT 112.735 80.090 113.025 80.135 ;
        RECT 111.800 79.950 113.025 80.090 ;
        RECT 111.800 79.890 112.120 79.950 ;
        RECT 112.735 79.905 113.025 79.950 ;
        RECT 115.020 80.090 115.340 80.150 ;
        RECT 116.415 80.090 116.705 80.135 ;
        RECT 115.020 79.950 116.705 80.090 ;
        RECT 115.020 79.890 115.340 79.950 ;
        RECT 116.415 79.905 116.705 79.950 ;
        RECT 117.780 79.890 118.100 80.150 ;
        RECT 124.680 80.090 125.000 80.150 ;
        RECT 125.615 80.090 125.905 80.135 ;
        RECT 124.680 79.950 125.905 80.090 ;
        RECT 124.680 79.890 125.000 79.950 ;
        RECT 125.615 79.905 125.905 79.950 ;
        RECT 127.900 80.090 128.220 80.150 ;
        RECT 129.295 80.090 129.585 80.135 ;
        RECT 127.900 79.950 129.585 80.090 ;
        RECT 127.900 79.890 128.220 79.950 ;
        RECT 129.295 79.905 129.585 79.950 ;
        RECT 131.120 80.090 131.440 80.150 ;
        RECT 132.515 80.090 132.805 80.135 ;
        RECT 131.120 79.950 132.805 80.090 ;
        RECT 131.120 79.890 131.440 79.950 ;
        RECT 132.515 79.905 132.805 79.950 ;
        RECT 134.340 80.090 134.660 80.150 ;
        RECT 135.275 80.090 135.565 80.135 ;
        RECT 134.340 79.950 135.565 80.090 ;
        RECT 134.340 79.890 134.660 79.950 ;
        RECT 135.275 79.905 135.565 79.950 ;
        RECT 17.430 79.270 143.010 79.750 ;
        RECT 12.750 48.490 48.630 48.970 ;
        RECT 21.575 48.290 21.865 48.335 ;
        RECT 26.620 48.290 26.940 48.350 ;
        RECT 21.575 48.150 26.940 48.290 ;
        RECT 21.575 48.105 21.865 48.150 ;
        RECT 26.620 48.090 26.940 48.150 ;
        RECT 32.155 48.290 32.445 48.335 ;
        RECT 33.060 48.290 33.380 48.350 ;
        RECT 32.155 48.150 33.380 48.290 ;
        RECT 32.155 48.105 32.445 48.150 ;
        RECT 33.060 48.090 33.380 48.150 ;
        RECT 39.500 48.290 39.820 48.350 ;
        RECT 40.435 48.290 40.725 48.335 ;
        RECT 39.500 48.150 40.725 48.290 ;
        RECT 39.500 48.090 39.820 48.150 ;
        RECT 40.435 48.105 40.725 48.150 ;
        RECT 23.875 47.950 24.165 47.995 ;
        RECT 31.220 47.950 31.540 48.010 ;
        RECT 38.120 47.950 38.440 48.010 ;
        RECT 23.875 47.810 31.540 47.950 ;
        RECT 23.875 47.765 24.165 47.810 ;
        RECT 31.220 47.750 31.540 47.810 ;
        RECT 32.690 47.810 38.440 47.950 ;
        RECT 27.095 47.610 27.385 47.655 ;
        RECT 20.730 47.470 27.385 47.610 ;
        RECT 18.340 47.270 18.660 47.330 ;
        RECT 20.730 47.315 20.870 47.470 ;
        RECT 27.095 47.425 27.385 47.470 ;
        RECT 20.655 47.270 20.945 47.315 ;
        RECT 18.340 47.130 20.945 47.270 ;
        RECT 18.340 47.070 18.660 47.130 ;
        RECT 20.655 47.085 20.945 47.130 ;
        RECT 22.940 47.070 23.260 47.330 ;
        RECT 23.400 47.070 23.720 47.330 ;
        RECT 24.335 47.270 24.625 47.315 ;
        RECT 32.690 47.270 32.830 47.810 ;
        RECT 38.120 47.750 38.440 47.810 ;
        RECT 24.335 47.130 32.830 47.270 ;
        RECT 33.075 47.270 33.365 47.315 ;
        RECT 33.520 47.270 33.840 47.330 ;
        RECT 33.075 47.130 33.840 47.270 ;
        RECT 24.335 47.085 24.625 47.130 ;
        RECT 33.075 47.085 33.365 47.130 ;
        RECT 33.520 47.070 33.840 47.130 ;
        RECT 36.280 47.270 36.600 47.330 ;
        RECT 37.215 47.270 37.505 47.315 ;
        RECT 36.280 47.130 37.505 47.270 ;
        RECT 36.280 47.070 36.600 47.130 ;
        RECT 37.215 47.085 37.505 47.130 ;
        RECT 41.340 47.070 41.660 47.330 ;
        RECT 44.100 47.070 44.420 47.330 ;
        RECT 45.480 47.070 45.800 47.330 ;
        RECT 46.860 47.070 47.180 47.330 ;
        RECT 25.240 46.390 25.560 46.650 ;
        RECT 30.300 46.390 30.620 46.650 ;
        RECT 33.980 46.590 34.300 46.650 ;
        RECT 36.755 46.590 37.045 46.635 ;
        RECT 33.980 46.450 37.045 46.590 ;
        RECT 33.980 46.390 34.300 46.450 ;
        RECT 36.755 46.405 37.045 46.450 ;
        RECT 39.960 46.590 40.280 46.650 ;
        RECT 43.195 46.590 43.485 46.635 ;
        RECT 39.960 46.450 43.485 46.590 ;
        RECT 39.960 46.390 40.280 46.450 ;
        RECT 43.195 46.405 43.485 46.450 ;
        RECT 43.640 46.590 43.960 46.650 ;
        RECT 44.575 46.590 44.865 46.635 ;
        RECT 43.640 46.450 44.865 46.590 ;
        RECT 43.640 46.390 43.960 46.450 ;
        RECT 44.575 46.405 44.865 46.450 ;
        RECT 45.955 46.590 46.245 46.635 ;
        RECT 46.400 46.590 46.720 46.650 ;
        RECT 45.955 46.450 46.720 46.590 ;
        RECT 45.955 46.405 46.245 46.450 ;
        RECT 46.400 46.390 46.720 46.450 ;
        RECT 12.750 45.770 48.630 46.250 ;
        RECT 18.340 45.370 18.660 45.630 ;
        RECT 22.940 45.570 23.260 45.630 ;
        RECT 32.615 45.570 32.905 45.615 ;
        RECT 33.520 45.570 33.840 45.630 ;
        RECT 22.940 45.430 28.230 45.570 ;
        RECT 22.940 45.370 23.260 45.430 ;
        RECT 25.240 45.230 25.560 45.290 ;
        RECT 26.940 45.230 27.230 45.275 ;
        RECT 25.240 45.090 27.230 45.230 ;
        RECT 28.090 45.230 28.230 45.430 ;
        RECT 32.615 45.430 33.840 45.570 ;
        RECT 32.615 45.385 32.905 45.430 ;
        RECT 33.520 45.370 33.840 45.430 ;
        RECT 33.075 45.230 33.365 45.275 ;
        RECT 28.090 45.090 33.365 45.230 ;
        RECT 25.240 45.030 25.560 45.090 ;
        RECT 26.940 45.045 27.230 45.090 ;
        RECT 33.075 45.045 33.365 45.090 ;
        RECT 33.980 45.030 34.300 45.290 ;
        RECT 23.975 44.890 24.265 44.935 ;
        RECT 26.160 44.890 26.480 44.950 ;
        RECT 23.975 44.750 26.480 44.890 ;
        RECT 23.975 44.705 24.265 44.750 ;
        RECT 26.160 44.690 26.480 44.750 ;
        RECT 34.900 44.690 35.220 44.950 ;
        RECT 35.375 44.705 35.665 44.935 ;
        RECT 36.280 44.890 36.600 44.950 ;
        RECT 37.215 44.890 37.505 44.935 ;
        RECT 36.280 44.750 37.505 44.890 ;
        RECT 20.665 44.550 20.955 44.595 ;
        RECT 23.185 44.550 23.475 44.595 ;
        RECT 24.375 44.550 24.665 44.595 ;
        RECT 20.665 44.410 24.665 44.550 ;
        RECT 20.665 44.365 20.955 44.410 ;
        RECT 23.185 44.365 23.475 44.410 ;
        RECT 24.375 44.365 24.665 44.410 ;
        RECT 25.255 44.550 25.545 44.595 ;
        RECT 25.715 44.550 26.005 44.595 ;
        RECT 25.255 44.410 26.005 44.550 ;
        RECT 25.255 44.365 25.545 44.410 ;
        RECT 25.715 44.365 26.005 44.410 ;
        RECT 26.595 44.550 26.885 44.595 ;
        RECT 27.785 44.550 28.075 44.595 ;
        RECT 30.305 44.550 30.595 44.595 ;
        RECT 26.595 44.410 30.595 44.550 ;
        RECT 26.595 44.365 26.885 44.410 ;
        RECT 27.785 44.365 28.075 44.410 ;
        RECT 30.305 44.365 30.595 44.410 ;
        RECT 31.680 44.550 32.000 44.610 ;
        RECT 35.450 44.550 35.590 44.705 ;
        RECT 36.280 44.690 36.600 44.750 ;
        RECT 37.215 44.705 37.505 44.750 ;
        RECT 38.120 44.890 38.440 44.950 ;
        RECT 39.975 44.890 40.265 44.935 ;
        RECT 38.120 44.750 40.265 44.890 ;
        RECT 38.120 44.690 38.440 44.750 ;
        RECT 39.975 44.705 40.265 44.750 ;
        RECT 40.880 44.690 41.200 44.950 ;
        RECT 41.355 44.890 41.645 44.935 ;
        RECT 44.100 44.890 44.420 44.950 ;
        RECT 41.355 44.750 44.420 44.890 ;
        RECT 41.355 44.705 41.645 44.750 ;
        RECT 44.100 44.690 44.420 44.750 ;
        RECT 46.860 44.690 47.180 44.950 ;
        RECT 31.680 44.410 35.590 44.550 ;
        RECT 35.820 44.550 36.140 44.610 ;
        RECT 38.210 44.550 38.350 44.690 ;
        RECT 35.820 44.410 38.350 44.550 ;
        RECT 21.100 44.210 21.390 44.255 ;
        RECT 22.670 44.210 22.960 44.255 ;
        RECT 24.770 44.210 25.060 44.255 ;
        RECT 21.100 44.070 25.060 44.210 ;
        RECT 21.100 44.025 21.390 44.070 ;
        RECT 22.670 44.025 22.960 44.070 ;
        RECT 24.770 44.025 25.060 44.070 ;
        RECT 23.860 43.870 24.180 43.930 ;
        RECT 25.790 43.870 25.930 44.365 ;
        RECT 31.680 44.350 32.000 44.410 ;
        RECT 35.820 44.350 36.140 44.410 ;
        RECT 42.275 44.365 42.565 44.595 ;
        RECT 26.200 44.210 26.490 44.255 ;
        RECT 28.300 44.210 28.590 44.255 ;
        RECT 29.870 44.210 30.160 44.255 ;
        RECT 26.200 44.070 30.160 44.210 ;
        RECT 26.200 44.025 26.490 44.070 ;
        RECT 28.300 44.025 28.590 44.070 ;
        RECT 29.870 44.025 30.160 44.070 ;
        RECT 30.760 44.210 31.080 44.270 ;
        RECT 36.295 44.210 36.585 44.255 ;
        RECT 30.760 44.070 36.585 44.210 ;
        RECT 30.760 44.010 31.080 44.070 ;
        RECT 36.295 44.025 36.585 44.070 ;
        RECT 37.675 44.210 37.965 44.255 ;
        RECT 40.435 44.210 40.725 44.255 ;
        RECT 37.675 44.070 40.725 44.210 ;
        RECT 37.675 44.025 37.965 44.070 ;
        RECT 40.435 44.025 40.725 44.070 ;
        RECT 41.340 44.210 41.660 44.270 ;
        RECT 42.350 44.210 42.490 44.365 ;
        RECT 41.340 44.070 42.490 44.210 ;
        RECT 44.560 44.210 44.880 44.270 ;
        RECT 45.955 44.210 46.245 44.255 ;
        RECT 44.560 44.070 46.245 44.210 ;
        RECT 41.340 44.010 41.660 44.070 ;
        RECT 44.560 44.010 44.880 44.070 ;
        RECT 45.955 44.025 46.245 44.070 ;
        RECT 34.440 43.870 34.760 43.930 ;
        RECT 23.860 43.730 34.760 43.870 ;
        RECT 23.860 43.670 24.180 43.730 ;
        RECT 34.440 43.670 34.760 43.730 ;
        RECT 37.200 43.870 37.520 43.930 ;
        RECT 39.055 43.870 39.345 43.915 ;
        RECT 37.200 43.730 39.345 43.870 ;
        RECT 37.200 43.670 37.520 43.730 ;
        RECT 39.055 43.685 39.345 43.730 ;
        RECT 43.180 43.870 43.500 43.930 ;
        RECT 45.495 43.870 45.785 43.915 ;
        RECT 43.180 43.730 45.785 43.870 ;
        RECT 43.180 43.670 43.500 43.730 ;
        RECT 45.495 43.685 45.785 43.730 ;
        RECT 12.750 43.050 48.630 43.530 ;
        RECT 26.160 42.650 26.480 42.910 ;
        RECT 31.220 42.850 31.540 42.910 ;
        RECT 33.535 42.850 33.825 42.895 ;
        RECT 36.280 42.850 36.600 42.910 ;
        RECT 31.220 42.710 33.825 42.850 ;
        RECT 31.220 42.650 31.540 42.710 ;
        RECT 33.535 42.665 33.825 42.710 ;
        RECT 34.530 42.710 39.730 42.850 ;
        RECT 14.700 42.510 14.990 42.555 ;
        RECT 16.800 42.510 17.090 42.555 ;
        RECT 18.370 42.510 18.660 42.555 ;
        RECT 34.530 42.510 34.670 42.710 ;
        RECT 36.280 42.650 36.600 42.710 ;
        RECT 14.700 42.370 18.660 42.510 ;
        RECT 14.700 42.325 14.990 42.370 ;
        RECT 16.800 42.325 17.090 42.370 ;
        RECT 18.370 42.325 18.660 42.370 ;
        RECT 29.470 42.370 34.670 42.510 ;
        RECT 34.940 42.510 35.230 42.555 ;
        RECT 37.040 42.510 37.330 42.555 ;
        RECT 38.610 42.510 38.900 42.555 ;
        RECT 34.940 42.370 38.900 42.510 ;
        RECT 29.470 42.215 29.610 42.370 ;
        RECT 34.940 42.325 35.230 42.370 ;
        RECT 37.040 42.325 37.330 42.370 ;
        RECT 38.610 42.325 38.900 42.370 ;
        RECT 15.095 42.170 15.385 42.215 ;
        RECT 16.285 42.170 16.575 42.215 ;
        RECT 18.805 42.170 19.095 42.215 ;
        RECT 15.095 42.030 19.095 42.170 ;
        RECT 15.095 41.985 15.385 42.030 ;
        RECT 16.285 41.985 16.575 42.030 ;
        RECT 18.805 41.985 19.095 42.030 ;
        RECT 29.395 41.985 29.685 42.215 ;
        RECT 34.440 41.970 34.760 42.230 ;
        RECT 35.335 42.170 35.625 42.215 ;
        RECT 36.525 42.170 36.815 42.215 ;
        RECT 39.045 42.170 39.335 42.215 ;
        RECT 35.335 42.030 39.335 42.170 ;
        RECT 35.335 41.985 35.625 42.030 ;
        RECT 36.525 41.985 36.815 42.030 ;
        RECT 39.045 41.985 39.335 42.030 ;
        RECT 14.215 41.830 14.505 41.875 ;
        RECT 23.860 41.830 24.180 41.890 ;
        RECT 14.215 41.690 24.180 41.830 ;
        RECT 14.215 41.645 14.505 41.690 ;
        RECT 23.860 41.630 24.180 41.690 ;
        RECT 24.335 41.645 24.625 41.875 ;
        RECT 28.015 41.830 28.305 41.875 ;
        RECT 30.300 41.830 30.620 41.890 ;
        RECT 28.015 41.690 30.620 41.830 ;
        RECT 28.015 41.645 28.305 41.690 ;
        RECT 15.550 41.490 15.840 41.535 ;
        RECT 16.040 41.490 16.360 41.550 ;
        RECT 24.410 41.490 24.550 41.645 ;
        RECT 30.300 41.630 30.620 41.690 ;
        RECT 30.760 41.630 31.080 41.890 ;
        RECT 31.680 41.830 32.000 41.890 ;
        RECT 33.520 41.830 33.840 41.890 ;
        RECT 31.680 41.690 33.840 41.830 ;
        RECT 31.680 41.630 32.000 41.690 ;
        RECT 33.520 41.630 33.840 41.690 ;
        RECT 33.980 41.830 34.300 41.890 ;
        RECT 34.900 41.830 35.220 41.890 ;
        RECT 33.980 41.690 35.220 41.830 ;
        RECT 33.980 41.630 34.300 41.690 ;
        RECT 34.900 41.630 35.220 41.690 ;
        RECT 35.790 41.830 36.080 41.875 ;
        RECT 37.200 41.830 37.520 41.890 ;
        RECT 35.790 41.690 37.520 41.830 ;
        RECT 39.590 41.830 39.730 42.710 ;
        RECT 41.340 42.650 41.660 42.910 ;
        RECT 44.100 42.650 44.420 42.910 ;
        RECT 42.275 41.830 42.565 41.875 ;
        RECT 39.590 41.690 42.565 41.830 ;
        RECT 35.790 41.645 36.080 41.690 ;
        RECT 37.200 41.630 37.520 41.690 ;
        RECT 42.275 41.645 42.565 41.690 ;
        RECT 43.180 41.630 43.500 41.890 ;
        RECT 44.560 41.630 44.880 41.890 ;
        RECT 46.860 41.630 47.180 41.890 ;
        RECT 15.550 41.350 16.360 41.490 ;
        RECT 15.550 41.305 15.840 41.350 ;
        RECT 16.040 41.290 16.360 41.350 ;
        RECT 21.190 41.350 24.550 41.490 ;
        RECT 28.475 41.490 28.765 41.535 ;
        RECT 36.280 41.490 36.600 41.550 ;
        RECT 28.475 41.350 36.600 41.490 ;
        RECT 21.190 41.210 21.330 41.350 ;
        RECT 28.475 41.305 28.765 41.350 ;
        RECT 36.280 41.290 36.600 41.350 ;
        RECT 21.100 40.950 21.420 41.210 ;
        RECT 21.560 40.950 21.880 41.210 ;
        RECT 30.300 41.150 30.620 41.210 ;
        RECT 32.615 41.150 32.905 41.195 ;
        RECT 30.300 41.010 32.905 41.150 ;
        RECT 30.300 40.950 30.620 41.010 ;
        RECT 32.615 40.965 32.905 41.010 ;
        RECT 45.480 40.950 45.800 41.210 ;
        RECT 45.940 40.950 46.260 41.210 ;
        RECT 12.750 40.330 48.630 40.810 ;
        RECT 13.740 40.130 14.060 40.190 ;
        RECT 14.675 40.130 14.965 40.175 ;
        RECT 13.740 39.990 14.965 40.130 ;
        RECT 13.740 39.930 14.060 39.990 ;
        RECT 14.675 39.945 14.965 39.990 ;
        RECT 16.040 39.930 16.360 40.190 ;
        RECT 17.895 40.130 18.185 40.175 ;
        RECT 21.560 40.130 21.880 40.190 ;
        RECT 17.895 39.990 21.880 40.130 ;
        RECT 17.895 39.945 18.185 39.990 ;
        RECT 21.560 39.930 21.880 39.990 ;
        RECT 23.860 40.130 24.180 40.190 ;
        RECT 26.160 40.130 26.480 40.190 ;
        RECT 23.860 39.990 26.480 40.130 ;
        RECT 23.860 39.930 24.180 39.990 ;
        RECT 26.160 39.930 26.480 39.990 ;
        RECT 27.080 40.130 27.400 40.190 ;
        RECT 30.760 40.130 31.080 40.190 ;
        RECT 43.640 40.130 43.960 40.190 ;
        RECT 27.080 39.990 31.080 40.130 ;
        RECT 27.080 39.930 27.400 39.990 ;
        RECT 30.760 39.930 31.080 39.990 ;
        RECT 37.290 39.990 43.960 40.130 ;
        RECT 35.820 39.590 36.140 39.850 ;
        RECT 15.595 39.450 15.885 39.495 ;
        RECT 21.100 39.450 21.420 39.510 ;
        RECT 15.595 39.310 21.420 39.450 ;
        RECT 15.595 39.265 15.885 39.310 ;
        RECT 21.100 39.250 21.420 39.310 ;
        RECT 30.315 39.450 30.605 39.495 ;
        RECT 30.760 39.450 31.080 39.510 ;
        RECT 37.290 39.495 37.430 39.990 ;
        RECT 43.640 39.930 43.960 39.990 ;
        RECT 45.940 39.930 46.260 40.190 ;
        RECT 39.055 39.790 39.345 39.835 ;
        RECT 40.420 39.790 40.740 39.850 ;
        RECT 39.055 39.650 40.740 39.790 ;
        RECT 39.055 39.605 39.345 39.650 ;
        RECT 40.420 39.590 40.740 39.650 ;
        RECT 40.880 39.790 41.200 39.850 ;
        RECT 46.030 39.790 46.170 39.930 ;
        RECT 40.880 39.650 46.170 39.790 ;
        RECT 40.880 39.590 41.200 39.650 ;
        RECT 30.315 39.310 31.080 39.450 ;
        RECT 30.315 39.265 30.605 39.310 ;
        RECT 30.760 39.250 31.080 39.310 ;
        RECT 37.215 39.265 37.505 39.495 ;
        RECT 39.960 39.250 40.280 39.510 ;
        RECT 42.350 39.495 42.490 39.650 ;
        RECT 41.355 39.265 41.645 39.495 ;
        RECT 42.275 39.265 42.565 39.495 ;
        RECT 18.355 38.925 18.645 39.155 ;
        RECT 19.275 39.110 19.565 39.155 ;
        RECT 19.720 39.110 20.040 39.170 ;
        RECT 19.275 38.970 20.040 39.110 ;
        RECT 19.275 38.925 19.565 38.970 ;
        RECT 16.500 38.770 16.820 38.830 ;
        RECT 18.430 38.770 18.570 38.925 ;
        RECT 19.720 38.910 20.040 38.970 ;
        RECT 33.995 39.110 34.285 39.155 ;
        RECT 34.440 39.110 34.760 39.170 ;
        RECT 33.995 38.970 34.760 39.110 ;
        RECT 33.995 38.925 34.285 38.970 ;
        RECT 34.440 38.910 34.760 38.970 ;
        RECT 36.755 39.110 37.045 39.155 ;
        RECT 40.050 39.110 40.190 39.250 ;
        RECT 36.755 38.970 40.190 39.110 ;
        RECT 41.430 39.110 41.570 39.265 ;
        RECT 43.640 39.250 43.960 39.510 ;
        RECT 45.020 39.250 45.340 39.510 ;
        RECT 45.955 39.450 46.245 39.495 ;
        RECT 46.400 39.450 46.720 39.510 ;
        RECT 45.955 39.310 46.720 39.450 ;
        RECT 45.955 39.265 46.245 39.310 ;
        RECT 46.400 39.250 46.720 39.310 ;
        RECT 42.735 39.110 43.025 39.155 ;
        RECT 41.430 38.970 43.025 39.110 ;
        RECT 36.755 38.925 37.045 38.970 ;
        RECT 42.735 38.925 43.025 38.970 ;
        RECT 36.280 38.770 36.600 38.830 ;
        RECT 40.880 38.770 41.200 38.830 ;
        RECT 16.500 38.630 36.600 38.770 ;
        RECT 16.500 38.570 16.820 38.630 ;
        RECT 36.280 38.570 36.600 38.630 ;
        RECT 37.290 38.630 41.200 38.770 ;
        RECT 30.775 38.430 31.065 38.475 ;
        RECT 31.220 38.430 31.540 38.490 ;
        RECT 37.290 38.475 37.430 38.630 ;
        RECT 40.880 38.570 41.200 38.630 ;
        RECT 30.775 38.290 31.540 38.430 ;
        RECT 30.775 38.245 31.065 38.290 ;
        RECT 31.220 38.230 31.540 38.290 ;
        RECT 37.215 38.245 37.505 38.475 ;
        RECT 38.120 38.230 38.440 38.490 ;
        RECT 12.750 37.610 48.630 38.090 ;
        RECT 27.080 37.410 27.400 37.470 ;
        RECT 18.430 37.270 27.400 37.410 ;
        RECT 16.500 36.530 16.820 36.790 ;
        RECT 17.435 36.730 17.725 36.775 ;
        RECT 18.430 36.730 18.570 37.270 ;
        RECT 27.080 37.210 27.400 37.270 ;
        RECT 33.075 37.410 33.365 37.455 ;
        RECT 33.520 37.410 33.840 37.470 ;
        RECT 33.075 37.270 33.840 37.410 ;
        RECT 33.075 37.225 33.365 37.270 ;
        RECT 33.520 37.210 33.840 37.270 ;
        RECT 43.195 37.410 43.485 37.455 ;
        RECT 45.020 37.410 45.340 37.470 ;
        RECT 43.195 37.270 45.340 37.410 ;
        RECT 43.195 37.225 43.485 37.270 ;
        RECT 45.020 37.210 45.340 37.270 ;
        RECT 18.840 37.070 19.130 37.115 ;
        RECT 20.940 37.070 21.230 37.115 ;
        RECT 22.510 37.070 22.800 37.115 ;
        RECT 18.840 36.930 22.800 37.070 ;
        RECT 18.840 36.885 19.130 36.930 ;
        RECT 20.940 36.885 21.230 36.930 ;
        RECT 22.510 36.885 22.800 36.930 ;
        RECT 25.255 36.885 25.545 37.115 ;
        RECT 26.660 37.070 26.950 37.115 ;
        RECT 28.760 37.070 29.050 37.115 ;
        RECT 30.330 37.070 30.620 37.115 ;
        RECT 26.660 36.930 30.620 37.070 ;
        RECT 26.660 36.885 26.950 36.930 ;
        RECT 28.760 36.885 29.050 36.930 ;
        RECT 30.330 36.885 30.620 36.930 ;
        RECT 17.435 36.590 18.570 36.730 ;
        RECT 19.235 36.730 19.525 36.775 ;
        RECT 20.425 36.730 20.715 36.775 ;
        RECT 22.945 36.730 23.235 36.775 ;
        RECT 19.235 36.590 23.235 36.730 ;
        RECT 17.435 36.545 17.725 36.590 ;
        RECT 19.235 36.545 19.525 36.590 ;
        RECT 20.425 36.545 20.715 36.590 ;
        RECT 22.945 36.545 23.235 36.590 ;
        RECT 18.355 36.390 18.645 36.435 ;
        RECT 21.100 36.390 21.420 36.450 ;
        RECT 23.860 36.390 24.180 36.450 ;
        RECT 18.355 36.250 24.180 36.390 ;
        RECT 25.330 36.390 25.470 36.885 ;
        RECT 34.900 36.870 35.220 37.130 ;
        RECT 41.800 37.070 42.120 37.130 ;
        RECT 46.400 37.070 46.720 37.130 ;
        RECT 39.590 36.930 46.720 37.070 ;
        RECT 26.160 36.530 26.480 36.790 ;
        RECT 39.590 36.775 39.730 36.930 ;
        RECT 41.800 36.870 42.120 36.930 ;
        RECT 46.400 36.870 46.720 36.930 ;
        RECT 27.055 36.730 27.345 36.775 ;
        RECT 28.245 36.730 28.535 36.775 ;
        RECT 30.765 36.730 31.055 36.775 ;
        RECT 27.055 36.590 31.055 36.730 ;
        RECT 27.055 36.545 27.345 36.590 ;
        RECT 28.245 36.545 28.535 36.590 ;
        RECT 30.765 36.545 31.055 36.590 ;
        RECT 39.515 36.545 39.805 36.775 ;
        RECT 39.975 36.730 40.265 36.775 ;
        RECT 42.720 36.730 43.040 36.790 ;
        RECT 39.975 36.590 43.040 36.730 ;
        RECT 39.975 36.545 40.265 36.590 ;
        RECT 42.720 36.530 43.040 36.590 ;
        RECT 34.440 36.390 34.760 36.450 ;
        RECT 25.330 36.250 35.590 36.390 ;
        RECT 18.355 36.205 18.645 36.250 ;
        RECT 21.100 36.190 21.420 36.250 ;
        RECT 23.860 36.190 24.180 36.250 ;
        RECT 34.440 36.190 34.760 36.250 ;
        RECT 35.450 36.110 35.590 36.250 ;
        RECT 39.055 36.205 39.345 36.435 ;
        RECT 40.435 36.205 40.725 36.435 ;
        RECT 40.880 36.390 41.200 36.450 ;
        RECT 41.355 36.390 41.645 36.435 ;
        RECT 40.880 36.250 41.645 36.390 ;
        RECT 19.720 36.095 20.040 36.110 ;
        RECT 19.690 36.050 20.040 36.095 ;
        RECT 27.510 36.050 27.800 36.095 ;
        RECT 33.980 36.050 34.300 36.110 ;
        RECT 19.285 35.910 27.310 36.050 ;
        RECT 19.690 35.865 20.040 35.910 ;
        RECT 19.720 35.850 20.040 35.865 ;
        RECT 14.200 35.510 14.520 35.770 ;
        RECT 16.055 35.710 16.345 35.755 ;
        RECT 18.800 35.710 19.120 35.770 ;
        RECT 16.055 35.570 19.120 35.710 ;
        RECT 27.170 35.710 27.310 35.910 ;
        RECT 27.510 35.910 34.300 36.050 ;
        RECT 27.510 35.865 27.800 35.910 ;
        RECT 33.980 35.850 34.300 35.910 ;
        RECT 35.360 36.050 35.680 36.110 ;
        RECT 36.755 36.050 37.045 36.095 ;
        RECT 35.360 35.910 37.045 36.050 ;
        RECT 39.130 36.050 39.270 36.205 ;
        RECT 40.510 36.050 40.650 36.205 ;
        RECT 40.880 36.190 41.200 36.250 ;
        RECT 41.355 36.205 41.645 36.250 ;
        RECT 42.275 36.390 42.565 36.435 ;
        RECT 43.640 36.390 43.960 36.450 ;
        RECT 42.275 36.250 43.960 36.390 ;
        RECT 42.275 36.205 42.565 36.250 ;
        RECT 43.640 36.190 43.960 36.250 ;
        RECT 44.100 36.190 44.420 36.450 ;
        RECT 45.480 36.190 45.800 36.450 ;
        RECT 45.940 36.390 46.260 36.450 ;
        RECT 46.415 36.390 46.705 36.435 ;
        RECT 45.940 36.250 46.705 36.390 ;
        RECT 45.940 36.190 46.260 36.250 ;
        RECT 46.415 36.205 46.705 36.250 ;
        RECT 41.815 36.050 42.105 36.095 ;
        RECT 39.130 35.910 39.730 36.050 ;
        RECT 40.510 35.910 42.105 36.050 ;
        RECT 35.360 35.850 35.680 35.910 ;
        RECT 36.755 35.865 37.045 35.910 ;
        RECT 33.520 35.710 33.840 35.770 ;
        RECT 34.455 35.710 34.745 35.755 ;
        RECT 27.170 35.570 34.745 35.710 ;
        RECT 16.055 35.525 16.345 35.570 ;
        RECT 18.800 35.510 19.120 35.570 ;
        RECT 33.520 35.510 33.840 35.570 ;
        RECT 34.455 35.525 34.745 35.570 ;
        RECT 38.135 35.710 38.425 35.755 ;
        RECT 39.040 35.710 39.360 35.770 ;
        RECT 38.135 35.570 39.360 35.710 ;
        RECT 39.590 35.710 39.730 35.910 ;
        RECT 41.815 35.865 42.105 35.910 ;
        RECT 44.190 35.710 44.330 36.190 ;
        RECT 39.590 35.570 44.330 35.710 ;
        RECT 38.135 35.525 38.425 35.570 ;
        RECT 39.040 35.510 39.360 35.570 ;
        RECT 12.750 34.890 48.630 35.370 ;
        RECT 33.980 34.490 34.300 34.750 ;
        RECT 36.280 34.690 36.600 34.750 ;
        RECT 40.895 34.690 41.185 34.735 ;
        RECT 36.280 34.550 41.185 34.690 ;
        RECT 36.280 34.490 36.600 34.550 ;
        RECT 40.895 34.505 41.185 34.550 ;
        RECT 45.955 34.505 46.245 34.735 ;
        RECT 14.200 34.350 14.520 34.410 ;
        RECT 19.780 34.350 20.070 34.395 ;
        RECT 14.200 34.210 20.070 34.350 ;
        RECT 14.200 34.150 14.520 34.210 ;
        RECT 19.780 34.165 20.070 34.210 ;
        RECT 24.780 34.150 25.100 34.410 ;
        RECT 46.030 34.350 46.170 34.505 ;
        RECT 44.650 34.210 46.170 34.350 ;
        RECT 44.650 34.070 44.790 34.210 ;
        RECT 21.100 33.810 21.420 34.070 ;
        RECT 39.040 33.810 39.360 34.070 ;
        RECT 39.960 33.810 40.280 34.070 ;
        RECT 44.560 33.810 44.880 34.070 ;
        RECT 45.495 34.010 45.785 34.055 ;
        RECT 45.940 34.010 46.260 34.070 ;
        RECT 45.495 33.870 46.260 34.010 ;
        RECT 45.495 33.825 45.785 33.870 ;
        RECT 45.940 33.810 46.260 33.870 ;
        RECT 46.860 33.810 47.180 34.070 ;
        RECT 16.525 33.670 16.815 33.715 ;
        RECT 19.045 33.670 19.335 33.715 ;
        RECT 20.235 33.670 20.525 33.715 ;
        RECT 16.525 33.530 20.525 33.670 ;
        RECT 16.525 33.485 16.815 33.530 ;
        RECT 19.045 33.485 19.335 33.530 ;
        RECT 20.235 33.485 20.525 33.530 ;
        RECT 31.220 33.670 31.540 33.730 ;
        RECT 36.755 33.670 37.045 33.715 ;
        RECT 31.220 33.530 37.045 33.670 ;
        RECT 31.220 33.470 31.540 33.530 ;
        RECT 36.755 33.485 37.045 33.530 ;
        RECT 16.960 33.330 17.250 33.375 ;
        RECT 18.530 33.330 18.820 33.375 ;
        RECT 20.630 33.330 20.920 33.375 ;
        RECT 16.960 33.190 20.920 33.330 ;
        RECT 16.960 33.145 17.250 33.190 ;
        RECT 18.530 33.145 18.820 33.190 ;
        RECT 20.630 33.145 20.920 33.190 ;
        RECT 14.200 32.790 14.520 33.050 ;
        RECT 30.760 32.990 31.080 33.050 ;
        RECT 31.235 32.990 31.525 33.035 ;
        RECT 30.760 32.850 31.525 32.990 ;
        RECT 30.760 32.790 31.080 32.850 ;
        RECT 31.235 32.805 31.525 32.850 ;
        RECT 35.820 32.990 36.140 33.050 ;
        RECT 39.055 32.990 39.345 33.035 ;
        RECT 35.820 32.850 39.345 32.990 ;
        RECT 35.820 32.790 36.140 32.850 ;
        RECT 39.055 32.805 39.345 32.850 ;
        RECT 42.260 32.990 42.580 33.050 ;
        RECT 45.495 32.990 45.785 33.035 ;
        RECT 42.260 32.850 45.785 32.990 ;
        RECT 42.260 32.790 42.580 32.850 ;
        RECT 45.495 32.805 45.785 32.850 ;
        RECT 12.750 32.170 48.630 32.650 ;
        RECT 18.800 31.770 19.120 32.030 ;
        RECT 27.080 31.770 27.400 32.030 ;
        RECT 27.540 31.970 27.860 32.030 ;
        RECT 29.395 31.970 29.685 32.015 ;
        RECT 27.540 31.830 29.685 31.970 ;
        RECT 27.540 31.770 27.860 31.830 ;
        RECT 29.395 31.785 29.685 31.830 ;
        RECT 38.120 31.770 38.440 32.030 ;
        RECT 45.480 31.970 45.800 32.030 ;
        RECT 46.415 31.970 46.705 32.015 ;
        RECT 45.480 31.830 46.705 31.970 ;
        RECT 45.480 31.770 45.800 31.830 ;
        RECT 46.415 31.785 46.705 31.830 ;
        RECT 28.475 31.630 28.765 31.675 ;
        RECT 31.680 31.630 32.000 31.690 ;
        RECT 35.820 31.630 36.140 31.690 ;
        RECT 28.475 31.490 32.000 31.630 ;
        RECT 28.475 31.445 28.765 31.490 ;
        RECT 14.200 31.290 14.520 31.350 ;
        RECT 15.595 31.290 15.885 31.335 ;
        RECT 28.550 31.290 28.690 31.445 ;
        RECT 31.680 31.430 32.000 31.490 ;
        RECT 34.530 31.490 36.140 31.630 ;
        RECT 14.200 31.150 15.885 31.290 ;
        RECT 14.200 31.090 14.520 31.150 ;
        RECT 15.595 31.105 15.885 31.150 ;
        RECT 27.170 31.150 28.690 31.290 ;
        RECT 28.935 31.290 29.225 31.335 ;
        RECT 34.530 31.290 34.670 31.490 ;
        RECT 35.820 31.430 36.140 31.490 ;
        RECT 44.100 31.430 44.420 31.690 ;
        RECT 28.935 31.150 34.670 31.290 ;
        RECT 22.020 30.750 22.340 31.010 ;
        RECT 27.170 30.995 27.310 31.150 ;
        RECT 28.935 31.105 29.225 31.150 ;
        RECT 34.900 31.090 35.220 31.350 ;
        RECT 44.190 31.290 44.330 31.430 ;
        RECT 37.750 31.150 44.330 31.290 ;
        RECT 26.175 30.765 26.465 30.995 ;
        RECT 27.095 30.765 27.385 30.995 ;
        RECT 26.250 30.610 26.390 30.765 ;
        RECT 27.540 30.750 27.860 31.010 ;
        RECT 29.855 30.950 30.145 30.995 ;
        RECT 30.300 30.950 30.620 31.010 ;
        RECT 29.855 30.810 30.620 30.950 ;
        RECT 29.855 30.765 30.145 30.810 ;
        RECT 30.300 30.750 30.620 30.810 ;
        RECT 31.220 30.750 31.540 31.010 ;
        RECT 37.750 30.995 37.890 31.150 ;
        RECT 37.675 30.765 37.965 30.995 ;
        RECT 38.595 30.950 38.885 30.995 ;
        RECT 40.435 30.950 40.725 30.995 ;
        RECT 40.880 30.950 41.200 31.010 ;
        RECT 41.430 30.995 41.570 31.150 ;
        RECT 38.595 30.810 41.200 30.950 ;
        RECT 38.595 30.765 38.885 30.810 ;
        RECT 40.435 30.765 40.725 30.810 ;
        RECT 40.880 30.750 41.200 30.810 ;
        RECT 41.355 30.765 41.645 30.995 ;
        RECT 41.800 30.750 42.120 31.010 ;
        RECT 43.195 30.765 43.485 30.995 ;
        RECT 31.695 30.610 31.985 30.655 ;
        RECT 26.250 30.470 31.985 30.610 ;
        RECT 31.695 30.425 31.985 30.470 ;
        RECT 39.975 30.610 40.265 30.655 ;
        RECT 42.260 30.610 42.580 30.670 ;
        RECT 43.270 30.610 43.410 30.765 ;
        RECT 44.100 30.750 44.420 31.010 ;
        RECT 44.560 30.950 44.880 31.010 ;
        RECT 45.495 30.950 45.785 30.995 ;
        RECT 44.560 30.810 45.785 30.950 ;
        RECT 44.560 30.750 44.880 30.810 ;
        RECT 45.495 30.765 45.785 30.810 ;
        RECT 45.020 30.610 45.340 30.670 ;
        RECT 39.975 30.470 42.580 30.610 ;
        RECT 39.975 30.425 40.265 30.470 ;
        RECT 42.260 30.410 42.580 30.470 ;
        RECT 42.810 30.470 45.340 30.610 ;
        RECT 19.260 30.070 19.580 30.330 ;
        RECT 36.755 30.270 37.045 30.315 ;
        RECT 37.660 30.270 37.980 30.330 ;
        RECT 36.755 30.130 37.980 30.270 ;
        RECT 36.755 30.085 37.045 30.130 ;
        RECT 37.660 30.070 37.980 30.130 ;
        RECT 40.420 30.270 40.740 30.330 ;
        RECT 42.810 30.315 42.950 30.470 ;
        RECT 45.020 30.410 45.340 30.470 ;
        RECT 40.895 30.270 41.185 30.315 ;
        RECT 40.420 30.130 41.185 30.270 ;
        RECT 40.420 30.070 40.740 30.130 ;
        RECT 40.895 30.085 41.185 30.130 ;
        RECT 42.735 30.085 43.025 30.315 ;
        RECT 12.750 29.450 48.630 29.930 ;
        RECT 13.740 29.250 14.060 29.310 ;
        RECT 14.675 29.250 14.965 29.295 ;
        RECT 13.740 29.110 14.965 29.250 ;
        RECT 13.740 29.050 14.060 29.110 ;
        RECT 14.675 29.065 14.965 29.110 ;
        RECT 18.355 29.250 18.645 29.295 ;
        RECT 19.260 29.250 19.580 29.310 ;
        RECT 18.355 29.110 19.580 29.250 ;
        RECT 18.355 29.065 18.645 29.110 ;
        RECT 19.260 29.050 19.580 29.110 ;
        RECT 27.540 29.250 27.860 29.310 ;
        RECT 34.440 29.250 34.760 29.310 ;
        RECT 27.540 29.110 34.760 29.250 ;
        RECT 27.540 29.050 27.860 29.110 ;
        RECT 34.440 29.050 34.760 29.110 ;
        RECT 44.100 29.250 44.420 29.310 ;
        RECT 46.415 29.250 46.705 29.295 ;
        RECT 44.100 29.110 46.705 29.250 ;
        RECT 44.100 29.050 44.420 29.110 ;
        RECT 46.415 29.065 46.705 29.110 ;
        RECT 21.990 28.910 22.280 28.955 ;
        RECT 25.700 28.910 26.020 28.970 ;
        RECT 27.080 28.910 27.400 28.970 ;
        RECT 42.260 28.910 42.580 28.970 ;
        RECT 21.990 28.770 27.400 28.910 ;
        RECT 21.990 28.725 22.280 28.770 ;
        RECT 25.700 28.710 26.020 28.770 ;
        RECT 27.080 28.710 27.400 28.770 ;
        RECT 40.050 28.770 42.580 28.910 ;
        RECT 14.200 28.570 14.520 28.630 ;
        RECT 15.595 28.570 15.885 28.615 ;
        RECT 14.200 28.430 15.885 28.570 ;
        RECT 14.200 28.370 14.520 28.430 ;
        RECT 15.595 28.385 15.885 28.430 ;
        RECT 29.855 28.570 30.145 28.615 ;
        RECT 32.155 28.570 32.445 28.615 ;
        RECT 29.855 28.430 32.445 28.570 ;
        RECT 29.855 28.385 30.145 28.430 ;
        RECT 32.155 28.385 32.445 28.430 ;
        RECT 38.120 28.570 38.440 28.630 ;
        RECT 40.050 28.615 40.190 28.770 ;
        RECT 42.260 28.710 42.580 28.770 ;
        RECT 39.515 28.570 39.805 28.615 ;
        RECT 38.120 28.430 39.805 28.570 ;
        RECT 38.120 28.370 38.440 28.430 ;
        RECT 39.515 28.385 39.805 28.430 ;
        RECT 39.975 28.385 40.265 28.615 ;
        RECT 40.420 28.370 40.740 28.630 ;
        RECT 43.195 28.570 43.485 28.615 ;
        RECT 43.640 28.570 43.960 28.630 ;
        RECT 43.195 28.430 43.960 28.570 ;
        RECT 43.195 28.385 43.485 28.430 ;
        RECT 43.640 28.370 43.960 28.430 ;
        RECT 44.100 28.370 44.420 28.630 ;
        RECT 45.495 28.570 45.785 28.615 ;
        RECT 45.940 28.570 46.260 28.630 ;
        RECT 45.495 28.430 46.260 28.570 ;
        RECT 45.495 28.385 45.785 28.430 ;
        RECT 45.940 28.370 46.260 28.430 ;
        RECT 18.815 28.230 19.105 28.275 ;
        RECT 19.260 28.230 19.580 28.290 ;
        RECT 18.815 28.090 19.580 28.230 ;
        RECT 18.815 28.045 19.105 28.090 ;
        RECT 19.260 28.030 19.580 28.090 ;
        RECT 19.720 28.030 20.040 28.290 ;
        RECT 20.655 28.045 20.945 28.275 ;
        RECT 21.535 28.230 21.825 28.275 ;
        RECT 22.725 28.230 23.015 28.275 ;
        RECT 25.245 28.230 25.535 28.275 ;
        RECT 21.535 28.090 25.535 28.230 ;
        RECT 21.535 28.045 21.825 28.090 ;
        RECT 22.725 28.045 23.015 28.090 ;
        RECT 25.245 28.045 25.535 28.090 ;
        RECT 30.315 28.045 30.605 28.275 ;
        RECT 31.235 28.230 31.525 28.275 ;
        RECT 33.520 28.230 33.840 28.290 ;
        RECT 31.235 28.090 33.840 28.230 ;
        RECT 31.235 28.045 31.525 28.090 ;
        RECT 14.200 27.890 14.520 27.950 ;
        RECT 20.730 27.890 20.870 28.045 ;
        RECT 14.200 27.750 20.870 27.890 ;
        RECT 21.140 27.890 21.430 27.935 ;
        RECT 23.240 27.890 23.530 27.935 ;
        RECT 24.810 27.890 25.100 27.935 ;
        RECT 21.140 27.750 25.100 27.890 ;
        RECT 14.200 27.690 14.520 27.750 ;
        RECT 21.140 27.705 21.430 27.750 ;
        RECT 23.240 27.705 23.530 27.750 ;
        RECT 24.810 27.705 25.100 27.750 ;
        RECT 27.080 27.890 27.400 27.950 ;
        RECT 28.015 27.890 28.305 27.935 ;
        RECT 27.080 27.750 28.305 27.890 ;
        RECT 30.390 27.890 30.530 28.045 ;
        RECT 33.520 28.030 33.840 28.090 ;
        RECT 33.980 28.230 34.300 28.290 ;
        RECT 34.915 28.230 35.205 28.275 ;
        RECT 33.980 28.090 35.205 28.230 ;
        RECT 33.980 28.030 34.300 28.090 ;
        RECT 34.915 28.045 35.205 28.090 ;
        RECT 40.895 28.230 41.185 28.275 ;
        RECT 44.560 28.230 44.880 28.290 ;
        RECT 40.895 28.090 44.880 28.230 ;
        RECT 40.895 28.045 41.185 28.090 ;
        RECT 44.560 28.030 44.880 28.090 ;
        RECT 35.820 27.890 36.140 27.950 ;
        RECT 41.815 27.890 42.105 27.935 ;
        RECT 30.390 27.750 42.105 27.890 ;
        RECT 27.080 27.690 27.400 27.750 ;
        RECT 28.015 27.705 28.305 27.750 ;
        RECT 35.820 27.690 36.140 27.750 ;
        RECT 41.815 27.705 42.105 27.750 ;
        RECT 16.500 27.350 16.820 27.610 ;
        RECT 12.750 26.730 48.630 27.210 ;
        RECT 21.115 26.530 21.405 26.575 ;
        RECT 22.020 26.530 22.340 26.590 ;
        RECT 21.115 26.390 22.340 26.530 ;
        RECT 21.115 26.345 21.405 26.390 ;
        RECT 22.020 26.330 22.340 26.390 ;
        RECT 35.835 26.530 36.125 26.575 ;
        RECT 36.740 26.530 37.060 26.590 ;
        RECT 35.835 26.390 37.060 26.530 ;
        RECT 35.835 26.345 36.125 26.390 ;
        RECT 36.740 26.330 37.060 26.390 ;
        RECT 42.720 26.530 43.040 26.590 ;
        RECT 43.655 26.530 43.945 26.575 ;
        RECT 42.720 26.390 43.945 26.530 ;
        RECT 42.720 26.330 43.040 26.390 ;
        RECT 43.655 26.345 43.945 26.390 ;
        RECT 14.700 26.190 14.990 26.235 ;
        RECT 16.800 26.190 17.090 26.235 ;
        RECT 18.370 26.190 18.660 26.235 ;
        RECT 14.700 26.050 18.660 26.190 ;
        RECT 14.700 26.005 14.990 26.050 ;
        RECT 16.800 26.005 17.090 26.050 ;
        RECT 18.370 26.005 18.660 26.050 ;
        RECT 26.660 26.190 26.950 26.235 ;
        RECT 28.760 26.190 29.050 26.235 ;
        RECT 30.330 26.190 30.620 26.235 ;
        RECT 26.660 26.050 30.620 26.190 ;
        RECT 26.660 26.005 26.950 26.050 ;
        RECT 28.760 26.005 29.050 26.050 ;
        RECT 30.330 26.005 30.620 26.050 ;
        RECT 35.360 25.990 35.680 26.250 ;
        RECT 14.200 25.650 14.520 25.910 ;
        RECT 15.095 25.850 15.385 25.895 ;
        RECT 16.285 25.850 16.575 25.895 ;
        RECT 18.805 25.850 19.095 25.895 ;
        RECT 15.095 25.710 19.095 25.850 ;
        RECT 15.095 25.665 15.385 25.710 ;
        RECT 16.285 25.665 16.575 25.710 ;
        RECT 18.805 25.665 19.095 25.710 ;
        RECT 27.055 25.850 27.345 25.895 ;
        RECT 28.245 25.850 28.535 25.895 ;
        RECT 30.765 25.850 31.055 25.895 ;
        RECT 27.055 25.710 31.055 25.850 ;
        RECT 27.055 25.665 27.345 25.710 ;
        RECT 28.245 25.665 28.535 25.710 ;
        RECT 30.765 25.665 31.055 25.710 ;
        RECT 33.535 25.850 33.825 25.895 ;
        RECT 34.440 25.850 34.760 25.910 ;
        RECT 33.535 25.710 34.760 25.850 ;
        RECT 33.535 25.665 33.825 25.710 ;
        RECT 34.440 25.650 34.760 25.710 ;
        RECT 42.260 25.850 42.580 25.910 ;
        RECT 42.260 25.710 46.170 25.850 ;
        RECT 42.260 25.650 42.580 25.710 ;
        RECT 14.290 25.510 14.430 25.650 ;
        RECT 21.100 25.510 21.420 25.570 ;
        RECT 26.175 25.510 26.465 25.555 ;
        RECT 14.290 25.370 26.465 25.510 ;
        RECT 21.100 25.310 21.420 25.370 ;
        RECT 26.175 25.325 26.465 25.370 ;
        RECT 27.510 25.325 27.800 25.555 ;
        RECT 15.550 25.170 15.840 25.215 ;
        RECT 16.500 25.170 16.820 25.230 ;
        RECT 15.550 25.030 16.820 25.170 ;
        RECT 15.550 24.985 15.840 25.030 ;
        RECT 16.500 24.970 16.820 25.030 ;
        RECT 26.250 24.830 26.390 25.325 ;
        RECT 27.080 25.170 27.400 25.230 ;
        RECT 27.630 25.170 27.770 25.325 ;
        RECT 39.960 25.310 40.280 25.570 ;
        RECT 42.720 25.510 43.040 25.570 ;
        RECT 44.575 25.510 44.865 25.555 ;
        RECT 42.720 25.370 44.865 25.510 ;
        RECT 42.720 25.310 43.040 25.370 ;
        RECT 44.575 25.325 44.865 25.370 ;
        RECT 45.020 25.310 45.340 25.570 ;
        RECT 45.480 25.310 45.800 25.570 ;
        RECT 46.030 25.555 46.170 25.710 ;
        RECT 45.955 25.325 46.245 25.555 ;
        RECT 27.080 25.030 27.770 25.170 ;
        RECT 27.080 24.970 27.400 25.030 ;
        RECT 31.220 24.830 31.540 24.890 ;
        RECT 26.250 24.690 31.540 24.830 ;
        RECT 31.220 24.630 31.540 24.690 ;
        RECT 33.075 24.830 33.365 24.875 ;
        RECT 33.980 24.830 34.300 24.890 ;
        RECT 33.075 24.690 34.300 24.830 ;
        RECT 33.075 24.645 33.365 24.690 ;
        RECT 33.980 24.630 34.300 24.690 ;
        RECT 40.880 24.830 41.200 24.890 ;
        RECT 43.195 24.830 43.485 24.875 ;
        RECT 40.880 24.690 43.485 24.830 ;
        RECT 40.880 24.630 41.200 24.690 ;
        RECT 43.195 24.645 43.485 24.690 ;
        RECT 12.750 24.010 48.630 24.490 ;
        RECT 40.880 23.610 41.200 23.870 ;
        RECT 44.560 23.610 44.880 23.870 ;
        RECT 35.820 23.470 36.140 23.530 ;
        RECT 30.850 23.330 36.140 23.470 ;
        RECT 15.595 23.130 15.885 23.175 ;
        RECT 22.020 23.130 22.340 23.190 ;
        RECT 15.595 22.990 22.340 23.130 ;
        RECT 15.595 22.945 15.885 22.990 ;
        RECT 22.020 22.930 22.340 22.990 ;
        RECT 24.795 23.130 25.085 23.175 ;
        RECT 27.095 23.130 27.385 23.175 ;
        RECT 24.795 22.990 27.385 23.130 ;
        RECT 24.795 22.945 25.085 22.990 ;
        RECT 27.095 22.945 27.385 22.990 ;
        RECT 14.200 22.790 14.520 22.850 ;
        RECT 16.975 22.790 17.265 22.835 ;
        RECT 14.200 22.650 17.265 22.790 ;
        RECT 14.200 22.590 14.520 22.650 ;
        RECT 16.975 22.605 17.265 22.650 ;
        RECT 21.560 22.590 21.880 22.850 ;
        RECT 25.700 22.590 26.020 22.850 ;
        RECT 26.635 22.790 26.925 22.835 ;
        RECT 30.850 22.790 30.990 23.330 ;
        RECT 35.820 23.270 36.140 23.330 ;
        RECT 45.020 23.470 45.340 23.530 ;
        RECT 46.875 23.470 47.165 23.515 ;
        RECT 45.020 23.330 47.165 23.470 ;
        RECT 45.020 23.270 45.340 23.330 ;
        RECT 46.875 23.285 47.165 23.330 ;
        RECT 31.220 22.930 31.540 23.190 ;
        RECT 32.570 23.130 32.860 23.175 ;
        RECT 36.740 23.130 37.060 23.190 ;
        RECT 32.570 22.990 36.510 23.130 ;
        RECT 32.570 22.945 32.860 22.990 ;
        RECT 26.635 22.650 30.990 22.790 ;
        RECT 32.115 22.790 32.405 22.835 ;
        RECT 33.305 22.790 33.595 22.835 ;
        RECT 35.825 22.790 36.115 22.835 ;
        RECT 32.115 22.650 36.115 22.790 ;
        RECT 26.635 22.605 26.925 22.650 ;
        RECT 32.115 22.605 32.405 22.650 ;
        RECT 33.305 22.605 33.595 22.650 ;
        RECT 35.825 22.605 36.115 22.650 ;
        RECT 13.740 22.450 14.060 22.510 ;
        RECT 14.675 22.450 14.965 22.495 ;
        RECT 13.740 22.310 14.965 22.450 ;
        RECT 13.740 22.250 14.060 22.310 ;
        RECT 14.675 22.265 14.965 22.310 ;
        RECT 19.260 22.450 19.580 22.510 ;
        RECT 31.720 22.450 32.010 22.495 ;
        RECT 33.820 22.450 34.110 22.495 ;
        RECT 35.390 22.450 35.680 22.495 ;
        RECT 19.260 22.310 31.450 22.450 ;
        RECT 19.260 22.250 19.580 22.310 ;
        RECT 18.800 22.110 19.120 22.170 ;
        RECT 20.195 22.110 20.485 22.155 ;
        RECT 18.800 21.970 20.485 22.110 ;
        RECT 18.800 21.910 19.120 21.970 ;
        RECT 20.195 21.925 20.485 21.970 ;
        RECT 28.935 22.110 29.225 22.155 ;
        RECT 30.300 22.110 30.620 22.170 ;
        RECT 28.935 21.970 30.620 22.110 ;
        RECT 31.310 22.110 31.450 22.310 ;
        RECT 31.720 22.310 35.680 22.450 ;
        RECT 36.370 22.450 36.510 22.990 ;
        RECT 36.740 22.990 42.030 23.130 ;
        RECT 36.740 22.930 37.060 22.990 ;
        RECT 37.660 22.790 37.980 22.850 ;
        RECT 41.890 22.835 42.030 22.990 ;
        RECT 43.180 22.930 43.500 23.190 ;
        RECT 44.560 23.130 44.880 23.190 ;
        RECT 45.495 23.130 45.785 23.175 ;
        RECT 44.560 22.990 45.785 23.130 ;
        RECT 44.560 22.930 44.880 22.990 ;
        RECT 45.495 22.945 45.785 22.990 ;
        RECT 41.355 22.790 41.645 22.835 ;
        RECT 37.660 22.650 41.645 22.790 ;
        RECT 37.660 22.590 37.980 22.650 ;
        RECT 41.355 22.605 41.645 22.650 ;
        RECT 41.815 22.605 42.105 22.835 ;
        RECT 42.720 22.790 43.040 22.850 ;
        RECT 45.940 22.790 46.260 22.850 ;
        RECT 42.720 22.650 46.260 22.790 ;
        RECT 42.720 22.590 43.040 22.650 ;
        RECT 45.940 22.590 46.260 22.650 ;
        RECT 39.055 22.450 39.345 22.495 ;
        RECT 36.370 22.310 39.345 22.450 ;
        RECT 31.720 22.265 32.010 22.310 ;
        RECT 33.820 22.265 34.110 22.310 ;
        RECT 35.390 22.265 35.680 22.310 ;
        RECT 39.055 22.265 39.345 22.310 ;
        RECT 44.115 22.450 44.405 22.495 ;
        RECT 46.860 22.450 47.180 22.510 ;
        RECT 44.115 22.310 47.180 22.450 ;
        RECT 44.115 22.265 44.405 22.310 ;
        RECT 46.860 22.250 47.180 22.310 ;
        RECT 37.660 22.110 37.980 22.170 ;
        RECT 31.310 21.970 37.980 22.110 ;
        RECT 28.935 21.925 29.225 21.970 ;
        RECT 30.300 21.910 30.620 21.970 ;
        RECT 37.660 21.910 37.980 21.970 ;
        RECT 38.135 22.110 38.425 22.155 ;
        RECT 39.960 22.110 40.280 22.170 ;
        RECT 38.135 21.970 40.280 22.110 ;
        RECT 38.135 21.925 38.425 21.970 ;
        RECT 39.960 21.910 40.280 21.970 ;
        RECT 43.640 22.110 43.960 22.170 ;
        RECT 45.495 22.110 45.785 22.155 ;
        RECT 43.640 21.970 45.785 22.110 ;
        RECT 43.640 21.910 43.960 21.970 ;
        RECT 45.495 21.925 45.785 21.970 ;
        RECT 12.750 21.290 48.630 21.770 ;
        RECT 14.200 20.890 14.520 21.150 ;
        RECT 31.220 21.090 31.540 21.150 ;
        RECT 32.615 21.090 32.905 21.135 ;
        RECT 31.220 20.950 32.905 21.090 ;
        RECT 31.220 20.890 31.540 20.950 ;
        RECT 32.615 20.905 32.905 20.950 ;
        RECT 40.435 21.090 40.725 21.135 ;
        RECT 42.720 21.090 43.040 21.150 ;
        RECT 40.435 20.950 43.040 21.090 ;
        RECT 40.435 20.905 40.725 20.950 ;
        RECT 42.720 20.890 43.040 20.950 ;
        RECT 43.655 21.090 43.945 21.135 ;
        RECT 44.100 21.090 44.420 21.150 ;
        RECT 43.655 20.950 44.420 21.090 ;
        RECT 43.655 20.905 43.945 20.950 ;
        RECT 44.100 20.890 44.420 20.950 ;
        RECT 16.960 20.750 17.250 20.795 ;
        RECT 18.530 20.750 18.820 20.795 ;
        RECT 20.630 20.750 20.920 20.795 ;
        RECT 16.960 20.610 20.920 20.750 ;
        RECT 16.960 20.565 17.250 20.610 ;
        RECT 18.530 20.565 18.820 20.610 ;
        RECT 20.630 20.565 20.920 20.610 ;
        RECT 37.675 20.750 37.965 20.795 ;
        RECT 43.180 20.750 43.500 20.810 ;
        RECT 37.675 20.610 43.500 20.750 ;
        RECT 37.675 20.565 37.965 20.610 ;
        RECT 43.180 20.550 43.500 20.610 ;
        RECT 16.525 20.410 16.815 20.455 ;
        RECT 19.045 20.410 19.335 20.455 ;
        RECT 20.235 20.410 20.525 20.455 ;
        RECT 16.525 20.270 20.525 20.410 ;
        RECT 16.525 20.225 16.815 20.270 ;
        RECT 19.045 20.225 19.335 20.270 ;
        RECT 20.235 20.225 20.525 20.270 ;
        RECT 21.100 20.210 21.420 20.470 ;
        RECT 46.400 20.410 46.720 20.470 ;
        RECT 36.830 20.270 46.720 20.410 ;
        RECT 26.175 20.070 26.465 20.115 ;
        RECT 30.760 20.070 31.080 20.130 ;
        RECT 36.830 20.115 36.970 20.270 ;
        RECT 46.400 20.210 46.720 20.270 ;
        RECT 26.175 19.930 31.080 20.070 ;
        RECT 26.175 19.885 26.465 19.930 ;
        RECT 30.760 19.870 31.080 19.930 ;
        RECT 36.755 19.885 37.045 20.115 ;
        RECT 38.120 19.870 38.440 20.130 ;
        RECT 39.500 19.870 39.820 20.130 ;
        RECT 40.880 19.870 41.200 20.130 ;
        RECT 42.275 19.885 42.565 20.115 ;
        RECT 43.195 20.070 43.485 20.115 ;
        RECT 43.640 20.070 43.960 20.130 ;
        RECT 43.195 19.930 43.960 20.070 ;
        RECT 43.195 19.885 43.485 19.930 ;
        RECT 16.960 19.730 17.280 19.790 ;
        RECT 19.780 19.730 20.070 19.775 ;
        RECT 42.350 19.730 42.490 19.885 ;
        RECT 43.640 19.870 43.960 19.930 ;
        RECT 44.560 19.870 44.880 20.130 ;
        RECT 45.940 19.870 46.260 20.130 ;
        RECT 46.860 19.870 47.180 20.130 ;
        RECT 44.650 19.730 44.790 19.870 ;
        RECT 16.960 19.590 20.070 19.730 ;
        RECT 16.960 19.530 17.280 19.590 ;
        RECT 19.780 19.545 20.070 19.590 ;
        RECT 39.130 19.590 44.790 19.730 ;
        RECT 39.130 19.435 39.270 19.590 ;
        RECT 39.055 19.205 39.345 19.435 ;
        RECT 41.815 19.390 42.105 19.435 ;
        RECT 42.260 19.390 42.580 19.450 ;
        RECT 41.815 19.250 42.580 19.390 ;
        RECT 41.815 19.205 42.105 19.250 ;
        RECT 42.260 19.190 42.580 19.250 ;
        RECT 42.720 19.190 43.040 19.450 ;
        RECT 12.750 18.570 48.630 19.050 ;
        RECT 16.960 18.170 17.280 18.430 ;
        RECT 18.800 18.170 19.120 18.430 ;
        RECT 19.260 18.170 19.580 18.430 ;
        RECT 21.560 18.370 21.880 18.430 ;
        RECT 23.860 18.370 24.180 18.430 ;
        RECT 26.175 18.370 26.465 18.415 ;
        RECT 21.560 18.230 26.465 18.370 ;
        RECT 21.560 18.170 21.880 18.230 ;
        RECT 23.860 18.170 24.180 18.230 ;
        RECT 26.175 18.185 26.465 18.230 ;
        RECT 30.300 18.170 30.620 18.430 ;
        RECT 35.820 18.170 36.140 18.430 ;
        RECT 45.480 18.370 45.800 18.430 ;
        RECT 45.955 18.370 46.245 18.415 ;
        RECT 45.480 18.230 46.245 18.370 ;
        RECT 45.480 18.170 45.800 18.230 ;
        RECT 45.955 18.185 46.245 18.230 ;
        RECT 14.200 17.690 14.520 17.750 ;
        RECT 15.595 17.690 15.885 17.735 ;
        RECT 14.200 17.550 15.885 17.690 ;
        RECT 30.390 17.690 30.530 18.170 ;
        RECT 31.220 18.030 31.540 18.090 ;
        RECT 31.220 17.890 33.290 18.030 ;
        RECT 31.220 17.830 31.540 17.890 ;
        RECT 33.150 17.735 33.290 17.890 ;
        RECT 31.740 17.690 32.030 17.735 ;
        RECT 30.390 17.550 32.030 17.690 ;
        RECT 14.200 17.490 14.520 17.550 ;
        RECT 15.595 17.505 15.885 17.550 ;
        RECT 31.740 17.505 32.030 17.550 ;
        RECT 33.075 17.505 33.365 17.735 ;
        RECT 35.375 17.690 35.665 17.735 ;
        RECT 39.055 17.690 39.345 17.735 ;
        RECT 35.375 17.550 39.345 17.690 ;
        RECT 35.375 17.505 35.665 17.550 ;
        RECT 39.055 17.505 39.345 17.550 ;
        RECT 42.720 17.690 43.040 17.750 ;
        RECT 45.035 17.690 45.325 17.735 ;
        RECT 42.720 17.550 45.325 17.690 ;
        RECT 42.720 17.490 43.040 17.550 ;
        RECT 45.035 17.505 45.325 17.550 ;
        RECT 20.195 17.350 20.485 17.395 ;
        RECT 25.700 17.350 26.020 17.410 ;
        RECT 20.195 17.210 26.020 17.350 ;
        RECT 20.195 17.165 20.485 17.210 ;
        RECT 25.700 17.150 26.020 17.210 ;
        RECT 28.485 17.350 28.775 17.395 ;
        RECT 31.005 17.350 31.295 17.395 ;
        RECT 32.195 17.350 32.485 17.395 ;
        RECT 28.485 17.210 32.485 17.350 ;
        RECT 28.485 17.165 28.775 17.210 ;
        RECT 31.005 17.165 31.295 17.210 ;
        RECT 32.195 17.165 32.485 17.210 ;
        RECT 36.740 17.150 37.060 17.410 ;
        RECT 37.200 17.350 37.520 17.410 ;
        RECT 41.815 17.350 42.105 17.395 ;
        RECT 37.200 17.210 42.105 17.350 ;
        RECT 37.200 17.150 37.520 17.210 ;
        RECT 41.815 17.165 42.105 17.210 ;
        RECT 42.260 17.350 42.580 17.410 ;
        RECT 43.655 17.350 43.945 17.395 ;
        RECT 42.260 17.210 43.945 17.350 ;
        RECT 42.260 17.150 42.580 17.210 ;
        RECT 43.655 17.165 43.945 17.210 ;
        RECT 44.115 17.350 44.405 17.395 ;
        RECT 46.860 17.350 47.180 17.410 ;
        RECT 44.115 17.210 47.180 17.350 ;
        RECT 44.115 17.165 44.405 17.210 ;
        RECT 46.860 17.150 47.180 17.210 ;
        RECT 11.440 17.010 11.760 17.070 ;
        RECT 14.675 17.010 14.965 17.055 ;
        RECT 11.440 16.870 14.965 17.010 ;
        RECT 11.440 16.810 11.760 16.870 ;
        RECT 14.675 16.825 14.965 16.870 ;
        RECT 28.920 17.010 29.210 17.055 ;
        RECT 30.490 17.010 30.780 17.055 ;
        RECT 32.590 17.010 32.880 17.055 ;
        RECT 28.920 16.870 32.880 17.010 ;
        RECT 28.920 16.825 29.210 16.870 ;
        RECT 30.490 16.825 30.780 16.870 ;
        RECT 32.590 16.825 32.880 16.870 ;
        RECT 31.220 16.670 31.540 16.730 ;
        RECT 33.535 16.670 33.825 16.715 ;
        RECT 31.220 16.530 33.825 16.670 ;
        RECT 31.220 16.470 31.540 16.530 ;
        RECT 33.535 16.485 33.825 16.530 ;
        RECT 12.750 15.850 48.630 16.330 ;
        RECT 33.980 15.650 34.300 15.710 ;
        RECT 28.090 15.510 34.300 15.650 ;
        RECT 23.860 14.430 24.180 14.690 ;
        RECT 28.090 14.675 28.230 15.510 ;
        RECT 33.980 15.450 34.300 15.510 ;
        RECT 41.815 15.650 42.105 15.695 ;
        RECT 43.640 15.650 43.960 15.710 ;
        RECT 41.815 15.510 43.960 15.650 ;
        RECT 41.815 15.465 42.105 15.510 ;
        RECT 43.640 15.450 43.960 15.510 ;
        RECT 45.940 15.650 46.260 15.710 ;
        RECT 46.415 15.650 46.705 15.695 ;
        RECT 45.940 15.510 46.705 15.650 ;
        RECT 45.940 15.450 46.260 15.510 ;
        RECT 46.415 15.465 46.705 15.510 ;
        RECT 28.960 15.310 29.250 15.355 ;
        RECT 31.060 15.310 31.350 15.355 ;
        RECT 32.630 15.310 32.920 15.355 ;
        RECT 28.960 15.170 32.920 15.310 ;
        RECT 28.960 15.125 29.250 15.170 ;
        RECT 31.060 15.125 31.350 15.170 ;
        RECT 32.630 15.125 32.920 15.170 ;
        RECT 35.375 15.310 35.665 15.355 ;
        RECT 37.200 15.310 37.520 15.370 ;
        RECT 35.375 15.170 37.520 15.310 ;
        RECT 35.375 15.125 35.665 15.170 ;
        RECT 37.200 15.110 37.520 15.170 ;
        RECT 43.180 15.310 43.500 15.370 ;
        RECT 45.495 15.310 45.785 15.355 ;
        RECT 43.180 15.170 45.785 15.310 ;
        RECT 43.180 15.110 43.500 15.170 ;
        RECT 45.495 15.125 45.785 15.170 ;
        RECT 29.355 14.970 29.645 15.015 ;
        RECT 30.545 14.970 30.835 15.015 ;
        RECT 33.065 14.970 33.355 15.015 ;
        RECT 29.355 14.830 33.355 14.970 ;
        RECT 29.355 14.785 29.645 14.830 ;
        RECT 30.545 14.785 30.835 14.830 ;
        RECT 33.065 14.785 33.355 14.830 ;
        RECT 42.260 14.970 42.580 15.030 ;
        RECT 44.115 14.970 44.405 15.015 ;
        RECT 42.260 14.830 44.405 14.970 ;
        RECT 42.260 14.770 42.580 14.830 ;
        RECT 44.115 14.785 44.405 14.830 ;
        RECT 28.015 14.445 28.305 14.675 ;
        RECT 28.475 14.630 28.765 14.675 ;
        RECT 28.920 14.630 29.240 14.690 ;
        RECT 28.475 14.490 29.240 14.630 ;
        RECT 28.475 14.445 28.765 14.490 ;
        RECT 28.920 14.430 29.240 14.490 ;
        RECT 37.200 14.430 37.520 14.690 ;
        RECT 39.960 14.430 40.280 14.690 ;
        RECT 42.720 14.430 43.040 14.690 ;
        RECT 29.810 14.290 30.100 14.335 ;
        RECT 31.220 14.290 31.540 14.350 ;
        RECT 29.810 14.150 31.540 14.290 ;
        RECT 29.810 14.105 30.100 14.150 ;
        RECT 31.220 14.090 31.540 14.150 ;
        RECT 33.610 14.150 36.510 14.290 ;
        RECT 33.610 14.010 33.750 14.150 ;
        RECT 24.795 13.950 25.085 13.995 ;
        RECT 26.620 13.950 26.940 14.010 ;
        RECT 24.795 13.810 26.940 13.950 ;
        RECT 24.795 13.765 25.085 13.810 ;
        RECT 26.620 13.750 26.940 13.810 ;
        RECT 27.095 13.950 27.385 13.995 ;
        RECT 29.380 13.950 29.700 14.010 ;
        RECT 27.095 13.810 29.700 13.950 ;
        RECT 27.095 13.765 27.385 13.810 ;
        RECT 29.380 13.750 29.700 13.810 ;
        RECT 33.520 13.750 33.840 14.010 ;
        RECT 36.370 13.995 36.510 14.150 ;
        RECT 36.295 13.765 36.585 13.995 ;
        RECT 39.500 13.950 39.820 14.010 ;
        RECT 40.895 13.950 41.185 13.995 ;
        RECT 39.500 13.810 41.185 13.950 ;
        RECT 39.500 13.750 39.820 13.810 ;
        RECT 40.895 13.765 41.185 13.810 ;
        RECT 12.750 13.130 48.630 13.610 ;
      LAYER met2 ;
        RECT 76.400 212.010 76.680 216.010 ;
        RECT 36.280 204.445 37.820 204.815 ;
        RECT 76.470 204.280 76.610 212.010 ;
        RECT 76.410 203.960 76.670 204.280 ;
        RECT 77.790 203.280 78.050 203.600 ;
        RECT 32.980 201.725 34.520 202.095 ;
        RECT 36.280 199.005 37.820 199.375 ;
        RECT 12.460 196.625 12.740 196.995 ;
        RECT 12.530 139.000 12.670 196.625 ;
        RECT 32.980 196.285 34.520 196.655 ;
        RECT 36.280 193.565 37.820 193.935 ;
        RECT 58.930 192.400 59.190 192.720 ;
        RECT 71.350 192.400 71.610 192.720 ;
        RECT 72.270 192.400 72.530 192.720 ;
        RECT 32.980 190.845 34.520 191.215 ;
        RECT 36.280 188.125 37.820 188.495 ;
        RECT 58.990 187.960 59.130 192.400 ;
        RECT 70.890 192.060 71.150 192.380 ;
        RECT 66.290 191.720 66.550 192.040 ;
        RECT 58.930 187.640 59.190 187.960 ;
        RECT 66.350 187.280 66.490 191.720 ;
        RECT 67.210 191.380 67.470 191.700 ;
        RECT 66.750 188.660 67.010 188.980 ;
        RECT 66.810 187.280 66.950 188.660 ;
        RECT 64.450 186.960 64.710 187.280 ;
        RECT 66.290 186.960 66.550 187.280 ;
        RECT 66.750 186.960 67.010 187.280 ;
        RECT 37.770 186.620 38.030 186.940 ;
        RECT 38.230 186.620 38.490 186.940 ;
        RECT 41.910 186.620 42.170 186.940 ;
        RECT 35.010 186.280 35.270 186.600 ;
        RECT 32.980 185.405 34.520 185.775 ;
        RECT 29.950 184.580 30.210 184.900 ;
        RECT 30.410 184.580 30.670 184.900 ;
        RECT 35.070 184.640 35.210 186.280 ;
        RECT 28.110 184.240 28.370 184.560 ;
        RECT 21.670 183.900 21.930 184.220 ;
        RECT 21.730 181.160 21.870 183.900 ;
        RECT 24.430 183.560 24.690 183.880 ;
        RECT 24.490 182.520 24.630 183.560 ;
        RECT 24.890 183.220 25.150 183.540 ;
        RECT 24.950 182.520 25.090 183.220 ;
        RECT 28.170 182.600 28.310 184.240 ;
        RECT 24.430 182.200 24.690 182.520 ;
        RECT 24.890 182.200 25.150 182.520 ;
        RECT 27.710 182.460 28.310 182.600 ;
        RECT 21.670 180.840 21.930 181.160 ;
        RECT 16.150 176.080 16.410 176.400 ;
        RECT 16.210 175.235 16.350 176.080 ;
        RECT 21.730 176.060 21.870 180.840 ;
        RECT 24.430 179.100 24.690 179.120 ;
        RECT 24.950 179.100 25.090 182.200 ;
        RECT 27.710 181.500 27.850 182.460 ;
        RECT 30.010 181.840 30.150 184.580 ;
        RECT 29.950 181.520 30.210 181.840 ;
        RECT 25.810 181.180 26.070 181.500 ;
        RECT 27.650 181.180 27.910 181.500 ;
        RECT 25.870 179.460 26.010 181.180 ;
        RECT 25.810 179.140 26.070 179.460 ;
        RECT 24.430 178.960 25.090 179.100 ;
        RECT 24.430 178.800 24.690 178.960 ;
        RECT 23.970 178.690 24.230 178.780 ;
        RECT 23.570 178.550 24.230 178.690 ;
        RECT 22.590 177.780 22.850 178.100 ;
        RECT 22.650 176.740 22.790 177.780 ;
        RECT 22.590 176.420 22.850 176.740 ;
        RECT 21.670 175.740 21.930 176.060 ;
        RECT 16.140 174.865 16.420 175.235 ;
        RECT 21.730 173.340 21.870 175.740 ;
        RECT 21.670 173.020 21.930 173.340 ;
        RECT 22.590 172.680 22.850 173.000 ;
        RECT 22.650 171.640 22.790 172.680 ;
        RECT 23.570 171.640 23.710 178.550 ;
        RECT 23.970 178.460 24.230 178.550 ;
        RECT 23.970 173.020 24.230 173.340 ;
        RECT 24.030 171.640 24.170 173.020 ;
        RECT 22.590 171.320 22.850 171.640 ;
        RECT 23.510 171.320 23.770 171.640 ;
        RECT 23.970 171.320 24.230 171.640 ;
        RECT 21.670 170.640 21.930 170.960 ;
        RECT 21.730 168.920 21.870 170.640 ;
        RECT 23.050 169.620 23.310 169.940 ;
        RECT 21.670 168.600 21.930 168.920 ;
        RECT 23.110 167.220 23.250 169.620 ;
        RECT 23.050 166.900 23.310 167.220 ;
        RECT 23.110 165.520 23.250 166.900 ;
        RECT 23.570 165.860 23.710 171.320 ;
        RECT 23.510 165.540 23.770 165.860 ;
        RECT 23.050 165.200 23.310 165.520 ;
        RECT 16.150 162.140 16.410 162.460 ;
        RECT 16.210 161.635 16.350 162.140 ;
        RECT 16.140 161.265 16.420 161.635 ;
        RECT 21.670 161.460 21.930 161.780 ;
        RECT 21.730 156.680 21.870 161.460 ;
        RECT 23.110 160.760 23.250 165.200 ;
        RECT 23.570 162.460 23.710 165.540 ;
        RECT 23.510 162.140 23.770 162.460 ;
        RECT 23.050 160.440 23.310 160.760 ;
        RECT 24.030 160.080 24.170 171.320 ;
        RECT 24.490 170.960 24.630 178.800 ;
        RECT 27.710 178.780 27.850 181.180 ;
        RECT 30.010 180.820 30.150 181.520 ;
        RECT 29.950 180.500 30.210 180.820 ;
        RECT 30.010 179.800 30.150 180.500 ;
        RECT 29.950 179.480 30.210 179.800 ;
        RECT 30.470 179.460 30.610 184.580 ;
        RECT 34.150 184.560 35.210 184.640 ;
        RECT 37.830 184.640 37.970 186.620 ;
        RECT 38.290 185.240 38.430 186.620 ;
        RECT 39.150 185.940 39.410 186.260 ;
        RECT 39.610 185.940 39.870 186.260 ;
        RECT 38.230 184.920 38.490 185.240 ;
        RECT 34.090 184.500 35.210 184.560 ;
        RECT 34.090 184.240 34.350 184.500 ;
        RECT 35.470 184.240 35.730 184.560 ;
        RECT 37.830 184.500 38.430 184.640 ;
        RECT 35.010 183.560 35.270 183.880 ;
        RECT 35.070 181.500 35.210 183.560 ;
        RECT 30.870 181.180 31.130 181.500 ;
        RECT 35.010 181.180 35.270 181.500 ;
        RECT 30.930 179.460 31.070 181.180 ;
        RECT 35.010 180.500 35.270 180.820 ;
        RECT 32.980 179.965 34.520 180.335 ;
        RECT 34.550 179.480 34.810 179.800 ;
        RECT 30.410 179.140 30.670 179.460 ;
        RECT 30.870 179.140 31.130 179.460 ;
        RECT 34.610 179.315 34.750 179.480 ;
        RECT 25.350 178.460 25.610 178.780 ;
        RECT 27.650 178.460 27.910 178.780 ;
        RECT 25.410 170.960 25.550 178.460 ;
        RECT 29.950 178.120 30.210 178.440 ;
        RECT 30.010 177.080 30.150 178.120 ;
        RECT 29.950 176.760 30.210 177.080 ;
        RECT 30.930 176.400 31.070 179.140 ;
        RECT 34.540 178.945 34.820 179.315 ;
        RECT 28.570 176.080 28.830 176.400 ;
        RECT 30.870 176.080 31.130 176.400 ;
        RECT 28.110 175.060 28.370 175.380 ;
        RECT 28.170 173.680 28.310 175.060 ;
        RECT 28.630 174.360 28.770 176.080 ;
        RECT 29.030 175.060 29.290 175.380 ;
        RECT 28.570 174.040 28.830 174.360 ;
        RECT 28.110 173.360 28.370 173.680 ;
        RECT 29.090 173.340 29.230 175.060 ;
        RECT 26.270 173.020 26.530 173.340 ;
        RECT 29.030 173.020 29.290 173.340 ;
        RECT 25.810 170.980 26.070 171.300 ;
        RECT 24.430 170.640 24.690 170.960 ;
        RECT 25.350 170.640 25.610 170.960 ;
        RECT 24.490 162.800 24.630 170.640 ;
        RECT 24.890 164.180 25.150 164.500 ;
        RECT 24.950 162.800 25.090 164.180 ;
        RECT 25.410 163.140 25.550 170.640 ;
        RECT 25.870 167.900 26.010 170.980 ;
        RECT 26.330 170.280 26.470 173.020 ;
        RECT 28.110 172.340 28.370 172.660 ;
        RECT 28.170 171.300 28.310 172.340 ;
        RECT 28.110 170.980 28.370 171.300 ;
        RECT 26.270 169.960 26.530 170.280 ;
        RECT 28.170 168.920 28.310 170.980 ;
        RECT 29.090 170.620 29.230 173.020 ;
        RECT 30.930 171.300 31.070 176.080 ;
        RECT 34.610 175.800 34.750 178.945 ;
        RECT 35.070 178.780 35.210 180.500 ;
        RECT 35.530 179.800 35.670 184.240 ;
        RECT 37.830 183.880 37.970 184.500 ;
        RECT 37.770 183.560 38.030 183.880 ;
        RECT 36.390 183.450 36.650 183.540 ;
        RECT 35.990 183.310 36.650 183.450 ;
        RECT 35.990 182.180 36.130 183.310 ;
        RECT 36.390 183.220 36.650 183.310 ;
        RECT 36.280 182.685 37.820 183.055 ;
        RECT 38.290 182.520 38.430 184.500 ;
        RECT 36.850 182.430 37.110 182.520 ;
        RECT 36.450 182.290 37.110 182.430 ;
        RECT 35.930 181.860 36.190 182.180 ;
        RECT 36.450 180.820 36.590 182.290 ;
        RECT 36.850 182.200 37.110 182.290 ;
        RECT 38.230 182.200 38.490 182.520 ;
        RECT 36.390 180.500 36.650 180.820 ;
        RECT 38.690 180.500 38.950 180.820 ;
        RECT 35.470 179.480 35.730 179.800 ;
        RECT 36.450 178.780 36.590 180.500 ;
        RECT 37.300 178.945 37.580 179.315 ;
        RECT 37.770 179.140 38.030 179.460 ;
        RECT 37.370 178.780 37.510 178.945 ;
        RECT 37.830 178.780 37.970 179.140 ;
        RECT 35.010 178.460 35.270 178.780 ;
        RECT 36.390 178.460 36.650 178.780 ;
        RECT 37.310 178.460 37.570 178.780 ;
        RECT 37.770 178.460 38.030 178.780 ;
        RECT 38.750 178.100 38.890 180.500 ;
        RECT 39.210 179.800 39.350 185.940 ;
        RECT 39.670 184.220 39.810 185.940 ;
        RECT 39.610 183.900 39.870 184.220 ;
        RECT 39.150 179.480 39.410 179.800 ;
        RECT 41.970 179.120 42.110 186.620 ;
        RECT 55.250 185.940 55.510 186.260 ;
        RECT 54.330 184.920 54.590 185.240 ;
        RECT 53.410 183.900 53.670 184.220 ;
        RECT 46.970 183.560 47.230 183.880 ;
        RECT 43.750 183.220 44.010 183.540 ;
        RECT 45.130 183.220 45.390 183.540 ;
        RECT 43.810 179.460 43.950 183.220 ;
        RECT 45.190 182.180 45.330 183.220 ;
        RECT 47.030 182.520 47.170 183.560 ;
        RECT 46.970 182.200 47.230 182.520 ;
        RECT 45.130 181.860 45.390 182.180 ;
        RECT 51.570 181.860 51.830 182.180 ;
        RECT 43.750 179.140 44.010 179.460 ;
        RECT 41.910 178.800 42.170 179.120 ;
        RECT 43.810 178.780 43.950 179.140 ;
        RECT 41.450 178.460 41.710 178.780 ;
        RECT 43.750 178.460 44.010 178.780 ;
        RECT 41.510 178.100 41.650 178.460 ;
        RECT 38.690 177.780 38.950 178.100 ;
        RECT 41.450 177.780 41.710 178.100 ;
        RECT 36.280 177.245 37.820 177.615 ;
        RECT 34.610 175.660 35.210 175.800 ;
        RECT 32.980 174.525 34.520 174.895 ;
        RECT 32.250 173.020 32.510 173.340 ;
        RECT 35.070 173.080 35.210 175.660 ;
        RECT 38.750 174.360 38.890 177.780 ;
        RECT 38.690 174.040 38.950 174.360 ;
        RECT 40.530 173.700 40.790 174.020 ;
        RECT 40.990 173.700 41.250 174.020 ;
        RECT 32.310 171.300 32.450 173.020 ;
        RECT 34.610 172.940 35.210 173.080 ;
        RECT 30.870 170.980 31.130 171.300 ;
        RECT 32.250 170.980 32.510 171.300 ;
        RECT 29.950 170.640 30.210 170.960 ;
        RECT 29.030 170.300 29.290 170.620 ;
        RECT 28.110 168.600 28.370 168.920 ;
        RECT 28.170 167.900 28.310 168.600 ;
        RECT 30.010 168.240 30.150 170.640 ;
        RECT 30.870 168.600 31.130 168.920 ;
        RECT 29.950 167.920 30.210 168.240 ;
        RECT 25.810 167.580 26.070 167.900 ;
        RECT 28.110 167.580 28.370 167.900 ;
        RECT 25.870 165.180 26.010 167.580 ;
        RECT 27.650 165.540 27.910 165.860 ;
        RECT 25.810 164.860 26.070 165.180 ;
        RECT 25.350 162.820 25.610 163.140 ;
        RECT 24.430 162.480 24.690 162.800 ;
        RECT 24.890 162.480 25.150 162.800 ;
        RECT 25.870 162.120 26.010 164.860 ;
        RECT 27.710 162.800 27.850 165.540 ;
        RECT 30.930 165.520 31.070 168.600 ;
        RECT 32.310 168.240 32.450 170.980 ;
        RECT 34.610 170.960 34.750 172.940 ;
        RECT 35.930 172.680 36.190 173.000 ;
        RECT 35.010 172.340 35.270 172.660 ;
        RECT 35.070 170.960 35.210 172.340 ;
        RECT 34.550 170.640 34.810 170.960 ;
        RECT 35.010 170.640 35.270 170.960 ;
        RECT 35.470 170.640 35.730 170.960 ;
        RECT 32.980 169.085 34.520 169.455 ;
        RECT 32.250 167.920 32.510 168.240 ;
        RECT 31.330 167.580 31.590 167.900 ;
        RECT 30.870 165.200 31.130 165.520 ;
        RECT 31.390 165.180 31.530 167.580 ;
        RECT 32.310 165.520 32.450 167.920 ;
        RECT 35.070 167.900 35.210 170.640 ;
        RECT 35.010 167.580 35.270 167.900 ;
        RECT 35.530 166.110 35.670 170.640 ;
        RECT 35.070 165.970 35.670 166.110 ;
        RECT 32.250 165.200 32.510 165.520 ;
        RECT 35.070 165.180 35.210 165.970 ;
        RECT 35.470 165.200 35.730 165.520 ;
        RECT 31.330 164.860 31.590 165.180 ;
        RECT 35.010 164.860 35.270 165.180 ;
        RECT 27.650 162.480 27.910 162.800 ;
        RECT 30.870 162.140 31.130 162.460 ;
        RECT 25.810 161.800 26.070 162.120 ;
        RECT 23.970 159.760 24.230 160.080 ;
        RECT 24.030 159.480 24.170 159.760 ;
        RECT 23.570 159.340 24.170 159.480 ;
        RECT 23.570 157.020 23.710 159.340 ;
        RECT 25.870 158.040 26.010 161.800 ;
        RECT 26.270 161.460 26.530 161.780 ;
        RECT 26.330 159.990 26.470 161.460 ;
        RECT 26.730 159.990 26.990 160.080 ;
        RECT 26.330 159.850 26.990 159.990 ;
        RECT 26.730 159.760 26.990 159.850 ;
        RECT 25.810 157.720 26.070 158.040 ;
        RECT 23.510 156.700 23.770 157.020 ;
        RECT 21.670 156.360 21.930 156.680 ;
        RECT 19.830 150.580 20.090 150.900 ;
        RECT 19.890 149.880 20.030 150.580 ;
        RECT 19.830 149.560 20.090 149.880 ;
        RECT 20.750 149.220 21.010 149.540 ;
        RECT 16.150 148.880 16.410 149.200 ;
        RECT 16.210 148.035 16.350 148.880 ;
        RECT 16.140 147.665 16.420 148.035 ;
        RECT 20.810 147.160 20.950 149.220 ;
        RECT 23.570 149.200 23.710 156.700 ;
        RECT 30.930 155.320 31.070 162.140 ;
        RECT 30.870 155.000 31.130 155.320 ;
        RECT 30.930 154.640 31.070 155.000 ;
        RECT 30.870 154.320 31.130 154.640 ;
        RECT 31.390 154.300 31.530 164.860 ;
        RECT 32.980 163.645 34.520 164.015 ;
        RECT 32.710 163.160 32.970 163.480 ;
        RECT 32.250 162.140 32.510 162.460 ;
        RECT 32.310 160.760 32.450 162.140 ;
        RECT 32.250 160.440 32.510 160.760 ;
        RECT 31.790 159.760 32.050 160.080 ;
        RECT 32.250 159.990 32.510 160.080 ;
        RECT 32.770 159.990 32.910 163.160 ;
        RECT 34.090 161.460 34.350 161.780 ;
        RECT 34.150 160.080 34.290 161.460 ;
        RECT 32.250 159.850 32.910 159.990 ;
        RECT 32.250 159.760 32.510 159.850 ;
        RECT 34.090 159.760 34.350 160.080 ;
        RECT 31.850 158.040 31.990 159.760 ;
        RECT 31.790 157.720 32.050 158.040 ;
        RECT 31.850 157.020 31.990 157.720 ;
        RECT 32.310 157.610 32.450 159.760 ;
        RECT 32.980 158.205 34.520 158.575 ;
        RECT 32.710 157.610 32.970 157.700 ;
        RECT 32.310 157.470 32.970 157.610 ;
        RECT 32.710 157.380 32.970 157.470 ;
        RECT 31.790 156.700 32.050 157.020 ;
        RECT 32.770 156.680 32.910 157.380 ;
        RECT 32.710 156.360 32.970 156.680 ;
        RECT 34.090 156.020 34.350 156.340 ;
        RECT 34.150 154.640 34.290 156.020 ;
        RECT 35.070 155.320 35.210 164.860 ;
        RECT 35.530 162.460 35.670 165.200 ;
        RECT 35.990 165.035 36.130 172.680 ;
        RECT 40.070 172.340 40.330 172.660 ;
        RECT 36.280 171.805 37.820 172.175 ;
        RECT 37.310 170.300 37.570 170.620 ;
        RECT 37.370 167.900 37.510 170.300 ;
        RECT 37.770 169.620 38.030 169.940 ;
        RECT 37.830 167.900 37.970 169.620 ;
        RECT 40.130 167.900 40.270 172.340 ;
        RECT 40.590 167.900 40.730 173.700 ;
        RECT 41.050 173.340 41.190 173.700 ;
        RECT 43.810 173.680 43.950 178.460 ;
        RECT 45.190 175.380 45.330 181.860 ;
        RECT 51.110 181.520 51.370 181.840 ;
        RECT 46.050 181.180 46.310 181.500 ;
        RECT 50.650 181.180 50.910 181.500 ;
        RECT 46.110 178.100 46.250 181.180 ;
        RECT 47.430 178.460 47.690 178.780 ;
        RECT 46.050 177.780 46.310 178.100 ;
        RECT 46.110 177.160 46.250 177.780 ;
        RECT 46.110 177.080 46.710 177.160 ;
        RECT 46.110 177.020 46.770 177.080 ;
        RECT 46.510 176.760 46.770 177.020 ;
        RECT 46.970 176.080 47.230 176.400 ;
        RECT 45.590 175.740 45.850 176.060 ;
        RECT 44.210 175.060 44.470 175.380 ;
        RECT 45.130 175.060 45.390 175.380 ;
        RECT 44.270 173.680 44.410 175.060 ;
        RECT 45.130 173.700 45.390 174.020 ;
        RECT 43.750 173.360 44.010 173.680 ;
        RECT 44.210 173.360 44.470 173.680 ;
        RECT 40.990 173.020 41.250 173.340 ;
        RECT 41.910 173.250 42.170 173.340 ;
        RECT 41.910 173.110 43.490 173.250 ;
        RECT 41.910 173.020 42.170 173.110 ;
        RECT 43.350 173.080 43.490 173.110 ;
        RECT 44.270 173.080 44.410 173.360 ;
        RECT 43.350 172.940 44.410 173.080 ;
        RECT 44.670 173.020 44.930 173.340 ;
        RECT 37.310 167.580 37.570 167.900 ;
        RECT 37.770 167.580 38.030 167.900 ;
        RECT 40.070 167.580 40.330 167.900 ;
        RECT 40.530 167.580 40.790 167.900 ;
        RECT 40.070 166.900 40.330 167.220 ;
        RECT 40.990 166.900 41.250 167.220 ;
        RECT 41.450 166.900 41.710 167.220 ;
        RECT 36.280 166.365 37.820 166.735 ;
        RECT 35.920 164.665 36.200 165.035 ;
        RECT 35.930 164.180 36.190 164.500 ;
        RECT 35.990 162.460 36.130 164.180 ;
        RECT 37.310 163.160 37.570 163.480 ;
        RECT 37.370 162.460 37.510 163.160 ;
        RECT 40.130 162.800 40.270 166.900 ;
        RECT 41.050 165.860 41.190 166.900 ;
        RECT 40.990 165.540 41.250 165.860 ;
        RECT 41.510 165.520 41.650 166.900 ;
        RECT 44.730 166.110 44.870 173.020 ;
        RECT 43.810 165.970 44.870 166.110 ;
        RECT 41.450 165.200 41.710 165.520 ;
        RECT 41.910 165.200 42.170 165.520 ;
        RECT 41.970 164.920 42.110 165.200 ;
        RECT 41.510 164.780 42.110 164.920 ;
        RECT 40.070 162.480 40.330 162.800 ;
        RECT 40.530 162.480 40.790 162.800 ;
        RECT 35.470 162.140 35.730 162.460 ;
        RECT 35.930 162.140 36.190 162.460 ;
        RECT 37.310 162.370 37.570 162.460 ;
        RECT 37.310 162.230 38.430 162.370 ;
        RECT 37.310 162.140 37.570 162.230 ;
        RECT 36.280 160.925 37.820 161.295 ;
        RECT 38.290 160.760 38.430 162.230 ;
        RECT 38.690 162.140 38.950 162.460 ;
        RECT 38.230 160.440 38.490 160.760 ;
        RECT 38.750 158.040 38.890 162.140 ;
        RECT 39.610 161.800 39.870 162.120 ;
        RECT 39.670 160.760 39.810 161.800 ;
        RECT 39.610 160.440 39.870 160.760 ;
        RECT 40.590 160.420 40.730 162.480 ;
        RECT 40.990 162.370 41.250 162.460 ;
        RECT 41.510 162.370 41.650 164.780 ;
        RECT 41.910 164.180 42.170 164.500 ;
        RECT 40.990 162.230 41.650 162.370 ;
        RECT 40.990 162.140 41.250 162.230 ;
        RECT 40.530 160.100 40.790 160.420 ;
        RECT 41.050 159.480 41.190 162.140 ;
        RECT 41.450 161.460 41.710 161.780 ;
        RECT 41.510 160.080 41.650 161.460 ;
        RECT 41.970 160.080 42.110 164.180 ;
        RECT 43.290 161.460 43.550 161.780 ;
        RECT 41.450 159.760 41.710 160.080 ;
        RECT 41.910 159.760 42.170 160.080 ;
        RECT 41.050 159.340 41.650 159.480 ;
        RECT 38.690 157.720 38.950 158.040 ;
        RECT 40.990 156.700 41.250 157.020 ;
        RECT 36.280 155.485 37.820 155.855 ;
        RECT 35.010 155.000 35.270 155.320 ;
        RECT 34.090 154.320 34.350 154.640 ;
        RECT 31.330 153.980 31.590 154.300 ;
        RECT 31.390 149.200 31.530 153.980 ;
        RECT 32.980 152.765 34.520 153.135 ;
        RECT 35.070 149.880 35.210 155.000 ;
        RECT 40.070 151.940 40.330 152.260 ;
        RECT 36.280 150.045 37.820 150.415 ;
        RECT 35.010 149.560 35.270 149.880 ;
        RECT 39.610 149.220 39.870 149.540 ;
        RECT 23.510 148.880 23.770 149.200 ;
        RECT 23.970 148.880 24.230 149.200 ;
        RECT 31.330 148.880 31.590 149.200 ;
        RECT 35.930 148.880 36.190 149.200 ;
        RECT 24.030 147.160 24.170 148.880 ;
        RECT 32.250 147.860 32.510 148.180 ;
        RECT 35.470 147.860 35.730 148.180 ;
        RECT 20.750 146.840 21.010 147.160 ;
        RECT 23.970 146.840 24.230 147.160 ;
        RECT 24.890 146.840 25.150 147.160 ;
        RECT 19.370 145.480 19.630 145.800 ;
        RECT 19.430 143.955 19.570 145.480 ;
        RECT 19.360 143.585 19.640 143.955 ;
        RECT 24.950 143.760 25.090 146.840 ;
        RECT 28.110 146.160 28.370 146.480 ;
        RECT 28.570 146.160 28.830 146.480 ;
        RECT 26.270 145.820 26.530 146.140 ;
        RECT 25.350 145.480 25.610 145.800 ;
        RECT 24.890 143.440 25.150 143.760 ;
        RECT 21.210 142.420 21.470 142.740 ;
        RECT 19.830 140.380 20.090 140.700 ;
        RECT 12.470 138.680 12.730 139.000 ;
        RECT 19.890 138.320 20.030 140.380 ;
        RECT 21.270 138.320 21.410 142.420 ;
        RECT 22.590 140.040 22.850 140.360 ;
        RECT 19.830 138.000 20.090 138.320 ;
        RECT 21.210 138.000 21.470 138.320 ;
        RECT 22.650 136.280 22.790 140.040 ;
        RECT 24.950 136.280 25.090 143.440 ;
        RECT 25.410 143.080 25.550 145.480 ;
        RECT 26.330 143.760 26.470 145.820 ;
        RECT 26.730 145.140 26.990 145.460 ;
        RECT 27.650 145.140 27.910 145.460 ;
        RECT 26.270 143.440 26.530 143.760 ;
        RECT 25.350 142.760 25.610 143.080 ;
        RECT 22.590 135.960 22.850 136.280 ;
        RECT 24.890 135.960 25.150 136.280 ;
        RECT 24.950 130.840 25.090 135.960 ;
        RECT 25.410 134.920 25.550 142.760 ;
        RECT 26.270 142.420 26.530 142.740 ;
        RECT 26.330 137.980 26.470 142.420 ;
        RECT 26.790 138.320 26.930 145.140 ;
        RECT 27.710 144.440 27.850 145.140 ;
        RECT 27.650 144.120 27.910 144.440 ;
        RECT 27.650 143.440 27.910 143.760 ;
        RECT 27.190 143.100 27.450 143.420 ;
        RECT 27.250 140.700 27.390 143.100 ;
        RECT 27.710 141.040 27.850 143.440 ;
        RECT 28.170 141.720 28.310 146.160 ;
        RECT 28.630 145.800 28.770 146.160 ;
        RECT 32.310 146.140 32.450 147.860 ;
        RECT 32.980 147.325 34.520 147.695 ;
        RECT 29.950 145.820 30.210 146.140 ;
        RECT 32.250 145.880 32.510 146.140 ;
        RECT 32.250 145.820 32.910 145.880 ;
        RECT 28.570 145.480 28.830 145.800 ;
        RECT 28.630 142.740 28.770 145.480 ;
        RECT 28.570 142.420 28.830 142.740 ;
        RECT 30.010 142.480 30.150 145.820 ;
        RECT 31.790 145.480 32.050 145.800 ;
        RECT 32.310 145.740 32.910 145.820 ;
        RECT 30.870 145.140 31.130 145.460 ;
        RECT 30.410 142.480 30.670 142.740 ;
        RECT 30.010 142.420 30.670 142.480 ;
        RECT 28.630 141.800 28.770 142.420 ;
        RECT 30.010 142.340 30.610 142.420 ;
        RECT 28.630 141.720 29.230 141.800 ;
        RECT 28.110 141.400 28.370 141.720 ;
        RECT 28.630 141.660 29.290 141.720 ;
        RECT 29.030 141.400 29.290 141.660 ;
        RECT 28.570 141.060 28.830 141.380 ;
        RECT 27.650 140.720 27.910 141.040 ;
        RECT 27.190 140.380 27.450 140.700 ;
        RECT 26.730 138.000 26.990 138.320 ;
        RECT 26.270 137.660 26.530 137.980 ;
        RECT 25.350 134.600 25.610 134.920 ;
        RECT 24.890 130.520 25.150 130.840 ;
        RECT 24.950 129.560 25.090 130.520 ;
        RECT 18.910 129.160 19.170 129.480 ;
        RECT 24.490 129.420 25.090 129.560 ;
        RECT 25.410 129.480 25.550 134.600 ;
        RECT 26.270 132.560 26.530 132.880 ;
        RECT 26.330 130.160 26.470 132.560 ;
        RECT 26.270 129.840 26.530 130.160 ;
        RECT 18.970 127.440 19.110 129.160 ;
        RECT 24.490 129.140 24.630 129.420 ;
        RECT 25.350 129.160 25.610 129.480 ;
        RECT 21.670 128.820 21.930 129.140 ;
        RECT 23.970 128.820 24.230 129.140 ;
        RECT 24.430 128.820 24.690 129.140 ;
        RECT 21.730 127.440 21.870 128.820 ;
        RECT 24.030 128.120 24.170 128.820 ;
        RECT 26.330 128.120 26.470 129.840 ;
        RECT 26.730 129.160 26.990 129.480 ;
        RECT 23.970 127.800 24.230 128.120 ;
        RECT 26.270 127.800 26.530 128.120 ;
        RECT 18.910 127.120 19.170 127.440 ;
        RECT 21.670 127.120 21.930 127.440 ;
        RECT 26.790 126.420 26.930 129.160 ;
        RECT 27.250 127.780 27.390 140.380 ;
        RECT 28.110 138.230 28.370 138.320 ;
        RECT 28.630 138.230 28.770 141.060 ;
        RECT 30.010 140.700 30.150 142.340 ;
        RECT 30.410 141.400 30.670 141.720 ;
        RECT 30.470 140.700 30.610 141.400 ;
        RECT 29.950 140.380 30.210 140.700 ;
        RECT 30.410 140.380 30.670 140.700 ;
        RECT 30.930 138.320 31.070 145.140 ;
        RECT 31.850 144.440 31.990 145.480 ;
        RECT 31.790 144.120 32.050 144.440 ;
        RECT 31.850 140.700 31.990 144.120 ;
        RECT 32.770 143.760 32.910 145.740 ;
        RECT 32.710 143.440 32.970 143.760 ;
        RECT 32.980 141.885 34.520 142.255 ;
        RECT 35.530 140.700 35.670 147.860 ;
        RECT 35.990 145.460 36.130 148.880 ;
        RECT 35.930 145.140 36.190 145.460 ;
        RECT 38.690 145.140 38.950 145.460 ;
        RECT 35.990 141.720 36.130 145.140 ;
        RECT 36.280 144.605 37.820 144.975 ;
        RECT 38.750 144.100 38.890 145.140 ;
        RECT 39.670 144.440 39.810 149.220 ;
        RECT 39.610 144.120 39.870 144.440 ;
        RECT 38.690 143.780 38.950 144.100 ;
        RECT 36.850 142.420 37.110 142.740 ;
        RECT 35.930 141.400 36.190 141.720 ;
        RECT 36.910 140.700 37.050 142.420 ;
        RECT 37.370 141.720 38.430 141.800 ;
        RECT 37.310 141.660 38.430 141.720 ;
        RECT 37.310 141.400 37.570 141.660 ;
        RECT 38.290 141.380 38.430 141.660 ;
        RECT 38.230 141.060 38.490 141.380 ;
        RECT 38.690 140.720 38.950 141.040 ;
        RECT 31.790 140.380 32.050 140.700 ;
        RECT 32.250 140.555 32.510 140.700 ;
        RECT 32.240 140.185 32.520 140.555 ;
        RECT 35.470 140.380 35.730 140.700 ;
        RECT 35.930 140.380 36.190 140.700 ;
        RECT 36.850 140.380 37.110 140.700 ;
        RECT 35.990 138.320 36.130 140.380 ;
        RECT 36.280 139.165 37.820 139.535 ;
        RECT 38.230 138.340 38.490 138.660 ;
        RECT 28.110 138.090 28.770 138.230 ;
        RECT 28.110 138.000 28.370 138.090 ;
        RECT 30.870 138.000 31.130 138.320 ;
        RECT 35.930 138.000 36.190 138.320 ;
        RECT 27.650 137.660 27.910 137.980 ;
        RECT 27.710 129.480 27.850 137.660 ;
        RECT 28.570 136.980 28.830 137.300 ;
        RECT 36.850 136.980 37.110 137.300 ;
        RECT 28.630 134.580 28.770 136.980 ;
        RECT 32.980 136.445 34.520 136.815 ;
        RECT 36.910 135.260 37.050 136.980 ;
        RECT 38.290 136.280 38.430 138.340 ;
        RECT 38.750 138.320 38.890 140.720 ;
        RECT 39.670 140.700 39.810 144.120 ;
        RECT 40.130 142.740 40.270 151.940 ;
        RECT 41.050 149.880 41.190 156.700 ;
        RECT 41.510 153.960 41.650 159.340 ;
        RECT 43.350 157.360 43.490 161.460 ;
        RECT 43.290 157.040 43.550 157.360 ;
        RECT 43.810 154.640 43.950 165.970 ;
        RECT 44.670 165.200 44.930 165.520 ;
        RECT 44.730 162.460 44.870 165.200 ;
        RECT 44.670 162.140 44.930 162.460 ;
        RECT 44.210 161.800 44.470 162.120 ;
        RECT 44.270 160.420 44.410 161.800 ;
        RECT 44.210 160.100 44.470 160.420 ;
        RECT 44.670 156.700 44.930 157.020 ;
        RECT 43.290 154.320 43.550 154.640 ;
        RECT 43.750 154.320 44.010 154.640 ;
        RECT 42.830 153.980 43.090 154.300 ;
        RECT 41.450 153.640 41.710 153.960 ;
        RECT 42.890 151.580 43.030 153.980 ;
        RECT 42.830 151.260 43.090 151.580 ;
        RECT 43.350 151.490 43.490 154.320 ;
        RECT 44.730 153.620 44.870 156.700 ;
        RECT 44.670 153.300 44.930 153.620 ;
        RECT 45.190 152.260 45.330 173.700 ;
        RECT 45.650 173.000 45.790 175.740 ;
        RECT 47.030 175.120 47.170 176.080 ;
        RECT 47.490 175.720 47.630 178.460 ;
        RECT 47.430 175.400 47.690 175.720 ;
        RECT 47.030 174.980 47.630 175.120 ;
        RECT 45.590 172.680 45.850 173.000 ;
        RECT 46.050 172.340 46.310 172.660 ;
        RECT 46.110 168.920 46.250 172.340 ;
        RECT 46.050 168.600 46.310 168.920 ;
        RECT 46.110 167.560 46.250 168.600 ;
        RECT 46.050 167.240 46.310 167.560 ;
        RECT 46.510 166.900 46.770 167.220 ;
        RECT 46.570 165.520 46.710 166.900 ;
        RECT 46.510 165.200 46.770 165.520 ;
        RECT 46.970 164.180 47.230 164.500 ;
        RECT 45.590 162.480 45.850 162.800 ;
        RECT 45.130 151.940 45.390 152.260 ;
        RECT 43.750 151.490 44.010 151.580 ;
        RECT 43.350 151.350 44.010 151.490 ;
        RECT 43.750 151.260 44.010 151.350 ;
        RECT 40.990 149.560 41.250 149.880 ;
        RECT 40.530 145.820 40.790 146.140 ;
        RECT 40.590 143.420 40.730 145.820 ;
        RECT 41.050 144.100 41.190 149.560 ;
        RECT 42.890 149.540 43.030 151.260 ;
        RECT 42.830 149.220 43.090 149.540 ;
        RECT 43.810 149.200 43.950 151.260 ;
        RECT 43.750 148.880 44.010 149.200 ;
        RECT 41.450 148.200 41.710 148.520 ;
        RECT 41.510 146.480 41.650 148.200 ;
        RECT 44.670 147.860 44.930 148.180 ;
        RECT 41.450 146.160 41.710 146.480 ;
        RECT 40.990 143.780 41.250 144.100 ;
        RECT 40.530 143.100 40.790 143.420 ;
        RECT 40.070 142.420 40.330 142.740 ;
        RECT 39.610 140.380 39.870 140.700 ;
        RECT 40.130 140.020 40.270 142.420 ;
        RECT 41.510 140.555 41.650 146.160 ;
        RECT 44.730 146.140 44.870 147.860 ;
        RECT 45.650 147.160 45.790 162.480 ;
        RECT 46.510 159.760 46.770 160.080 ;
        RECT 46.570 158.040 46.710 159.760 ;
        RECT 47.030 159.740 47.170 164.180 ;
        RECT 47.490 159.740 47.630 174.980 ;
        RECT 48.810 172.340 49.070 172.660 ;
        RECT 48.870 171.640 49.010 172.340 ;
        RECT 48.810 171.320 49.070 171.640 ;
        RECT 48.870 162.460 49.010 171.320 ;
        RECT 50.710 168.240 50.850 181.180 ;
        RECT 51.170 178.100 51.310 181.520 ;
        RECT 51.630 178.100 51.770 181.860 ;
        RECT 51.110 177.780 51.370 178.100 ;
        RECT 51.570 177.780 51.830 178.100 ;
        RECT 52.950 177.780 53.210 178.100 ;
        RECT 50.650 167.920 50.910 168.240 ;
        RECT 49.270 164.520 49.530 164.840 ;
        RECT 48.810 162.140 49.070 162.460 ;
        RECT 48.810 160.440 49.070 160.760 ;
        RECT 48.350 160.100 48.610 160.420 ;
        RECT 47.890 159.760 48.150 160.080 ;
        RECT 46.970 159.420 47.230 159.740 ;
        RECT 47.430 159.420 47.690 159.740 ;
        RECT 46.050 157.720 46.310 158.040 ;
        RECT 46.510 157.720 46.770 158.040 ;
        RECT 46.110 157.440 46.250 157.720 ;
        RECT 46.110 157.300 47.170 157.440 ;
        RECT 46.050 153.300 46.310 153.620 ;
        RECT 45.590 147.070 45.850 147.160 ;
        RECT 45.190 146.930 45.850 147.070 ;
        RECT 44.670 145.820 44.930 146.140 ;
        RECT 45.190 143.760 45.330 146.930 ;
        RECT 45.590 146.840 45.850 146.930 ;
        RECT 45.590 145.140 45.850 145.460 ;
        RECT 41.910 143.440 42.170 143.760 ;
        RECT 45.130 143.440 45.390 143.760 ;
        RECT 40.990 140.040 41.250 140.360 ;
        RECT 41.440 140.185 41.720 140.555 ;
        RECT 39.150 139.700 39.410 140.020 ;
        RECT 40.070 139.700 40.330 140.020 ;
        RECT 38.690 138.000 38.950 138.320 ;
        RECT 38.690 137.320 38.950 137.640 ;
        RECT 38.230 135.960 38.490 136.280 ;
        RECT 36.850 134.940 37.110 135.260 ;
        RECT 38.750 135.170 38.890 137.320 ;
        RECT 39.210 135.940 39.350 139.700 ;
        RECT 39.610 138.000 39.870 138.320 ;
        RECT 39.150 135.620 39.410 135.940 ;
        RECT 38.750 135.030 39.350 135.170 ;
        RECT 28.570 134.260 28.830 134.580 ;
        RECT 36.280 133.725 37.820 134.095 ;
        RECT 39.210 132.880 39.350 135.030 ;
        RECT 35.010 132.560 35.270 132.880 ;
        RECT 39.150 132.560 39.410 132.880 ;
        RECT 29.030 131.540 29.290 131.860 ;
        RECT 29.090 129.480 29.230 131.540 ;
        RECT 32.980 131.005 34.520 131.375 ;
        RECT 29.950 130.180 30.210 130.500 ;
        RECT 27.650 129.160 27.910 129.480 ;
        RECT 29.030 129.160 29.290 129.480 ;
        RECT 28.110 128.820 28.370 129.140 ;
        RECT 27.190 127.460 27.450 127.780 ;
        RECT 26.730 126.100 26.990 126.420 ;
        RECT 27.250 124.380 27.390 127.460 ;
        RECT 27.190 124.060 27.450 124.380 ;
        RECT 27.250 122.340 27.390 124.060 ;
        RECT 28.170 124.040 28.310 128.820 ;
        RECT 29.030 127.460 29.290 127.780 ;
        RECT 29.090 125.400 29.230 127.460 ;
        RECT 30.010 126.760 30.150 130.180 ;
        RECT 34.090 129.500 34.350 129.820 ;
        RECT 30.410 128.820 30.670 129.140 ;
        RECT 30.870 128.820 31.130 129.140 ;
        RECT 32.250 128.820 32.510 129.140 ;
        RECT 30.470 128.120 30.610 128.820 ;
        RECT 30.410 127.800 30.670 128.120 ;
        RECT 29.950 126.440 30.210 126.760 ;
        RECT 29.030 125.080 29.290 125.400 ;
        RECT 28.110 123.720 28.370 124.040 ;
        RECT 30.010 122.680 30.150 126.440 ;
        RECT 30.930 124.040 31.070 128.820 ;
        RECT 31.790 127.800 32.050 128.120 ;
        RECT 31.330 127.460 31.590 127.780 ;
        RECT 31.390 126.420 31.530 127.460 ;
        RECT 31.850 127.440 31.990 127.800 ;
        RECT 31.790 127.120 32.050 127.440 ;
        RECT 31.330 126.100 31.590 126.420 ;
        RECT 32.310 124.800 32.450 128.820 ;
        RECT 34.150 127.780 34.290 129.500 ;
        RECT 34.090 127.460 34.350 127.780 ;
        RECT 35.070 126.420 35.210 132.560 ;
        RECT 35.930 132.220 36.190 132.540 ;
        RECT 35.470 131.540 35.730 131.860 ;
        RECT 35.530 127.440 35.670 131.540 ;
        RECT 35.990 128.120 36.130 132.220 ;
        RECT 39.210 129.820 39.350 132.560 ;
        RECT 39.670 132.200 39.810 138.000 ;
        RECT 40.130 137.640 40.270 139.700 ;
        RECT 41.050 138.320 41.190 140.040 ;
        RECT 40.990 138.000 41.250 138.320 ;
        RECT 40.070 137.320 40.330 137.640 ;
        RECT 41.050 137.300 41.190 138.000 ;
        RECT 40.990 136.980 41.250 137.300 ;
        RECT 40.070 134.940 40.330 135.260 ;
        RECT 40.530 134.940 40.790 135.260 ;
        RECT 39.610 131.880 39.870 132.200 ;
        RECT 40.130 130.840 40.270 134.940 ;
        RECT 40.590 132.880 40.730 134.940 ;
        RECT 40.990 132.900 41.250 133.220 ;
        RECT 40.530 132.560 40.790 132.880 ;
        RECT 40.070 130.520 40.330 130.840 ;
        RECT 40.070 129.840 40.330 130.160 ;
        RECT 39.150 129.500 39.410 129.820 ;
        RECT 38.230 129.160 38.490 129.480 ;
        RECT 36.280 128.285 37.820 128.655 ;
        RECT 38.290 128.120 38.430 129.160 ;
        RECT 38.690 128.820 38.950 129.140 ;
        RECT 35.930 127.800 36.190 128.120 ;
        RECT 38.230 127.800 38.490 128.120 ;
        RECT 35.470 127.120 35.730 127.440 ;
        RECT 35.920 127.265 36.200 127.635 ;
        RECT 37.760 127.265 38.040 127.635 ;
        RECT 38.750 127.520 38.890 128.820 ;
        RECT 38.290 127.440 38.890 127.520 ;
        RECT 38.230 127.380 38.890 127.440 ;
        RECT 35.990 127.100 36.130 127.265 ;
        RECT 37.770 127.120 38.030 127.265 ;
        RECT 38.230 127.120 38.490 127.380 ;
        RECT 35.930 127.010 36.190 127.100 ;
        RECT 35.930 126.870 36.590 127.010 ;
        RECT 35.930 126.780 36.190 126.870 ;
        RECT 35.470 126.440 35.730 126.760 ;
        RECT 35.010 126.100 35.270 126.420 ;
        RECT 32.980 125.565 34.520 125.935 ;
        RECT 32.310 124.660 33.370 124.800 ;
        RECT 35.530 124.720 35.670 126.440 ;
        RECT 35.930 126.100 36.190 126.420 ;
        RECT 35.990 125.400 36.130 126.100 ;
        RECT 35.930 125.080 36.190 125.400 ;
        RECT 36.450 124.800 36.590 126.870 ;
        RECT 33.230 124.380 33.370 124.660 ;
        RECT 35.470 124.400 35.730 124.720 ;
        RECT 35.990 124.660 36.590 124.800 ;
        RECT 33.170 124.060 33.430 124.380 ;
        RECT 30.870 123.720 31.130 124.040 ;
        RECT 33.630 123.720 33.890 124.040 ;
        RECT 30.930 122.680 31.070 123.720 ;
        RECT 32.710 123.380 32.970 123.700 ;
        RECT 29.950 122.360 30.210 122.680 ;
        RECT 30.870 122.360 31.130 122.680 ;
        RECT 27.190 122.020 27.450 122.340 ;
        RECT 27.250 118.940 27.390 122.020 ;
        RECT 32.770 122.000 32.910 123.380 ;
        RECT 33.690 122.340 33.830 123.720 ;
        RECT 33.630 122.020 33.890 122.340 ;
        RECT 32.710 121.680 32.970 122.000 ;
        RECT 32.980 120.125 34.520 120.495 ;
        RECT 27.190 118.620 27.450 118.940 ;
        RECT 35.470 118.620 35.730 118.940 ;
        RECT 20.750 116.580 21.010 116.900 ;
        RECT 20.810 111.800 20.950 116.580 ;
        RECT 24.890 115.900 25.150 116.220 ;
        RECT 21.670 114.200 21.930 114.520 ;
        RECT 20.750 111.480 21.010 111.800 ;
        RECT 21.730 111.460 21.870 114.200 ;
        RECT 24.950 111.800 25.090 115.900 ;
        RECT 26.730 115.560 26.990 115.880 ;
        RECT 25.810 115.220 26.070 115.540 ;
        RECT 25.870 113.500 26.010 115.220 ;
        RECT 26.790 113.500 26.930 115.560 ;
        RECT 28.570 115.220 28.830 115.540 ;
        RECT 29.030 115.220 29.290 115.540 ;
        RECT 25.810 113.180 26.070 113.500 ;
        RECT 26.730 113.180 26.990 113.500 ;
        RECT 24.890 111.480 25.150 111.800 ;
        RECT 21.670 111.140 21.930 111.460 ;
        RECT 21.670 109.780 21.930 110.100 ;
        RECT 21.730 105.340 21.870 109.780 ;
        RECT 24.950 107.720 25.090 111.480 ;
        RECT 26.790 111.120 26.930 113.180 ;
        RECT 27.190 111.200 27.450 111.460 ;
        RECT 28.110 111.200 28.370 111.460 ;
        RECT 27.190 111.140 28.370 111.200 ;
        RECT 26.730 110.800 26.990 111.120 ;
        RECT 27.250 111.060 28.310 111.140 ;
        RECT 25.810 110.520 26.070 110.780 ;
        RECT 25.810 110.460 28.310 110.520 ;
        RECT 25.870 110.380 28.310 110.460 ;
        RECT 28.170 110.100 28.310 110.380 ;
        RECT 27.650 109.780 27.910 110.100 ;
        RECT 28.110 109.780 28.370 110.100 ;
        RECT 27.710 109.080 27.850 109.780 ;
        RECT 25.810 108.760 26.070 109.080 ;
        RECT 27.650 108.760 27.910 109.080 ;
        RECT 24.890 107.400 25.150 107.720 ;
        RECT 23.510 107.060 23.770 107.380 ;
        RECT 23.570 105.680 23.710 107.060 ;
        RECT 23.510 105.360 23.770 105.680 ;
        RECT 21.670 105.020 21.930 105.340 ;
        RECT 21.730 102.960 21.870 105.020 ;
        RECT 24.950 103.200 25.090 107.400 ;
        RECT 24.490 103.060 25.090 103.200 ;
        RECT 21.670 102.640 21.930 102.960 ;
        RECT 21.730 95.480 21.870 102.640 ;
        RECT 23.510 101.960 23.770 102.280 ;
        RECT 22.590 101.620 22.850 101.940 ;
        RECT 22.650 100.580 22.790 101.620 ;
        RECT 23.570 100.920 23.710 101.960 ;
        RECT 23.510 100.600 23.770 100.920 ;
        RECT 22.590 100.260 22.850 100.580 ;
        RECT 24.490 99.220 24.630 103.060 ;
        RECT 25.870 100.920 26.010 108.760 ;
        RECT 28.630 108.740 28.770 115.220 ;
        RECT 29.090 112.820 29.230 115.220 ;
        RECT 32.980 114.685 34.520 115.055 ;
        RECT 29.490 114.200 29.750 114.520 ;
        RECT 29.030 112.500 29.290 112.820 ;
        RECT 28.570 108.420 28.830 108.740 ;
        RECT 29.090 105.340 29.230 112.500 ;
        RECT 29.550 108.060 29.690 114.200 ;
        RECT 29.950 113.860 30.210 114.180 ;
        RECT 30.010 111.460 30.150 113.860 ;
        RECT 35.530 113.500 35.670 118.620 ;
        RECT 35.990 115.540 36.130 124.660 ;
        RECT 38.290 124.380 38.430 127.120 ;
        RECT 38.690 126.840 38.950 127.100 ;
        RECT 39.210 126.840 39.350 129.500 ;
        RECT 38.690 126.780 39.350 126.840 ;
        RECT 38.750 126.700 39.350 126.780 ;
        RECT 38.230 124.060 38.490 124.380 ;
        RECT 38.750 123.440 38.890 126.700 ;
        RECT 40.130 126.420 40.270 129.840 ;
        RECT 40.590 128.120 40.730 132.560 ;
        RECT 41.050 129.140 41.190 132.900 ;
        RECT 40.990 128.820 41.250 129.140 ;
        RECT 40.530 127.800 40.790 128.120 ;
        RECT 40.070 126.100 40.330 126.420 ;
        RECT 39.610 125.080 39.870 125.400 ;
        RECT 38.290 123.300 38.890 123.440 ;
        RECT 36.280 122.845 37.820 123.215 ;
        RECT 36.280 117.405 37.820 117.775 ;
        RECT 36.390 115.560 36.650 115.880 ;
        RECT 35.930 115.220 36.190 115.540 ;
        RECT 34.540 112.985 34.820 113.355 ;
        RECT 35.470 113.180 35.730 113.500 ;
        RECT 36.450 113.240 36.590 115.560 ;
        RECT 35.990 113.160 36.590 113.240 ;
        RECT 34.610 111.460 34.750 112.985 ;
        RECT 35.010 112.840 35.270 113.160 ;
        RECT 35.990 113.100 36.650 113.160 ;
        RECT 29.950 111.140 30.210 111.460 ;
        RECT 34.550 111.140 34.810 111.460 ;
        RECT 30.010 108.060 30.150 111.140 ;
        RECT 35.070 110.100 35.210 112.840 ;
        RECT 35.470 112.500 35.730 112.820 ;
        RECT 30.870 109.780 31.130 110.100 ;
        RECT 35.010 109.780 35.270 110.100 ;
        RECT 29.490 107.740 29.750 108.060 ;
        RECT 29.950 107.740 30.210 108.060 ;
        RECT 29.550 107.380 29.690 107.740 ;
        RECT 29.490 107.060 29.750 107.380 ;
        RECT 29.030 105.020 29.290 105.340 ;
        RECT 29.550 104.660 29.690 107.060 ;
        RECT 30.010 106.020 30.150 107.740 ;
        RECT 30.930 106.360 31.070 109.780 ;
        RECT 32.980 109.245 34.520 109.615 ;
        RECT 31.330 107.740 31.590 108.060 ;
        RECT 32.250 107.740 32.510 108.060 ;
        RECT 30.870 106.040 31.130 106.360 ;
        RECT 29.950 105.700 30.210 106.020 ;
        RECT 28.110 104.340 28.370 104.660 ;
        RECT 29.490 104.340 29.750 104.660 ;
        RECT 28.170 102.620 28.310 104.340 ;
        RECT 30.010 102.960 30.150 105.700 ;
        RECT 29.950 102.640 30.210 102.960 ;
        RECT 31.390 102.620 31.530 107.740 ;
        RECT 28.110 102.300 28.370 102.620 ;
        RECT 31.330 102.300 31.590 102.620 ;
        RECT 27.650 101.960 27.910 102.280 ;
        RECT 25.810 100.600 26.070 100.920 ;
        RECT 27.710 100.240 27.850 101.960 ;
        RECT 28.170 100.240 28.310 102.300 ;
        RECT 30.410 101.620 30.670 101.940 ;
        RECT 30.470 100.240 30.610 101.620 ;
        RECT 32.310 100.920 32.450 107.740 ;
        RECT 33.630 107.400 33.890 107.720 ;
        RECT 33.690 106.360 33.830 107.400 ;
        RECT 35.070 107.380 35.210 109.780 ;
        RECT 35.530 108.060 35.670 112.500 ;
        RECT 35.990 111.120 36.130 113.100 ;
        RECT 36.390 112.840 36.650 113.100 ;
        RECT 36.280 111.965 37.820 112.335 ;
        RECT 38.290 111.460 38.430 123.300 ;
        RECT 39.670 122.340 39.810 125.080 ;
        RECT 39.610 122.020 39.870 122.340 ;
        RECT 40.130 120.980 40.270 126.100 ;
        RECT 40.530 123.720 40.790 124.040 ;
        RECT 40.590 122.680 40.730 123.720 ;
        RECT 40.530 122.360 40.790 122.680 ;
        RECT 40.070 120.660 40.330 120.980 ;
        RECT 41.510 117.000 41.650 140.185 ;
        RECT 41.970 138.320 42.110 143.440 ;
        RECT 45.190 143.080 45.330 143.440 ;
        RECT 45.130 142.760 45.390 143.080 ;
        RECT 42.370 142.420 42.630 142.740 ;
        RECT 44.670 142.420 44.930 142.740 ;
        RECT 42.430 141.040 42.570 142.420 ;
        RECT 42.370 140.720 42.630 141.040 ;
        RECT 44.730 140.700 44.870 142.420 ;
        RECT 42.830 140.380 43.090 140.700 ;
        RECT 44.670 140.380 44.930 140.700 ;
        RECT 45.130 140.380 45.390 140.700 ;
        RECT 41.910 138.000 42.170 138.320 ;
        RECT 41.970 137.640 42.110 138.000 ;
        RECT 41.910 137.320 42.170 137.640 ;
        RECT 42.890 135.940 43.030 140.380 ;
        RECT 44.210 139.700 44.470 140.020 ;
        RECT 44.270 138.660 44.410 139.700 ;
        RECT 43.290 138.340 43.550 138.660 ;
        RECT 44.210 138.340 44.470 138.660 ;
        RECT 43.350 136.280 43.490 138.340 ;
        RECT 45.190 137.980 45.330 140.380 ;
        RECT 45.130 137.660 45.390 137.980 ;
        RECT 45.650 137.210 45.790 145.140 ;
        RECT 45.190 137.070 45.790 137.210 ;
        RECT 43.290 135.960 43.550 136.280 ;
        RECT 42.830 135.620 43.090 135.940 ;
        RECT 42.890 133.560 43.030 135.620 ;
        RECT 42.830 133.240 43.090 133.560 ;
        RECT 40.590 116.860 41.650 117.000 ;
        RECT 39.150 114.200 39.410 114.520 ;
        RECT 39.210 113.500 39.350 114.200 ;
        RECT 40.590 113.500 40.730 116.860 ;
        RECT 44.670 115.220 44.930 115.540 ;
        RECT 44.210 114.200 44.470 114.520 ;
        RECT 41.450 114.090 41.710 114.180 ;
        RECT 42.830 114.090 43.090 114.180 ;
        RECT 41.450 113.950 43.090 114.090 ;
        RECT 41.450 113.860 41.710 113.950 ;
        RECT 42.830 113.860 43.090 113.950 ;
        RECT 44.270 113.500 44.410 114.200 ;
        RECT 44.730 113.840 44.870 115.220 ;
        RECT 44.670 113.520 44.930 113.840 ;
        RECT 39.150 113.180 39.410 113.500 ;
        RECT 38.230 111.140 38.490 111.460 ;
        RECT 35.930 110.800 36.190 111.120 ;
        RECT 38.290 108.060 38.430 111.140 ;
        RECT 39.210 110.100 39.350 113.180 ;
        RECT 39.610 112.840 39.870 113.160 ;
        RECT 40.060 112.985 40.340 113.355 ;
        RECT 40.530 113.180 40.790 113.500 ;
        RECT 40.070 112.840 40.330 112.985 ;
        RECT 41.450 112.840 41.710 113.160 ;
        RECT 42.820 112.985 43.100 113.355 ;
        RECT 44.210 113.180 44.470 113.500 ;
        RECT 39.150 109.780 39.410 110.100 ;
        RECT 39.670 108.740 39.810 112.840 ;
        RECT 40.530 112.500 40.790 112.820 ;
        RECT 40.070 110.800 40.330 111.120 ;
        RECT 40.130 109.080 40.270 110.800 ;
        RECT 40.070 108.760 40.330 109.080 ;
        RECT 39.610 108.420 39.870 108.740 ;
        RECT 40.590 108.400 40.730 112.500 ;
        RECT 40.990 111.480 41.250 111.800 ;
        RECT 41.050 109.080 41.190 111.480 ;
        RECT 40.990 108.760 41.250 109.080 ;
        RECT 40.530 108.080 40.790 108.400 ;
        RECT 40.990 108.080 41.250 108.400 ;
        RECT 35.470 107.740 35.730 108.060 ;
        RECT 38.230 107.740 38.490 108.060 ;
        RECT 41.050 107.380 41.190 108.080 ;
        RECT 41.510 108.060 41.650 112.840 ;
        RECT 42.890 111.800 43.030 112.985 ;
        RECT 42.830 111.480 43.090 111.800 ;
        RECT 43.750 109.780 44.010 110.100 ;
        RECT 44.210 109.780 44.470 110.100 ;
        RECT 42.370 108.420 42.630 108.740 ;
        RECT 41.450 107.740 41.710 108.060 ;
        RECT 35.010 107.060 35.270 107.380 ;
        RECT 39.610 107.060 39.870 107.380 ;
        RECT 40.990 107.060 41.250 107.380 ;
        RECT 35.070 106.360 35.210 107.060 ;
        RECT 36.280 106.525 37.820 106.895 ;
        RECT 33.630 106.040 33.890 106.360 ;
        RECT 35.010 106.040 35.270 106.360 ;
        RECT 39.670 106.020 39.810 107.060 ;
        RECT 39.610 105.700 39.870 106.020 ;
        RECT 35.010 105.360 35.270 105.680 ;
        RECT 32.980 103.805 34.520 104.175 ;
        RECT 35.070 102.620 35.210 105.360 ;
        RECT 41.050 102.620 41.190 107.060 ;
        RECT 32.710 102.300 32.970 102.620 ;
        RECT 35.010 102.300 35.270 102.620 ;
        RECT 40.990 102.300 41.250 102.620 ;
        RECT 32.250 100.600 32.510 100.920 ;
        RECT 24.890 99.920 25.150 100.240 ;
        RECT 27.650 99.920 27.910 100.240 ;
        RECT 28.110 99.920 28.370 100.240 ;
        RECT 29.030 99.920 29.290 100.240 ;
        RECT 30.410 99.920 30.670 100.240 ;
        RECT 24.950 99.640 25.090 99.920 ;
        RECT 24.950 99.500 25.550 99.640 ;
        RECT 24.430 98.900 24.690 99.220 ;
        RECT 24.890 98.900 25.150 99.220 ;
        RECT 24.490 98.200 24.630 98.900 ;
        RECT 24.430 97.880 24.690 98.200 ;
        RECT 21.670 95.160 21.930 95.480 ;
        RECT 21.730 92.080 21.870 95.160 ;
        RECT 24.490 94.120 24.630 97.880 ;
        RECT 24.950 96.840 25.090 98.900 ;
        RECT 25.410 97.180 25.550 99.500 ;
        RECT 27.710 97.180 27.850 99.920 ;
        RECT 29.090 99.560 29.230 99.920 ;
        RECT 32.770 99.560 32.910 102.300 ;
        RECT 35.010 101.620 35.270 101.940 ;
        RECT 35.070 100.580 35.210 101.620 ;
        RECT 36.280 101.085 37.820 101.455 ;
        RECT 35.010 100.260 35.270 100.580 ;
        RECT 38.230 100.260 38.490 100.580 ;
        RECT 29.030 99.240 29.290 99.560 ;
        RECT 32.710 99.240 32.970 99.560 ;
        RECT 32.980 98.365 34.520 98.735 ;
        RECT 34.090 98.110 34.350 98.200 ;
        RECT 35.070 98.110 35.210 100.260 ;
        RECT 38.290 98.200 38.430 100.260 ;
        RECT 39.610 98.900 39.870 99.220 ;
        RECT 40.530 98.900 40.790 99.220 ;
        RECT 39.670 98.200 39.810 98.900 ;
        RECT 34.090 97.970 35.210 98.110 ;
        RECT 34.090 97.880 34.350 97.970 ;
        RECT 38.230 97.880 38.490 98.200 ;
        RECT 39.610 97.880 39.870 98.200 ;
        RECT 25.350 96.860 25.610 97.180 ;
        RECT 27.650 96.860 27.910 97.180 ;
        RECT 24.890 96.520 25.150 96.840 ;
        RECT 24.950 94.120 25.090 96.520 ;
        RECT 25.410 94.800 25.550 96.860 ;
        RECT 28.110 96.180 28.370 96.500 ;
        RECT 28.170 95.480 28.310 96.180 ;
        RECT 28.110 95.160 28.370 95.480 ;
        RECT 25.350 94.480 25.610 94.800 ;
        RECT 24.430 93.800 24.690 94.120 ;
        RECT 24.890 93.800 25.150 94.120 ;
        RECT 23.050 93.460 23.310 93.780 ;
        RECT 21.670 91.760 21.930 92.080 ;
        RECT 23.110 91.740 23.250 93.460 ;
        RECT 25.410 92.840 25.550 94.480 ;
        RECT 34.150 93.780 34.290 97.880 ;
        RECT 38.230 96.860 38.490 97.180 ;
        RECT 36.280 95.645 37.820 96.015 ;
        RECT 35.010 94.820 35.270 95.140 ;
        RECT 35.070 94.120 35.210 94.820 ;
        RECT 38.290 94.800 38.430 96.860 ;
        RECT 39.610 96.520 39.870 96.840 ;
        RECT 39.670 95.480 39.810 96.520 ;
        RECT 39.610 95.160 39.870 95.480 ;
        RECT 38.230 94.480 38.490 94.800 ;
        RECT 35.010 93.800 35.270 94.120 ;
        RECT 40.590 93.780 40.730 98.900 ;
        RECT 41.050 95.480 41.190 102.300 ;
        RECT 42.430 100.240 42.570 108.420 ;
        RECT 43.810 107.720 43.950 109.780 ;
        RECT 43.750 107.400 44.010 107.720 ;
        RECT 44.270 100.920 44.410 109.780 ;
        RECT 45.190 108.060 45.330 137.070 ;
        RECT 46.110 135.260 46.250 153.300 ;
        RECT 47.030 136.280 47.170 157.300 ;
        RECT 47.490 154.640 47.630 159.420 ;
        RECT 47.950 157.700 48.090 159.760 ;
        RECT 47.890 157.380 48.150 157.700 ;
        RECT 48.410 157.020 48.550 160.100 ;
        RECT 48.870 157.360 49.010 160.440 ;
        RECT 49.330 159.060 49.470 164.520 ;
        RECT 49.730 161.460 49.990 161.780 ;
        RECT 49.270 158.740 49.530 159.060 ;
        RECT 48.810 157.040 49.070 157.360 ;
        RECT 47.890 156.700 48.150 157.020 ;
        RECT 48.350 156.700 48.610 157.020 ;
        RECT 47.950 156.340 48.090 156.700 ;
        RECT 47.890 156.020 48.150 156.340 ;
        RECT 47.950 154.640 48.090 156.020 ;
        RECT 47.430 154.320 47.690 154.640 ;
        RECT 47.890 154.320 48.150 154.640 ;
        RECT 48.870 146.140 49.010 157.040 ;
        RECT 49.790 156.340 49.930 161.460 ;
        RECT 50.710 159.740 50.850 167.920 ;
        RECT 51.170 165.860 51.310 177.780 ;
        RECT 51.110 165.540 51.370 165.860 ;
        RECT 51.630 164.840 51.770 177.780 ;
        RECT 53.010 176.400 53.150 177.780 ;
        RECT 53.470 176.740 53.610 183.900 ;
        RECT 54.390 181.840 54.530 184.920 ;
        RECT 55.310 182.180 55.450 185.940 ;
        RECT 64.510 185.240 64.650 186.960 ;
        RECT 64.450 184.920 64.710 185.240 ;
        RECT 66.350 184.560 66.490 186.960 ;
        RECT 66.290 184.240 66.550 184.560 ;
        RECT 67.270 183.880 67.410 191.380 ;
        RECT 69.050 189.340 69.310 189.660 ;
        RECT 70.430 189.340 70.690 189.660 ;
        RECT 67.670 186.620 67.930 186.940 ;
        RECT 68.130 186.620 68.390 186.940 ;
        RECT 67.730 184.075 67.870 186.620 ;
        RECT 55.710 183.560 55.970 183.880 ;
        RECT 67.210 183.560 67.470 183.880 ;
        RECT 67.660 183.705 67.940 184.075 ;
        RECT 67.670 183.560 67.930 183.705 ;
        RECT 55.250 181.860 55.510 182.180 ;
        RECT 54.330 181.520 54.590 181.840 ;
        RECT 54.790 181.520 55.050 181.840 ;
        RECT 53.410 176.420 53.670 176.740 ;
        RECT 52.950 176.080 53.210 176.400 ;
        RECT 53.470 173.000 53.610 176.420 ;
        RECT 53.410 172.680 53.670 173.000 ;
        RECT 53.870 172.680 54.130 173.000 ;
        RECT 53.470 171.300 53.610 172.680 ;
        RECT 53.410 170.980 53.670 171.300 ;
        RECT 53.930 168.920 54.070 172.680 ;
        RECT 53.870 168.600 54.130 168.920 ;
        RECT 54.390 168.580 54.530 181.520 ;
        RECT 53.410 168.260 53.670 168.580 ;
        RECT 54.330 168.260 54.590 168.580 ;
        RECT 52.950 165.540 53.210 165.860 ;
        RECT 51.570 164.520 51.830 164.840 ;
        RECT 52.490 164.520 52.750 164.840 ;
        RECT 51.110 162.820 51.370 163.140 ;
        RECT 51.170 160.080 51.310 162.820 ;
        RECT 52.550 160.760 52.690 164.520 ;
        RECT 53.010 160.955 53.150 165.540 ;
        RECT 52.490 160.440 52.750 160.760 ;
        RECT 52.940 160.585 53.220 160.955 ;
        RECT 51.570 160.100 51.830 160.420 ;
        RECT 51.110 159.760 51.370 160.080 ;
        RECT 50.650 159.420 50.910 159.740 ;
        RECT 50.710 157.700 50.850 159.420 ;
        RECT 50.650 157.380 50.910 157.700 ;
        RECT 51.630 157.020 51.770 160.100 ;
        RECT 53.010 159.740 53.150 160.585 ;
        RECT 52.950 159.420 53.210 159.740 ;
        RECT 53.470 157.360 53.610 168.260 ;
        RECT 54.330 167.580 54.590 167.900 ;
        RECT 53.870 165.200 54.130 165.520 ;
        RECT 53.930 162.800 54.070 165.200 ;
        RECT 54.390 165.180 54.530 167.580 ;
        RECT 54.850 166.960 54.990 181.520 ;
        RECT 55.310 179.460 55.450 181.860 ;
        RECT 55.770 181.160 55.910 183.560 ;
        RECT 57.090 183.220 57.350 183.540 ;
        RECT 55.710 180.840 55.970 181.160 ;
        RECT 55.250 179.140 55.510 179.460 ;
        RECT 57.150 173.000 57.290 183.220 ;
        RECT 67.270 181.500 67.410 183.560 ;
        RECT 67.210 181.180 67.470 181.500 ;
        RECT 67.670 179.100 67.930 179.120 ;
        RECT 68.190 179.100 68.330 186.620 ;
        RECT 68.590 185.940 68.850 186.260 ;
        RECT 68.650 184.560 68.790 185.940 ;
        RECT 69.110 184.900 69.250 189.340 ;
        RECT 70.490 185.240 70.630 189.340 ;
        RECT 70.950 187.960 71.090 192.060 ;
        RECT 71.410 189.320 71.550 192.400 ;
        RECT 71.350 189.000 71.610 189.320 ;
        RECT 71.410 187.960 71.550 189.000 ;
        RECT 70.890 187.640 71.150 187.960 ;
        RECT 71.350 187.640 71.610 187.960 ;
        RECT 70.430 184.920 70.690 185.240 ;
        RECT 71.810 184.920 72.070 185.240 ;
        RECT 69.050 184.580 69.310 184.900 ;
        RECT 69.970 184.580 70.230 184.900 ;
        RECT 68.590 184.240 68.850 184.560 ;
        RECT 70.030 182.520 70.170 184.580 ;
        RECT 69.970 182.200 70.230 182.520 ;
        RECT 71.870 181.840 72.010 184.920 ;
        RECT 72.330 184.900 72.470 192.400 ;
        RECT 77.850 192.040 77.990 203.280 ;
        RECT 81.470 192.400 81.730 192.720 ;
        RECT 120.570 192.400 120.830 192.720 ;
        RECT 78.710 192.060 78.970 192.380 ;
        RECT 77.790 191.720 78.050 192.040 ;
        RECT 74.570 190.020 74.830 190.340 ;
        RECT 73.650 189.340 73.910 189.660 ;
        RECT 73.190 188.660 73.450 188.980 ;
        RECT 72.730 186.960 72.990 187.280 ;
        RECT 72.790 185.240 72.930 186.960 ;
        RECT 72.730 184.920 72.990 185.240 ;
        RECT 72.270 184.580 72.530 184.900 ;
        RECT 72.270 183.900 72.530 184.220 ;
        RECT 71.810 181.520 72.070 181.840 ;
        RECT 72.330 181.500 72.470 183.900 ;
        RECT 73.250 181.750 73.390 188.660 ;
        RECT 73.710 187.620 73.850 189.340 ;
        RECT 74.110 187.640 74.370 187.960 ;
        RECT 73.650 187.300 73.910 187.620 ;
        RECT 73.710 184.220 73.850 187.300 ;
        RECT 74.170 185.240 74.310 187.640 ;
        RECT 74.630 187.280 74.770 190.020 ;
        RECT 77.850 189.320 77.990 191.720 ;
        RECT 78.250 191.380 78.510 191.700 ;
        RECT 78.310 190.680 78.450 191.380 ;
        RECT 78.250 190.360 78.510 190.680 ;
        RECT 77.790 189.000 78.050 189.320 ;
        RECT 78.770 188.980 78.910 192.060 ;
        RECT 78.710 188.660 78.970 188.980 ;
        RECT 74.570 186.960 74.830 187.280 ;
        RECT 74.110 184.920 74.370 185.240 ;
        RECT 73.650 183.900 73.910 184.220 ;
        RECT 74.170 182.180 74.310 184.920 ;
        RECT 74.630 184.220 74.770 186.960 ;
        RECT 78.770 186.940 78.910 188.660 ;
        RECT 78.710 186.620 78.970 186.940 ;
        RECT 79.630 186.620 79.890 186.940 ;
        RECT 76.870 185.940 77.130 186.260 ;
        RECT 77.330 185.940 77.590 186.260 ;
        RECT 76.930 184.220 77.070 185.940 ;
        RECT 77.390 184.560 77.530 185.940 ;
        RECT 77.330 184.240 77.590 184.560 ;
        RECT 78.770 184.220 78.910 186.620 ;
        RECT 79.690 186.115 79.830 186.620 ;
        RECT 79.620 185.745 79.900 186.115 ;
        RECT 81.010 185.940 81.270 186.260 ;
        RECT 80.550 184.920 80.810 185.240 ;
        RECT 80.610 184.220 80.750 184.920 ;
        RECT 81.070 184.560 81.210 185.940 ;
        RECT 81.010 184.240 81.270 184.560 ;
        RECT 74.570 183.900 74.830 184.220 ;
        RECT 75.490 184.075 75.750 184.220 ;
        RECT 75.480 183.705 75.760 184.075 ;
        RECT 76.870 183.900 77.130 184.220 ;
        RECT 78.710 183.900 78.970 184.220 ;
        RECT 80.550 183.900 80.810 184.220 ;
        RECT 77.790 183.560 78.050 183.880 ;
        RECT 77.850 182.520 77.990 183.560 ;
        RECT 78.770 183.540 78.910 183.900 ;
        RECT 78.710 183.220 78.970 183.540 ;
        RECT 80.550 183.280 80.810 183.540 ;
        RECT 81.530 183.280 81.670 192.400 ;
        RECT 83.310 191.380 83.570 191.700 ;
        RECT 117.810 191.380 118.070 191.700 ;
        RECT 81.930 186.960 82.190 187.280 ;
        RECT 81.990 185.240 82.130 186.960 ;
        RECT 81.930 184.920 82.190 185.240 ;
        RECT 83.370 184.075 83.510 191.380 ;
        RECT 108.150 189.680 108.410 190.000 ;
        RECT 99.870 189.570 100.130 189.660 ;
        RECT 99.870 189.430 100.530 189.570 ;
        RECT 99.870 189.340 100.130 189.430 ;
        RECT 84.230 188.660 84.490 188.980 ;
        RECT 94.810 188.660 95.070 188.980 ;
        RECT 95.730 188.660 95.990 188.980 ;
        RECT 84.290 187.620 84.430 188.660 ;
        RECT 84.230 187.300 84.490 187.620 ;
        RECT 94.350 187.300 94.610 187.620 ;
        RECT 84.690 186.960 84.950 187.280 ;
        RECT 85.610 186.960 85.870 187.280 ;
        RECT 83.300 183.705 83.580 184.075 ;
        RECT 80.550 183.220 81.670 183.280 ;
        RECT 80.610 183.140 81.670 183.220 ;
        RECT 77.790 182.200 78.050 182.520 ;
        RECT 74.110 181.860 74.370 182.180 ;
        RECT 73.250 181.610 73.850 181.750 ;
        RECT 69.050 181.180 69.310 181.500 ;
        RECT 72.270 181.180 72.530 181.500 ;
        RECT 67.670 178.960 68.330 179.100 ;
        RECT 67.670 178.800 67.930 178.960 ;
        RECT 57.550 178.460 57.810 178.780 ;
        RECT 57.610 177.080 57.750 178.460 ;
        RECT 67.730 178.100 67.870 178.800 ;
        RECT 69.110 178.780 69.250 181.180 ;
        RECT 70.430 180.500 70.690 180.820 ;
        RECT 71.350 180.500 71.610 180.820 ;
        RECT 71.810 180.500 72.070 180.820 ;
        RECT 68.130 178.460 68.390 178.780 ;
        RECT 69.050 178.460 69.310 178.780 ;
        RECT 62.610 177.780 62.870 178.100 ;
        RECT 67.670 177.780 67.930 178.100 ;
        RECT 57.550 176.760 57.810 177.080 ;
        RECT 56.630 172.680 56.890 173.000 ;
        RECT 57.090 172.680 57.350 173.000 ;
        RECT 55.250 169.620 55.510 169.940 ;
        RECT 55.310 167.900 55.450 169.620 ;
        RECT 56.690 168.240 56.830 172.680 ;
        RECT 57.610 171.300 57.750 176.760 ;
        RECT 59.850 175.740 60.110 176.060 ;
        RECT 59.390 175.060 59.650 175.380 ;
        RECT 59.450 174.020 59.590 175.060 ;
        RECT 59.390 173.700 59.650 174.020 ;
        RECT 59.910 173.340 60.050 175.740 ;
        RECT 62.670 173.340 62.810 177.780 ;
        RECT 68.190 174.360 68.330 178.460 ;
        RECT 70.490 178.440 70.630 180.500 ;
        RECT 71.410 178.780 71.550 180.500 ;
        RECT 71.350 178.690 71.610 178.780 ;
        RECT 70.950 178.550 71.610 178.690 ;
        RECT 70.430 178.120 70.690 178.440 ;
        RECT 70.490 176.400 70.630 178.120 ;
        RECT 70.950 177.080 71.090 178.550 ;
        RECT 71.350 178.460 71.610 178.550 ;
        RECT 71.350 177.780 71.610 178.100 ;
        RECT 71.410 177.080 71.550 177.780 ;
        RECT 70.890 176.760 71.150 177.080 ;
        RECT 71.350 176.760 71.610 177.080 ;
        RECT 71.870 176.400 72.010 180.500 ;
        RECT 72.330 176.400 72.470 181.180 ;
        RECT 73.190 180.840 73.450 181.160 ;
        RECT 73.250 179.460 73.390 180.840 ;
        RECT 73.190 179.140 73.450 179.460 ;
        RECT 73.250 177.080 73.390 179.140 ;
        RECT 73.710 178.780 73.850 181.610 ;
        RECT 81.070 180.820 81.210 183.140 ;
        RECT 81.470 181.860 81.730 182.180 ;
        RECT 81.010 180.500 81.270 180.820 ;
        RECT 73.650 178.460 73.910 178.780 ;
        RECT 74.570 178.460 74.830 178.780 ;
        RECT 75.950 178.460 76.210 178.780 ;
        RECT 79.630 178.460 79.890 178.780 ;
        RECT 73.190 176.760 73.450 177.080 ;
        RECT 70.430 176.080 70.690 176.400 ;
        RECT 71.810 176.080 72.070 176.400 ;
        RECT 72.270 176.080 72.530 176.400 ;
        RECT 71.870 174.360 72.010 176.080 ;
        RECT 68.130 174.040 68.390 174.360 ;
        RECT 71.810 174.040 72.070 174.360 ;
        RECT 59.850 173.020 60.110 173.340 ;
        RECT 62.610 173.020 62.870 173.340 ;
        RECT 58.470 172.340 58.730 172.660 ;
        RECT 69.510 172.340 69.770 172.660 ;
        RECT 71.350 172.340 71.610 172.660 ;
        RECT 58.530 171.640 58.670 172.340 ;
        RECT 58.470 171.320 58.730 171.640 ;
        RECT 57.090 170.980 57.350 171.300 ;
        RECT 57.550 170.980 57.810 171.300 ;
        RECT 69.570 171.155 69.710 172.340 ;
        RECT 56.630 167.920 56.890 168.240 ;
        RECT 57.150 167.900 57.290 170.980 ;
        RECT 69.500 170.785 69.780 171.155 ;
        RECT 64.450 170.300 64.710 170.620 ;
        RECT 64.510 167.900 64.650 170.300 ;
        RECT 55.250 167.580 55.510 167.900 ;
        RECT 57.090 167.580 57.350 167.900 ;
        RECT 64.450 167.580 64.710 167.900 ;
        RECT 67.210 167.580 67.470 167.900 ;
        RECT 69.510 167.580 69.770 167.900 ;
        RECT 55.250 166.960 55.510 167.220 ;
        RECT 54.850 166.900 55.510 166.960 ;
        RECT 54.850 166.820 55.450 166.900 ;
        RECT 55.310 165.180 55.450 166.820 ;
        RECT 54.330 164.860 54.590 165.180 ;
        RECT 55.250 164.860 55.510 165.180 ;
        RECT 54.390 163.140 54.530 164.860 ;
        RECT 54.330 162.820 54.590 163.140 ;
        RECT 53.870 162.480 54.130 162.800 ;
        RECT 53.930 161.780 54.070 162.480 ;
        RECT 53.870 161.460 54.130 161.780 ;
        RECT 53.930 160.760 54.070 161.460 ;
        RECT 53.870 160.440 54.130 160.760 ;
        RECT 54.790 159.760 55.050 160.080 ;
        RECT 54.330 158.740 54.590 159.060 ;
        RECT 53.410 157.040 53.670 157.360 ;
        RECT 51.570 156.700 51.830 157.020 ;
        RECT 49.730 156.020 49.990 156.340 ;
        RECT 50.190 156.020 50.450 156.340 ;
        RECT 49.790 154.640 49.930 156.020 ;
        RECT 49.730 154.320 49.990 154.640 ;
        RECT 50.250 153.620 50.390 156.020 ;
        RECT 54.390 154.300 54.530 158.740 ;
        RECT 54.850 155.320 54.990 159.760 ;
        RECT 55.310 156.680 55.450 164.860 ;
        RECT 63.990 164.520 64.250 164.840 ;
        RECT 63.530 164.180 63.790 164.500 ;
        RECT 56.630 162.140 56.890 162.460 ;
        RECT 63.070 162.140 63.330 162.460 ;
        RECT 55.710 161.460 55.970 161.780 ;
        RECT 55.770 157.360 55.910 161.460 ;
        RECT 56.160 160.585 56.440 160.955 ;
        RECT 56.170 160.440 56.430 160.585 ;
        RECT 56.690 157.700 56.830 162.140 ;
        RECT 60.310 161.800 60.570 162.120 ;
        RECT 60.370 158.040 60.510 161.800 ;
        RECT 62.610 159.650 62.870 159.740 ;
        RECT 63.130 159.650 63.270 162.140 ;
        RECT 63.590 160.420 63.730 164.180 ;
        RECT 64.050 160.420 64.190 164.520 ;
        RECT 65.830 164.180 66.090 164.500 ;
        RECT 64.450 163.160 64.710 163.480 ;
        RECT 63.530 160.100 63.790 160.420 ;
        RECT 63.990 160.100 64.250 160.420 ;
        RECT 64.510 159.740 64.650 163.160 ;
        RECT 65.890 163.140 66.030 164.180 ;
        RECT 65.830 162.820 66.090 163.140 ;
        RECT 62.610 159.510 63.270 159.650 ;
        RECT 62.610 159.420 62.870 159.510 ;
        RECT 62.150 158.740 62.410 159.060 ;
        RECT 60.310 157.720 60.570 158.040 ;
        RECT 56.630 157.380 56.890 157.700 ;
        RECT 55.710 157.040 55.970 157.360 ;
        RECT 55.250 156.360 55.510 156.680 ;
        RECT 54.790 155.000 55.050 155.320 ;
        RECT 56.690 154.640 56.830 157.380 ;
        RECT 62.210 157.020 62.350 158.740 ;
        RECT 63.130 157.020 63.270 159.510 ;
        RECT 64.450 159.420 64.710 159.740 ;
        RECT 62.150 156.700 62.410 157.020 ;
        RECT 63.070 156.700 63.330 157.020 ;
        RECT 67.270 156.680 67.410 167.580 ;
        RECT 69.050 167.240 69.310 167.560 ;
        RECT 69.110 165.520 69.250 167.240 ;
        RECT 69.570 165.520 69.710 167.580 ;
        RECT 71.410 167.560 71.550 172.340 ;
        RECT 72.330 167.900 72.470 176.080 ;
        RECT 73.710 175.970 73.850 178.460 ;
        RECT 72.790 175.830 73.850 175.970 ;
        RECT 72.790 173.340 72.930 175.830 ;
        RECT 73.190 175.060 73.450 175.380 ;
        RECT 72.730 173.020 72.990 173.340 ;
        RECT 72.270 167.580 72.530 167.900 ;
        RECT 71.350 167.240 71.610 167.560 ;
        RECT 69.050 165.200 69.310 165.520 ;
        RECT 69.510 165.200 69.770 165.520 ;
        RECT 73.250 162.120 73.390 175.060 ;
        RECT 74.110 173.020 74.370 173.340 ;
        RECT 74.170 171.300 74.310 173.020 ;
        RECT 74.630 171.640 74.770 178.460 ;
        RECT 76.010 177.080 76.150 178.460 ;
        RECT 77.790 177.780 78.050 178.100 ;
        RECT 75.950 176.760 76.210 177.080 ;
        RECT 75.490 176.420 75.750 176.740 ;
        RECT 75.550 174.360 75.690 176.420 ;
        RECT 76.010 174.360 76.150 176.760 ;
        RECT 76.410 176.080 76.670 176.400 ;
        RECT 75.490 174.040 75.750 174.360 ;
        RECT 75.950 174.040 76.210 174.360 ;
        RECT 75.030 173.700 75.290 174.020 ;
        RECT 74.570 171.320 74.830 171.640 ;
        RECT 75.090 171.300 75.230 173.700 ;
        RECT 75.480 173.505 75.760 173.875 ;
        RECT 75.490 173.360 75.750 173.505 ;
        RECT 75.950 173.020 76.210 173.340 ;
        RECT 76.010 171.835 76.150 173.020 ;
        RECT 75.940 171.465 76.220 171.835 ;
        RECT 76.470 171.640 76.610 176.080 ;
        RECT 76.870 173.360 77.130 173.680 ;
        RECT 77.320 173.505 77.600 173.875 ;
        RECT 76.410 171.320 76.670 171.640 ;
        RECT 74.110 170.980 74.370 171.300 ;
        RECT 75.030 170.980 75.290 171.300 ;
        RECT 74.170 166.200 74.310 170.980 ;
        RECT 76.410 170.300 76.670 170.620 ;
        RECT 74.570 169.620 74.830 169.940 ;
        RECT 74.110 165.880 74.370 166.200 ;
        RECT 74.170 165.600 74.310 165.880 ;
        RECT 73.710 165.460 74.310 165.600 ;
        RECT 73.710 162.800 73.850 165.460 ;
        RECT 74.630 163.480 74.770 169.620 ;
        RECT 76.470 167.900 76.610 170.300 ;
        RECT 76.930 169.940 77.070 173.360 ;
        RECT 76.870 169.620 77.130 169.940 ;
        RECT 76.410 167.580 76.670 167.900 ;
        RECT 77.390 165.300 77.530 173.505 ;
        RECT 77.850 170.960 77.990 177.780 ;
        RECT 79.690 177.080 79.830 178.460 ;
        RECT 79.630 176.760 79.890 177.080 ;
        RECT 79.170 176.420 79.430 176.740 ;
        RECT 79.230 174.360 79.370 176.420 ;
        RECT 80.090 175.060 80.350 175.380 ;
        RECT 81.010 175.060 81.270 175.380 ;
        RECT 79.170 174.040 79.430 174.360 ;
        RECT 79.230 173.680 79.830 173.760 ;
        RECT 80.150 173.680 80.290 175.060 ;
        RECT 79.170 173.620 79.830 173.680 ;
        RECT 79.170 173.360 79.430 173.620 ;
        RECT 77.790 170.640 78.050 170.960 ;
        RECT 79.160 170.785 79.440 171.155 ;
        RECT 79.690 170.960 79.830 173.620 ;
        RECT 80.090 173.360 80.350 173.680 ;
        RECT 80.540 173.505 80.820 173.875 ;
        RECT 79.170 170.640 79.430 170.785 ;
        RECT 79.630 170.640 79.890 170.960 ;
        RECT 79.690 170.360 79.830 170.640 ;
        RECT 78.770 170.280 79.830 170.360 ;
        RECT 78.710 170.220 79.830 170.280 ;
        RECT 78.710 169.960 78.970 170.220 ;
        RECT 79.170 169.620 79.430 169.940 ;
        RECT 77.390 165.160 77.990 165.300 ;
        RECT 74.570 163.160 74.830 163.480 ;
        RECT 74.110 162.820 74.370 163.140 ;
        RECT 73.650 162.480 73.910 162.800 ;
        RECT 72.270 161.800 72.530 162.120 ;
        RECT 73.190 161.800 73.450 162.120 ;
        RECT 70.430 161.460 70.690 161.780 ;
        RECT 71.350 161.460 71.610 161.780 ;
        RECT 66.750 156.360 67.010 156.680 ;
        RECT 67.210 156.360 67.470 156.680 ;
        RECT 56.630 154.320 56.890 154.640 ;
        RECT 66.810 154.300 66.950 156.360 ;
        RECT 67.270 155.320 67.410 156.360 ;
        RECT 67.210 155.000 67.470 155.320 ;
        RECT 51.570 153.980 51.830 154.300 ;
        RECT 54.330 153.980 54.590 154.300 ;
        RECT 66.750 153.980 67.010 154.300 ;
        RECT 50.190 153.300 50.450 153.620 ;
        RECT 48.810 145.820 49.070 146.140 ;
        RECT 50.190 143.440 50.450 143.760 ;
        RECT 49.270 139.700 49.530 140.020 ;
        RECT 49.330 138.320 49.470 139.700 ;
        RECT 50.250 138.320 50.390 143.440 ;
        RECT 49.270 138.000 49.530 138.320 ;
        RECT 50.190 138.000 50.450 138.320 ;
        RECT 50.650 138.000 50.910 138.320 ;
        RECT 48.350 137.320 48.610 137.640 ;
        RECT 46.970 135.960 47.230 136.280 ;
        RECT 46.050 134.940 46.310 135.260 ;
        RECT 46.110 132.540 46.250 134.940 ;
        RECT 46.050 132.220 46.310 132.540 ;
        RECT 48.410 131.860 48.550 137.320 ;
        RECT 49.330 136.280 49.470 138.000 ;
        RECT 49.270 135.960 49.530 136.280 ;
        RECT 49.270 134.940 49.530 135.260 ;
        RECT 48.350 131.540 48.610 131.860 ;
        RECT 47.890 129.840 48.150 130.160 ;
        RECT 45.590 128.820 45.850 129.140 ;
        RECT 45.650 127.440 45.790 128.820 ;
        RECT 45.590 127.120 45.850 127.440 ;
        RECT 45.650 125.400 45.790 127.120 ;
        RECT 45.590 125.080 45.850 125.400 ;
        RECT 45.650 124.040 45.790 125.080 ;
        RECT 47.950 124.040 48.090 129.840 ;
        RECT 48.410 125.400 48.550 131.540 ;
        RECT 48.350 125.080 48.610 125.400 ;
        RECT 45.590 123.720 45.850 124.040 ;
        RECT 47.890 123.720 48.150 124.040 ;
        RECT 48.800 123.865 49.080 124.235 ;
        RECT 48.810 123.720 49.070 123.865 ;
        RECT 47.430 122.250 47.690 122.340 ;
        RECT 47.950 122.250 48.090 123.720 ;
        RECT 49.330 122.680 49.470 134.940 ;
        RECT 50.710 133.220 50.850 138.000 ;
        RECT 51.110 136.980 51.370 137.300 ;
        RECT 51.170 135.260 51.310 136.980 ;
        RECT 51.110 134.940 51.370 135.260 ;
        RECT 51.170 133.560 51.310 134.940 ;
        RECT 51.110 133.240 51.370 133.560 ;
        RECT 50.650 132.900 50.910 133.220 ;
        RECT 51.110 127.120 51.370 127.440 ;
        RECT 50.190 126.780 50.450 127.100 ;
        RECT 50.250 124.040 50.390 126.780 ;
        RECT 51.170 125.400 51.310 127.120 ;
        RECT 51.110 125.080 51.370 125.400 ;
        RECT 50.190 123.720 50.450 124.040 ;
        RECT 50.250 122.680 50.390 123.720 ;
        RECT 49.270 122.360 49.530 122.680 ;
        RECT 50.190 122.360 50.450 122.680 ;
        RECT 47.430 122.110 48.090 122.250 ;
        RECT 47.430 122.020 47.690 122.110 ;
        RECT 45.590 121.340 45.850 121.660 ;
        RECT 45.650 112.820 45.790 121.340 ;
        RECT 51.630 114.180 51.770 153.980 ;
        RECT 66.810 148.860 66.950 153.980 ;
        RECT 69.970 150.580 70.230 150.900 ;
        RECT 66.750 148.540 67.010 148.860 ;
        RECT 54.790 145.820 55.050 146.140 ;
        RECT 52.490 141.400 52.750 141.720 ;
        RECT 52.030 140.380 52.290 140.700 ;
        RECT 52.090 138.660 52.230 140.380 ;
        RECT 52.030 138.340 52.290 138.660 ;
        RECT 52.030 137.660 52.290 137.980 ;
        RECT 52.090 136.280 52.230 137.660 ;
        RECT 52.550 137.640 52.690 141.400 ;
        RECT 54.850 140.700 54.990 145.820 ;
        RECT 57.090 145.480 57.350 145.800 ;
        RECT 59.850 145.480 60.110 145.800 ;
        RECT 56.630 145.140 56.890 145.460 ;
        RECT 54.790 140.380 55.050 140.700 ;
        RECT 53.410 138.570 53.670 138.660 ;
        RECT 53.410 138.430 54.070 138.570 ;
        RECT 53.410 138.340 53.670 138.430 ;
        RECT 52.490 137.320 52.750 137.640 ;
        RECT 53.410 136.980 53.670 137.300 ;
        RECT 52.030 135.960 52.290 136.280 ;
        RECT 53.470 135.600 53.610 136.980 ;
        RECT 53.410 135.280 53.670 135.600 ;
        RECT 52.490 134.940 52.750 135.260 ;
        RECT 52.030 134.260 52.290 134.580 ;
        RECT 52.090 132.880 52.230 134.260 ;
        RECT 52.550 133.560 52.690 134.940 ;
        RECT 52.950 134.600 53.210 134.920 ;
        RECT 52.490 133.240 52.750 133.560 ;
        RECT 52.030 132.560 52.290 132.880 ;
        RECT 52.030 127.120 52.290 127.440 ;
        RECT 52.090 124.720 52.230 127.120 ;
        RECT 53.010 127.100 53.150 134.600 ;
        RECT 53.930 133.560 54.070 138.430 ;
        RECT 54.330 137.660 54.590 137.980 ;
        RECT 54.390 134.580 54.530 137.660 ;
        RECT 54.330 134.260 54.590 134.580 ;
        RECT 53.870 133.240 54.130 133.560 ;
        RECT 54.850 133.220 54.990 140.380 ;
        RECT 55.710 138.340 55.970 138.660 ;
        RECT 55.770 136.280 55.910 138.340 ;
        RECT 56.170 138.230 56.430 138.320 ;
        RECT 56.690 138.230 56.830 145.140 ;
        RECT 56.170 138.090 56.830 138.230 ;
        RECT 56.170 138.000 56.430 138.090 ;
        RECT 55.710 135.960 55.970 136.280 ;
        RECT 55.250 134.600 55.510 134.920 ;
        RECT 55.310 133.560 55.450 134.600 ;
        RECT 55.250 133.240 55.510 133.560 ;
        RECT 54.790 132.900 55.050 133.220 ;
        RECT 54.330 132.560 54.590 132.880 ;
        RECT 54.390 129.820 54.530 132.560 ;
        RECT 53.410 129.500 53.670 129.820 ;
        RECT 54.330 129.500 54.590 129.820 ;
        RECT 52.950 126.780 53.210 127.100 ;
        RECT 53.470 125.400 53.610 129.500 ;
        RECT 54.390 128.120 54.530 129.500 ;
        RECT 54.330 127.800 54.590 128.120 ;
        RECT 53.410 125.080 53.670 125.400 ;
        RECT 52.030 124.400 52.290 124.720 ;
        RECT 52.090 123.700 52.230 124.400 ;
        RECT 53.470 124.380 53.610 125.080 ;
        RECT 54.330 124.740 54.590 125.060 ;
        RECT 52.950 124.235 53.210 124.380 ;
        RECT 52.940 123.865 53.220 124.235 ;
        RECT 53.410 124.060 53.670 124.380 ;
        RECT 52.030 123.380 52.290 123.700 ;
        RECT 54.390 122.340 54.530 124.740 ;
        RECT 54.850 124.720 54.990 132.900 ;
        RECT 55.710 129.500 55.970 129.820 ;
        RECT 55.250 128.820 55.510 129.140 ;
        RECT 54.790 124.400 55.050 124.720 ;
        RECT 55.310 124.040 55.450 128.820 ;
        RECT 55.770 127.780 55.910 129.500 ;
        RECT 56.230 128.030 56.370 138.000 ;
        RECT 57.150 137.300 57.290 145.480 ;
        RECT 57.550 143.440 57.810 143.760 ;
        RECT 58.010 143.440 58.270 143.760 ;
        RECT 57.610 138.320 57.750 143.440 ;
        RECT 57.550 138.000 57.810 138.320 ;
        RECT 57.090 136.980 57.350 137.300 ;
        RECT 56.630 132.900 56.890 133.220 ;
        RECT 56.690 130.840 56.830 132.900 ;
        RECT 56.630 130.520 56.890 130.840 ;
        RECT 57.150 130.160 57.290 136.980 ;
        RECT 57.610 135.600 57.750 138.000 ;
        RECT 58.070 137.300 58.210 143.440 ;
        RECT 59.910 141.720 60.050 145.480 ;
        RECT 63.070 145.140 63.330 145.460 ;
        RECT 63.130 143.760 63.270 145.140 ;
        RECT 66.810 144.100 66.950 148.540 ;
        RECT 66.750 143.780 67.010 144.100 ;
        RECT 70.030 143.760 70.170 150.580 ;
        RECT 70.490 149.540 70.630 161.460 ;
        RECT 71.410 159.060 71.550 161.460 ;
        RECT 71.350 158.740 71.610 159.060 ;
        RECT 72.330 157.700 72.470 161.800 ;
        RECT 74.170 160.760 74.310 162.820 ;
        RECT 73.190 160.440 73.450 160.760 ;
        RECT 74.110 160.440 74.370 160.760 ;
        RECT 73.250 160.080 73.390 160.440 ;
        RECT 74.630 160.160 74.770 163.160 ;
        RECT 77.330 162.140 77.590 162.460 ;
        RECT 76.870 161.460 77.130 161.780 ;
        RECT 73.190 159.760 73.450 160.080 ;
        RECT 73.710 160.020 74.770 160.160 ;
        RECT 76.930 160.080 77.070 161.460 ;
        RECT 77.390 160.760 77.530 162.140 ;
        RECT 77.330 160.440 77.590 160.760 ;
        RECT 77.850 160.080 77.990 165.160 ;
        RECT 78.250 164.860 78.510 165.180 ;
        RECT 73.710 159.740 73.850 160.020 ;
        RECT 73.650 159.420 73.910 159.740 ;
        RECT 74.630 159.060 74.770 160.020 ;
        RECT 76.870 159.760 77.130 160.080 ;
        RECT 77.790 159.760 78.050 160.080 ;
        RECT 75.030 159.420 75.290 159.740 ;
        RECT 74.570 158.740 74.830 159.060 ;
        RECT 74.630 158.040 74.770 158.740 ;
        RECT 75.090 158.040 75.230 159.420 ;
        RECT 76.410 159.080 76.670 159.400 ;
        RECT 74.570 157.720 74.830 158.040 ;
        RECT 75.030 157.720 75.290 158.040 ;
        RECT 72.270 157.380 72.530 157.700 ;
        RECT 74.110 156.020 74.370 156.340 ;
        RECT 70.890 154.320 71.150 154.640 ;
        RECT 70.950 152.600 71.090 154.320 ;
        RECT 73.190 153.300 73.450 153.620 ;
        RECT 70.890 152.280 71.150 152.600 ;
        RECT 73.250 151.920 73.390 153.300 ;
        RECT 74.170 151.920 74.310 156.020 ;
        RECT 76.470 154.640 76.610 159.080 ;
        RECT 76.410 154.320 76.670 154.640 ;
        RECT 76.470 153.620 76.610 154.320 ;
        RECT 76.410 153.300 76.670 153.620 ;
        RECT 73.190 151.600 73.450 151.920 ;
        RECT 74.110 151.600 74.370 151.920 ;
        RECT 74.170 149.880 74.310 151.600 ;
        RECT 76.870 150.920 77.130 151.240 ;
        RECT 75.950 150.580 76.210 150.900 ;
        RECT 76.410 150.580 76.670 150.900 ;
        RECT 74.110 149.560 74.370 149.880 ;
        RECT 70.430 149.220 70.690 149.540 ;
        RECT 70.490 147.160 70.630 149.220 ;
        RECT 72.270 148.880 72.530 149.200 ;
        RECT 70.890 147.860 71.150 148.180 ;
        RECT 70.430 146.840 70.690 147.160 ;
        RECT 70.950 143.760 71.090 147.860 ;
        RECT 72.330 147.160 72.470 148.880 ;
        RECT 73.190 147.860 73.450 148.180 ;
        RECT 72.270 146.840 72.530 147.160 ;
        RECT 73.250 146.140 73.390 147.860 ;
        RECT 76.010 146.820 76.150 150.580 ;
        RECT 75.950 146.500 76.210 146.820 ;
        RECT 76.470 146.480 76.610 150.580 ;
        RECT 76.410 146.160 76.670 146.480 ;
        RECT 73.190 145.820 73.450 146.140 ;
        RECT 73.650 145.820 73.910 146.140 ;
        RECT 73.710 144.100 73.850 145.820 ;
        RECT 73.650 143.780 73.910 144.100 ;
        RECT 60.770 143.440 61.030 143.760 ;
        RECT 63.070 143.440 63.330 143.760 ;
        RECT 69.970 143.440 70.230 143.760 ;
        RECT 70.890 143.440 71.150 143.760 ;
        RECT 59.850 141.400 60.110 141.720 ;
        RECT 60.830 140.700 60.970 143.440 ;
        RECT 68.590 142.420 68.850 142.740 ;
        RECT 68.650 141.040 68.790 142.420 ;
        RECT 70.030 141.720 70.170 143.440 ;
        RECT 69.970 141.400 70.230 141.720 ;
        RECT 68.590 140.720 68.850 141.040 ;
        RECT 70.950 140.700 71.090 143.440 ;
        RECT 71.810 141.060 72.070 141.380 ;
        RECT 71.870 140.700 72.010 141.060 ;
        RECT 76.930 141.040 77.070 150.920 ;
        RECT 77.790 145.880 78.050 146.140 ;
        RECT 77.390 145.820 78.050 145.880 ;
        RECT 77.390 145.740 77.990 145.820 ;
        RECT 77.390 143.760 77.530 145.740 ;
        RECT 78.310 144.440 78.450 164.860 ;
        RECT 78.710 162.480 78.970 162.800 ;
        RECT 78.770 158.040 78.910 162.480 ;
        RECT 79.230 160.420 79.370 169.620 ;
        RECT 80.150 165.180 80.290 173.360 ;
        RECT 80.610 173.340 80.750 173.505 ;
        RECT 80.550 173.020 80.810 173.340 ;
        RECT 81.070 171.640 81.210 175.060 ;
        RECT 81.010 171.320 81.270 171.640 ;
        RECT 81.010 166.900 81.270 167.220 ;
        RECT 80.090 164.860 80.350 165.180 ;
        RECT 80.150 162.460 80.290 164.860 ;
        RECT 81.070 164.840 81.210 166.900 ;
        RECT 81.530 166.200 81.670 181.860 ;
        RECT 82.390 174.040 82.650 174.360 ;
        RECT 81.920 171.465 82.200 171.835 ;
        RECT 81.930 171.320 82.190 171.465 ;
        RECT 82.450 171.300 82.590 174.040 ;
        RECT 83.370 173.680 83.510 183.705 ;
        RECT 84.750 183.540 84.890 186.960 ;
        RECT 85.150 184.580 85.410 184.900 ;
        RECT 84.690 183.220 84.950 183.540 ;
        RECT 85.210 178.100 85.350 184.580 ;
        RECT 85.670 182.520 85.810 186.960 ;
        RECT 92.970 186.620 93.230 186.940 ;
        RECT 89.750 185.940 90.010 186.260 ;
        RECT 89.810 184.220 89.950 185.940 ;
        RECT 89.750 183.900 90.010 184.220 ;
        RECT 90.210 183.900 90.470 184.220 ;
        RECT 85.610 182.200 85.870 182.520 ;
        RECT 89.750 181.180 90.010 181.500 ;
        RECT 89.290 180.500 89.550 180.820 ;
        RECT 84.230 177.780 84.490 178.100 ;
        RECT 85.150 177.780 85.410 178.100 ;
        RECT 83.770 173.700 84.030 174.020 ;
        RECT 83.310 173.360 83.570 173.680 ;
        RECT 82.390 170.980 82.650 171.300 ;
        RECT 82.450 167.900 82.590 170.980 ;
        RECT 83.370 169.940 83.510 173.360 ;
        RECT 83.830 170.960 83.970 173.700 ;
        RECT 84.290 173.680 84.430 177.780 ;
        RECT 86.070 176.080 86.330 176.400 ;
        RECT 86.130 174.360 86.270 176.080 ;
        RECT 86.070 174.040 86.330 174.360 ;
        RECT 84.230 173.360 84.490 173.680 ;
        RECT 86.990 173.020 87.250 173.340 ;
        RECT 87.050 171.300 87.190 173.020 ;
        RECT 87.910 172.340 88.170 172.660 ;
        RECT 87.970 171.640 88.110 172.340 ;
        RECT 87.910 171.320 88.170 171.640 ;
        RECT 86.990 170.980 87.250 171.300 ;
        RECT 83.770 170.640 84.030 170.960 ;
        RECT 88.830 170.640 89.090 170.960 ;
        RECT 83.310 169.620 83.570 169.940 ;
        RECT 82.390 167.580 82.650 167.900 ;
        RECT 81.470 165.880 81.730 166.200 ;
        RECT 82.390 165.200 82.650 165.520 ;
        RECT 81.010 164.520 81.270 164.840 ;
        RECT 81.930 164.180 82.190 164.500 ;
        RECT 81.010 163.160 81.270 163.480 ;
        RECT 80.090 162.140 80.350 162.460 ;
        RECT 79.620 160.585 79.900 160.955 ;
        RECT 79.630 160.440 79.890 160.585 ;
        RECT 79.170 160.100 79.430 160.420 ;
        RECT 80.150 159.740 80.290 162.140 ;
        RECT 81.070 160.760 81.210 163.160 ;
        RECT 81.010 160.440 81.270 160.760 ;
        RECT 81.990 160.080 82.130 164.180 ;
        RECT 81.930 159.760 82.190 160.080 ;
        RECT 80.090 159.420 80.350 159.740 ;
        RECT 82.450 158.040 82.590 165.200 ;
        RECT 83.830 160.080 83.970 170.640 ;
        RECT 84.230 170.300 84.490 170.620 ;
        RECT 84.290 168.920 84.430 170.300 ;
        RECT 88.370 169.960 88.630 170.280 ;
        RECT 87.910 169.620 88.170 169.940 ;
        RECT 84.230 168.600 84.490 168.920 ;
        RECT 84.290 166.200 84.430 168.600 ;
        RECT 86.070 167.240 86.330 167.560 ;
        RECT 86.130 166.200 86.270 167.240 ;
        RECT 84.230 165.880 84.490 166.200 ;
        RECT 86.070 165.880 86.330 166.200 ;
        RECT 87.970 162.800 88.110 169.620 ;
        RECT 88.430 165.180 88.570 169.960 ;
        RECT 88.370 164.860 88.630 165.180 ;
        RECT 87.910 162.480 88.170 162.800 ;
        RECT 84.230 162.140 84.490 162.460 ;
        RECT 84.690 162.140 84.950 162.460 ;
        RECT 84.290 160.760 84.430 162.140 ;
        RECT 84.230 160.440 84.490 160.760 ;
        RECT 83.770 159.760 84.030 160.080 ;
        RECT 78.710 157.720 78.970 158.040 ;
        RECT 82.390 157.720 82.650 158.040 ;
        RECT 84.750 156.680 84.890 162.140 ;
        RECT 87.970 158.040 88.110 162.480 ;
        RECT 87.910 157.720 88.170 158.040 ;
        RECT 84.690 156.360 84.950 156.680 ;
        RECT 84.750 153.620 84.890 156.360 ;
        RECT 85.610 155.000 85.870 155.320 ;
        RECT 84.690 153.300 84.950 153.620 ;
        RECT 80.090 151.600 80.350 151.920 ;
        RECT 78.710 148.880 78.970 149.200 ;
        RECT 78.770 147.160 78.910 148.880 ;
        RECT 80.150 148.860 80.290 151.600 ;
        RECT 80.090 148.540 80.350 148.860 ;
        RECT 78.710 146.840 78.970 147.160 ;
        RECT 80.150 146.480 80.290 148.540 ;
        RECT 80.090 146.160 80.350 146.480 ;
        RECT 80.090 145.480 80.350 145.800 ;
        RECT 78.710 145.140 78.970 145.460 ;
        RECT 78.770 144.440 78.910 145.140 ;
        RECT 78.250 144.120 78.510 144.440 ;
        RECT 78.710 144.120 78.970 144.440 ;
        RECT 78.770 143.760 78.910 144.120 ;
        RECT 77.330 143.440 77.590 143.760 ;
        RECT 78.710 143.440 78.970 143.760 ;
        RECT 72.730 140.720 72.990 141.040 ;
        RECT 76.870 140.720 77.130 141.040 ;
        RECT 60.770 140.380 61.030 140.700 ;
        RECT 70.890 140.380 71.150 140.700 ;
        RECT 71.810 140.380 72.070 140.700 ;
        RECT 58.470 139.700 58.730 140.020 ;
        RECT 59.850 139.700 60.110 140.020 ;
        RECT 58.530 138.320 58.670 139.700 ;
        RECT 58.930 138.340 59.190 138.660 ;
        RECT 59.390 138.340 59.650 138.660 ;
        RECT 58.470 138.000 58.730 138.320 ;
        RECT 58.010 136.980 58.270 137.300 ;
        RECT 57.550 135.280 57.810 135.600 ;
        RECT 58.470 134.490 58.730 134.580 ;
        RECT 58.990 134.490 59.130 138.340 ;
        RECT 59.450 135.260 59.590 138.340 ;
        RECT 59.910 137.300 60.050 139.700 ;
        RECT 70.950 138.320 71.090 140.380 ;
        RECT 71.870 139.080 72.010 140.380 ;
        RECT 71.870 138.940 72.470 139.080 ;
        RECT 62.150 138.000 62.410 138.320 ;
        RECT 70.890 138.230 71.150 138.320 ;
        RECT 70.890 138.090 72.010 138.230 ;
        RECT 70.890 138.000 71.150 138.090 ;
        RECT 59.850 136.980 60.110 137.300 ;
        RECT 59.390 134.940 59.650 135.260 ;
        RECT 58.470 134.350 59.130 134.490 ;
        RECT 58.470 134.260 58.730 134.350 ;
        RECT 58.530 131.860 58.670 134.260 ;
        RECT 58.470 131.540 58.730 131.860 ;
        RECT 57.090 129.840 57.350 130.160 ;
        RECT 58.530 129.820 58.670 131.540 ;
        RECT 59.450 130.160 59.590 134.940 ;
        RECT 59.910 134.920 60.050 136.980 ;
        RECT 62.210 136.280 62.350 138.000 ;
        RECT 71.350 136.980 71.610 137.300 ;
        RECT 62.150 135.960 62.410 136.280 ;
        RECT 59.850 134.600 60.110 134.920 ;
        RECT 66.750 132.220 67.010 132.540 ;
        RECT 66.810 130.160 66.950 132.220 ;
        RECT 59.390 129.840 59.650 130.160 ;
        RECT 66.750 129.840 67.010 130.160 ;
        RECT 58.470 129.500 58.730 129.820 ;
        RECT 56.230 127.890 56.830 128.030 ;
        RECT 55.710 127.460 55.970 127.780 ;
        RECT 56.170 127.120 56.430 127.440 ;
        RECT 56.230 125.400 56.370 127.120 ;
        RECT 56.690 126.420 56.830 127.890 ;
        RECT 66.810 127.440 66.950 129.840 ;
        RECT 66.750 127.120 67.010 127.440 ;
        RECT 70.890 127.120 71.150 127.440 ;
        RECT 56.630 126.100 56.890 126.420 ;
        RECT 56.170 125.080 56.430 125.400 ;
        RECT 56.690 125.060 56.830 126.100 ;
        RECT 56.630 124.740 56.890 125.060 ;
        RECT 55.250 123.720 55.510 124.040 ;
        RECT 66.810 122.340 66.950 127.120 ;
        RECT 70.950 125.400 71.090 127.120 ;
        RECT 70.890 125.080 71.150 125.400 ;
        RECT 54.330 122.020 54.590 122.340 ;
        RECT 66.750 122.020 67.010 122.340 ;
        RECT 60.310 121.680 60.570 122.000 ;
        RECT 60.370 118.260 60.510 121.680 ;
        RECT 66.810 118.940 66.950 122.020 ;
        RECT 68.130 121.680 68.390 122.000 ;
        RECT 68.190 119.280 68.330 121.680 ;
        RECT 68.130 118.960 68.390 119.280 ;
        RECT 66.750 118.620 67.010 118.940 ;
        RECT 60.310 117.940 60.570 118.260 ;
        RECT 61.690 117.940 61.950 118.260 ;
        RECT 59.850 115.900 60.110 116.220 ;
        RECT 47.890 113.860 48.150 114.180 ;
        RECT 51.570 113.860 51.830 114.180 ;
        RECT 46.050 113.180 46.310 113.500 ;
        RECT 45.590 112.500 45.850 112.820 ;
        RECT 46.110 110.780 46.250 113.180 ;
        RECT 46.050 110.460 46.310 110.780 ;
        RECT 46.050 109.780 46.310 110.100 ;
        RECT 44.670 107.740 44.930 108.060 ;
        RECT 45.130 107.740 45.390 108.060 ;
        RECT 46.110 107.970 46.250 109.780 ;
        RECT 47.950 108.060 48.090 113.860 ;
        RECT 58.470 113.180 58.730 113.500 ;
        RECT 57.090 112.500 57.350 112.820 ;
        RECT 57.150 111.800 57.290 112.500 ;
        RECT 55.710 111.480 55.970 111.800 ;
        RECT 57.090 111.480 57.350 111.800 ;
        RECT 48.810 111.140 49.070 111.460 ;
        RECT 48.350 109.780 48.610 110.100 ;
        RECT 46.510 107.970 46.770 108.060 ;
        RECT 46.110 107.830 46.770 107.970 ;
        RECT 46.510 107.740 46.770 107.830 ;
        RECT 47.890 107.740 48.150 108.060 ;
        RECT 44.730 100.920 44.870 107.740 ;
        RECT 45.190 106.360 45.330 107.740 ;
        RECT 47.430 107.060 47.690 107.380 ;
        RECT 45.130 106.040 45.390 106.360 ;
        RECT 47.490 105.680 47.630 107.060 ;
        RECT 48.410 105.680 48.550 109.780 ;
        RECT 48.870 109.080 49.010 111.140 ;
        RECT 52.030 110.460 52.290 110.780 ;
        RECT 48.810 108.760 49.070 109.080 ;
        RECT 48.870 106.360 49.010 108.760 ;
        RECT 52.090 107.380 52.230 110.460 ;
        RECT 55.770 107.380 55.910 111.480 ;
        RECT 58.530 111.120 58.670 113.180 ;
        RECT 58.470 110.800 58.730 111.120 ;
        RECT 59.910 110.440 60.050 115.900 ;
        RECT 60.370 111.460 60.510 117.940 ;
        RECT 61.750 114.520 61.890 117.940 ;
        RECT 66.810 116.560 66.950 118.620 ;
        RECT 67.210 118.280 67.470 118.600 ;
        RECT 63.070 116.240 63.330 116.560 ;
        RECT 66.750 116.240 67.010 116.560 ;
        RECT 61.690 114.200 61.950 114.520 ;
        RECT 63.130 112.820 63.270 116.240 ;
        RECT 67.270 115.540 67.410 118.280 ;
        RECT 67.210 115.220 67.470 115.540 ;
        RECT 64.450 112.840 64.710 113.160 ;
        RECT 63.070 112.500 63.330 112.820 ;
        RECT 60.310 111.140 60.570 111.460 ;
        RECT 63.130 110.440 63.270 112.500 ;
        RECT 64.510 110.780 64.650 112.840 ;
        RECT 64.450 110.460 64.710 110.780 ;
        RECT 59.850 110.120 60.110 110.440 ;
        RECT 63.070 110.120 63.330 110.440 ;
        RECT 63.990 108.080 64.250 108.400 ;
        RECT 57.550 107.400 57.810 107.720 ;
        RECT 52.030 107.060 52.290 107.380 ;
        RECT 55.710 107.060 55.970 107.380 ;
        RECT 52.090 106.360 52.230 107.060 ;
        RECT 57.610 106.360 57.750 107.400 ;
        RECT 48.810 106.040 49.070 106.360 ;
        RECT 52.030 106.040 52.290 106.360 ;
        RECT 57.550 106.040 57.810 106.360 ;
        RECT 64.050 105.680 64.190 108.080 ;
        RECT 64.510 108.060 64.650 110.460 ;
        RECT 66.740 109.585 67.020 109.955 ;
        RECT 66.810 108.400 66.950 109.585 ;
        RECT 67.270 108.740 67.410 115.220 ;
        RECT 68.190 112.820 68.330 118.960 ;
        RECT 69.510 113.180 69.770 113.500 ;
        RECT 68.130 112.500 68.390 112.820 ;
        RECT 68.590 112.500 68.850 112.820 ;
        RECT 68.190 110.780 68.330 112.500 ;
        RECT 68.650 111.800 68.790 112.500 ;
        RECT 69.570 111.800 69.710 113.180 ;
        RECT 68.590 111.480 68.850 111.800 ;
        RECT 69.510 111.480 69.770 111.800 ;
        RECT 68.130 110.460 68.390 110.780 ;
        RECT 67.210 108.420 67.470 108.740 ;
        RECT 66.750 108.080 67.010 108.400 ;
        RECT 68.190 108.060 68.330 110.460 ;
        RECT 69.570 109.080 69.710 111.480 ;
        RECT 69.970 110.800 70.230 111.120 ;
        RECT 69.510 108.760 69.770 109.080 ;
        RECT 64.450 107.740 64.710 108.060 ;
        RECT 68.130 107.740 68.390 108.060 ;
        RECT 47.430 105.360 47.690 105.680 ;
        RECT 48.350 105.360 48.610 105.680 ;
        RECT 51.110 105.360 51.370 105.680 ;
        RECT 51.570 105.360 51.830 105.680 ;
        RECT 52.490 105.360 52.750 105.680 ;
        RECT 54.330 105.360 54.590 105.680 ;
        RECT 63.990 105.360 64.250 105.680 ;
        RECT 51.170 103.640 51.310 105.360 ;
        RECT 51.630 105.000 51.770 105.360 ;
        RECT 51.570 104.680 51.830 105.000 ;
        RECT 51.110 103.320 51.370 103.640 ;
        RECT 50.650 101.620 50.910 101.940 ;
        RECT 44.210 100.600 44.470 100.920 ;
        RECT 44.670 100.600 44.930 100.920 ;
        RECT 44.270 100.240 44.410 100.600 ;
        RECT 42.370 99.920 42.630 100.240 ;
        RECT 44.210 99.920 44.470 100.240 ;
        RECT 42.430 97.180 42.570 99.920 ;
        RECT 42.370 96.860 42.630 97.180 ;
        RECT 42.430 95.480 42.570 96.860 ;
        RECT 44.270 96.500 44.410 99.920 ;
        RECT 44.730 97.860 44.870 100.600 ;
        RECT 50.710 100.240 50.850 101.620 ;
        RECT 51.630 100.580 51.770 104.680 ;
        RECT 52.550 101.940 52.690 105.360 ;
        RECT 54.390 104.660 54.530 105.360 ;
        RECT 54.330 104.340 54.590 104.660 ;
        RECT 52.490 101.620 52.750 101.940 ;
        RECT 52.550 100.920 52.690 101.620 ;
        RECT 52.490 100.600 52.750 100.920 ;
        RECT 51.570 100.260 51.830 100.580 ;
        RECT 53.410 100.260 53.670 100.580 ;
        RECT 49.270 99.920 49.530 100.240 ;
        RECT 50.650 99.920 50.910 100.240 ;
        RECT 44.670 97.540 44.930 97.860 ;
        RECT 44.210 96.180 44.470 96.500 ;
        RECT 44.730 95.560 44.870 97.540 ;
        RECT 45.130 96.180 45.390 96.500 ;
        RECT 40.990 95.160 41.250 95.480 ;
        RECT 42.370 95.160 42.630 95.480 ;
        RECT 44.270 95.420 44.870 95.560 ;
        RECT 44.270 95.140 44.410 95.420 ;
        RECT 44.210 94.820 44.470 95.140 ;
        RECT 45.190 93.780 45.330 96.180 ;
        RECT 49.330 95.140 49.470 99.920 ;
        RECT 50.710 96.840 50.850 99.920 ;
        RECT 50.650 96.520 50.910 96.840 ;
        RECT 51.630 95.140 51.770 100.260 ;
        RECT 53.470 99.220 53.610 100.260 ;
        RECT 54.390 100.240 54.530 104.340 ;
        RECT 55.710 102.300 55.970 102.620 ;
        RECT 53.870 99.920 54.130 100.240 ;
        RECT 54.330 99.920 54.590 100.240 ;
        RECT 53.930 99.560 54.070 99.920 ;
        RECT 53.870 99.240 54.130 99.560 ;
        RECT 53.410 98.900 53.670 99.220 ;
        RECT 53.470 97.860 53.610 98.900 ;
        RECT 53.410 97.540 53.670 97.860 ;
        RECT 49.270 94.820 49.530 95.140 ;
        RECT 51.570 94.820 51.830 95.140 ;
        RECT 51.630 94.120 51.770 94.820 ;
        RECT 51.570 93.800 51.830 94.120 ;
        RECT 34.090 93.460 34.350 93.780 ;
        RECT 40.530 93.460 40.790 93.780 ;
        RECT 45.130 93.460 45.390 93.780 ;
        RECT 32.980 92.925 34.520 93.295 ;
        RECT 25.410 92.760 26.010 92.840 ;
        RECT 25.410 92.700 26.070 92.760 ;
        RECT 25.810 92.440 26.070 92.700 ;
        RECT 53.470 91.740 53.610 97.540 ;
        RECT 53.930 92.760 54.070 99.240 ;
        RECT 53.870 92.440 54.130 92.760 ;
        RECT 54.390 92.080 54.530 99.920 ;
        RECT 54.790 97.880 55.050 98.200 ;
        RECT 54.850 95.480 54.990 97.880 ;
        RECT 55.770 97.520 55.910 102.300 ;
        RECT 56.170 101.960 56.430 102.280 ;
        RECT 56.230 100.920 56.370 101.960 ;
        RECT 56.170 100.600 56.430 100.920 ;
        RECT 56.630 99.920 56.890 100.240 ;
        RECT 58.470 99.920 58.730 100.240 ;
        RECT 56.690 98.200 56.830 99.920 ;
        RECT 56.630 97.880 56.890 98.200 ;
        RECT 55.710 97.200 55.970 97.520 ;
        RECT 55.250 96.180 55.510 96.500 ;
        RECT 54.790 95.160 55.050 95.480 ;
        RECT 55.310 94.800 55.450 96.180 ;
        RECT 55.770 95.140 55.910 97.200 ;
        RECT 58.530 96.840 58.670 99.920 ;
        RECT 59.390 98.900 59.650 99.220 ;
        RECT 59.450 96.840 59.590 98.900 ;
        RECT 58.470 96.520 58.730 96.840 ;
        RECT 59.390 96.520 59.650 96.840 ;
        RECT 55.710 94.820 55.970 95.140 ;
        RECT 55.250 94.480 55.510 94.800 ;
        RECT 54.330 91.760 54.590 92.080 ;
        RECT 23.050 91.420 23.310 91.740 ;
        RECT 53.410 91.420 53.670 91.740 ;
        RECT 36.280 90.205 37.820 90.575 ;
        RECT 32.980 87.485 34.520 87.855 ;
        RECT 36.280 84.765 37.820 85.135 ;
        RECT 32.980 82.045 34.520 82.415 ;
        RECT 64.050 81.880 64.190 105.360 ;
        RECT 64.510 102.280 64.650 107.740 ;
        RECT 66.750 107.400 67.010 107.720 ;
        RECT 66.290 105.590 66.550 105.680 ;
        RECT 66.810 105.590 66.950 107.400 ;
        RECT 69.050 107.060 69.310 107.380 ;
        RECT 66.290 105.450 66.950 105.590 ;
        RECT 66.290 105.360 66.550 105.450 ;
        RECT 68.590 104.680 68.850 105.000 ;
        RECT 67.210 102.980 67.470 103.300 ;
        RECT 66.750 102.640 67.010 102.960 ;
        RECT 64.450 101.960 64.710 102.280 ;
        RECT 64.510 97.180 64.650 101.960 ;
        RECT 66.810 100.920 66.950 102.640 ;
        RECT 66.750 100.600 67.010 100.920 ;
        RECT 66.750 100.150 67.010 100.240 ;
        RECT 67.270 100.150 67.410 102.980 ;
        RECT 68.650 102.620 68.790 104.680 ;
        RECT 69.110 103.640 69.250 107.060 ;
        RECT 69.570 105.680 69.710 108.760 ;
        RECT 70.030 106.360 70.170 110.800 ;
        RECT 70.890 109.780 71.150 110.100 ;
        RECT 70.950 109.080 71.090 109.780 ;
        RECT 70.890 108.760 71.150 109.080 ;
        RECT 70.430 108.080 70.690 108.400 ;
        RECT 69.970 106.040 70.230 106.360 ;
        RECT 70.490 105.680 70.630 108.080 ;
        RECT 69.510 105.360 69.770 105.680 ;
        RECT 70.430 105.360 70.690 105.680 ;
        RECT 71.410 105.340 71.550 136.980 ;
        RECT 71.870 105.930 72.010 138.090 ;
        RECT 72.330 137.300 72.470 138.940 ;
        RECT 72.790 138.660 72.930 140.720 ;
        RECT 75.030 140.040 75.290 140.360 ;
        RECT 73.650 139.700 73.910 140.020 ;
        RECT 72.730 138.340 72.990 138.660 ;
        RECT 72.270 136.980 72.530 137.300 ;
        RECT 73.710 137.040 73.850 139.700 ;
        RECT 75.090 137.980 75.230 140.040 ;
        RECT 77.390 138.320 77.530 143.440 ;
        RECT 75.950 138.000 76.210 138.320 ;
        RECT 77.330 138.000 77.590 138.320 ;
        RECT 75.030 137.660 75.290 137.980 ;
        RECT 74.110 137.040 74.370 137.300 ;
        RECT 73.710 136.980 74.370 137.040 ;
        RECT 73.710 136.900 74.310 136.980 ;
        RECT 72.270 134.260 72.530 134.580 ;
        RECT 72.330 124.040 72.470 134.260 ;
        RECT 72.270 123.720 72.530 124.040 ;
        RECT 73.710 122.680 73.850 136.900 ;
        RECT 74.110 134.940 74.370 135.260 ;
        RECT 74.170 128.120 74.310 134.940 ;
        RECT 74.110 127.800 74.370 128.120 ;
        RECT 75.030 124.060 75.290 124.380 ;
        RECT 74.110 123.720 74.370 124.040 ;
        RECT 73.650 122.360 73.910 122.680 ;
        RECT 74.170 122.000 74.310 123.720 ;
        RECT 75.090 122.000 75.230 124.060 ;
        RECT 73.190 121.680 73.450 122.000 ;
        RECT 74.110 121.680 74.370 122.000 ;
        RECT 75.030 121.680 75.290 122.000 ;
        RECT 72.270 121.000 72.530 121.320 ;
        RECT 72.330 111.460 72.470 121.000 ;
        RECT 72.730 120.660 72.990 120.980 ;
        RECT 72.790 116.900 72.930 120.660 ;
        RECT 73.250 119.960 73.390 121.680 ;
        RECT 73.190 119.640 73.450 119.960 ;
        RECT 74.170 118.600 74.310 121.680 ;
        RECT 74.110 118.280 74.370 118.600 ;
        RECT 72.730 116.580 72.990 116.900 ;
        RECT 72.730 115.220 72.990 115.540 ;
        RECT 72.790 113.840 72.930 115.220 ;
        RECT 72.730 113.520 72.990 113.840 ;
        RECT 74.170 112.820 74.310 118.280 ;
        RECT 73.650 112.500 73.910 112.820 ;
        RECT 74.110 112.500 74.370 112.820 ;
        RECT 74.570 112.500 74.830 112.820 ;
        RECT 72.270 111.140 72.530 111.460 ;
        RECT 72.330 107.720 72.470 111.140 ;
        RECT 72.730 109.955 72.990 110.100 ;
        RECT 72.720 109.585 73.000 109.955 ;
        RECT 73.710 107.720 73.850 112.500 ;
        RECT 74.110 109.780 74.370 110.100 ;
        RECT 74.170 107.800 74.310 109.780 ;
        RECT 74.630 108.400 74.770 112.500 ;
        RECT 75.490 111.480 75.750 111.800 ;
        RECT 75.550 110.100 75.690 111.480 ;
        RECT 75.490 109.780 75.750 110.100 ;
        RECT 74.570 108.080 74.830 108.400 ;
        RECT 74.170 107.720 74.770 107.800 ;
        RECT 75.030 107.740 75.290 108.060 ;
        RECT 72.270 107.400 72.530 107.720 ;
        RECT 73.650 107.400 73.910 107.720 ;
        RECT 74.170 107.660 74.830 107.720 ;
        RECT 74.570 107.400 74.830 107.660 ;
        RECT 74.110 107.060 74.370 107.380 ;
        RECT 74.170 106.020 74.310 107.060 ;
        RECT 71.870 105.790 72.470 105.930 ;
        RECT 72.330 105.340 72.470 105.790 ;
        RECT 74.110 105.700 74.370 106.020 ;
        RECT 69.960 104.825 70.240 105.195 ;
        RECT 71.350 105.020 71.610 105.340 ;
        RECT 72.270 105.020 72.530 105.340 ;
        RECT 74.110 105.195 74.370 105.340 ;
        RECT 69.970 104.680 70.230 104.825 ;
        RECT 69.050 103.320 69.310 103.640 ;
        RECT 68.590 102.300 68.850 102.620 ;
        RECT 71.410 102.280 71.550 105.020 ;
        RECT 71.810 104.340 72.070 104.660 ;
        RECT 71.870 103.640 72.010 104.340 ;
        RECT 71.810 103.320 72.070 103.640 ;
        RECT 71.350 101.960 71.610 102.280 ;
        RECT 68.590 101.620 68.850 101.940 ;
        RECT 66.750 100.010 67.410 100.150 ;
        RECT 66.750 99.920 67.010 100.010 ;
        RECT 68.650 99.900 68.790 101.620 ;
        RECT 72.330 100.580 72.470 105.020 ;
        RECT 74.100 104.825 74.380 105.195 ;
        RECT 75.090 103.640 75.230 107.740 ;
        RECT 75.550 105.680 75.690 109.780 ;
        RECT 75.490 105.360 75.750 105.680 ;
        RECT 75.030 103.320 75.290 103.640 ;
        RECT 72.270 100.260 72.530 100.580 ;
        RECT 68.590 99.580 68.850 99.900 ;
        RECT 71.810 99.580 72.070 99.900 ;
        RECT 65.830 98.900 66.090 99.220 ;
        RECT 65.890 97.180 66.030 98.900 ;
        RECT 64.450 96.860 64.710 97.180 ;
        RECT 65.830 96.860 66.090 97.180 ;
        RECT 71.870 96.500 72.010 99.580 ;
        RECT 71.810 96.180 72.070 96.500 ;
        RECT 63.990 81.560 64.250 81.880 ;
        RECT 71.870 80.860 72.010 96.180 ;
        RECT 74.570 91.420 74.830 91.740 ;
        RECT 74.630 89.020 74.770 91.420 ;
        RECT 76.010 91.060 76.150 138.000 ;
        RECT 78.770 135.600 78.910 143.440 ;
        RECT 79.630 139.700 79.890 140.020 ;
        RECT 78.710 135.280 78.970 135.600 ;
        RECT 79.690 135.260 79.830 139.700 ;
        RECT 80.150 137.980 80.290 145.480 ;
        RECT 81.930 143.440 82.190 143.760 ;
        RECT 81.470 142.420 81.730 142.740 ;
        RECT 81.530 141.040 81.670 142.420 ;
        RECT 81.470 140.720 81.730 141.040 ;
        RECT 80.090 137.660 80.350 137.980 ;
        RECT 81.990 136.280 82.130 143.440 ;
        RECT 85.670 139.000 85.810 155.000 ;
        RECT 87.970 151.920 88.110 157.720 ;
        RECT 87.910 151.600 88.170 151.920 ;
        RECT 88.370 151.600 88.630 151.920 ;
        RECT 88.430 148.180 88.570 151.600 ;
        RECT 88.370 147.860 88.630 148.180 ;
        RECT 88.430 146.480 88.570 147.860 ;
        RECT 88.890 146.480 89.030 170.640 ;
        RECT 89.350 165.180 89.490 180.500 ;
        RECT 89.810 178.780 89.950 181.180 ;
        RECT 89.750 178.460 90.010 178.780 ;
        RECT 89.290 164.860 89.550 165.180 ;
        RECT 89.810 164.240 89.950 178.460 ;
        RECT 90.270 176.400 90.410 183.900 ;
        RECT 92.050 183.220 92.310 183.540 ;
        RECT 92.110 181.840 92.250 183.220 ;
        RECT 93.030 182.520 93.170 186.620 ;
        RECT 94.410 184.560 94.550 187.300 ;
        RECT 94.350 184.240 94.610 184.560 ;
        RECT 94.870 184.220 95.010 188.660 ;
        RECT 95.270 185.940 95.530 186.260 ;
        RECT 94.810 183.900 95.070 184.220 ;
        RECT 92.970 182.200 93.230 182.520 ;
        RECT 92.050 181.520 92.310 181.840 ;
        RECT 92.510 181.520 92.770 181.840 ;
        RECT 92.570 179.120 92.710 181.520 ;
        RECT 95.330 181.500 95.470 185.940 ;
        RECT 95.790 185.240 95.930 188.660 ;
        RECT 95.730 184.920 95.990 185.240 ;
        RECT 95.270 181.180 95.530 181.500 ;
        RECT 95.330 179.120 95.470 181.180 ;
        RECT 92.510 178.800 92.770 179.120 ;
        RECT 95.270 178.800 95.530 179.120 ;
        RECT 95.790 178.440 95.930 184.920 ;
        RECT 97.110 183.220 97.370 183.540 ;
        RECT 97.170 181.500 97.310 183.220 ;
        RECT 98.030 181.920 98.290 182.180 ;
        RECT 98.030 181.860 98.690 181.920 ;
        RECT 98.090 181.780 98.690 181.860 ;
        RECT 97.110 181.180 97.370 181.500 ;
        RECT 97.170 178.780 97.310 181.180 ;
        RECT 98.550 179.460 98.690 181.780 ;
        RECT 99.870 181.180 100.130 181.500 ;
        RECT 98.490 179.140 98.750 179.460 ;
        RECT 97.110 178.460 97.370 178.780 ;
        RECT 98.030 178.460 98.290 178.780 ;
        RECT 95.730 178.120 95.990 178.440 ;
        RECT 98.090 178.100 98.230 178.460 ;
        RECT 98.030 177.780 98.290 178.100 ;
        RECT 90.210 176.080 90.470 176.400 ;
        RECT 90.270 168.240 90.410 176.080 ;
        RECT 98.550 173.340 98.690 179.140 ;
        RECT 99.930 178.780 100.070 181.180 ;
        RECT 100.390 181.160 100.530 189.430 ;
        RECT 102.630 189.340 102.890 189.660 ;
        RECT 105.390 189.340 105.650 189.660 ;
        RECT 101.250 188.660 101.510 188.980 ;
        RECT 100.790 185.940 101.050 186.260 ;
        RECT 100.850 184.220 100.990 185.940 ;
        RECT 100.790 183.900 101.050 184.220 ;
        RECT 100.330 180.840 100.590 181.160 ;
        RECT 101.310 180.820 101.450 188.660 ;
        RECT 102.690 187.620 102.830 189.340 ;
        RECT 103.550 189.000 103.810 189.320 ;
        RECT 102.630 187.300 102.890 187.620 ;
        RECT 101.710 187.190 101.970 187.280 ;
        RECT 101.710 187.050 102.370 187.190 ;
        RECT 101.710 186.960 101.970 187.050 ;
        RECT 101.710 183.220 101.970 183.540 ;
        RECT 101.770 182.180 101.910 183.220 ;
        RECT 102.230 182.520 102.370 187.050 ;
        RECT 102.170 182.200 102.430 182.520 ;
        RECT 101.710 181.860 101.970 182.180 ;
        RECT 101.250 180.500 101.510 180.820 ;
        RECT 101.310 179.800 101.450 180.500 ;
        RECT 101.250 179.480 101.510 179.800 ;
        RECT 101.770 179.100 101.910 181.860 ;
        RECT 103.610 181.840 103.750 189.000 ;
        RECT 105.450 187.190 105.590 189.340 ;
        RECT 105.450 187.050 106.970 187.190 ;
        RECT 105.390 185.940 105.650 186.260 ;
        RECT 104.930 183.560 105.190 183.880 ;
        RECT 104.990 182.180 105.130 183.560 ;
        RECT 104.930 181.860 105.190 182.180 ;
        RECT 105.450 181.840 105.590 185.940 ;
        RECT 106.830 184.220 106.970 187.050 ;
        RECT 107.690 186.960 107.950 187.280 ;
        RECT 107.750 185.240 107.890 186.960 ;
        RECT 107.690 184.920 107.950 185.240 ;
        RECT 107.690 184.240 107.950 184.560 ;
        RECT 106.770 183.900 107.030 184.220 ;
        RECT 106.830 181.840 106.970 183.900 ;
        RECT 107.230 183.220 107.490 183.540 ;
        RECT 103.550 181.520 103.810 181.840 ;
        RECT 105.390 181.520 105.650 181.840 ;
        RECT 106.770 181.520 107.030 181.840 ;
        RECT 106.830 179.800 106.970 181.520 ;
        RECT 106.770 179.480 107.030 179.800 ;
        RECT 102.170 179.100 102.430 179.120 ;
        RECT 101.770 178.960 102.430 179.100 ;
        RECT 102.170 178.800 102.430 178.960 ;
        RECT 107.290 178.780 107.430 183.220 ;
        RECT 107.750 181.840 107.890 184.240 ;
        RECT 107.690 181.520 107.950 181.840 ;
        RECT 108.210 181.750 108.350 189.680 ;
        RECT 110.450 189.340 110.710 189.660 ;
        RECT 109.990 189.000 110.250 189.320 ;
        RECT 109.070 188.660 109.330 188.980 ;
        RECT 109.130 184.220 109.270 188.660 ;
        RECT 110.050 185.240 110.190 189.000 ;
        RECT 109.990 184.920 110.250 185.240 ;
        RECT 109.070 183.900 109.330 184.220 ;
        RECT 110.050 182.180 110.190 184.920 ;
        RECT 110.510 184.900 110.650 189.340 ;
        RECT 117.350 189.000 117.610 189.320 ;
        RECT 112.750 188.660 113.010 188.980 ;
        RECT 110.450 184.580 110.710 184.900 ;
        RECT 109.990 181.860 110.250 182.180 ;
        RECT 108.610 181.750 108.870 181.840 ;
        RECT 108.210 181.610 108.870 181.750 ;
        RECT 108.610 181.520 108.870 181.610 ;
        RECT 109.070 181.180 109.330 181.500 ;
        RECT 107.690 180.500 107.950 180.820 ;
        RECT 99.870 178.460 100.130 178.780 ;
        RECT 107.230 178.460 107.490 178.780 ;
        RECT 107.290 173.680 107.430 178.460 ;
        RECT 107.750 175.380 107.890 180.500 ;
        RECT 108.610 179.480 108.870 179.800 ;
        RECT 108.670 179.100 108.810 179.480 ;
        RECT 109.130 179.460 109.270 181.180 ;
        RECT 109.530 180.500 109.790 180.820 ;
        RECT 109.070 179.140 109.330 179.460 ;
        RECT 108.210 178.960 108.810 179.100 ;
        RECT 107.690 175.060 107.950 175.380 ;
        RECT 98.950 173.360 99.210 173.680 ;
        RECT 107.230 173.360 107.490 173.680 ;
        RECT 98.490 173.020 98.750 173.340 ;
        RECT 95.270 172.340 95.530 172.660 ;
        RECT 90.210 167.920 90.470 168.240 ;
        RECT 90.270 165.180 90.410 167.920 ;
        RECT 95.330 167.900 95.470 172.340 ;
        RECT 99.010 171.640 99.150 173.360 ;
        RECT 99.410 173.020 99.670 173.340 ;
        RECT 98.950 171.320 99.210 171.640 ;
        RECT 98.490 170.640 98.750 170.960 ;
        RECT 97.570 168.600 97.830 168.920 ;
        RECT 95.270 167.580 95.530 167.900 ;
        RECT 95.270 165.200 95.530 165.520 ;
        RECT 90.210 164.860 90.470 165.180 ;
        RECT 89.350 164.100 89.950 164.240 ;
        RECT 89.350 159.480 89.490 164.100 ;
        RECT 89.750 161.460 90.010 161.780 ;
        RECT 89.810 160.420 89.950 161.460 ;
        RECT 89.750 160.100 90.010 160.420 ;
        RECT 90.270 159.990 90.410 164.860 ;
        RECT 95.330 163.480 95.470 165.200 ;
        RECT 95.270 163.160 95.530 163.480 ;
        RECT 97.630 162.800 97.770 168.600 ;
        RECT 98.030 165.200 98.290 165.520 ;
        RECT 97.570 162.480 97.830 162.800 ;
        RECT 96.190 162.140 96.450 162.460 ;
        RECT 92.050 161.460 92.310 161.780 ;
        RECT 90.670 159.990 90.930 160.080 ;
        RECT 90.270 159.850 90.930 159.990 ;
        RECT 90.670 159.760 90.930 159.850 ;
        RECT 89.350 159.340 89.950 159.480 ;
        RECT 89.290 156.700 89.550 157.020 ;
        RECT 89.350 154.640 89.490 156.700 ;
        RECT 89.290 154.320 89.550 154.640 ;
        RECT 88.370 146.160 88.630 146.480 ;
        RECT 88.830 146.160 89.090 146.480 ;
        RECT 86.070 145.140 86.330 145.460 ;
        RECT 86.130 142.740 86.270 145.140 ;
        RECT 87.910 143.100 88.170 143.420 ;
        RECT 88.890 143.160 89.030 146.160 ;
        RECT 86.070 142.420 86.330 142.740 ;
        RECT 87.970 140.360 88.110 143.100 ;
        RECT 88.430 143.020 89.030 143.160 ;
        RECT 89.810 143.080 89.950 159.340 ;
        RECT 91.590 156.020 91.850 156.340 ;
        RECT 91.650 152.600 91.790 156.020 ;
        RECT 92.110 154.640 92.250 161.460 ;
        RECT 96.250 159.060 96.390 162.140 ;
        RECT 97.570 161.460 97.830 161.780 ;
        RECT 96.190 158.740 96.450 159.060 ;
        RECT 92.510 157.040 92.770 157.360 ;
        RECT 92.050 154.320 92.310 154.640 ;
        RECT 92.570 154.300 92.710 157.040 ;
        RECT 94.810 156.700 95.070 157.020 ;
        RECT 94.870 155.320 95.010 156.700 ;
        RECT 94.810 155.000 95.070 155.320 ;
        RECT 92.510 153.980 92.770 154.300 ;
        RECT 91.590 152.280 91.850 152.600 ;
        RECT 96.250 151.920 96.390 158.740 ;
        RECT 96.650 154.660 96.910 154.980 ;
        RECT 96.710 151.920 96.850 154.660 ;
        RECT 96.190 151.600 96.450 151.920 ;
        RECT 96.650 151.600 96.910 151.920 ;
        RECT 91.130 150.580 91.390 150.900 ;
        RECT 90.670 143.780 90.930 144.100 ;
        RECT 87.910 140.040 88.170 140.360 ;
        RECT 88.430 140.020 88.570 143.020 ;
        RECT 89.750 142.760 90.010 143.080 ;
        RECT 88.830 142.420 89.090 142.740 ;
        RECT 88.890 140.020 89.030 142.420 ;
        RECT 90.210 140.380 90.470 140.700 ;
        RECT 88.370 139.700 88.630 140.020 ;
        RECT 88.830 139.700 89.090 140.020 ;
        RECT 85.610 138.680 85.870 139.000 ;
        RECT 81.930 135.960 82.190 136.280 ;
        RECT 79.630 134.940 79.890 135.260 ;
        RECT 76.870 134.600 77.130 134.920 ;
        RECT 83.310 134.600 83.570 134.920 ;
        RECT 76.410 132.560 76.670 132.880 ;
        RECT 76.470 125.400 76.610 132.560 ;
        RECT 76.930 127.440 77.070 134.600 ;
        RECT 78.250 131.540 78.510 131.860 ;
        RECT 77.330 129.840 77.590 130.160 ;
        RECT 77.390 128.120 77.530 129.840 ;
        RECT 77.330 127.800 77.590 128.120 ;
        RECT 76.870 127.120 77.130 127.440 ;
        RECT 76.410 125.080 76.670 125.400 ;
        RECT 77.390 125.060 77.530 127.800 ;
        RECT 78.310 127.440 78.450 131.540 ;
        RECT 78.710 129.500 78.970 129.820 ;
        RECT 78.250 127.120 78.510 127.440 ;
        RECT 77.790 126.440 78.050 126.760 ;
        RECT 77.330 124.740 77.590 125.060 ;
        RECT 77.850 124.380 77.990 126.440 ;
        RECT 78.310 124.720 78.450 127.120 ;
        RECT 78.250 124.400 78.510 124.720 ;
        RECT 77.790 124.060 78.050 124.380 ;
        RECT 78.770 124.120 78.910 129.500 ;
        RECT 82.850 128.820 83.110 129.140 ;
        RECT 80.090 127.460 80.350 127.780 ;
        RECT 80.150 124.380 80.290 127.460 ;
        RECT 81.470 127.120 81.730 127.440 ;
        RECT 77.850 122.680 77.990 124.060 ;
        RECT 78.310 123.980 78.910 124.120 ;
        RECT 80.090 124.060 80.350 124.380 ;
        RECT 77.790 122.360 78.050 122.680 ;
        RECT 76.410 115.220 76.670 115.540 ;
        RECT 76.470 114.520 76.610 115.220 ;
        RECT 76.410 114.200 76.670 114.520 ;
        RECT 78.310 113.240 78.450 123.980 ;
        RECT 80.550 121.340 80.810 121.660 ;
        RECT 80.610 118.940 80.750 121.340 ;
        RECT 78.710 118.620 78.970 118.940 ;
        RECT 80.550 118.850 80.810 118.940 ;
        RECT 80.150 118.710 80.810 118.850 ;
        RECT 77.850 113.100 78.450 113.240 ;
        RECT 77.850 94.800 77.990 113.100 ;
        RECT 78.250 112.500 78.510 112.820 ;
        RECT 78.310 111.120 78.450 112.500 ;
        RECT 78.250 110.800 78.510 111.120 ;
        RECT 78.310 108.400 78.450 110.800 ;
        RECT 78.770 110.440 78.910 118.620 ;
        RECT 79.170 117.940 79.430 118.260 ;
        RECT 78.710 110.120 78.970 110.440 ;
        RECT 79.230 108.400 79.370 117.940 ;
        RECT 80.150 114.520 80.290 118.710 ;
        RECT 80.550 118.620 80.810 118.710 ;
        RECT 80.550 115.220 80.810 115.540 ;
        RECT 80.090 114.200 80.350 114.520 ;
        RECT 80.090 113.180 80.350 113.500 ;
        RECT 79.630 112.840 79.890 113.160 ;
        RECT 79.690 111.120 79.830 112.840 ;
        RECT 79.630 110.800 79.890 111.120 ;
        RECT 80.150 110.780 80.290 113.180 ;
        RECT 80.610 110.780 80.750 115.220 ;
        RECT 81.010 113.180 81.270 113.500 ;
        RECT 81.070 111.800 81.210 113.180 ;
        RECT 81.010 111.480 81.270 111.800 ;
        RECT 80.090 110.460 80.350 110.780 ;
        RECT 80.550 110.460 80.810 110.780 ;
        RECT 78.250 108.080 78.510 108.400 ;
        RECT 79.170 108.080 79.430 108.400 ;
        RECT 79.230 105.340 79.370 108.080 ;
        RECT 81.530 107.290 81.670 127.120 ;
        RECT 82.910 127.100 83.050 128.820 ;
        RECT 82.850 126.780 83.110 127.100 ;
        RECT 82.850 126.100 83.110 126.420 ;
        RECT 82.910 125.400 83.050 126.100 ;
        RECT 82.850 125.080 83.110 125.400 ;
        RECT 82.910 119.960 83.050 125.080 ;
        RECT 82.850 119.640 83.110 119.960 ;
        RECT 82.390 115.220 82.650 115.540 ;
        RECT 82.450 111.120 82.590 115.220 ;
        RECT 82.850 111.140 83.110 111.460 ;
        RECT 82.390 110.800 82.650 111.120 ;
        RECT 82.910 108.060 83.050 111.140 ;
        RECT 82.850 107.740 83.110 108.060 ;
        RECT 81.530 107.150 82.130 107.290 ;
        RECT 79.170 105.020 79.430 105.340 ;
        RECT 81.010 102.300 81.270 102.620 ;
        RECT 81.070 97.860 81.210 102.300 ;
        RECT 81.470 98.900 81.730 99.220 ;
        RECT 81.010 97.540 81.270 97.860 ;
        RECT 81.010 96.520 81.270 96.840 ;
        RECT 77.790 94.480 78.050 94.800 ;
        RECT 78.250 93.460 78.510 93.780 ;
        RECT 78.310 91.740 78.450 93.460 ;
        RECT 81.070 92.760 81.210 96.520 ;
        RECT 81.010 92.440 81.270 92.760 ;
        RECT 78.250 91.420 78.510 91.740 ;
        RECT 75.950 90.740 76.210 91.060 ;
        RECT 74.570 88.700 74.830 89.020 ;
        RECT 76.010 82.500 76.150 90.740 ;
        RECT 81.070 88.340 81.210 92.440 ;
        RECT 80.550 88.020 80.810 88.340 ;
        RECT 81.010 88.020 81.270 88.340 ;
        RECT 80.610 86.300 80.750 88.020 ;
        RECT 80.550 85.980 80.810 86.300 ;
        RECT 80.610 83.920 80.750 85.980 ;
        RECT 80.550 83.600 80.810 83.920 ;
        RECT 75.090 82.360 76.150 82.500 ;
        RECT 75.090 81.200 75.230 82.360 ;
        RECT 75.030 80.880 75.290 81.200 ;
        RECT 81.070 80.860 81.210 88.020 ;
        RECT 81.530 80.860 81.670 98.900 ;
        RECT 81.990 97.520 82.130 107.150 ;
        RECT 83.370 103.640 83.510 134.600 ;
        RECT 85.670 130.800 85.810 138.680 ;
        RECT 87.440 138.145 87.720 138.515 ;
        RECT 88.830 138.340 89.090 138.660 ;
        RECT 90.270 138.515 90.410 140.380 ;
        RECT 87.450 138.000 87.710 138.145 ;
        RECT 88.890 136.280 89.030 138.340 ;
        RECT 90.200 138.145 90.480 138.515 ;
        RECT 88.830 135.960 89.090 136.280 ;
        RECT 88.370 134.600 88.630 134.920 ;
        RECT 85.210 130.660 85.810 130.800 ;
        RECT 84.690 129.160 84.950 129.480 ;
        RECT 84.230 128.820 84.490 129.140 ;
        RECT 84.290 127.440 84.430 128.820 ;
        RECT 84.750 128.120 84.890 129.160 ;
        RECT 84.690 127.800 84.950 128.120 ;
        RECT 84.230 127.120 84.490 127.440 ;
        RECT 84.690 123.720 84.950 124.040 ;
        RECT 84.750 122.000 84.890 123.720 ;
        RECT 85.210 122.340 85.350 130.660 ;
        RECT 85.610 129.500 85.870 129.820 ;
        RECT 86.070 129.500 86.330 129.820 ;
        RECT 85.670 127.440 85.810 129.500 ;
        RECT 85.610 127.120 85.870 127.440 ;
        RECT 85.670 124.720 85.810 127.120 ;
        RECT 86.130 125.400 86.270 129.500 ;
        RECT 86.070 125.080 86.330 125.400 ;
        RECT 86.530 124.800 86.790 125.060 ;
        RECT 86.130 124.740 86.790 124.800 ;
        RECT 85.610 124.400 85.870 124.720 ;
        RECT 86.130 124.660 86.730 124.740 ;
        RECT 85.150 122.020 85.410 122.340 ;
        RECT 84.690 121.680 84.950 122.000 ;
        RECT 84.750 119.960 84.890 121.680 ;
        RECT 84.690 119.640 84.950 119.960 ;
        RECT 84.750 118.940 84.890 119.640 ;
        RECT 84.690 118.620 84.950 118.940 ;
        RECT 85.150 117.940 85.410 118.260 ;
        RECT 85.210 116.220 85.350 117.940 ;
        RECT 85.670 116.560 85.810 124.400 ;
        RECT 86.130 122.000 86.270 124.660 ;
        RECT 86.530 123.380 86.790 123.700 ;
        RECT 86.590 122.680 86.730 123.380 ;
        RECT 86.530 122.360 86.790 122.680 ;
        RECT 86.070 121.680 86.330 122.000 ;
        RECT 87.910 118.280 88.170 118.600 ;
        RECT 87.450 116.810 87.710 116.900 ;
        RECT 87.970 116.810 88.110 118.280 ;
        RECT 87.450 116.670 88.110 116.810 ;
        RECT 87.450 116.580 87.710 116.670 ;
        RECT 85.610 116.240 85.870 116.560 ;
        RECT 84.690 115.900 84.950 116.220 ;
        RECT 85.150 115.900 85.410 116.220 ;
        RECT 84.750 111.120 84.890 115.900 ;
        RECT 85.670 113.840 85.810 116.240 ;
        RECT 85.610 113.520 85.870 113.840 ;
        RECT 85.670 111.460 85.810 113.520 ;
        RECT 85.610 111.140 85.870 111.460 ;
        RECT 84.690 111.030 84.950 111.120 ;
        RECT 83.830 110.890 84.950 111.030 ;
        RECT 83.310 103.320 83.570 103.640 ;
        RECT 83.310 101.960 83.570 102.280 ;
        RECT 82.850 100.600 83.110 100.920 ;
        RECT 82.390 99.920 82.650 100.240 ;
        RECT 82.450 98.200 82.590 99.920 ;
        RECT 82.390 97.880 82.650 98.200 ;
        RECT 82.910 97.860 83.050 100.600 ;
        RECT 83.370 99.220 83.510 101.960 ;
        RECT 83.310 98.900 83.570 99.220 ;
        RECT 82.850 97.540 83.110 97.860 ;
        RECT 81.930 97.200 82.190 97.520 ;
        RECT 82.390 96.520 82.650 96.840 ;
        RECT 82.450 94.800 82.590 96.520 ;
        RECT 82.390 94.480 82.650 94.800 ;
        RECT 82.450 94.200 82.590 94.480 ;
        RECT 81.990 94.060 82.590 94.200 ;
        RECT 82.910 94.120 83.050 97.540 ;
        RECT 81.990 91.060 82.130 94.060 ;
        RECT 82.850 93.800 83.110 94.120 ;
        RECT 83.830 91.740 83.970 110.890 ;
        RECT 84.690 110.800 84.950 110.890 ;
        RECT 87.970 109.080 88.110 116.670 ;
        RECT 87.910 108.760 88.170 109.080 ;
        RECT 85.150 102.300 85.410 102.620 ;
        RECT 87.450 102.300 87.710 102.620 ;
        RECT 84.690 101.620 84.950 101.940 ;
        RECT 84.230 99.240 84.490 99.560 ;
        RECT 84.290 97.180 84.430 99.240 ;
        RECT 84.750 97.180 84.890 101.620 ;
        RECT 84.230 96.860 84.490 97.180 ;
        RECT 84.690 96.860 84.950 97.180 ;
        RECT 84.290 95.480 84.430 96.860 ;
        RECT 84.690 96.180 84.950 96.500 ;
        RECT 84.230 95.160 84.490 95.480 ;
        RECT 84.290 91.740 84.430 95.160 ;
        RECT 84.750 91.740 84.890 96.180 ;
        RECT 85.210 95.140 85.350 102.300 ;
        RECT 85.610 99.580 85.870 99.900 ;
        RECT 85.670 97.860 85.810 99.580 ;
        RECT 85.610 97.540 85.870 97.860 ;
        RECT 85.670 97.180 85.810 97.540 ;
        RECT 87.510 97.180 87.650 102.300 ;
        RECT 88.430 98.200 88.570 134.600 ;
        RECT 89.750 128.820 90.010 129.140 ;
        RECT 89.810 127.440 89.950 128.820 ;
        RECT 89.750 127.120 90.010 127.440 ;
        RECT 90.210 126.100 90.470 126.420 ;
        RECT 88.830 123.720 89.090 124.040 ;
        RECT 88.890 122.680 89.030 123.720 ;
        RECT 88.830 122.360 89.090 122.680 ;
        RECT 90.270 121.660 90.410 126.100 ;
        RECT 90.210 121.340 90.470 121.660 ;
        RECT 90.270 118.600 90.410 121.340 ;
        RECT 90.210 118.280 90.470 118.600 ;
        RECT 88.830 117.940 89.090 118.260 ;
        RECT 88.890 116.900 89.030 117.940 ;
        RECT 88.830 116.580 89.090 116.900 ;
        RECT 89.750 107.400 90.010 107.720 ;
        RECT 89.810 106.020 89.950 107.400 ;
        RECT 89.750 105.700 90.010 106.020 ;
        RECT 88.830 105.360 89.090 105.680 ;
        RECT 88.890 100.920 89.030 105.360 ;
        RECT 89.290 102.300 89.550 102.620 ;
        RECT 88.830 100.600 89.090 100.920 ;
        RECT 89.350 100.580 89.490 102.300 ;
        RECT 89.810 102.280 89.950 105.700 ;
        RECT 89.750 101.960 90.010 102.280 ;
        RECT 89.290 100.260 89.550 100.580 ;
        RECT 89.810 100.240 89.950 101.960 ;
        RECT 89.750 99.920 90.010 100.240 ;
        RECT 88.370 97.880 88.630 98.200 ;
        RECT 88.820 97.345 89.100 97.715 ;
        RECT 89.810 97.520 89.950 99.920 ;
        RECT 88.890 97.180 89.030 97.345 ;
        RECT 89.750 97.200 90.010 97.520 ;
        RECT 85.610 96.860 85.870 97.180 ;
        RECT 87.450 96.860 87.710 97.180 ;
        RECT 88.830 96.860 89.090 97.180 ;
        RECT 85.150 94.820 85.410 95.140 ;
        RECT 85.150 94.140 85.410 94.460 ;
        RECT 85.210 92.760 85.350 94.140 ;
        RECT 85.670 92.760 85.810 96.860 ;
        RECT 87.510 94.800 87.650 96.860 ;
        RECT 88.820 95.985 89.100 96.355 ;
        RECT 87.450 94.480 87.710 94.800 ;
        RECT 88.890 93.780 89.030 95.985 ;
        RECT 89.290 94.480 89.550 94.800 ;
        RECT 88.830 93.460 89.090 93.780 ;
        RECT 85.150 92.440 85.410 92.760 ;
        RECT 85.610 92.440 85.870 92.760 ;
        RECT 85.670 91.740 85.810 92.440 ;
        RECT 83.770 91.420 84.030 91.740 ;
        RECT 84.230 91.420 84.490 91.740 ;
        RECT 84.690 91.420 84.950 91.740 ;
        RECT 85.610 91.420 85.870 91.740 ;
        RECT 81.930 90.740 82.190 91.060 ;
        RECT 82.390 90.740 82.650 91.060 ;
        RECT 81.990 80.860 82.130 90.740 ;
        RECT 82.450 89.360 82.590 90.740 ;
        RECT 83.830 89.360 83.970 91.420 ;
        RECT 85.670 90.040 85.810 91.420 ;
        RECT 85.610 89.720 85.870 90.040 ;
        RECT 88.890 89.360 89.030 93.460 ;
        RECT 89.350 92.760 89.490 94.480 ;
        RECT 89.290 92.440 89.550 92.760 ;
        RECT 89.810 92.160 89.950 97.200 ;
        RECT 90.210 96.860 90.470 97.180 ;
        RECT 89.350 92.020 89.950 92.160 ;
        RECT 82.390 89.040 82.650 89.360 ;
        RECT 83.770 89.040 84.030 89.360 ;
        RECT 88.830 89.040 89.090 89.360 ;
        RECT 88.370 88.700 88.630 89.020 ;
        RECT 83.770 88.020 84.030 88.340 ;
        RECT 87.450 88.020 87.710 88.340 ;
        RECT 83.830 85.960 83.970 88.020 ;
        RECT 83.770 85.640 84.030 85.960 ;
        RECT 87.510 84.260 87.650 88.020 ;
        RECT 88.430 84.260 88.570 88.700 ;
        RECT 89.350 86.300 89.490 92.020 ;
        RECT 89.750 89.040 90.010 89.360 ;
        RECT 89.290 85.980 89.550 86.300 ;
        RECT 89.810 84.600 89.950 89.040 ;
        RECT 90.270 88.680 90.410 96.860 ;
        RECT 90.730 94.800 90.870 143.780 ;
        RECT 91.190 139.000 91.330 150.580 ;
        RECT 96.710 149.200 96.850 151.600 ;
        RECT 96.650 148.880 96.910 149.200 ;
        RECT 91.590 145.140 91.850 145.460 ;
        RECT 91.650 144.440 91.790 145.140 ;
        RECT 91.590 144.120 91.850 144.440 ;
        RECT 95.730 143.100 95.990 143.420 ;
        RECT 95.270 142.420 95.530 142.740 ;
        RECT 95.330 140.360 95.470 142.420 ;
        RECT 95.270 140.040 95.530 140.360 ;
        RECT 91.130 138.680 91.390 139.000 ;
        RECT 92.970 138.680 93.230 139.000 ;
        RECT 93.030 135.600 93.170 138.680 ;
        RECT 92.970 135.280 93.230 135.600 ;
        RECT 92.050 128.820 92.310 129.140 ;
        RECT 94.810 128.820 95.070 129.140 ;
        RECT 92.110 126.420 92.250 128.820 ;
        RECT 94.870 126.420 95.010 128.820 ;
        RECT 92.050 126.100 92.310 126.420 ;
        RECT 94.810 126.100 95.070 126.420 ;
        RECT 91.590 123.380 91.850 123.700 ;
        RECT 91.650 121.660 91.790 123.380 ;
        RECT 94.350 122.360 94.610 122.680 ;
        RECT 91.590 121.340 91.850 121.660 ;
        RECT 93.890 120.660 94.150 120.980 ;
        RECT 93.950 116.900 94.090 120.660 ;
        RECT 94.410 118.260 94.550 122.360 ;
        RECT 95.270 122.020 95.530 122.340 ;
        RECT 94.350 117.940 94.610 118.260 ;
        RECT 93.890 116.580 94.150 116.900 ;
        RECT 94.410 116.220 94.550 117.940 ;
        RECT 94.350 115.960 94.610 116.220 ;
        RECT 93.950 115.900 94.610 115.960 ;
        RECT 93.950 115.820 94.550 115.900 ;
        RECT 91.130 107.060 91.390 107.380 ;
        RECT 91.190 100.240 91.330 107.060 ;
        RECT 92.510 103.320 92.770 103.640 ;
        RECT 91.590 101.620 91.850 101.940 ;
        RECT 92.050 101.620 92.310 101.940 ;
        RECT 91.650 100.920 91.790 101.620 ;
        RECT 91.590 100.600 91.850 100.920 ;
        RECT 92.110 100.240 92.250 101.620 ;
        RECT 91.130 99.920 91.390 100.240 ;
        RECT 91.590 99.920 91.850 100.240 ;
        RECT 92.050 99.920 92.310 100.240 ;
        RECT 91.190 98.200 91.330 99.920 ;
        RECT 91.650 99.220 91.790 99.920 ;
        RECT 91.590 98.900 91.850 99.220 ;
        RECT 91.130 97.880 91.390 98.200 ;
        RECT 91.130 96.520 91.390 96.840 ;
        RECT 91.190 95.480 91.330 96.520 ;
        RECT 92.570 96.500 92.710 103.320 ;
        RECT 93.950 100.320 94.090 115.820 ;
        RECT 94.810 115.560 95.070 115.880 ;
        RECT 94.350 115.220 94.610 115.540 ;
        RECT 94.410 113.500 94.550 115.220 ;
        RECT 94.870 114.520 95.010 115.560 ;
        RECT 94.810 114.200 95.070 114.520 ;
        RECT 94.350 113.180 94.610 113.500 ;
        RECT 95.330 111.120 95.470 122.020 ;
        RECT 95.270 110.800 95.530 111.120 ;
        RECT 94.810 107.060 95.070 107.380 ;
        RECT 94.870 106.360 95.010 107.060 ;
        RECT 94.810 106.040 95.070 106.360 ;
        RECT 95.330 105.875 95.470 110.800 ;
        RECT 95.790 106.360 95.930 143.100 ;
        RECT 96.710 140.700 96.850 148.880 ;
        RECT 97.630 144.100 97.770 161.460 ;
        RECT 98.090 157.700 98.230 165.200 ;
        RECT 98.550 162.800 98.690 170.640 ;
        RECT 99.470 168.920 99.610 173.020 ;
        RECT 107.750 173.000 107.890 175.060 ;
        RECT 107.690 172.680 107.950 173.000 ;
        RECT 105.390 172.340 105.650 172.660 ;
        RECT 105.450 170.960 105.590 172.340 ;
        RECT 105.390 170.640 105.650 170.960 ;
        RECT 102.170 170.300 102.430 170.620 ;
        RECT 99.410 168.600 99.670 168.920 ;
        RECT 102.230 167.900 102.370 170.300 ;
        RECT 107.230 167.920 107.490 168.240 ;
        RECT 102.170 167.580 102.430 167.900 ;
        RECT 102.230 165.180 102.370 167.580 ;
        RECT 103.550 166.900 103.810 167.220 ;
        RECT 102.170 164.860 102.430 165.180 ;
        RECT 98.490 162.480 98.750 162.800 ;
        RECT 98.030 157.380 98.290 157.700 ;
        RECT 98.550 157.020 98.690 162.480 ;
        RECT 101.250 161.800 101.510 162.120 ;
        RECT 101.310 158.040 101.450 161.800 ;
        RECT 102.230 159.990 102.370 164.860 ;
        RECT 102.630 159.990 102.890 160.080 ;
        RECT 102.230 159.850 102.890 159.990 ;
        RECT 102.630 159.760 102.890 159.850 ;
        RECT 101.250 157.720 101.510 158.040 ;
        RECT 103.610 157.360 103.750 166.900 ;
        RECT 107.290 166.200 107.430 167.920 ;
        RECT 107.230 165.880 107.490 166.200 ;
        RECT 104.930 161.460 105.190 161.780 ;
        RECT 104.990 160.080 105.130 161.460 ;
        RECT 107.290 160.080 107.430 165.880 ;
        RECT 104.930 159.760 105.190 160.080 ;
        RECT 107.230 159.760 107.490 160.080 ;
        RECT 103.550 157.040 103.810 157.360 ;
        RECT 98.490 156.700 98.750 157.020 ;
        RECT 101.250 156.700 101.510 157.020 ;
        RECT 99.870 156.360 100.130 156.680 ;
        RECT 99.930 154.980 100.070 156.360 ;
        RECT 99.870 154.660 100.130 154.980 ;
        RECT 101.310 154.640 101.450 156.700 ;
        RECT 103.090 156.020 103.350 156.340 ;
        RECT 101.250 154.320 101.510 154.640 ;
        RECT 101.310 148.180 101.450 154.320 ;
        RECT 101.250 147.860 101.510 148.180 ;
        RECT 101.310 146.560 101.450 147.860 ;
        RECT 101.310 146.480 101.910 146.560 ;
        RECT 101.310 146.420 101.970 146.480 ;
        RECT 101.710 146.160 101.970 146.420 ;
        RECT 97.570 143.780 97.830 144.100 ;
        RECT 97.630 141.380 97.770 143.780 ;
        RECT 98.490 142.760 98.750 143.080 ;
        RECT 98.550 141.720 98.690 142.760 ;
        RECT 98.490 141.400 98.750 141.720 ;
        RECT 97.570 141.060 97.830 141.380 ;
        RECT 96.650 140.380 96.910 140.700 ;
        RECT 96.710 138.320 96.850 140.380 ;
        RECT 96.190 138.000 96.450 138.320 ;
        RECT 96.650 138.000 96.910 138.320 ;
        RECT 96.250 130.160 96.390 138.000 ;
        RECT 96.710 135.600 96.850 138.000 ;
        RECT 103.150 136.280 103.290 156.020 ;
        RECT 104.010 154.660 104.270 154.980 ;
        RECT 103.550 153.980 103.810 154.300 ;
        RECT 103.610 151.920 103.750 153.980 ;
        RECT 103.550 151.600 103.810 151.920 ;
        RECT 103.610 149.880 103.750 151.600 ;
        RECT 103.550 149.560 103.810 149.880 ;
        RECT 103.550 137.320 103.810 137.640 ;
        RECT 103.090 135.960 103.350 136.280 ;
        RECT 103.610 135.680 103.750 137.320 ;
        RECT 96.650 135.280 96.910 135.600 ;
        RECT 103.150 135.540 103.750 135.680 ;
        RECT 103.150 135.260 103.290 135.540 ;
        RECT 103.090 134.940 103.350 135.260 ;
        RECT 101.250 134.600 101.510 134.920 ;
        RECT 101.310 133.560 101.450 134.600 ;
        RECT 101.250 133.240 101.510 133.560 ;
        RECT 103.150 132.540 103.290 134.940 ;
        RECT 103.090 132.220 103.350 132.540 ;
        RECT 96.190 129.840 96.450 130.160 ;
        RECT 98.490 128.820 98.750 129.140 ;
        RECT 100.790 128.820 101.050 129.140 ;
        RECT 98.550 127.780 98.690 128.820 ;
        RECT 98.490 127.460 98.750 127.780 ;
        RECT 97.110 127.120 97.370 127.440 ;
        RECT 97.170 124.720 97.310 127.120 ;
        RECT 98.950 126.160 99.210 126.420 ;
        RECT 98.950 126.100 99.610 126.160 ;
        RECT 99.010 126.020 99.610 126.100 ;
        RECT 97.110 124.400 97.370 124.720 ;
        RECT 98.950 123.720 99.210 124.040 ;
        RECT 97.570 123.380 97.830 123.700 ;
        RECT 97.630 122.000 97.770 123.380 ;
        RECT 97.570 121.680 97.830 122.000 ;
        RECT 96.190 110.800 96.450 111.120 ;
        RECT 95.730 106.040 95.990 106.360 ;
        RECT 95.260 105.505 95.540 105.875 ;
        RECT 96.250 105.680 96.390 110.800 ;
        RECT 97.110 108.080 97.370 108.400 ;
        RECT 95.330 102.620 95.470 105.505 ;
        RECT 96.190 105.360 96.450 105.680 ;
        RECT 96.650 105.360 96.910 105.680 ;
        RECT 96.250 102.960 96.390 105.360 ;
        RECT 96.710 104.660 96.850 105.360 ;
        RECT 96.650 104.340 96.910 104.660 ;
        RECT 96.190 102.640 96.450 102.960 ;
        RECT 95.270 102.300 95.530 102.620 ;
        RECT 96.190 102.190 96.450 102.280 ;
        RECT 96.710 102.190 96.850 104.340 ;
        RECT 96.190 102.050 96.850 102.190 ;
        RECT 96.190 101.960 96.450 102.050 ;
        RECT 93.950 100.180 94.550 100.320 ;
        RECT 93.890 99.580 94.150 99.900 ;
        RECT 92.970 99.240 93.230 99.560 ;
        RECT 92.510 96.180 92.770 96.500 ;
        RECT 91.130 95.160 91.390 95.480 ;
        RECT 92.570 95.390 92.710 96.180 ;
        RECT 92.110 95.250 92.710 95.390 ;
        RECT 92.110 94.800 92.250 95.250 ;
        RECT 90.670 94.480 90.930 94.800 ;
        RECT 92.050 94.480 92.310 94.800 ;
        RECT 91.130 94.140 91.390 94.460 ;
        RECT 91.190 89.360 91.330 94.140 ;
        RECT 92.050 91.420 92.310 91.740 ;
        RECT 92.110 89.360 92.250 91.420 ;
        RECT 93.030 91.400 93.170 99.240 ;
        RECT 93.950 94.800 94.090 99.580 ;
        RECT 93.890 94.480 94.150 94.800 ;
        RECT 92.510 91.080 92.770 91.400 ;
        RECT 92.970 91.080 93.230 91.400 ;
        RECT 91.130 89.040 91.390 89.360 ;
        RECT 92.050 89.040 92.310 89.360 ;
        RECT 91.590 88.700 91.850 89.020 ;
        RECT 90.210 88.360 90.470 88.680 ;
        RECT 89.750 84.280 90.010 84.600 ;
        RECT 87.450 83.940 87.710 84.260 ;
        RECT 88.370 83.940 88.630 84.260 ;
        RECT 91.650 83.580 91.790 88.700 ;
        RECT 92.570 87.320 92.710 91.080 ;
        RECT 93.030 89.360 93.170 91.080 ;
        RECT 92.970 89.040 93.230 89.360 ;
        RECT 93.890 89.040 94.150 89.360 ;
        RECT 93.950 87.400 94.090 89.040 ;
        RECT 94.410 88.340 94.550 100.180 ;
        RECT 95.730 99.920 95.990 100.240 ;
        RECT 95.790 97.520 95.930 99.920 ;
        RECT 95.730 97.200 95.990 97.520 ;
        RECT 95.790 92.080 95.930 97.200 ;
        RECT 95.730 91.760 95.990 92.080 ;
        RECT 95.730 89.380 95.990 89.700 ;
        RECT 94.810 88.360 95.070 88.680 ;
        RECT 94.350 88.020 94.610 88.340 ;
        RECT 93.950 87.320 94.550 87.400 ;
        RECT 92.510 87.000 92.770 87.320 ;
        RECT 93.950 87.260 94.610 87.320 ;
        RECT 94.350 87.000 94.610 87.260 ;
        RECT 92.570 84.260 92.710 87.000 ;
        RECT 94.870 84.260 95.010 88.360 ;
        RECT 95.270 85.640 95.530 85.960 ;
        RECT 95.330 84.600 95.470 85.640 ;
        RECT 95.790 84.600 95.930 89.380 ;
        RECT 95.270 84.280 95.530 84.600 ;
        RECT 95.730 84.280 95.990 84.600 ;
        RECT 92.510 83.940 92.770 84.260 ;
        RECT 94.810 83.940 95.070 84.260 ;
        RECT 91.590 83.260 91.850 83.580 ;
        RECT 87.910 82.920 88.170 83.240 ;
        RECT 87.970 80.860 88.110 82.920 ;
        RECT 92.570 80.860 92.710 83.940 ;
        RECT 96.250 80.860 96.390 101.960 ;
        RECT 97.170 100.240 97.310 108.080 ;
        RECT 96.650 99.920 96.910 100.240 ;
        RECT 97.110 99.920 97.370 100.240 ;
        RECT 96.710 97.860 96.850 99.920 ;
        RECT 96.650 97.540 96.910 97.860 ;
        RECT 97.110 96.180 97.370 96.500 ;
        RECT 97.170 95.140 97.310 96.180 ;
        RECT 97.110 94.820 97.370 95.140 ;
        RECT 97.110 90.740 97.370 91.060 ;
        RECT 96.650 89.040 96.910 89.360 ;
        RECT 96.710 85.620 96.850 89.040 ;
        RECT 96.650 85.300 96.910 85.620 ;
        RECT 96.640 83.745 96.920 84.115 ;
        RECT 96.650 83.600 96.910 83.745 ;
        RECT 97.170 83.240 97.310 90.740 ;
        RECT 97.630 84.115 97.770 121.680 ;
        RECT 99.010 109.080 99.150 123.720 ;
        RECT 99.470 118.600 99.610 126.020 ;
        RECT 99.870 118.620 100.130 118.940 ;
        RECT 99.410 118.280 99.670 118.600 ;
        RECT 98.950 108.760 99.210 109.080 ;
        RECT 99.010 99.220 99.150 108.760 ;
        RECT 98.950 98.900 99.210 99.220 ;
        RECT 98.030 97.540 98.290 97.860 ;
        RECT 98.090 96.840 98.230 97.540 ;
        RECT 98.030 96.520 98.290 96.840 ;
        RECT 98.950 96.520 99.210 96.840 ;
        RECT 97.560 83.745 97.840 84.115 ;
        RECT 97.110 82.920 97.370 83.240 ;
        RECT 98.090 80.860 98.230 96.520 ;
        RECT 99.010 90.040 99.150 96.520 ;
        RECT 98.950 89.720 99.210 90.040 ;
        RECT 98.490 89.040 98.750 89.360 ;
        RECT 98.550 84.600 98.690 89.040 ;
        RECT 98.490 84.280 98.750 84.600 ;
        RECT 99.010 83.920 99.150 89.720 ;
        RECT 99.470 89.360 99.610 118.280 ;
        RECT 99.930 116.220 100.070 118.620 ;
        RECT 99.870 115.900 100.130 116.220 ;
        RECT 99.930 111.460 100.070 115.900 ;
        RECT 100.850 115.540 100.990 128.820 ;
        RECT 104.070 125.400 104.210 154.660 ;
        RECT 104.470 153.640 104.730 153.960 ;
        RECT 104.530 152.600 104.670 153.640 ;
        RECT 105.390 153.300 105.650 153.620 ;
        RECT 104.470 152.280 104.730 152.600 ;
        RECT 104.530 146.820 104.670 152.280 ;
        RECT 105.450 151.580 105.590 153.300 ;
        RECT 105.390 151.260 105.650 151.580 ;
        RECT 107.750 151.240 107.890 172.680 ;
        RECT 108.210 170.960 108.350 178.960 ;
        RECT 109.070 172.340 109.330 172.660 ;
        RECT 109.130 171.300 109.270 172.340 ;
        RECT 109.070 170.980 109.330 171.300 ;
        RECT 108.150 170.640 108.410 170.960 ;
        RECT 108.610 170.640 108.870 170.960 ;
        RECT 108.670 168.580 108.810 170.640 ;
        RECT 109.130 168.920 109.270 170.980 ;
        RECT 109.070 168.600 109.330 168.920 ;
        RECT 108.610 168.260 108.870 168.580 ;
        RECT 108.150 167.580 108.410 167.900 ;
        RECT 108.210 167.220 108.350 167.580 ;
        RECT 108.150 166.900 108.410 167.220 ;
        RECT 109.130 165.860 109.270 168.600 ;
        RECT 109.070 165.540 109.330 165.860 ;
        RECT 108.150 165.200 108.410 165.520 ;
        RECT 108.210 157.020 108.350 165.200 ;
        RECT 108.610 160.440 108.870 160.760 ;
        RECT 108.670 158.040 108.810 160.440 ;
        RECT 109.070 159.420 109.330 159.740 ;
        RECT 108.610 157.720 108.870 158.040 ;
        RECT 108.150 156.700 108.410 157.020 ;
        RECT 109.130 154.980 109.270 159.420 ;
        RECT 109.590 157.360 109.730 180.500 ;
        RECT 110.050 179.800 110.190 181.860 ;
        RECT 109.990 179.480 110.250 179.800 ;
        RECT 110.510 178.440 110.650 184.580 ;
        RECT 112.810 184.220 112.950 188.660 ;
        RECT 115.050 186.960 115.310 187.280 ;
        RECT 116.890 186.960 117.150 187.280 ;
        RECT 113.210 185.940 113.470 186.260 ;
        RECT 110.910 183.900 111.170 184.220 ;
        RECT 112.750 183.900 113.010 184.220 ;
        RECT 110.970 180.820 111.110 183.900 ;
        RECT 110.910 180.500 111.170 180.820 ;
        RECT 111.830 180.500 112.090 180.820 ;
        RECT 110.450 178.120 110.710 178.440 ;
        RECT 110.510 173.340 110.650 178.120 ;
        RECT 110.910 177.780 111.170 178.100 ;
        RECT 111.370 177.780 111.630 178.100 ;
        RECT 110.970 177.275 111.110 177.780 ;
        RECT 110.900 176.905 111.180 177.275 ;
        RECT 111.430 176.060 111.570 177.780 ;
        RECT 111.890 176.400 112.030 180.500 ;
        RECT 112.810 179.800 112.950 183.900 ;
        RECT 113.270 183.880 113.410 185.940 ;
        RECT 114.590 184.240 114.850 184.560 ;
        RECT 113.210 183.560 113.470 183.880 ;
        RECT 113.270 182.090 113.410 183.560 ;
        RECT 113.670 182.090 113.930 182.180 ;
        RECT 113.270 181.950 113.930 182.090 ;
        RECT 113.670 181.860 113.930 181.950 ;
        RECT 113.730 181.160 113.870 181.860 ;
        RECT 113.670 180.840 113.930 181.160 ;
        RECT 112.750 179.480 113.010 179.800 ;
        RECT 113.730 179.120 113.870 180.840 ;
        RECT 113.670 178.800 113.930 179.120 ;
        RECT 114.650 176.990 114.790 184.240 ;
        RECT 115.110 183.880 115.250 186.960 ;
        RECT 116.950 184.560 117.090 186.960 ;
        RECT 117.410 185.240 117.550 189.000 ;
        RECT 117.870 186.940 118.010 191.380 ;
        RECT 119.190 189.000 119.450 189.320 ;
        RECT 119.250 187.960 119.390 189.000 ;
        RECT 120.630 188.980 120.770 192.400 ;
        RECT 128.850 189.340 129.110 189.660 ;
        RECT 120.570 188.660 120.830 188.980 ;
        RECT 119.190 187.640 119.450 187.960 ;
        RECT 117.810 186.620 118.070 186.940 ;
        RECT 117.350 184.920 117.610 185.240 ;
        RECT 116.890 184.240 117.150 184.560 ;
        RECT 117.870 184.220 118.010 186.620 ;
        RECT 119.650 184.920 119.910 185.240 ;
        RECT 118.270 184.580 118.530 184.900 ;
        RECT 118.330 184.220 118.470 184.580 ;
        RECT 117.810 184.075 118.070 184.220 ;
        RECT 115.050 183.560 115.310 183.880 ;
        RECT 115.970 183.560 116.230 183.880 ;
        RECT 117.800 183.705 118.080 184.075 ;
        RECT 118.270 183.900 118.530 184.220 ;
        RECT 115.040 183.025 115.320 183.395 ;
        RECT 115.110 178.780 115.250 183.025 ;
        RECT 116.030 182.520 116.170 183.560 ;
        RECT 117.810 183.220 118.070 183.540 ;
        RECT 115.970 182.200 116.230 182.520 ;
        RECT 115.970 181.520 116.230 181.840 ;
        RECT 115.510 180.500 115.770 180.820 ;
        RECT 115.570 179.460 115.710 180.500 ;
        RECT 115.510 179.140 115.770 179.460 ;
        RECT 115.050 178.460 115.310 178.780 ;
        RECT 114.190 176.850 114.790 176.990 ;
        RECT 111.830 176.080 112.090 176.400 ;
        RECT 111.370 175.740 111.630 176.060 ;
        RECT 113.670 175.740 113.930 176.060 ;
        RECT 111.830 175.400 112.090 175.720 ;
        RECT 111.890 174.360 112.030 175.400 ;
        RECT 112.750 175.060 113.010 175.380 ;
        RECT 111.830 174.040 112.090 174.360 ;
        RECT 112.810 173.340 112.950 175.060 ;
        RECT 113.730 173.340 113.870 175.740 ;
        RECT 110.450 173.020 110.710 173.340 ;
        RECT 111.370 173.020 111.630 173.340 ;
        RECT 112.750 173.020 113.010 173.340 ;
        RECT 113.670 173.195 113.930 173.340 ;
        RECT 110.510 170.960 110.650 173.020 ;
        RECT 110.910 172.340 111.170 172.660 ;
        RECT 110.970 171.640 111.110 172.340 ;
        RECT 111.430 171.835 111.570 173.020 ;
        RECT 110.910 171.320 111.170 171.640 ;
        RECT 111.360 171.465 111.640 171.835 ;
        RECT 110.450 170.640 110.710 170.960 ;
        RECT 111.430 170.620 111.570 171.465 ;
        RECT 112.810 170.960 112.950 173.020 ;
        RECT 113.660 172.825 113.940 173.195 ;
        RECT 112.750 170.640 113.010 170.960 ;
        RECT 111.370 170.300 111.630 170.620 ;
        RECT 110.910 169.960 111.170 170.280 ;
        RECT 109.990 161.460 110.250 161.780 ;
        RECT 110.050 160.080 110.190 161.460 ;
        RECT 109.990 159.760 110.250 160.080 ;
        RECT 110.970 158.040 111.110 169.960 ;
        RECT 111.430 167.900 111.570 170.300 ;
        RECT 113.670 169.620 113.930 169.940 ;
        RECT 111.370 167.580 111.630 167.900 ;
        RECT 111.430 160.275 111.570 167.580 ;
        RECT 113.210 161.460 113.470 161.780 ;
        RECT 111.360 159.905 111.640 160.275 ;
        RECT 111.370 159.760 111.630 159.905 ;
        RECT 112.750 159.760 113.010 160.080 ;
        RECT 112.290 159.080 112.550 159.400 ;
        RECT 110.910 157.720 111.170 158.040 ;
        RECT 109.530 157.040 109.790 157.360 ;
        RECT 110.450 156.020 110.710 156.340 ;
        RECT 110.510 154.980 110.650 156.020 ;
        RECT 109.070 154.660 109.330 154.980 ;
        RECT 110.450 154.660 110.710 154.980 ;
        RECT 111.830 151.500 112.090 151.580 ;
        RECT 112.350 151.500 112.490 159.080 ;
        RECT 111.830 151.360 112.490 151.500 ;
        RECT 111.830 151.260 112.090 151.360 ;
        RECT 107.690 150.920 107.950 151.240 ;
        RECT 110.450 150.920 110.710 151.240 ;
        RECT 110.510 149.200 110.650 150.920 ;
        RECT 110.450 148.880 110.710 149.200 ;
        RECT 105.390 147.860 105.650 148.180 ;
        RECT 104.470 146.500 104.730 146.820 ;
        RECT 105.450 146.140 105.590 147.860 ;
        RECT 112.810 146.140 112.950 159.760 ;
        RECT 113.270 159.740 113.410 161.460 ;
        RECT 113.210 159.420 113.470 159.740 ;
        RECT 113.210 154.320 113.470 154.640 ;
        RECT 113.270 152.600 113.410 154.320 ;
        RECT 113.210 152.280 113.470 152.600 ;
        RECT 113.730 152.000 113.870 169.620 ;
        RECT 114.190 159.990 114.330 176.850 ;
        RECT 114.590 176.080 114.850 176.400 ;
        RECT 114.650 170.280 114.790 176.080 ;
        RECT 115.570 176.060 115.710 179.140 ;
        RECT 116.030 178.780 116.170 181.520 ;
        RECT 117.350 180.840 117.610 181.160 ;
        RECT 116.890 180.500 117.150 180.820 ;
        RECT 115.970 178.460 116.230 178.780 ;
        RECT 116.950 178.350 117.090 180.500 ;
        RECT 117.410 179.370 117.550 180.840 ;
        RECT 117.870 180.820 118.010 183.220 ;
        RECT 117.810 180.500 118.070 180.820 ;
        RECT 117.810 179.370 118.070 179.460 ;
        RECT 117.410 179.230 118.070 179.370 ;
        RECT 117.810 179.140 118.070 179.230 ;
        RECT 116.950 178.210 117.550 178.350 ;
        RECT 115.970 177.780 116.230 178.100 ;
        RECT 115.040 175.545 115.320 175.915 ;
        RECT 115.510 175.740 115.770 176.060 ;
        RECT 116.030 175.800 116.170 177.780 ;
        RECT 116.880 176.905 117.160 177.275 ;
        RECT 116.950 176.740 117.090 176.905 ;
        RECT 116.890 176.420 117.150 176.740 ;
        RECT 117.410 175.800 117.550 178.210 ;
        RECT 117.870 178.100 118.010 179.140 ;
        RECT 118.330 179.120 118.470 183.900 ;
        RECT 118.730 180.500 118.990 180.820 ;
        RECT 119.190 180.500 119.450 180.820 ;
        RECT 118.790 179.800 118.930 180.500 ;
        RECT 118.730 179.480 118.990 179.800 ;
        RECT 118.270 178.800 118.530 179.120 ;
        RECT 118.730 178.120 118.990 178.440 ;
        RECT 117.810 177.780 118.070 178.100 ;
        RECT 117.870 176.400 118.010 177.780 ;
        RECT 117.810 176.080 118.070 176.400 ;
        RECT 118.270 176.080 118.530 176.400 ;
        RECT 118.330 175.800 118.470 176.080 ;
        RECT 116.030 175.660 116.630 175.800 ;
        RECT 115.110 174.020 115.250 175.545 ;
        RECT 115.970 175.060 116.230 175.380 ;
        RECT 115.510 174.040 115.770 174.360 ;
        RECT 115.050 173.700 115.310 174.020 ;
        RECT 115.050 173.020 115.310 173.340 ;
        RECT 115.110 171.640 115.250 173.020 ;
        RECT 115.570 173.000 115.710 174.040 ;
        RECT 116.030 173.340 116.170 175.060 ;
        RECT 115.970 173.020 116.230 173.340 ;
        RECT 115.510 172.680 115.770 173.000 ;
        RECT 115.050 171.320 115.310 171.640 ;
        RECT 115.570 170.620 115.710 172.680 ;
        RECT 115.510 170.300 115.770 170.620 ;
        RECT 114.590 169.960 114.850 170.280 ;
        RECT 116.030 168.920 116.170 173.020 ;
        RECT 115.970 168.600 116.230 168.920 ;
        RECT 115.510 162.140 115.770 162.460 ;
        RECT 115.050 160.440 115.310 160.760 ;
        RECT 114.590 159.990 114.850 160.080 ;
        RECT 114.190 159.850 114.850 159.990 ;
        RECT 114.190 159.060 114.330 159.850 ;
        RECT 114.590 159.760 114.850 159.850 ;
        RECT 114.130 158.740 114.390 159.060 ;
        RECT 114.590 157.720 114.850 158.040 ;
        RECT 114.650 153.960 114.790 157.720 ;
        RECT 115.110 154.640 115.250 160.440 ;
        RECT 115.570 160.275 115.710 162.140 ;
        RECT 115.500 159.905 115.780 160.275 ;
        RECT 116.490 160.080 116.630 175.660 ;
        RECT 116.950 175.660 117.550 175.800 ;
        RECT 117.870 175.720 118.470 175.800 ;
        RECT 117.810 175.660 118.470 175.720 ;
        RECT 116.950 173.340 117.090 175.660 ;
        RECT 117.810 175.400 118.070 175.660 ;
        RECT 117.350 175.060 117.610 175.380 ;
        RECT 118.270 175.060 118.530 175.380 ;
        RECT 116.890 173.020 117.150 173.340 ;
        RECT 116.950 168.580 117.090 173.020 ;
        RECT 117.410 170.620 117.550 175.060 ;
        RECT 117.810 174.040 118.070 174.360 ;
        RECT 117.350 170.300 117.610 170.620 ;
        RECT 116.890 168.260 117.150 168.580 ;
        RECT 116.890 167.580 117.150 167.900 ;
        RECT 116.950 166.200 117.090 167.580 ;
        RECT 116.890 165.880 117.150 166.200 ;
        RECT 116.950 162.995 117.090 165.880 ;
        RECT 117.410 164.920 117.550 170.300 ;
        RECT 117.870 168.240 118.010 174.040 ;
        RECT 118.330 173.340 118.470 175.060 ;
        RECT 118.790 174.020 118.930 178.120 ;
        RECT 118.730 173.700 118.990 174.020 ;
        RECT 118.270 173.020 118.530 173.340 ;
        RECT 118.730 173.020 118.990 173.340 ;
        RECT 118.330 170.280 118.470 173.020 ;
        RECT 118.790 172.515 118.930 173.020 ;
        RECT 118.720 172.145 119.000 172.515 ;
        RECT 118.720 171.465 119.000 171.835 ;
        RECT 118.730 171.320 118.990 171.465 ;
        RECT 118.270 169.960 118.530 170.280 ;
        RECT 118.790 168.580 118.930 171.320 ;
        RECT 118.730 168.260 118.990 168.580 ;
        RECT 117.810 167.920 118.070 168.240 ;
        RECT 118.730 167.580 118.990 167.900 ;
        RECT 118.270 166.900 118.530 167.220 ;
        RECT 117.410 164.780 118.010 164.920 ;
        RECT 117.870 164.500 118.010 164.780 ;
        RECT 117.350 164.180 117.610 164.500 ;
        RECT 117.810 164.180 118.070 164.500 ;
        RECT 116.880 162.625 117.160 162.995 ;
        RECT 115.510 159.760 115.770 159.905 ;
        RECT 116.430 159.760 116.690 160.080 ;
        RECT 116.490 157.360 116.630 159.760 ;
        RECT 116.950 158.040 117.090 162.625 ;
        RECT 116.890 157.720 117.150 158.040 ;
        RECT 116.430 157.040 116.690 157.360 ;
        RECT 116.490 154.640 116.630 157.040 ;
        RECT 116.890 156.700 117.150 157.020 ;
        RECT 116.950 154.720 117.090 156.700 ;
        RECT 117.410 155.320 117.550 164.180 ;
        RECT 117.800 161.265 118.080 161.635 ;
        RECT 117.870 159.740 118.010 161.265 ;
        RECT 117.810 159.420 118.070 159.740 ;
        RECT 117.870 156.680 118.010 159.420 ;
        RECT 118.330 159.060 118.470 166.900 ;
        RECT 118.790 161.780 118.930 167.580 ;
        RECT 119.250 162.460 119.390 180.500 ;
        RECT 119.710 179.800 119.850 184.920 ;
        RECT 120.110 183.900 120.370 184.220 ;
        RECT 120.170 181.500 120.310 183.900 ;
        RECT 120.630 183.880 120.770 188.660 ;
        RECT 128.910 186.000 129.050 189.340 ;
        RECT 128.910 185.860 129.510 186.000 ;
        RECT 122.870 184.580 123.130 184.900 ;
        RECT 121.030 183.900 121.290 184.220 ;
        RECT 120.570 183.560 120.830 183.880 ;
        RECT 120.630 183.395 120.770 183.560 ;
        RECT 120.560 183.025 120.840 183.395 ;
        RECT 120.110 181.180 120.370 181.500 ;
        RECT 119.650 179.480 119.910 179.800 ;
        RECT 119.650 178.350 119.910 178.670 ;
        RECT 119.710 173.000 119.850 178.350 ;
        RECT 120.170 176.060 120.310 181.180 ;
        RECT 120.570 176.310 120.830 176.400 ;
        RECT 121.090 176.310 121.230 183.900 ;
        RECT 121.490 183.220 121.750 183.540 ;
        RECT 121.550 182.520 121.690 183.220 ;
        RECT 121.490 182.200 121.750 182.520 ;
        RECT 121.490 179.480 121.750 179.800 ;
        RECT 121.550 179.100 121.690 179.480 ;
        RECT 122.410 179.100 122.670 179.120 ;
        RECT 122.930 179.100 123.070 184.580 ;
        RECT 129.370 181.840 129.510 185.860 ;
        RECT 138.050 183.900 138.310 184.220 ;
        RECT 141.270 183.900 141.530 184.220 ;
        RECT 138.110 181.840 138.250 183.900 ;
        RECT 139.890 183.220 140.150 183.540 ;
        RECT 139.950 181.840 140.090 183.220 ;
        RECT 129.310 181.520 129.570 181.840 ;
        RECT 133.910 181.520 134.170 181.840 ;
        RECT 138.050 181.520 138.310 181.840 ;
        RECT 139.890 181.520 140.150 181.840 ;
        RECT 129.370 181.240 129.510 181.520 ;
        RECT 129.370 181.100 129.970 181.240 ;
        RECT 121.550 178.960 122.150 179.100 ;
        RECT 122.010 178.520 122.150 178.960 ;
        RECT 122.410 178.960 123.070 179.100 ;
        RECT 122.410 178.800 122.670 178.960 ;
        RECT 122.010 178.380 122.610 178.520 ;
        RECT 121.950 177.780 122.210 178.100 ;
        RECT 122.010 176.400 122.150 177.780 ;
        RECT 120.570 176.170 121.230 176.310 ;
        RECT 120.570 176.080 120.830 176.170 ;
        RECT 120.110 175.740 120.370 176.060 ;
        RECT 121.090 175.720 121.230 176.170 ;
        RECT 121.490 176.080 121.750 176.400 ;
        RECT 121.950 176.080 122.210 176.400 ;
        RECT 121.030 175.400 121.290 175.720 ;
        RECT 120.110 173.700 120.370 174.020 ;
        RECT 119.650 172.680 119.910 173.000 ;
        RECT 120.170 170.960 120.310 173.700 ;
        RECT 120.570 173.195 120.830 173.340 ;
        RECT 120.560 172.825 120.840 173.195 ;
        RECT 121.020 171.465 121.300 171.835 ;
        RECT 120.110 170.640 120.370 170.960 ;
        RECT 120.170 167.900 120.310 170.640 ;
        RECT 120.110 167.580 120.370 167.900 ;
        RECT 120.170 165.860 120.310 167.580 ;
        RECT 121.090 167.220 121.230 171.465 ;
        RECT 121.550 170.960 121.690 176.080 ;
        RECT 121.950 172.515 122.210 172.660 ;
        RECT 121.940 172.145 122.220 172.515 ;
        RECT 121.940 171.465 122.220 171.835 ;
        RECT 122.010 171.040 122.150 171.465 ;
        RECT 122.470 171.040 122.610 178.380 ;
        RECT 122.930 177.080 123.070 178.960 ;
        RECT 125.630 178.800 125.890 179.120 ;
        RECT 129.310 178.800 129.570 179.120 ;
        RECT 123.790 177.780 124.050 178.100 ;
        RECT 122.870 176.760 123.130 177.080 ;
        RECT 122.930 171.300 123.070 176.760 ;
        RECT 123.330 176.420 123.590 176.740 ;
        RECT 123.390 174.360 123.530 176.420 ;
        RECT 123.850 175.915 123.990 177.780 ;
        RECT 123.780 175.545 124.060 175.915 ;
        RECT 123.330 174.040 123.590 174.360 ;
        RECT 123.330 172.680 123.590 173.000 ;
        RECT 122.010 170.960 122.610 171.040 ;
        RECT 122.870 170.980 123.130 171.300 ;
        RECT 121.490 170.640 121.750 170.960 ;
        RECT 122.010 170.900 122.670 170.960 ;
        RECT 122.410 170.640 122.670 170.900 ;
        RECT 121.550 168.920 121.690 170.640 ;
        RECT 122.870 170.300 123.130 170.620 ;
        RECT 121.950 169.960 122.210 170.280 ;
        RECT 121.490 168.600 121.750 168.920 ;
        RECT 121.030 166.900 121.290 167.220 ;
        RECT 120.110 165.540 120.370 165.860 ;
        RECT 121.550 165.520 121.690 168.600 ;
        RECT 121.490 165.200 121.750 165.520 ;
        RECT 119.650 164.180 119.910 164.500 ;
        RECT 119.710 162.460 119.850 164.180 ;
        RECT 119.190 162.315 119.450 162.460 ;
        RECT 119.180 161.945 119.460 162.315 ;
        RECT 119.650 162.140 119.910 162.460 ;
        RECT 118.730 161.460 118.990 161.780 ;
        RECT 119.190 159.760 119.450 160.080 ;
        RECT 118.730 159.080 118.990 159.400 ;
        RECT 118.270 158.740 118.530 159.060 ;
        RECT 118.270 157.720 118.530 158.040 ;
        RECT 118.330 156.680 118.470 157.720 ;
        RECT 117.810 156.360 118.070 156.680 ;
        RECT 118.270 156.360 118.530 156.680 ;
        RECT 117.350 155.000 117.610 155.320 ;
        RECT 115.050 154.320 115.310 154.640 ;
        RECT 115.510 154.320 115.770 154.640 ;
        RECT 116.430 154.320 116.690 154.640 ;
        RECT 116.950 154.580 117.550 154.720 ;
        RECT 118.330 154.640 118.470 156.360 ;
        RECT 118.790 155.320 118.930 159.080 ;
        RECT 118.730 155.000 118.990 155.320 ;
        RECT 114.590 153.640 114.850 153.960 ;
        RECT 113.730 151.860 114.330 152.000 ;
        RECT 113.670 151.260 113.930 151.580 ;
        RECT 113.730 148.180 113.870 151.260 ;
        RECT 113.210 147.860 113.470 148.180 ;
        RECT 113.670 147.860 113.930 148.180 ;
        RECT 105.390 145.820 105.650 146.140 ;
        RECT 112.750 145.820 113.010 146.140 ;
        RECT 113.270 145.800 113.410 147.860 ;
        RECT 113.730 146.820 113.870 147.860 ;
        RECT 113.670 146.500 113.930 146.820 ;
        RECT 104.470 145.480 104.730 145.800 ;
        RECT 113.210 145.480 113.470 145.800 ;
        RECT 104.530 140.700 104.670 145.480 ;
        RECT 104.930 145.140 105.190 145.460 ;
        RECT 104.990 141.720 105.130 145.140 ;
        RECT 114.190 143.420 114.330 151.860 ;
        RECT 114.650 151.580 114.790 153.640 ;
        RECT 114.590 151.260 114.850 151.580 ;
        RECT 115.570 146.140 115.710 154.320 ;
        RECT 117.410 154.300 117.550 154.580 ;
        RECT 118.270 154.320 118.530 154.640 ;
        RECT 117.350 153.980 117.610 154.300 ;
        RECT 115.970 153.300 116.230 153.620 ;
        RECT 116.430 153.300 116.690 153.620 ;
        RECT 116.030 149.880 116.170 153.300 ;
        RECT 116.490 151.920 116.630 153.300 ;
        RECT 116.430 151.600 116.690 151.920 ;
        RECT 116.430 150.920 116.690 151.240 ;
        RECT 115.970 149.560 116.230 149.880 ;
        RECT 116.490 149.200 116.630 150.920 ;
        RECT 117.410 150.900 117.550 153.980 ;
        RECT 118.330 151.240 118.470 154.320 ;
        RECT 118.730 153.980 118.990 154.300 ;
        RECT 118.270 150.920 118.530 151.240 ;
        RECT 117.350 150.580 117.610 150.900 ;
        RECT 116.430 148.880 116.690 149.200 ;
        RECT 118.790 147.160 118.930 153.980 ;
        RECT 118.730 146.840 118.990 147.160 ;
        RECT 115.510 145.820 115.770 146.140 ;
        RECT 116.890 145.140 117.150 145.460 ;
        RECT 114.130 143.100 114.390 143.420 ;
        RECT 104.930 141.400 105.190 141.720 ;
        RECT 113.210 141.400 113.470 141.720 ;
        RECT 104.470 140.380 104.730 140.700 ;
        RECT 104.530 139.000 104.670 140.380 ;
        RECT 104.930 140.040 105.190 140.360 ;
        RECT 104.990 139.000 105.130 140.040 ;
        RECT 106.770 139.700 107.030 140.020 ;
        RECT 110.910 139.700 111.170 140.020 ;
        RECT 106.830 139.000 106.970 139.700 ;
        RECT 110.970 139.000 111.110 139.700 ;
        RECT 104.470 138.680 104.730 139.000 ;
        RECT 104.930 138.680 105.190 139.000 ;
        RECT 106.770 138.680 107.030 139.000 ;
        RECT 110.910 138.680 111.170 139.000 ;
        RECT 112.290 138.680 112.550 139.000 ;
        RECT 109.530 138.000 109.790 138.320 ;
        RECT 108.150 134.260 108.410 134.580 ;
        RECT 108.210 133.560 108.350 134.260 ;
        RECT 109.590 133.560 109.730 138.000 ;
        RECT 111.370 135.620 111.630 135.940 ;
        RECT 108.150 133.240 108.410 133.560 ;
        RECT 109.530 133.240 109.790 133.560 ;
        RECT 111.430 132.880 111.570 135.620 ;
        RECT 109.990 132.560 110.250 132.880 ;
        RECT 110.450 132.560 110.710 132.880 ;
        RECT 111.370 132.560 111.630 132.880 ;
        RECT 107.230 132.220 107.490 132.540 ;
        RECT 109.530 132.220 109.790 132.540 ;
        RECT 107.290 127.100 107.430 132.220 ;
        RECT 108.610 128.820 108.870 129.140 ;
        RECT 108.670 128.120 108.810 128.820 ;
        RECT 108.610 127.800 108.870 128.120 ;
        RECT 108.150 127.120 108.410 127.440 ;
        RECT 106.770 126.780 107.030 127.100 ;
        RECT 107.230 126.780 107.490 127.100 ;
        RECT 104.470 126.100 104.730 126.420 ;
        RECT 104.010 125.080 104.270 125.400 ;
        RECT 104.530 124.380 104.670 126.100 ;
        RECT 106.830 125.060 106.970 126.780 ;
        RECT 106.770 124.740 107.030 125.060 ;
        RECT 104.470 124.060 104.730 124.380 ;
        RECT 106.770 121.680 107.030 122.000 ;
        RECT 104.010 121.340 104.270 121.660 ;
        RECT 101.250 120.660 101.510 120.980 ;
        RECT 101.310 118.940 101.450 120.660 ;
        RECT 104.070 118.940 104.210 121.340 ;
        RECT 106.830 119.960 106.970 121.680 ;
        RECT 107.290 121.660 107.430 126.780 ;
        RECT 108.210 125.400 108.350 127.120 ;
        RECT 108.150 125.080 108.410 125.400 ;
        RECT 107.230 121.340 107.490 121.660 ;
        RECT 106.770 119.640 107.030 119.960 ;
        RECT 101.250 118.620 101.510 118.940 ;
        RECT 104.010 118.620 104.270 118.940 ;
        RECT 105.850 118.620 106.110 118.940 ;
        RECT 100.790 115.220 101.050 115.540 ;
        RECT 100.330 113.520 100.590 113.840 ;
        RECT 99.870 111.140 100.130 111.460 ;
        RECT 100.390 111.120 100.530 113.520 ;
        RECT 105.390 112.840 105.650 113.160 ;
        RECT 105.450 111.460 105.590 112.840 ;
        RECT 101.250 111.140 101.510 111.460 ;
        RECT 104.010 111.370 104.270 111.460 ;
        RECT 105.390 111.370 105.650 111.460 ;
        RECT 104.010 111.230 105.650 111.370 ;
        RECT 104.010 111.140 104.270 111.230 ;
        RECT 105.390 111.140 105.650 111.230 ;
        RECT 100.330 110.800 100.590 111.120 ;
        RECT 100.790 110.120 101.050 110.440 ;
        RECT 100.330 97.540 100.590 97.860 ;
        RECT 100.390 91.400 100.530 97.540 ;
        RECT 100.850 97.520 100.990 110.120 ;
        RECT 101.310 108.060 101.450 111.140 ;
        RECT 104.010 110.520 104.270 110.780 ;
        RECT 105.910 110.520 106.050 118.620 ;
        RECT 106.830 116.560 106.970 119.640 ;
        RECT 108.150 117.940 108.410 118.260 ;
        RECT 108.210 116.900 108.350 117.940 ;
        RECT 108.150 116.580 108.410 116.900 ;
        RECT 106.770 116.240 107.030 116.560 ;
        RECT 106.830 114.520 106.970 116.240 ;
        RECT 108.610 115.560 108.870 115.880 ;
        RECT 106.770 114.200 107.030 114.520 ;
        RECT 106.830 110.780 106.970 114.200 ;
        RECT 108.670 113.500 108.810 115.560 ;
        RECT 108.610 113.180 108.870 113.500 ;
        RECT 107.230 112.500 107.490 112.820 ;
        RECT 107.290 111.120 107.430 112.500 ;
        RECT 107.230 110.800 107.490 111.120 ;
        RECT 104.010 110.460 106.050 110.520 ;
        RECT 106.770 110.460 107.030 110.780 ;
        RECT 104.070 110.380 106.050 110.460 ;
        RECT 102.170 108.420 102.430 108.740 ;
        RECT 101.250 107.740 101.510 108.060 ;
        RECT 102.230 102.620 102.370 108.420 ;
        RECT 105.390 105.700 105.650 106.020 ;
        RECT 104.930 102.980 105.190 103.300 ;
        RECT 104.990 102.620 105.130 102.980 ;
        RECT 105.450 102.620 105.590 105.700 ;
        RECT 105.910 102.620 106.050 110.380 ;
        RECT 108.150 108.760 108.410 109.080 ;
        RECT 107.230 107.060 107.490 107.380 ;
        RECT 107.290 106.360 107.430 107.060 ;
        RECT 107.230 106.040 107.490 106.360 ;
        RECT 106.310 102.640 106.570 102.960 ;
        RECT 107.290 102.870 107.430 106.040 ;
        RECT 108.210 105.680 108.350 108.760 ;
        RECT 107.690 105.360 107.950 105.680 ;
        RECT 108.150 105.360 108.410 105.680 ;
        RECT 109.070 105.360 109.330 105.680 ;
        RECT 107.750 105.195 107.890 105.360 ;
        RECT 107.680 104.825 107.960 105.195 ;
        RECT 107.750 103.640 107.890 104.825 ;
        RECT 108.610 104.340 108.870 104.660 ;
        RECT 107.690 103.320 107.950 103.640 ;
        RECT 106.830 102.730 107.430 102.870 ;
        RECT 102.170 102.300 102.430 102.620 ;
        RECT 104.930 102.300 105.190 102.620 ;
        RECT 105.390 102.300 105.650 102.620 ;
        RECT 105.850 102.300 106.110 102.620 ;
        RECT 101.710 101.620 101.970 101.940 ;
        RECT 100.790 97.200 101.050 97.520 ;
        RECT 101.770 91.740 101.910 101.620 ;
        RECT 103.550 97.880 103.810 98.200 ;
        RECT 103.090 96.860 103.350 97.180 ;
        RECT 103.150 95.140 103.290 96.860 ;
        RECT 103.090 94.820 103.350 95.140 ;
        RECT 102.170 94.480 102.430 94.800 ;
        RECT 102.230 92.760 102.370 94.480 ;
        RECT 102.630 94.140 102.890 94.460 ;
        RECT 102.170 92.440 102.430 92.760 ;
        RECT 101.710 91.420 101.970 91.740 ;
        RECT 100.330 91.080 100.590 91.400 ;
        RECT 99.410 89.040 99.670 89.360 ;
        RECT 99.470 88.875 99.610 89.040 ;
        RECT 100.390 89.020 100.530 91.080 ;
        RECT 102.690 89.360 102.830 94.140 ;
        RECT 103.610 92.420 103.750 97.880 ;
        RECT 106.370 92.760 106.510 102.640 ;
        RECT 106.830 102.280 106.970 102.730 ;
        RECT 107.690 102.530 107.950 102.620 ;
        RECT 107.290 102.390 107.950 102.530 ;
        RECT 106.770 101.960 107.030 102.280 ;
        RECT 107.290 99.900 107.430 102.390 ;
        RECT 107.690 102.300 107.950 102.390 ;
        RECT 108.670 100.580 108.810 104.340 ;
        RECT 109.130 103.640 109.270 105.360 ;
        RECT 109.070 103.320 109.330 103.640 ;
        RECT 108.610 100.260 108.870 100.580 ;
        RECT 107.230 99.580 107.490 99.900 ;
        RECT 107.290 97.520 107.430 99.580 ;
        RECT 108.610 97.540 108.870 97.860 ;
        RECT 107.230 97.200 107.490 97.520 ;
        RECT 106.310 92.440 106.570 92.760 ;
        RECT 103.550 92.100 103.810 92.420 ;
        RECT 106.370 91.740 106.510 92.440 ;
        RECT 106.310 91.420 106.570 91.740 ;
        RECT 106.770 91.420 107.030 91.740 ;
        RECT 106.370 89.700 106.510 91.420 ;
        RECT 106.310 89.380 106.570 89.700 ;
        RECT 102.630 89.040 102.890 89.360 ;
        RECT 99.400 88.505 99.680 88.875 ;
        RECT 100.330 88.700 100.590 89.020 ;
        RECT 100.790 88.020 101.050 88.340 ;
        RECT 100.850 85.960 100.990 88.020 ;
        RECT 102.690 86.300 102.830 89.040 ;
        RECT 106.830 87.320 106.970 91.420 ;
        RECT 108.150 89.040 108.410 89.360 ;
        RECT 108.210 87.320 108.350 89.040 ;
        RECT 106.770 87.000 107.030 87.320 ;
        RECT 108.150 87.000 108.410 87.320 ;
        RECT 105.390 86.660 105.650 86.980 ;
        RECT 102.630 85.980 102.890 86.300 ;
        RECT 100.790 85.640 101.050 85.960 ;
        RECT 100.330 85.300 100.590 85.620 ;
        RECT 98.490 83.600 98.750 83.920 ;
        RECT 98.950 83.600 99.210 83.920 ;
        RECT 98.550 83.240 98.690 83.600 ;
        RECT 98.490 82.920 98.750 83.240 ;
        RECT 100.390 82.500 100.530 85.300 ;
        RECT 105.450 84.260 105.590 86.660 ;
        RECT 108.670 86.640 108.810 97.540 ;
        RECT 109.070 95.160 109.330 95.480 ;
        RECT 109.130 91.740 109.270 95.160 ;
        RECT 109.590 92.840 109.730 132.220 ;
        RECT 110.050 130.840 110.190 132.560 ;
        RECT 109.990 130.520 110.250 130.840 ;
        RECT 110.510 129.820 110.650 132.560 ;
        RECT 110.910 129.840 111.170 130.160 ;
        RECT 110.450 129.500 110.710 129.820 ;
        RECT 110.970 119.280 111.110 129.840 ;
        RECT 111.370 127.120 111.630 127.440 ;
        RECT 111.430 125.400 111.570 127.120 ;
        RECT 111.370 125.080 111.630 125.400 ;
        RECT 112.350 122.680 112.490 138.680 ;
        RECT 112.750 138.000 113.010 138.320 ;
        RECT 112.810 130.840 112.950 138.000 ;
        RECT 113.270 135.260 113.410 141.400 ;
        RECT 115.970 141.060 116.230 141.380 ;
        RECT 114.130 140.040 114.390 140.360 ;
        RECT 113.670 138.000 113.930 138.320 ;
        RECT 113.730 136.280 113.870 138.000 ;
        RECT 114.190 137.300 114.330 140.040 ;
        RECT 115.510 139.700 115.770 140.020 ;
        RECT 114.130 136.980 114.390 137.300 ;
        RECT 113.670 135.960 113.930 136.280 ;
        RECT 113.210 134.940 113.470 135.260 ;
        RECT 114.190 132.880 114.330 136.980 ;
        RECT 115.570 135.680 115.710 139.700 ;
        RECT 116.030 136.280 116.170 141.060 ;
        RECT 116.430 138.000 116.690 138.320 ;
        RECT 115.970 135.960 116.230 136.280 ;
        RECT 114.650 135.540 116.170 135.680 ;
        RECT 116.490 135.600 116.630 138.000 ;
        RECT 114.650 135.260 114.790 135.540 ;
        RECT 114.590 134.940 114.850 135.260 ;
        RECT 114.130 132.560 114.390 132.880 ;
        RECT 112.750 130.520 113.010 130.840 ;
        RECT 114.650 130.800 114.790 134.940 ;
        RECT 116.030 132.880 116.170 135.540 ;
        RECT 116.430 135.280 116.690 135.600 ;
        RECT 115.970 132.560 116.230 132.880 ;
        RECT 115.510 131.540 115.770 131.860 ;
        RECT 116.950 131.600 117.090 145.140 ;
        RECT 119.250 143.760 119.390 159.760 ;
        RECT 119.710 157.020 119.850 162.140 ;
        RECT 120.560 161.945 120.840 162.315 ;
        RECT 120.110 161.460 120.370 161.780 ;
        RECT 120.170 160.080 120.310 161.460 ;
        RECT 120.110 159.760 120.370 160.080 ;
        RECT 120.110 158.740 120.370 159.060 ;
        RECT 120.170 157.360 120.310 158.740 ;
        RECT 120.110 157.040 120.370 157.360 ;
        RECT 119.650 156.700 119.910 157.020 ;
        RECT 120.170 154.640 120.310 157.040 ;
        RECT 120.630 157.020 120.770 161.945 ;
        RECT 121.030 161.460 121.290 161.780 ;
        RECT 121.550 161.690 121.690 165.200 ;
        RECT 122.010 164.500 122.150 169.960 ;
        RECT 122.930 168.920 123.070 170.300 ;
        RECT 122.870 168.600 123.130 168.920 ;
        RECT 122.410 167.580 122.670 167.900 ;
        RECT 122.470 165.600 122.610 167.580 ;
        RECT 122.930 166.200 123.070 168.600 ;
        RECT 123.390 167.900 123.530 172.680 ;
        RECT 123.850 170.870 123.990 175.545 ;
        RECT 124.710 175.060 124.970 175.380 ;
        RECT 124.770 173.000 124.910 175.060 ;
        RECT 124.710 172.680 124.970 173.000 ;
        RECT 125.170 172.340 125.430 172.660 ;
        RECT 124.250 170.870 124.510 170.960 ;
        RECT 123.850 170.730 124.910 170.870 ;
        RECT 124.250 170.640 124.510 170.730 ;
        RECT 124.250 167.920 124.510 168.240 ;
        RECT 123.330 167.580 123.590 167.900 ;
        RECT 123.790 167.240 124.050 167.560 ;
        RECT 122.870 165.880 123.130 166.200 ;
        RECT 122.470 165.460 123.070 165.600 ;
        RECT 122.410 164.520 122.670 164.840 ;
        RECT 121.950 164.180 122.210 164.500 ;
        RECT 121.950 162.480 122.210 162.800 ;
        RECT 122.010 162.315 122.150 162.480 ;
        RECT 121.940 161.945 122.220 162.315 ;
        RECT 121.950 161.690 122.210 161.780 ;
        RECT 121.550 161.635 122.210 161.690 ;
        RECT 121.480 161.550 122.210 161.635 ;
        RECT 121.090 160.760 121.230 161.460 ;
        RECT 121.480 161.265 121.760 161.550 ;
        RECT 121.950 161.460 122.210 161.550 ;
        RECT 121.030 160.440 121.290 160.760 ;
        RECT 121.090 160.080 121.230 160.440 ;
        RECT 121.030 159.760 121.290 160.080 ;
        RECT 121.490 159.080 121.750 159.400 ;
        RECT 121.550 157.020 121.690 159.080 ;
        RECT 122.470 159.060 122.610 164.520 ;
        RECT 122.930 162.120 123.070 165.460 ;
        RECT 123.850 163.560 123.990 167.240 ;
        RECT 124.310 166.200 124.450 167.920 ;
        RECT 124.770 167.900 124.910 170.730 ;
        RECT 124.710 167.580 124.970 167.900 ;
        RECT 124.250 165.880 124.510 166.200 ;
        RECT 124.710 164.180 124.970 164.500 ;
        RECT 123.850 163.480 124.450 163.560 ;
        RECT 123.850 163.420 124.510 163.480 ;
        RECT 124.250 163.160 124.510 163.420 ;
        RECT 123.320 162.625 123.600 162.995 ;
        RECT 123.390 162.460 123.530 162.625 ;
        RECT 123.330 162.140 123.590 162.460 ;
        RECT 123.790 162.140 124.050 162.460 ;
        RECT 122.870 161.800 123.130 162.120 ;
        RECT 122.410 158.740 122.670 159.060 ;
        RECT 120.570 156.700 120.830 157.020 ;
        RECT 121.490 156.930 121.750 157.020 ;
        RECT 121.490 156.790 122.150 156.930 ;
        RECT 121.490 156.700 121.750 156.790 ;
        RECT 121.490 156.020 121.750 156.340 ;
        RECT 120.110 154.320 120.370 154.640 ;
        RECT 121.030 153.300 121.290 153.620 ;
        RECT 121.090 151.580 121.230 153.300 ;
        RECT 121.030 151.260 121.290 151.580 ;
        RECT 121.550 151.240 121.690 156.020 ;
        RECT 122.010 154.640 122.150 156.790 ;
        RECT 122.410 155.000 122.670 155.320 ;
        RECT 121.950 154.320 122.210 154.640 ;
        RECT 121.490 150.920 121.750 151.240 ;
        RECT 119.650 150.580 119.910 150.900 ;
        RECT 120.570 150.580 120.830 150.900 ;
        RECT 119.710 149.200 119.850 150.580 ;
        RECT 119.650 148.880 119.910 149.200 ;
        RECT 120.630 148.860 120.770 150.580 ;
        RECT 122.010 149.200 122.150 154.320 ;
        RECT 122.470 152.260 122.610 155.000 ;
        RECT 122.930 153.960 123.070 161.800 ;
        RECT 123.330 159.760 123.590 160.080 ;
        RECT 123.390 157.700 123.530 159.760 ;
        RECT 123.330 157.380 123.590 157.700 ;
        RECT 123.390 154.980 123.530 157.380 ;
        RECT 123.850 155.320 123.990 162.140 ;
        RECT 123.790 155.000 124.050 155.320 ;
        RECT 123.330 154.660 123.590 154.980 ;
        RECT 122.870 153.640 123.130 153.960 ;
        RECT 124.310 153.620 124.450 163.160 ;
        RECT 124.770 163.140 124.910 164.180 ;
        RECT 124.710 162.820 124.970 163.140 ;
        RECT 124.250 153.300 124.510 153.620 ;
        RECT 122.410 151.940 122.670 152.260 ;
        RECT 125.230 152.000 125.370 172.340 ;
        RECT 125.690 160.080 125.830 178.800 ;
        RECT 129.370 177.160 129.510 178.800 ;
        RECT 128.910 177.080 129.510 177.160 ;
        RECT 128.850 177.020 129.510 177.080 ;
        RECT 128.850 176.760 129.110 177.020 ;
        RECT 129.830 176.400 129.970 181.100 ;
        RECT 133.970 179.800 134.110 181.520 ;
        RECT 135.750 181.180 136.010 181.500 ;
        RECT 141.330 181.355 141.470 183.900 ;
        RECT 133.910 179.480 134.170 179.800 ;
        RECT 135.810 178.780 135.950 181.180 ;
        RECT 141.260 180.985 141.540 181.355 ;
        RECT 140.810 180.500 141.070 180.820 ;
        RECT 135.750 178.460 136.010 178.780 ;
        RECT 139.890 178.460 140.150 178.780 ;
        RECT 130.230 178.120 130.490 178.440 ;
        RECT 127.930 176.080 128.190 176.400 ;
        RECT 129.770 176.080 130.030 176.400 ;
        RECT 126.550 175.740 126.810 176.060 ;
        RECT 126.610 173.340 126.750 175.740 ;
        RECT 127.990 173.340 128.130 176.080 ;
        RECT 130.290 175.720 130.430 178.120 ;
        RECT 131.610 177.780 131.870 178.100 ;
        RECT 138.970 177.780 139.230 178.100 ;
        RECT 130.690 176.080 130.950 176.400 ;
        RECT 130.230 175.400 130.490 175.720 ;
        RECT 130.750 173.680 130.890 176.080 ;
        RECT 131.670 174.360 131.810 177.780 ;
        RECT 132.070 176.080 132.330 176.400 ;
        RECT 132.130 174.360 132.270 176.080 ;
        RECT 138.050 175.060 138.310 175.380 ;
        RECT 131.610 174.040 131.870 174.360 ;
        RECT 132.070 174.040 132.330 174.360 ;
        RECT 130.690 173.360 130.950 173.680 ;
        RECT 126.550 173.020 126.810 173.340 ;
        RECT 127.930 173.020 128.190 173.340 ;
        RECT 126.610 171.640 126.750 173.020 ;
        RECT 127.990 172.570 128.130 173.020 ;
        RECT 127.530 172.430 128.130 172.570 ;
        RECT 127.530 171.640 127.670 172.430 ;
        RECT 130.230 172.340 130.490 172.660 ;
        RECT 130.290 171.640 130.430 172.340 ;
        RECT 126.550 171.320 126.810 171.640 ;
        RECT 127.470 171.320 127.730 171.640 ;
        RECT 130.230 171.320 130.490 171.640 ;
        RECT 126.090 170.300 126.350 170.620 ;
        RECT 125.630 159.760 125.890 160.080 ;
        RECT 125.690 159.400 125.830 159.760 ;
        RECT 125.630 159.080 125.890 159.400 ;
        RECT 124.310 151.860 125.370 152.000 ;
        RECT 121.950 148.880 122.210 149.200 ;
        RECT 122.410 148.880 122.670 149.200 ;
        RECT 120.570 148.540 120.830 148.860 ;
        RECT 120.630 146.480 120.770 148.540 ;
        RECT 120.570 146.160 120.830 146.480 ;
        RECT 121.480 146.305 121.760 146.675 ;
        RECT 121.550 146.140 121.690 146.305 ;
        RECT 121.490 145.820 121.750 146.140 ;
        RECT 122.010 144.440 122.150 148.880 ;
        RECT 121.950 144.120 122.210 144.440 ;
        RECT 122.470 144.100 122.610 148.880 ;
        RECT 122.410 143.780 122.670 144.100 ;
        RECT 119.190 143.440 119.450 143.760 ;
        RECT 120.570 142.420 120.830 142.740 ;
        RECT 117.350 140.380 117.610 140.700 ;
        RECT 117.410 139.000 117.550 140.380 ;
        RECT 118.730 139.700 118.990 140.020 ;
        RECT 118.790 139.000 118.930 139.700 ;
        RECT 117.350 138.680 117.610 139.000 ;
        RECT 118.730 138.680 118.990 139.000 ;
        RECT 120.100 138.145 120.380 138.515 ;
        RECT 120.110 138.000 120.370 138.145 ;
        RECT 120.630 137.640 120.770 142.420 ;
        RECT 122.870 141.400 123.130 141.720 ;
        RECT 121.030 140.040 121.290 140.360 ;
        RECT 119.190 137.320 119.450 137.640 ;
        RECT 120.570 137.320 120.830 137.640 ;
        RECT 117.350 135.960 117.610 136.280 ;
        RECT 114.650 130.660 115.250 130.800 ;
        RECT 113.270 130.160 114.790 130.240 ;
        RECT 113.210 130.100 114.790 130.160 ;
        RECT 113.210 129.840 113.470 130.100 ;
        RECT 114.650 129.820 114.790 130.100 ;
        RECT 113.670 129.500 113.930 129.820 ;
        RECT 114.590 129.500 114.850 129.820 ;
        RECT 112.750 128.820 113.010 129.140 ;
        RECT 112.810 127.440 112.950 128.820 ;
        RECT 112.750 127.120 113.010 127.440 ;
        RECT 112.290 122.360 112.550 122.680 ;
        RECT 111.830 121.000 112.090 121.320 ;
        RECT 110.910 118.960 111.170 119.280 ;
        RECT 111.890 115.540 112.030 121.000 ;
        RECT 112.290 116.580 112.550 116.900 ;
        RECT 111.830 115.220 112.090 115.540 ;
        RECT 109.990 113.520 110.250 113.840 ;
        RECT 110.050 111.120 110.190 113.520 ;
        RECT 109.990 110.800 110.250 111.120 ;
        RECT 111.890 107.800 112.030 115.220 ;
        RECT 112.350 111.120 112.490 116.580 ;
        RECT 112.810 116.560 112.950 127.120 ;
        RECT 113.210 124.060 113.470 124.380 ;
        RECT 113.270 121.320 113.410 124.060 ;
        RECT 113.210 121.000 113.470 121.320 ;
        RECT 112.750 116.240 113.010 116.560 ;
        RECT 113.210 111.480 113.470 111.800 ;
        RECT 112.290 110.800 112.550 111.120 ;
        RECT 112.350 108.400 112.490 110.800 ;
        RECT 112.290 108.080 112.550 108.400 ;
        RECT 111.890 107.660 112.490 107.800 ;
        RECT 110.910 105.360 111.170 105.680 ;
        RECT 110.970 100.240 111.110 105.360 ;
        RECT 111.830 104.680 112.090 105.000 ;
        RECT 110.910 99.920 111.170 100.240 ;
        RECT 110.970 99.220 111.110 99.920 ;
        RECT 110.910 98.900 111.170 99.220 ;
        RECT 111.890 93.780 112.030 104.680 ;
        RECT 111.830 93.460 112.090 93.780 ;
        RECT 112.350 92.840 112.490 107.660 ;
        RECT 113.270 99.900 113.410 111.480 ;
        RECT 113.210 99.580 113.470 99.900 ;
        RECT 113.270 97.180 113.410 99.580 ;
        RECT 113.210 97.090 113.470 97.180 ;
        RECT 112.810 96.950 113.470 97.090 ;
        RECT 112.810 94.800 112.950 96.950 ;
        RECT 113.210 96.860 113.470 96.950 ;
        RECT 112.750 94.480 113.010 94.800 ;
        RECT 113.210 94.480 113.470 94.800 ;
        RECT 109.590 92.700 111.570 92.840 ;
        RECT 109.070 91.420 109.330 91.740 ;
        RECT 109.530 91.080 109.790 91.400 ;
        RECT 109.070 90.740 109.330 91.060 ;
        RECT 109.130 89.020 109.270 90.740 ;
        RECT 109.070 88.700 109.330 89.020 ;
        RECT 109.130 86.640 109.270 88.700 ;
        RECT 108.610 86.320 108.870 86.640 ;
        RECT 109.070 86.320 109.330 86.640 ;
        RECT 105.850 85.640 106.110 85.960 ;
        RECT 108.610 85.640 108.870 85.960 ;
        RECT 103.550 83.940 103.810 84.260 ;
        RECT 105.390 83.940 105.650 84.260 ;
        RECT 101.250 83.600 101.510 83.920 ;
        RECT 101.310 82.500 101.450 83.600 ;
        RECT 100.390 82.360 100.990 82.500 ;
        RECT 101.310 82.360 101.910 82.500 ;
        RECT 100.850 80.860 100.990 82.360 ;
        RECT 101.770 81.200 101.910 82.360 ;
        RECT 101.710 80.880 101.970 81.200 ;
        RECT 103.610 80.860 103.750 83.940 ;
        RECT 105.910 83.920 106.050 85.640 ;
        RECT 105.850 83.600 106.110 83.920 ;
        RECT 108.670 82.900 108.810 85.640 ;
        RECT 109.070 85.475 109.330 85.620 ;
        RECT 109.060 85.105 109.340 85.475 ;
        RECT 109.590 83.920 109.730 91.080 ;
        RECT 109.990 89.720 110.250 90.040 ;
        RECT 110.050 84.600 110.190 89.720 ;
        RECT 110.910 89.380 111.170 89.700 ;
        RECT 110.450 88.360 110.710 88.680 ;
        RECT 110.510 86.835 110.650 88.360 ;
        RECT 110.440 86.465 110.720 86.835 ;
        RECT 110.970 86.640 111.110 89.380 ;
        RECT 110.910 86.320 111.170 86.640 ;
        RECT 110.450 86.040 110.710 86.300 ;
        RECT 110.450 85.980 111.110 86.040 ;
        RECT 110.510 85.900 111.110 85.980 ;
        RECT 109.990 84.280 110.250 84.600 ;
        RECT 110.440 84.425 110.720 84.795 ;
        RECT 110.970 84.600 111.110 85.900 ;
        RECT 111.430 84.600 111.570 92.700 ;
        RECT 111.890 92.700 112.490 92.840 ;
        RECT 110.510 83.920 110.650 84.425 ;
        RECT 110.910 84.280 111.170 84.600 ;
        RECT 111.370 84.280 111.630 84.600 ;
        RECT 111.890 84.000 112.030 92.700 ;
        RECT 112.810 90.040 112.950 94.480 ;
        RECT 113.270 91.740 113.410 94.480 ;
        RECT 113.210 91.420 113.470 91.740 ;
        RECT 112.750 89.950 113.010 90.040 ;
        RECT 112.750 89.810 113.410 89.950 ;
        RECT 112.750 89.720 113.010 89.810 ;
        RECT 112.290 89.040 112.550 89.360 ;
        RECT 112.740 89.185 113.020 89.555 ;
        RECT 109.530 83.600 109.790 83.920 ;
        RECT 110.450 83.600 110.710 83.920 ;
        RECT 111.430 83.860 112.030 84.000 ;
        RECT 104.930 82.580 105.190 82.900 ;
        RECT 108.610 82.580 108.870 82.900 ;
        RECT 104.990 81.880 105.130 82.580 ;
        RECT 109.590 82.500 109.730 83.600 ;
        RECT 109.130 82.360 109.730 82.500 ;
        RECT 104.930 81.560 105.190 81.880 ;
        RECT 104.990 80.860 105.130 81.560 ;
        RECT 105.390 81.220 105.650 81.540 ;
        RECT 63.530 80.540 63.790 80.860 ;
        RECT 71.810 80.540 72.070 80.860 ;
        RECT 73.190 80.540 73.450 80.860 ;
        RECT 81.010 80.540 81.270 80.860 ;
        RECT 81.470 80.540 81.730 80.860 ;
        RECT 81.930 80.540 82.190 80.860 ;
        RECT 87.910 80.540 88.170 80.860 ;
        RECT 92.510 80.540 92.770 80.860 ;
        RECT 96.190 80.540 96.450 80.860 ;
        RECT 98.030 80.540 98.290 80.860 ;
        RECT 100.790 80.540 101.050 80.860 ;
        RECT 103.550 80.540 103.810 80.860 ;
        RECT 104.930 80.540 105.190 80.860 ;
        RECT 36.280 79.325 37.820 79.695 ;
        RECT 63.590 72.630 63.730 80.540 ;
        RECT 69.970 79.860 70.230 80.180 ;
        RECT 70.030 72.630 70.170 79.860 ;
        RECT 73.250 72.630 73.390 80.540 ;
        RECT 76.410 79.860 76.670 80.180 ;
        RECT 79.630 79.860 79.890 80.180 ;
        RECT 82.850 79.860 83.110 80.180 ;
        RECT 86.070 79.860 86.330 80.180 ;
        RECT 89.290 79.860 89.550 80.180 ;
        RECT 92.510 79.860 92.770 80.180 ;
        RECT 95.730 79.860 95.990 80.180 ;
        RECT 98.950 79.860 99.210 80.180 ;
        RECT 102.170 79.860 102.430 80.180 ;
        RECT 76.470 72.630 76.610 79.860 ;
        RECT 79.690 72.630 79.830 79.860 ;
        RECT 82.910 72.630 83.050 79.860 ;
        RECT 86.130 72.630 86.270 79.860 ;
        RECT 89.350 72.630 89.490 79.860 ;
        RECT 92.570 72.630 92.710 79.860 ;
        RECT 95.790 72.630 95.930 79.860 ;
        RECT 99.010 72.630 99.150 79.860 ;
        RECT 102.230 72.630 102.370 79.860 ;
        RECT 105.450 72.630 105.590 81.220 ;
        RECT 109.130 81.200 109.270 82.360 ;
        RECT 109.070 80.880 109.330 81.200 ;
        RECT 110.510 80.860 110.650 83.600 ;
        RECT 111.430 82.900 111.570 83.860 ;
        RECT 111.370 82.580 111.630 82.900 ;
        RECT 110.450 80.540 110.710 80.860 ;
        RECT 112.350 80.520 112.490 89.040 ;
        RECT 112.810 86.300 112.950 89.185 ;
        RECT 112.750 85.980 113.010 86.300 ;
        RECT 113.270 85.620 113.410 89.810 ;
        RECT 113.730 85.620 113.870 129.500 ;
        RECT 114.130 128.820 114.390 129.140 ;
        RECT 114.190 124.380 114.330 128.820 ;
        RECT 114.650 126.420 114.790 129.500 ;
        RECT 114.590 126.100 114.850 126.420 ;
        RECT 114.650 124.720 114.790 126.100 ;
        RECT 114.590 124.400 114.850 124.720 ;
        RECT 114.130 124.060 114.390 124.380 ;
        RECT 114.130 115.220 114.390 115.540 ;
        RECT 114.190 113.500 114.330 115.220 ;
        RECT 114.650 113.840 114.790 124.400 ;
        RECT 115.110 123.700 115.250 130.660 ;
        RECT 115.570 130.500 115.710 131.540 ;
        RECT 116.030 131.460 117.090 131.600 ;
        RECT 115.510 130.180 115.770 130.500 ;
        RECT 115.510 126.440 115.770 126.760 ;
        RECT 115.050 123.380 115.310 123.700 ;
        RECT 115.050 118.620 115.310 118.940 ;
        RECT 115.110 116.220 115.250 118.620 ;
        RECT 115.050 115.900 115.310 116.220 ;
        RECT 115.570 113.920 115.710 126.440 ;
        RECT 116.030 115.540 116.170 131.460 ;
        RECT 117.410 130.800 117.550 135.960 ;
        RECT 117.810 134.600 118.070 134.920 ;
        RECT 117.870 133.560 118.010 134.600 ;
        RECT 118.270 134.260 118.530 134.580 ;
        RECT 118.330 133.560 118.470 134.260 ;
        RECT 117.810 133.240 118.070 133.560 ;
        RECT 118.270 133.240 118.530 133.560 ;
        RECT 119.250 132.880 119.390 137.320 ;
        RECT 119.650 136.980 119.910 137.300 ;
        RECT 119.710 136.280 119.850 136.980 ;
        RECT 119.650 135.960 119.910 136.280 ;
        RECT 119.710 135.260 119.850 135.960 ;
        RECT 119.650 134.940 119.910 135.260 ;
        RECT 121.090 134.920 121.230 140.040 ;
        RECT 121.490 138.000 121.750 138.320 ;
        RECT 121.550 136.280 121.690 138.000 ;
        RECT 121.490 135.960 121.750 136.280 ;
        RECT 121.030 134.600 121.290 134.920 ;
        RECT 121.090 132.960 121.230 134.600 ;
        RECT 122.410 134.260 122.670 134.580 ;
        RECT 120.170 132.880 121.230 132.960 ;
        RECT 117.810 132.560 118.070 132.880 ;
        RECT 119.190 132.560 119.450 132.880 ;
        RECT 120.110 132.820 121.230 132.880 ;
        RECT 120.110 132.560 120.370 132.820 ;
        RECT 116.950 130.660 117.550 130.800 ;
        RECT 117.870 130.800 118.010 132.560 ;
        RECT 117.870 130.660 118.470 130.800 ;
        RECT 116.430 127.460 116.690 127.780 ;
        RECT 116.490 119.280 116.630 127.460 ;
        RECT 116.950 123.700 117.090 130.660 ;
        RECT 117.350 129.500 117.610 129.820 ;
        RECT 116.890 123.380 117.150 123.700 ;
        RECT 116.890 120.660 117.150 120.980 ;
        RECT 116.430 118.960 116.690 119.280 ;
        RECT 115.970 115.220 116.230 115.540 ;
        RECT 114.590 113.520 114.850 113.840 ;
        RECT 115.110 113.780 115.710 113.920 ;
        RECT 116.490 113.840 116.630 118.960 ;
        RECT 116.950 118.940 117.090 120.660 ;
        RECT 116.890 118.620 117.150 118.940 ;
        RECT 114.130 113.180 114.390 113.500 ;
        RECT 114.190 106.020 114.330 113.180 ;
        RECT 115.110 108.740 115.250 113.780 ;
        RECT 116.430 113.520 116.690 113.840 ;
        RECT 115.510 113.180 115.770 113.500 ;
        RECT 115.570 111.800 115.710 113.180 ;
        RECT 115.510 111.480 115.770 111.800 ;
        RECT 116.490 111.460 116.630 113.520 ;
        RECT 116.890 111.480 117.150 111.800 ;
        RECT 116.430 111.370 116.690 111.460 ;
        RECT 116.030 111.230 116.690 111.370 ;
        RECT 115.510 109.780 115.770 110.100 ;
        RECT 115.050 108.420 115.310 108.740 ;
        RECT 114.130 105.700 114.390 106.020 ;
        RECT 114.590 105.360 114.850 105.680 ;
        RECT 114.650 99.560 114.790 105.360 ;
        RECT 115.050 104.400 115.310 104.660 ;
        RECT 115.570 104.400 115.710 109.780 ;
        RECT 116.030 108.060 116.170 111.230 ;
        RECT 116.430 111.140 116.690 111.230 ;
        RECT 116.950 110.440 117.090 111.480 ;
        RECT 116.890 110.120 117.150 110.440 ;
        RECT 116.430 108.760 116.690 109.080 ;
        RECT 115.970 107.740 116.230 108.060 ;
        RECT 115.970 105.360 116.230 105.680 ;
        RECT 115.050 104.340 115.710 104.400 ;
        RECT 115.110 104.260 115.710 104.340 ;
        RECT 115.510 101.620 115.770 101.940 ;
        RECT 114.590 99.240 114.850 99.560 ;
        RECT 114.650 97.860 114.790 99.240 ;
        RECT 114.590 97.540 114.850 97.860 ;
        RECT 114.130 94.480 114.390 94.800 ;
        RECT 114.190 89.360 114.330 94.480 ;
        RECT 114.590 93.800 114.850 94.120 ;
        RECT 114.650 89.700 114.790 93.800 ;
        RECT 114.590 89.555 114.850 89.700 ;
        RECT 114.580 89.440 114.860 89.555 ;
        RECT 114.130 89.040 114.390 89.360 ;
        RECT 114.580 89.300 115.250 89.440 ;
        RECT 114.580 89.185 114.860 89.300 ;
        RECT 114.590 88.700 114.850 89.020 ;
        RECT 114.130 88.360 114.390 88.680 ;
        RECT 113.210 85.300 113.470 85.620 ;
        RECT 113.670 85.300 113.930 85.620 ;
        RECT 112.740 84.425 113.020 84.795 ;
        RECT 112.810 83.580 112.950 84.425 ;
        RECT 113.270 83.920 113.410 85.300 ;
        RECT 113.670 84.280 113.930 84.600 ;
        RECT 113.210 83.600 113.470 83.920 ;
        RECT 112.750 83.260 113.010 83.580 ;
        RECT 113.730 81.540 113.870 84.280 ;
        RECT 113.670 81.220 113.930 81.540 ;
        RECT 114.190 80.860 114.330 88.360 ;
        RECT 114.650 86.835 114.790 88.700 ;
        RECT 114.580 86.465 114.860 86.835 ;
        RECT 114.590 85.980 114.850 86.300 ;
        RECT 114.650 82.900 114.790 85.980 ;
        RECT 115.110 84.260 115.250 89.300 ;
        RECT 115.050 83.940 115.310 84.260 ;
        RECT 115.110 83.435 115.250 83.940 ;
        RECT 115.040 83.065 115.320 83.435 ;
        RECT 114.590 82.580 114.850 82.900 ;
        RECT 115.570 80.860 115.710 101.620 ;
        RECT 116.030 99.640 116.170 105.360 ;
        RECT 116.490 105.250 116.630 108.760 ;
        RECT 116.890 107.400 117.150 107.720 ;
        RECT 116.950 106.360 117.090 107.400 ;
        RECT 116.890 106.040 117.150 106.360 ;
        RECT 116.890 105.250 117.150 105.340 ;
        RECT 116.490 105.110 117.150 105.250 ;
        RECT 116.890 105.020 117.150 105.110 ;
        RECT 116.430 104.340 116.690 104.660 ;
        RECT 116.490 102.620 116.630 104.340 ;
        RECT 116.950 102.620 117.090 105.020 ;
        RECT 116.430 102.300 116.690 102.620 ;
        RECT 116.890 102.300 117.150 102.620 ;
        RECT 116.030 99.500 117.090 99.640 ;
        RECT 116.430 98.900 116.690 99.220 ;
        RECT 115.970 96.520 116.230 96.840 ;
        RECT 116.030 95.140 116.170 96.520 ;
        RECT 115.970 94.820 116.230 95.140 ;
        RECT 116.490 94.200 116.630 98.900 ;
        RECT 116.950 95.480 117.090 99.500 ;
        RECT 116.890 95.160 117.150 95.480 ;
        RECT 116.030 94.060 116.630 94.200 ;
        RECT 116.030 82.500 116.170 94.060 ;
        RECT 116.950 92.760 117.090 95.160 ;
        RECT 116.890 92.440 117.150 92.760 ;
        RECT 116.420 85.105 116.700 85.475 ;
        RECT 116.490 83.920 116.630 85.105 ;
        RECT 117.410 84.600 117.550 129.500 ;
        RECT 117.810 124.060 118.070 124.380 ;
        RECT 117.870 88.340 118.010 124.060 ;
        RECT 118.330 118.260 118.470 130.660 ;
        RECT 119.250 130.500 119.390 132.560 ;
        RECT 118.720 129.985 119.000 130.355 ;
        RECT 119.190 130.180 119.450 130.500 ;
        RECT 118.790 129.820 118.930 129.985 ;
        RECT 121.090 129.820 121.230 132.820 ;
        RECT 121.950 132.220 122.210 132.540 ;
        RECT 118.730 129.500 118.990 129.820 ;
        RECT 118.790 128.120 118.930 129.500 ;
        RECT 120.100 129.305 120.380 129.675 ;
        RECT 121.030 129.500 121.290 129.820 ;
        RECT 118.730 127.800 118.990 128.120 ;
        RECT 118.790 124.720 118.930 127.800 ;
        RECT 118.730 124.400 118.990 124.720 ;
        RECT 119.190 124.060 119.450 124.380 ;
        RECT 119.650 124.060 119.910 124.380 ;
        RECT 119.250 119.870 119.390 124.060 ;
        RECT 119.710 122.680 119.850 124.060 ;
        RECT 119.650 122.360 119.910 122.680 ;
        RECT 119.650 119.870 119.910 119.960 ;
        RECT 119.250 119.730 119.910 119.870 ;
        RECT 119.650 119.640 119.910 119.730 ;
        RECT 118.270 117.940 118.530 118.260 ;
        RECT 119.650 112.500 119.910 112.820 ;
        RECT 119.710 111.120 119.850 112.500 ;
        RECT 118.730 111.030 118.990 111.120 ;
        RECT 118.330 110.890 118.990 111.030 ;
        RECT 118.330 107.380 118.470 110.890 ;
        RECT 118.730 110.800 118.990 110.890 ;
        RECT 119.650 110.800 119.910 111.120 ;
        RECT 118.270 107.060 118.530 107.380 ;
        RECT 118.330 102.620 118.470 107.060 ;
        RECT 119.190 105.360 119.450 105.680 ;
        RECT 119.250 102.960 119.390 105.360 ;
        RECT 119.710 103.640 119.850 110.800 ;
        RECT 119.650 103.320 119.910 103.640 ;
        RECT 120.170 103.200 120.310 129.305 ;
        RECT 121.090 126.760 121.230 129.500 ;
        RECT 121.490 127.120 121.750 127.440 ;
        RECT 121.030 126.440 121.290 126.760 ;
        RECT 121.550 125.400 121.690 127.120 ;
        RECT 121.490 125.080 121.750 125.400 ;
        RECT 121.030 123.720 121.290 124.040 ;
        RECT 121.090 120.890 121.230 123.720 ;
        RECT 121.490 121.570 121.750 121.660 ;
        RECT 122.010 121.570 122.150 132.220 ;
        RECT 122.470 129.140 122.610 134.260 ;
        RECT 122.410 128.820 122.670 129.140 ;
        RECT 122.410 126.100 122.670 126.420 ;
        RECT 122.470 124.380 122.610 126.100 ;
        RECT 122.930 125.060 123.070 141.400 ;
        RECT 122.870 124.740 123.130 125.060 ;
        RECT 122.410 124.060 122.670 124.380 ;
        RECT 123.790 124.060 124.050 124.380 ;
        RECT 123.330 122.360 123.590 122.680 ;
        RECT 121.490 121.430 122.150 121.570 ;
        RECT 121.490 121.340 121.750 121.430 ;
        RECT 121.090 120.750 121.690 120.890 ;
        RECT 121.550 116.560 121.690 120.750 ;
        RECT 121.490 116.240 121.750 116.560 ;
        RECT 121.030 107.400 121.290 107.720 ;
        RECT 121.090 106.020 121.230 107.400 ;
        RECT 121.030 105.875 121.290 106.020 ;
        RECT 121.020 105.505 121.300 105.875 ;
        RECT 121.550 105.250 121.690 116.240 ;
        RECT 122.010 116.220 122.150 121.430 ;
        RECT 123.390 119.620 123.530 122.360 ;
        RECT 123.850 122.000 123.990 124.060 ;
        RECT 123.790 121.680 124.050 122.000 ;
        RECT 123.330 119.300 123.590 119.620 ;
        RECT 121.950 115.900 122.210 116.220 ;
        RECT 122.010 106.360 122.150 115.900 ;
        RECT 122.410 113.860 122.670 114.180 ;
        RECT 122.470 111.120 122.610 113.860 ;
        RECT 122.870 111.480 123.130 111.800 ;
        RECT 122.410 110.800 122.670 111.120 ;
        RECT 122.410 107.060 122.670 107.380 ;
        RECT 121.950 106.040 122.210 106.360 ;
        RECT 121.090 105.110 121.690 105.250 ;
        RECT 120.170 103.060 120.770 103.200 ;
        RECT 119.190 102.640 119.450 102.960 ;
        RECT 118.270 102.300 118.530 102.620 ;
        RECT 119.250 102.360 119.390 102.640 ;
        RECT 118.330 100.240 118.470 102.300 ;
        RECT 119.250 102.220 120.310 102.360 ;
        RECT 120.630 102.280 120.770 103.060 ;
        RECT 118.730 101.620 118.990 101.940 ;
        RECT 118.270 99.920 118.530 100.240 ;
        RECT 118.330 96.500 118.470 99.920 ;
        RECT 118.790 96.840 118.930 101.620 ;
        RECT 119.190 99.920 119.450 100.240 ;
        RECT 118.730 96.520 118.990 96.840 ;
        RECT 118.270 96.180 118.530 96.500 ;
        RECT 119.250 96.355 119.390 99.920 ;
        RECT 119.650 98.900 119.910 99.220 ;
        RECT 119.710 96.840 119.850 98.900 ;
        RECT 119.650 96.520 119.910 96.840 ;
        RECT 119.180 95.985 119.460 96.355 ;
        RECT 118.270 95.160 118.530 95.480 ;
        RECT 118.330 94.800 118.470 95.160 ;
        RECT 118.270 94.480 118.530 94.800 ;
        RECT 119.190 94.480 119.450 94.800 ;
        RECT 119.250 92.760 119.390 94.480 ;
        RECT 119.190 92.440 119.450 92.760 ;
        RECT 119.710 91.400 119.850 96.520 ;
        RECT 120.170 91.740 120.310 102.220 ;
        RECT 120.570 101.960 120.830 102.280 ;
        RECT 120.630 100.240 120.770 101.960 ;
        RECT 120.570 99.920 120.830 100.240 ;
        RECT 120.570 99.240 120.830 99.560 ;
        RECT 120.630 98.200 120.770 99.240 ;
        RECT 120.570 97.880 120.830 98.200 ;
        RECT 120.570 94.480 120.830 94.800 ;
        RECT 120.630 92.760 120.770 94.480 ;
        RECT 120.570 92.440 120.830 92.760 ;
        RECT 120.110 91.420 120.370 91.740 ;
        RECT 119.650 91.080 119.910 91.400 ;
        RECT 119.710 90.040 119.850 91.080 ;
        RECT 120.630 91.060 120.770 92.440 ;
        RECT 121.090 92.420 121.230 105.110 ;
        RECT 122.470 102.280 122.610 107.060 ;
        RECT 122.930 105.000 123.070 111.480 ;
        RECT 122.870 104.680 123.130 105.000 ;
        RECT 122.410 101.960 122.670 102.280 ;
        RECT 122.410 97.880 122.670 98.200 ;
        RECT 122.470 96.500 122.610 97.880 ;
        RECT 122.870 96.860 123.130 97.180 ;
        RECT 122.410 96.180 122.670 96.500 ;
        RECT 122.410 95.160 122.670 95.480 ;
        RECT 121.030 92.100 121.290 92.420 ;
        RECT 120.570 90.740 120.830 91.060 ;
        RECT 119.650 89.720 119.910 90.040 ;
        RECT 119.190 89.380 119.450 89.700 ;
        RECT 118.730 89.040 118.990 89.360 ;
        RECT 117.810 88.020 118.070 88.340 ;
        RECT 117.810 85.300 118.070 85.620 ;
        RECT 117.350 84.280 117.610 84.600 ;
        RECT 116.890 83.940 117.150 84.260 ;
        RECT 116.430 83.600 116.690 83.920 ;
        RECT 116.950 82.900 117.090 83.940 ;
        RECT 117.870 83.920 118.010 85.300 ;
        RECT 118.790 83.920 118.930 89.040 ;
        RECT 119.250 84.795 119.390 89.380 ;
        RECT 119.710 86.300 119.850 89.720 ;
        RECT 120.630 89.360 120.770 90.740 ;
        RECT 122.470 90.040 122.610 95.160 ;
        RECT 122.930 95.140 123.070 96.860 ;
        RECT 122.870 94.820 123.130 95.140 ;
        RECT 122.410 89.720 122.670 90.040 ;
        RECT 122.470 89.360 122.610 89.720 ;
        RECT 120.570 89.040 120.830 89.360 ;
        RECT 122.410 89.040 122.670 89.360 ;
        RECT 122.930 86.640 123.070 94.820 ;
        RECT 123.390 89.020 123.530 119.300 ;
        RECT 123.850 117.240 123.990 121.680 ;
        RECT 124.310 118.600 124.450 151.860 ;
        RECT 124.710 148.880 124.970 149.200 ;
        RECT 125.170 148.880 125.430 149.200 ;
        RECT 124.770 129.675 124.910 148.880 ;
        RECT 125.230 148.520 125.370 148.880 ;
        RECT 125.170 148.200 125.430 148.520 ;
        RECT 125.230 146.820 125.370 148.200 ;
        RECT 125.170 146.500 125.430 146.820 ;
        RECT 125.630 146.160 125.890 146.480 ;
        RECT 125.170 145.820 125.430 146.140 ;
        RECT 125.230 143.080 125.370 145.820 ;
        RECT 125.170 142.760 125.430 143.080 ;
        RECT 125.690 138.515 125.830 146.160 ;
        RECT 126.150 141.720 126.290 170.300 ;
        RECT 126.610 162.120 126.750 171.320 ;
        RECT 127.530 170.960 127.670 171.320 ;
        RECT 127.470 170.640 127.730 170.960 ;
        RECT 128.390 170.640 128.650 170.960 ;
        RECT 129.770 170.640 130.030 170.960 ;
        RECT 127.530 169.940 127.670 170.640 ;
        RECT 127.470 169.620 127.730 169.940 ;
        RECT 126.550 161.800 126.810 162.120 ;
        RECT 126.610 149.450 126.750 161.800 ;
        RECT 127.010 153.980 127.270 154.300 ;
        RECT 127.070 151.580 127.210 153.980 ;
        RECT 127.010 151.260 127.270 151.580 ;
        RECT 127.010 149.450 127.270 149.540 ;
        RECT 126.610 149.310 127.270 149.450 ;
        RECT 127.010 149.220 127.270 149.310 ;
        RECT 127.530 148.520 127.670 169.620 ;
        RECT 128.450 168.580 128.590 170.640 ;
        RECT 128.390 168.260 128.650 168.580 ;
        RECT 129.830 167.220 129.970 170.640 ;
        RECT 129.770 166.900 130.030 167.220 ;
        RECT 130.750 165.520 130.890 173.360 ;
        RECT 138.110 173.340 138.250 175.060 ;
        RECT 139.030 174.555 139.170 177.780 ;
        RECT 138.960 174.185 139.240 174.555 ;
        RECT 138.050 173.020 138.310 173.340 ;
        RECT 135.290 172.680 135.550 173.000 ;
        RECT 135.350 171.640 135.490 172.680 ;
        RECT 139.950 171.640 140.090 178.460 ;
        RECT 140.870 177.955 141.010 180.500 ;
        RECT 140.800 177.585 141.080 177.955 ;
        RECT 141.730 177.780 141.990 178.100 ;
        RECT 140.810 172.340 141.070 172.660 ;
        RECT 135.290 171.320 135.550 171.640 ;
        RECT 139.890 171.320 140.150 171.640 ;
        RECT 140.870 170.960 141.010 172.340 ;
        RECT 141.790 171.155 141.930 177.780 ;
        RECT 140.810 170.640 141.070 170.960 ;
        RECT 141.720 170.785 142.000 171.155 ;
        RECT 131.610 167.580 131.870 167.900 ;
        RECT 131.150 166.900 131.410 167.220 ;
        RECT 130.690 165.200 130.950 165.520 ;
        RECT 129.770 162.480 130.030 162.800 ;
        RECT 127.930 162.140 128.190 162.460 ;
        RECT 127.990 160.760 128.130 162.140 ;
        RECT 127.930 160.440 128.190 160.760 ;
        RECT 129.830 158.040 129.970 162.480 ;
        RECT 130.230 162.140 130.490 162.460 ;
        RECT 129.770 157.720 130.030 158.040 ;
        RECT 128.390 154.320 128.650 154.640 ;
        RECT 128.450 153.620 128.590 154.320 ;
        RECT 128.390 153.300 128.650 153.620 ;
        RECT 129.770 153.300 130.030 153.620 ;
        RECT 129.830 149.200 129.970 153.300 ;
        RECT 127.930 148.880 128.190 149.200 ;
        RECT 129.770 148.880 130.030 149.200 ;
        RECT 127.470 148.200 127.730 148.520 ;
        RECT 126.090 141.400 126.350 141.720 ;
        RECT 127.990 140.020 128.130 148.880 ;
        RECT 130.290 146.140 130.430 162.140 ;
        RECT 130.750 160.080 130.890 165.200 ;
        RECT 130.690 159.760 130.950 160.080 ;
        RECT 130.750 157.020 130.890 159.760 ;
        RECT 130.690 156.700 130.950 157.020 ;
        RECT 130.750 154.640 130.890 156.700 ;
        RECT 130.690 154.320 130.950 154.640 ;
        RECT 131.210 151.320 131.350 166.900 ;
        RECT 131.670 166.200 131.810 167.580 ;
        RECT 132.520 167.385 132.800 167.755 ;
        RECT 138.510 167.580 138.770 167.900 ;
        RECT 132.590 167.220 132.730 167.385 ;
        RECT 132.530 166.900 132.790 167.220 ;
        RECT 133.910 166.900 134.170 167.220 ;
        RECT 134.370 166.900 134.630 167.220 ;
        RECT 131.610 165.880 131.870 166.200 ;
        RECT 133.970 165.860 134.110 166.900 ;
        RECT 133.910 165.540 134.170 165.860 ;
        RECT 134.430 163.480 134.570 166.900 ;
        RECT 138.570 166.200 138.710 167.580 ;
        RECT 138.510 165.880 138.770 166.200 ;
        RECT 140.810 165.880 141.070 166.200 ;
        RECT 136.210 165.540 136.470 165.860 ;
        RECT 134.370 163.160 134.630 163.480 ;
        RECT 132.990 161.800 133.250 162.120 ;
        RECT 132.070 156.020 132.330 156.340 ;
        RECT 132.130 154.640 132.270 156.020 ;
        RECT 132.070 154.320 132.330 154.640 ;
        RECT 131.210 151.180 131.810 151.320 ;
        RECT 130.690 150.580 130.950 150.900 ;
        RECT 131.150 150.580 131.410 150.900 ;
        RECT 130.750 149.880 130.890 150.580 ;
        RECT 131.210 149.880 131.350 150.580 ;
        RECT 130.690 149.560 130.950 149.880 ;
        RECT 131.150 149.560 131.410 149.880 ;
        RECT 131.150 148.880 131.410 149.200 ;
        RECT 130.690 146.840 130.950 147.160 ;
        RECT 130.230 145.820 130.490 146.140 ;
        RECT 128.390 145.480 128.650 145.800 ;
        RECT 128.850 145.480 129.110 145.800 ;
        RECT 128.450 144.440 128.590 145.480 ;
        RECT 128.390 144.120 128.650 144.440 ;
        RECT 128.910 140.700 129.050 145.480 ;
        RECT 130.750 144.100 130.890 146.840 ;
        RECT 130.690 143.780 130.950 144.100 ;
        RECT 128.850 140.380 129.110 140.700 ;
        RECT 127.930 139.700 128.190 140.020 ;
        RECT 128.910 139.000 129.050 140.380 ;
        RECT 128.850 138.680 129.110 139.000 ;
        RECT 125.620 138.145 125.900 138.515 ;
        RECT 130.690 138.340 130.950 138.660 ;
        RECT 126.550 136.980 126.810 137.300 ;
        RECT 126.610 134.920 126.750 136.980 ;
        RECT 127.930 135.620 128.190 135.940 ;
        RECT 127.990 134.920 128.130 135.620 ;
        RECT 128.850 134.940 129.110 135.260 ;
        RECT 126.550 134.600 126.810 134.920 ;
        RECT 127.930 134.600 128.190 134.920 ;
        RECT 125.630 134.260 125.890 134.580 ;
        RECT 125.690 133.220 125.830 134.260 ;
        RECT 125.630 132.900 125.890 133.220 ;
        RECT 127.990 130.800 128.130 134.600 ;
        RECT 127.990 130.660 128.590 130.800 ;
        RECT 124.700 129.305 124.980 129.675 ;
        RECT 125.170 129.500 125.430 129.820 ;
        RECT 125.230 122.680 125.370 129.500 ;
        RECT 126.550 129.160 126.810 129.480 ;
        RECT 126.610 125.400 126.750 129.160 ;
        RECT 127.930 128.820 128.190 129.140 ;
        RECT 127.990 126.420 128.130 128.820 ;
        RECT 127.930 126.100 128.190 126.420 ;
        RECT 126.550 125.080 126.810 125.400 ;
        RECT 126.610 124.040 126.750 125.080 ;
        RECT 127.990 124.720 128.130 126.100 ;
        RECT 127.930 124.400 128.190 124.720 ;
        RECT 126.550 123.720 126.810 124.040 ;
        RECT 125.170 122.360 125.430 122.680 ;
        RECT 124.250 118.280 124.510 118.600 ;
        RECT 123.790 116.920 124.050 117.240 ;
        RECT 123.850 113.500 123.990 116.920 ;
        RECT 126.090 113.860 126.350 114.180 ;
        RECT 123.790 113.180 124.050 113.500 ;
        RECT 123.790 110.800 124.050 111.120 ;
        RECT 123.850 107.380 123.990 110.800 ;
        RECT 126.150 110.780 126.290 113.860 ;
        RECT 126.610 113.160 126.750 123.720 ;
        RECT 128.450 122.340 128.590 130.660 ;
        RECT 128.910 129.820 129.050 134.940 ;
        RECT 130.230 134.830 130.490 134.920 ;
        RECT 130.750 134.830 130.890 138.340 ;
        RECT 130.230 134.690 130.890 134.830 ;
        RECT 130.230 134.600 130.490 134.690 ;
        RECT 129.310 132.900 129.570 133.220 ;
        RECT 129.370 130.500 129.510 132.900 ;
        RECT 129.770 132.560 130.030 132.880 ;
        RECT 130.230 132.560 130.490 132.880 ;
        RECT 129.830 130.840 129.970 132.560 ;
        RECT 129.770 130.520 130.030 130.840 ;
        RECT 129.310 130.180 129.570 130.500 ;
        RECT 128.850 129.500 129.110 129.820 ;
        RECT 128.910 124.720 129.050 129.500 ;
        RECT 130.290 127.780 130.430 132.560 ;
        RECT 130.750 132.540 130.890 134.690 ;
        RECT 130.690 132.220 130.950 132.540 ;
        RECT 131.210 130.160 131.350 148.880 ;
        RECT 131.670 135.260 131.810 151.180 ;
        RECT 132.070 139.700 132.330 140.020 ;
        RECT 132.130 138.320 132.270 139.700 ;
        RECT 132.070 138.000 132.330 138.320 ;
        RECT 132.530 138.000 132.790 138.320 ;
        RECT 132.590 135.940 132.730 138.000 ;
        RECT 132.530 135.620 132.790 135.940 ;
        RECT 131.610 134.940 131.870 135.260 ;
        RECT 132.070 134.940 132.330 135.260 ;
        RECT 131.610 134.260 131.870 134.580 ;
        RECT 131.670 132.880 131.810 134.260 ;
        RECT 132.130 132.880 132.270 134.940 ;
        RECT 132.530 134.600 132.790 134.920 ;
        RECT 132.590 133.560 132.730 134.600 ;
        RECT 132.530 133.240 132.790 133.560 ;
        RECT 131.610 132.560 131.870 132.880 ;
        RECT 132.070 132.560 132.330 132.880 ;
        RECT 132.590 130.800 132.730 133.240 ;
        RECT 131.670 130.660 132.730 130.800 ;
        RECT 131.150 129.840 131.410 130.160 ;
        RECT 130.230 127.460 130.490 127.780 ;
        RECT 131.150 126.780 131.410 127.100 ;
        RECT 130.230 126.440 130.490 126.760 ;
        RECT 129.770 124.740 130.030 125.060 ;
        RECT 128.850 124.400 129.110 124.720 ;
        RECT 128.390 122.020 128.650 122.340 ;
        RECT 128.450 117.320 128.590 122.020 ;
        RECT 128.910 122.000 129.050 124.400 ;
        RECT 129.830 122.000 129.970 124.740 ;
        RECT 130.290 124.720 130.430 126.440 ;
        RECT 130.230 124.400 130.490 124.720 ;
        RECT 130.290 122.680 130.430 124.400 ;
        RECT 130.230 122.360 130.490 122.680 ;
        RECT 128.850 121.680 129.110 122.000 ;
        RECT 129.770 121.680 130.030 122.000 ;
        RECT 129.310 117.940 129.570 118.260 ;
        RECT 128.450 117.180 129.050 117.320 ;
        RECT 128.390 116.240 128.650 116.560 ;
        RECT 128.450 114.520 128.590 116.240 ;
        RECT 128.390 114.200 128.650 114.520 ;
        RECT 128.910 113.840 129.050 117.180 ;
        RECT 128.850 113.520 129.110 113.840 ;
        RECT 126.550 112.840 126.810 113.160 ;
        RECT 126.090 110.460 126.350 110.780 ;
        RECT 123.790 107.060 124.050 107.380 ;
        RECT 124.250 105.020 124.510 105.340 ;
        RECT 125.170 105.020 125.430 105.340 ;
        RECT 124.310 102.960 124.450 105.020 ;
        RECT 124.250 102.640 124.510 102.960 ;
        RECT 125.230 99.900 125.370 105.020 ;
        RECT 126.610 102.620 126.750 112.840 ;
        RECT 128.910 111.800 129.050 113.520 ;
        RECT 129.370 113.500 129.510 117.940 ;
        RECT 130.290 117.320 130.430 122.360 ;
        RECT 130.690 121.680 130.950 122.000 ;
        RECT 130.750 121.320 130.890 121.680 ;
        RECT 131.210 121.320 131.350 126.780 ;
        RECT 131.670 124.380 131.810 130.660 ;
        RECT 132.530 127.120 132.790 127.440 ;
        RECT 132.590 124.380 132.730 127.120 ;
        RECT 131.610 124.060 131.870 124.380 ;
        RECT 132.530 124.060 132.790 124.380 ;
        RECT 133.050 122.000 133.190 161.800 ;
        RECT 133.450 161.460 133.710 161.780 ;
        RECT 133.910 161.460 134.170 161.780 ;
        RECT 134.830 161.460 135.090 161.780 ;
        RECT 133.510 157.360 133.650 161.460 ;
        RECT 133.970 160.420 134.110 161.460 ;
        RECT 133.910 160.100 134.170 160.420 ;
        RECT 133.450 157.040 133.710 157.360 ;
        RECT 134.370 156.020 134.630 156.340 ;
        RECT 134.430 148.520 134.570 156.020 ;
        RECT 134.370 148.200 134.630 148.520 ;
        RECT 134.890 148.180 135.030 161.460 ;
        RECT 135.750 153.980 136.010 154.300 ;
        RECT 135.810 148.520 135.950 153.980 ;
        RECT 135.750 148.200 136.010 148.520 ;
        RECT 134.830 147.860 135.090 148.180 ;
        RECT 133.450 145.140 133.710 145.460 ;
        RECT 133.510 144.440 133.650 145.140 ;
        RECT 133.450 144.120 133.710 144.440 ;
        RECT 136.270 142.740 136.410 165.540 ;
        RECT 139.430 165.200 139.690 165.520 ;
        RECT 138.510 164.180 138.770 164.500 ;
        RECT 137.590 162.140 137.850 162.460 ;
        RECT 137.650 160.760 137.790 162.140 ;
        RECT 137.590 160.440 137.850 160.760 ;
        RECT 138.570 160.080 138.710 164.180 ;
        RECT 138.960 163.985 139.240 164.355 ;
        RECT 139.030 160.760 139.170 163.985 ;
        RECT 139.490 162.460 139.630 165.200 ;
        RECT 139.430 162.140 139.690 162.460 ;
        RECT 140.870 160.955 141.010 165.880 ;
        RECT 138.970 160.440 139.230 160.760 ;
        RECT 140.800 160.585 141.080 160.955 ;
        RECT 138.510 159.760 138.770 160.080 ;
        RECT 139.890 159.760 140.150 160.080 ;
        RECT 137.590 156.700 137.850 157.020 ;
        RECT 137.650 155.320 137.790 156.700 ;
        RECT 139.950 155.320 140.090 159.760 ;
        RECT 140.810 158.740 141.070 159.060 ;
        RECT 140.870 157.555 141.010 158.740 ;
        RECT 140.800 157.185 141.080 157.555 ;
        RECT 137.590 155.000 137.850 155.320 ;
        RECT 139.890 155.000 140.150 155.320 ;
        RECT 140.800 153.785 141.080 154.155 ;
        RECT 140.810 153.640 141.070 153.785 ;
        RECT 139.430 150.580 139.690 150.900 ;
        RECT 139.490 149.200 139.630 150.580 ;
        RECT 142.180 150.385 142.460 150.755 ;
        RECT 139.430 148.880 139.690 149.200 ;
        RECT 140.350 148.880 140.610 149.200 ;
        RECT 136.670 146.160 136.930 146.480 ;
        RECT 136.730 143.760 136.870 146.160 ;
        RECT 138.050 145.820 138.310 146.140 ;
        RECT 138.110 144.440 138.250 145.820 ;
        RECT 138.970 145.140 139.230 145.460 ;
        RECT 138.050 144.120 138.310 144.440 ;
        RECT 139.030 143.955 139.170 145.140 ;
        RECT 136.670 143.440 136.930 143.760 ;
        RECT 138.960 143.585 139.240 143.955 ;
        RECT 136.210 142.420 136.470 142.740 ;
        RECT 133.910 140.380 134.170 140.700 ;
        RECT 133.450 140.040 133.710 140.360 ;
        RECT 133.510 139.000 133.650 140.040 ;
        RECT 133.450 138.680 133.710 139.000 ;
        RECT 133.970 138.515 134.110 140.380 ;
        RECT 140.410 140.020 140.550 148.880 ;
        RECT 140.810 147.860 141.070 148.180 ;
        RECT 140.870 147.355 141.010 147.860 ;
        RECT 140.800 146.985 141.080 147.355 ;
        RECT 142.250 147.160 142.390 150.385 ;
        RECT 142.190 146.840 142.450 147.160 ;
        RECT 140.800 140.185 141.080 140.555 ;
        RECT 140.350 139.700 140.610 140.020 ;
        RECT 138.970 138.680 139.230 139.000 ;
        RECT 133.900 138.145 134.180 138.515 ;
        RECT 134.370 138.340 134.630 138.660 ;
        RECT 133.970 135.260 134.110 138.145 ;
        RECT 133.910 134.940 134.170 135.260 ;
        RECT 133.910 130.180 134.170 130.500 ;
        RECT 133.450 129.840 133.710 130.160 ;
        RECT 132.990 121.680 133.250 122.000 ;
        RECT 130.690 121.000 130.950 121.320 ;
        RECT 131.150 121.000 131.410 121.320 ;
        RECT 129.830 117.180 130.430 117.320 ;
        RECT 129.310 113.180 129.570 113.500 ;
        RECT 127.010 111.480 127.270 111.800 ;
        RECT 128.850 111.480 129.110 111.800 ;
        RECT 126.550 102.300 126.810 102.620 ;
        RECT 127.070 102.280 127.210 111.480 ;
        RECT 127.470 110.800 127.730 111.120 ;
        RECT 128.850 111.030 129.110 111.120 ;
        RECT 129.830 111.030 129.970 117.180 ;
        RECT 130.230 116.470 130.490 116.560 ;
        RECT 130.750 116.470 130.890 121.000 ;
        RECT 131.210 116.560 131.350 121.000 ;
        RECT 132.070 118.620 132.330 118.940 ;
        RECT 131.610 118.280 131.870 118.600 ;
        RECT 130.230 116.330 130.890 116.470 ;
        RECT 130.230 116.240 130.490 116.330 ;
        RECT 131.150 116.240 131.410 116.560 ;
        RECT 131.210 111.120 131.350 116.240 ;
        RECT 128.850 110.890 129.970 111.030 ;
        RECT 128.850 110.800 129.110 110.890 ;
        RECT 127.530 108.060 127.670 110.800 ;
        RECT 129.370 110.440 129.510 110.890 ;
        RECT 130.690 110.800 130.950 111.120 ;
        RECT 131.150 110.800 131.410 111.120 ;
        RECT 130.750 110.520 130.890 110.800 ;
        RECT 131.670 110.520 131.810 118.280 ;
        RECT 132.130 117.000 132.270 118.620 ;
        RECT 132.130 116.860 133.190 117.000 ;
        RECT 129.310 110.120 129.570 110.440 ;
        RECT 130.750 110.380 132.730 110.520 ;
        RECT 129.370 108.060 129.510 110.120 ;
        RECT 131.610 108.080 131.870 108.400 ;
        RECT 127.470 107.740 127.730 108.060 ;
        RECT 129.310 107.740 129.570 108.060 ;
        RECT 130.690 107.740 130.950 108.060 ;
        RECT 127.010 101.960 127.270 102.280 ;
        RECT 127.530 101.000 127.670 107.740 ;
        RECT 128.390 105.700 128.650 106.020 ;
        RECT 128.450 105.195 128.590 105.700 ;
        RECT 129.370 105.680 129.510 107.740 ;
        RECT 129.310 105.360 129.570 105.680 ;
        RECT 130.750 105.250 130.890 107.740 ;
        RECT 131.150 107.060 131.410 107.380 ;
        RECT 131.210 106.020 131.350 107.060 ;
        RECT 131.150 105.700 131.410 106.020 ;
        RECT 131.670 105.680 131.810 108.080 ;
        RECT 132.070 107.400 132.330 107.720 ;
        RECT 132.130 105.680 132.270 107.400 ;
        RECT 131.610 105.360 131.870 105.680 ;
        RECT 132.070 105.360 132.330 105.680 ;
        RECT 128.380 104.825 128.660 105.195 ;
        RECT 130.750 105.110 131.350 105.250 ;
        RECT 127.070 100.860 127.670 101.000 ;
        RECT 127.070 100.240 127.210 100.860 ;
        RECT 128.450 100.240 128.590 104.825 ;
        RECT 129.310 104.680 129.570 105.000 ;
        RECT 129.370 102.960 129.510 104.680 ;
        RECT 129.310 102.640 129.570 102.960 ;
        RECT 127.010 99.920 127.270 100.240 ;
        RECT 127.470 99.920 127.730 100.240 ;
        RECT 127.930 99.920 128.190 100.240 ;
        RECT 128.390 99.920 128.650 100.240 ;
        RECT 130.690 100.150 130.950 100.240 ;
        RECT 131.210 100.150 131.350 105.110 ;
        RECT 130.690 100.010 131.350 100.150 ;
        RECT 130.690 99.920 130.950 100.010 ;
        RECT 124.710 99.580 124.970 99.900 ;
        RECT 125.170 99.580 125.430 99.900 ;
        RECT 124.770 98.395 124.910 99.580 ;
        RECT 124.700 98.025 124.980 98.395 ;
        RECT 125.230 97.180 125.370 99.580 ;
        RECT 125.170 96.860 125.430 97.180 ;
        RECT 127.070 94.800 127.210 99.920 ;
        RECT 127.530 98.200 127.670 99.920 ;
        RECT 127.470 97.880 127.730 98.200 ;
        RECT 127.010 94.480 127.270 94.800 ;
        RECT 127.070 91.740 127.210 94.480 ;
        RECT 127.990 94.460 128.130 99.920 ;
        RECT 130.690 97.540 130.950 97.860 ;
        RECT 128.390 96.240 128.650 96.500 ;
        RECT 128.390 96.180 129.050 96.240 ;
        RECT 129.310 96.180 129.570 96.500 ;
        RECT 130.230 96.180 130.490 96.500 ;
        RECT 128.450 96.100 129.050 96.180 ;
        RECT 128.390 94.820 128.650 95.140 ;
        RECT 127.930 94.140 128.190 94.460 ;
        RECT 127.930 93.460 128.190 93.780 ;
        RECT 127.990 92.080 128.130 93.460 ;
        RECT 128.450 92.080 128.590 94.820 ;
        RECT 127.930 91.760 128.190 92.080 ;
        RECT 128.390 91.760 128.650 92.080 ;
        RECT 127.010 91.420 127.270 91.740 ;
        RECT 127.470 90.970 127.730 91.060 ;
        RECT 127.070 90.830 127.730 90.970 ;
        RECT 127.070 90.040 127.210 90.830 ;
        RECT 127.470 90.740 127.730 90.830 ;
        RECT 124.710 89.720 124.970 90.040 ;
        RECT 127.010 89.720 127.270 90.040 ;
        RECT 127.470 89.720 127.730 90.040 ;
        RECT 123.330 88.700 123.590 89.020 ;
        RECT 124.250 88.020 124.510 88.340 ;
        RECT 122.870 86.320 123.130 86.640 ;
        RECT 119.650 85.980 119.910 86.300 ;
        RECT 119.180 84.425 119.460 84.795 ;
        RECT 117.350 83.600 117.610 83.920 ;
        RECT 117.810 83.600 118.070 83.920 ;
        RECT 118.730 83.600 118.990 83.920 ;
        RECT 117.410 83.435 117.550 83.600 ;
        RECT 117.340 83.065 117.620 83.435 ;
        RECT 116.890 82.580 117.150 82.900 ;
        RECT 117.350 82.580 117.610 82.900 ;
        RECT 116.030 82.360 116.630 82.500 ;
        RECT 116.490 81.200 116.630 82.360 ;
        RECT 116.430 80.880 116.690 81.200 ;
        RECT 117.410 80.860 117.550 82.580 ;
        RECT 114.130 80.540 114.390 80.860 ;
        RECT 115.510 80.540 115.770 80.860 ;
        RECT 117.350 80.540 117.610 80.860 ;
        RECT 112.290 80.200 112.550 80.520 ;
        RECT 117.870 80.180 118.010 83.600 ;
        RECT 119.710 82.900 119.850 85.980 ;
        RECT 121.030 85.640 121.290 85.960 ;
        RECT 121.090 84.600 121.230 85.640 ;
        RECT 122.930 84.600 123.070 86.320 ;
        RECT 124.310 86.300 124.450 88.020 ;
        RECT 124.250 85.980 124.510 86.300 ;
        RECT 121.030 84.280 121.290 84.600 ;
        RECT 122.870 84.280 123.130 84.600 ;
        RECT 124.250 84.280 124.510 84.600 ;
        RECT 122.400 83.745 122.680 84.115 ;
        RECT 124.310 83.920 124.450 84.280 ;
        RECT 122.410 83.600 122.670 83.745 ;
        RECT 123.330 83.600 123.590 83.920 ;
        RECT 124.250 83.600 124.510 83.920 ;
        RECT 119.650 82.580 119.910 82.900 ;
        RECT 118.270 81.560 118.530 81.880 ;
        RECT 109.070 79.860 109.330 80.180 ;
        RECT 111.830 79.860 112.090 80.180 ;
        RECT 115.050 79.860 115.310 80.180 ;
        RECT 117.810 79.860 118.070 80.180 ;
        RECT 109.130 74.480 109.270 79.860 ;
        RECT 108.670 74.340 109.270 74.480 ;
        RECT 108.670 72.630 108.810 74.340 ;
        RECT 111.890 72.630 112.030 79.860 ;
        RECT 115.110 72.630 115.250 79.860 ;
        RECT 118.330 72.630 118.470 81.560 ;
        RECT 123.390 81.540 123.530 83.600 ;
        RECT 124.770 83.580 124.910 89.720 ;
        RECT 127.070 89.360 127.210 89.720 ;
        RECT 126.090 89.040 126.350 89.360 ;
        RECT 127.010 89.040 127.270 89.360 ;
        RECT 126.150 85.620 126.290 89.040 ;
        RECT 127.530 88.760 127.670 89.720 ;
        RECT 127.070 88.620 127.670 88.760 ;
        RECT 126.550 88.020 126.810 88.340 ;
        RECT 126.090 85.300 126.350 85.620 ;
        RECT 126.610 84.260 126.750 88.020 ;
        RECT 127.070 85.620 127.210 88.620 ;
        RECT 127.470 88.020 127.730 88.340 ;
        RECT 127.530 87.320 127.670 88.020 ;
        RECT 127.470 87.000 127.730 87.320 ;
        RECT 127.010 85.300 127.270 85.620 ;
        RECT 126.550 83.940 126.810 84.260 ;
        RECT 124.710 83.260 124.970 83.580 ;
        RECT 123.330 81.220 123.590 81.540 ;
        RECT 127.070 80.860 127.210 85.300 ;
        RECT 127.530 84.260 127.670 87.000 ;
        RECT 127.470 83.940 127.730 84.260 ;
        RECT 127.990 80.860 128.130 91.760 ;
        RECT 128.390 91.080 128.650 91.400 ;
        RECT 128.450 89.360 128.590 91.080 ;
        RECT 128.390 89.040 128.650 89.360 ;
        RECT 128.450 85.870 128.590 89.040 ;
        RECT 128.910 86.980 129.050 96.100 ;
        RECT 129.370 94.800 129.510 96.180 ;
        RECT 129.310 94.480 129.570 94.800 ;
        RECT 130.290 94.120 130.430 96.180 ;
        RECT 130.230 93.800 130.490 94.120 ;
        RECT 130.750 91.740 130.890 97.540 ;
        RECT 131.210 94.800 131.350 100.010 ;
        RECT 132.070 98.900 132.330 99.220 ;
        RECT 131.610 97.880 131.870 98.200 ;
        RECT 131.670 96.840 131.810 97.880 ;
        RECT 132.130 96.840 132.270 98.900 ;
        RECT 131.610 96.520 131.870 96.840 ;
        RECT 132.070 96.520 132.330 96.840 ;
        RECT 131.150 94.480 131.410 94.800 ;
        RECT 131.150 93.800 131.410 94.120 ;
        RECT 131.210 91.740 131.350 93.800 ;
        RECT 132.590 91.740 132.730 110.380 ;
        RECT 133.050 103.640 133.190 116.860 ;
        RECT 133.510 106.360 133.650 129.840 ;
        RECT 133.970 118.600 134.110 130.180 ;
        RECT 134.430 130.160 134.570 138.340 ;
        RECT 138.050 138.000 138.310 138.320 ;
        RECT 137.130 132.560 137.390 132.880 ;
        RECT 137.190 130.840 137.330 132.560 ;
        RECT 137.590 131.540 137.850 131.860 ;
        RECT 137.650 130.840 137.790 131.540 ;
        RECT 135.750 130.520 136.010 130.840 ;
        RECT 137.130 130.520 137.390 130.840 ;
        RECT 137.590 130.520 137.850 130.840 ;
        RECT 134.370 129.840 134.630 130.160 ;
        RECT 135.290 129.500 135.550 129.820 ;
        RECT 135.810 129.730 135.950 130.520 ;
        RECT 138.110 130.355 138.250 138.000 ;
        RECT 139.030 137.155 139.170 138.680 ;
        RECT 140.410 138.660 140.550 139.700 ;
        RECT 140.870 139.000 141.010 140.185 ;
        RECT 140.810 138.680 141.070 139.000 ;
        RECT 140.350 138.340 140.610 138.660 ;
        RECT 138.960 136.785 139.240 137.155 ;
        RECT 139.890 134.260 140.150 134.580 ;
        RECT 139.950 132.880 140.090 134.260 ;
        RECT 139.890 132.560 140.150 132.880 ;
        RECT 138.970 131.540 139.230 131.860 ;
        RECT 138.040 129.985 138.320 130.355 ;
        RECT 136.210 129.730 136.470 129.820 ;
        RECT 135.810 129.590 136.470 129.730 ;
        RECT 134.830 127.460 135.090 127.780 ;
        RECT 134.890 124.040 135.030 127.460 ;
        RECT 134.830 123.720 135.090 124.040 ;
        RECT 135.350 122.680 135.490 129.500 ;
        RECT 135.290 122.360 135.550 122.680 ;
        RECT 135.810 119.280 135.950 129.590 ;
        RECT 136.210 129.500 136.470 129.590 ;
        RECT 139.030 129.480 139.170 131.540 ;
        RECT 140.410 129.820 140.550 138.340 ;
        RECT 140.800 133.385 141.080 133.755 ;
        RECT 140.810 133.240 141.070 133.385 ;
        RECT 140.800 129.985 141.080 130.355 ;
        RECT 140.350 129.500 140.610 129.820 ;
        RECT 138.970 129.160 139.230 129.480 ;
        RECT 139.890 128.820 140.150 129.140 ;
        RECT 139.950 127.440 140.090 128.820 ;
        RECT 140.870 128.120 141.010 129.985 ;
        RECT 140.810 127.800 141.070 128.120 ;
        RECT 139.890 127.120 140.150 127.440 ;
        RECT 139.890 126.440 140.150 126.760 ;
        RECT 140.800 126.585 141.080 126.955 ;
        RECT 138.510 126.100 138.770 126.420 ;
        RECT 138.570 124.380 138.710 126.100 ;
        RECT 138.510 124.060 138.770 124.380 ;
        RECT 136.210 123.720 136.470 124.040 ;
        RECT 136.270 120.980 136.410 123.720 ;
        RECT 136.210 120.660 136.470 120.980 ;
        RECT 135.750 118.960 136.010 119.280 ;
        RECT 136.270 118.940 136.410 120.660 ;
        RECT 139.950 118.940 140.090 126.440 ;
        RECT 140.870 125.400 141.010 126.585 ;
        RECT 140.810 125.080 141.070 125.400 ;
        RECT 140.800 123.185 141.080 123.555 ;
        RECT 140.870 122.680 141.010 123.185 ;
        RECT 140.810 122.360 141.070 122.680 ;
        RECT 140.800 119.785 141.080 120.155 ;
        RECT 140.810 119.640 141.070 119.785 ;
        RECT 136.210 118.620 136.470 118.940 ;
        RECT 137.590 118.680 137.850 118.940 ;
        RECT 137.590 118.620 138.250 118.680 ;
        RECT 139.890 118.620 140.150 118.940 ;
        RECT 133.910 118.280 134.170 118.600 ;
        RECT 137.650 118.540 138.250 118.620 ;
        RECT 133.970 114.180 134.110 118.280 ;
        RECT 138.110 115.540 138.250 118.540 ;
        RECT 138.970 117.940 139.230 118.260 ;
        RECT 139.030 116.755 139.170 117.940 ;
        RECT 138.960 116.385 139.240 116.755 ;
        RECT 138.050 115.220 138.310 115.540 ;
        RECT 133.910 113.860 134.170 114.180 ;
        RECT 138.110 113.840 138.250 115.220 ;
        RECT 138.050 113.520 138.310 113.840 ;
        RECT 137.130 112.840 137.390 113.160 ;
        RECT 134.370 112.500 134.630 112.820 ;
        RECT 134.430 108.060 134.570 112.500 ;
        RECT 136.210 110.120 136.470 110.440 ;
        RECT 134.370 107.740 134.630 108.060 ;
        RECT 133.450 106.040 133.710 106.360 ;
        RECT 135.290 105.360 135.550 105.680 ;
        RECT 132.990 103.320 133.250 103.640 ;
        RECT 134.830 103.320 135.090 103.640 ;
        RECT 134.890 102.620 135.030 103.320 ;
        RECT 135.350 103.300 135.490 105.360 ;
        RECT 135.290 102.980 135.550 103.300 ;
        RECT 135.350 102.620 135.490 102.980 ;
        RECT 134.830 102.300 135.090 102.620 ;
        RECT 135.290 102.300 135.550 102.620 ;
        RECT 133.910 101.620 134.170 101.940 ;
        RECT 133.970 100.920 134.110 101.620 ;
        RECT 133.910 100.600 134.170 100.920 ;
        RECT 134.890 100.150 135.030 102.300 ;
        RECT 135.750 101.960 136.010 102.280 ;
        RECT 135.290 100.150 135.550 100.240 ;
        RECT 134.890 100.010 135.550 100.150 ;
        RECT 134.890 97.180 135.030 100.010 ;
        RECT 135.290 99.920 135.550 100.010 ;
        RECT 135.810 99.900 135.950 101.960 ;
        RECT 135.750 99.580 136.010 99.900 ;
        RECT 135.810 98.395 135.950 99.580 ;
        RECT 135.740 98.025 136.020 98.395 ;
        RECT 134.830 96.860 135.090 97.180 ;
        RECT 135.810 96.840 135.950 98.025 ;
        RECT 136.270 97.180 136.410 110.120 ;
        RECT 137.190 106.360 137.330 112.840 ;
        RECT 137.130 106.040 137.390 106.360 ;
        RECT 136.670 102.300 136.930 102.620 ;
        RECT 136.730 99.560 136.870 102.300 ;
        RECT 136.670 99.240 136.930 99.560 ;
        RECT 137.590 98.900 137.850 99.220 ;
        RECT 137.650 97.715 137.790 98.900 ;
        RECT 137.580 97.345 137.860 97.715 ;
        RECT 136.210 96.860 136.470 97.180 ;
        RECT 135.750 96.520 136.010 96.840 ;
        RECT 130.690 91.420 130.950 91.740 ;
        RECT 131.150 91.420 131.410 91.740 ;
        RECT 132.530 91.420 132.790 91.740 ;
        RECT 136.210 91.080 136.470 91.400 ;
        RECT 135.750 90.970 136.010 91.060 ;
        RECT 135.350 90.830 136.010 90.970 ;
        RECT 129.770 89.380 130.030 89.700 ;
        RECT 129.300 88.505 129.580 88.875 ;
        RECT 128.850 86.660 129.110 86.980 ;
        RECT 129.370 86.640 129.510 88.505 ;
        RECT 129.830 87.320 129.970 89.380 ;
        RECT 129.770 87.000 130.030 87.320 ;
        RECT 129.310 86.320 129.570 86.640 ;
        RECT 131.140 86.465 131.420 86.835 ;
        RECT 131.210 85.960 131.350 86.465 ;
        RECT 135.350 86.300 135.490 90.830 ;
        RECT 135.750 90.740 136.010 90.830 ;
        RECT 136.270 89.360 136.410 91.080 ;
        RECT 135.750 89.040 136.010 89.360 ;
        RECT 136.210 89.040 136.470 89.360 ;
        RECT 135.810 87.320 135.950 89.040 ;
        RECT 135.750 87.000 136.010 87.320 ;
        RECT 132.530 85.980 132.790 86.300 ;
        RECT 134.370 85.980 134.630 86.300 ;
        RECT 135.290 85.980 135.550 86.300 ;
        RECT 129.310 85.870 129.570 85.960 ;
        RECT 128.450 85.730 129.570 85.870 ;
        RECT 128.450 84.600 128.590 85.730 ;
        RECT 129.310 85.640 129.570 85.730 ;
        RECT 131.150 85.640 131.410 85.960 ;
        RECT 131.210 84.600 131.350 85.640 ;
        RECT 128.390 84.280 128.650 84.600 ;
        RECT 131.150 84.280 131.410 84.600 ;
        RECT 131.210 80.860 131.350 84.280 ;
        RECT 132.590 84.260 132.730 85.980 ;
        RECT 134.430 84.600 134.570 85.980 ;
        RECT 134.370 84.280 134.630 84.600 ;
        RECT 132.530 83.940 132.790 84.260 ;
        RECT 138.110 83.920 138.250 113.520 ;
        RECT 139.890 113.180 140.150 113.500 ;
        RECT 138.510 112.840 138.770 113.160 ;
        RECT 138.570 111.120 138.710 112.840 ;
        RECT 139.950 111.120 140.090 113.180 ;
        RECT 140.800 112.985 141.080 113.355 ;
        RECT 140.870 112.820 141.010 112.985 ;
        RECT 140.810 112.500 141.070 112.820 ;
        RECT 138.510 110.800 138.770 111.120 ;
        RECT 139.890 110.800 140.150 111.120 ;
        RECT 142.640 109.585 142.920 109.955 ;
        RECT 140.350 107.060 140.610 107.380 ;
        RECT 139.890 106.040 140.150 106.360 ;
        RECT 138.960 102.785 139.240 103.155 ;
        RECT 139.030 101.940 139.170 102.785 ;
        RECT 139.950 102.620 140.090 106.040 ;
        RECT 140.410 105.680 140.550 107.060 ;
        RECT 140.800 106.185 141.080 106.555 ;
        RECT 142.710 106.360 142.850 109.585 ;
        RECT 140.350 105.360 140.610 105.680 ;
        RECT 139.890 102.300 140.150 102.620 ;
        RECT 138.970 101.620 139.230 101.940 ;
        RECT 139.950 100.580 140.090 102.300 ;
        RECT 140.870 101.940 141.010 106.185 ;
        RECT 142.650 106.040 142.910 106.360 ;
        RECT 140.810 101.620 141.070 101.940 ;
        RECT 139.890 100.260 140.150 100.580 ;
        RECT 138.510 99.240 138.770 99.560 ;
        RECT 140.800 99.385 141.080 99.755 ;
        RECT 138.570 98.200 138.710 99.240 ;
        RECT 139.890 98.900 140.150 99.220 ;
        RECT 138.510 97.880 138.770 98.200 ;
        RECT 138.570 95.480 138.710 97.880 ;
        RECT 139.950 97.180 140.090 98.900 ;
        RECT 140.870 98.200 141.010 99.385 ;
        RECT 140.810 97.880 141.070 98.200 ;
        RECT 139.890 96.860 140.150 97.180 ;
        RECT 139.430 96.520 139.690 96.840 ;
        RECT 138.510 95.160 138.770 95.480 ;
        RECT 139.490 92.760 139.630 96.520 ;
        RECT 140.800 95.985 141.080 96.355 ;
        RECT 140.870 95.480 141.010 95.985 ;
        RECT 140.810 95.160 141.070 95.480 ;
        RECT 139.430 92.440 139.690 92.760 ;
        RECT 140.800 92.585 141.080 92.955 ;
        RECT 138.960 89.185 139.240 89.555 ;
        RECT 139.490 89.360 139.630 92.440 ;
        RECT 139.030 88.680 139.170 89.185 ;
        RECT 139.430 89.040 139.690 89.360 ;
        RECT 140.870 88.680 141.010 92.585 ;
        RECT 138.970 88.360 139.230 88.680 ;
        RECT 140.810 88.360 141.070 88.680 ;
        RECT 140.800 85.785 141.080 86.155 ;
        RECT 140.870 85.620 141.010 85.785 ;
        RECT 140.810 85.300 141.070 85.620 ;
        RECT 136.210 83.600 136.470 83.920 ;
        RECT 138.050 83.600 138.310 83.920 ;
        RECT 136.270 80.860 136.410 83.600 ;
        RECT 140.810 82.755 141.070 82.900 ;
        RECT 140.800 82.385 141.080 82.755 ;
        RECT 121.490 80.540 121.750 80.860 ;
        RECT 127.010 80.540 127.270 80.860 ;
        RECT 127.930 80.540 128.190 80.860 ;
        RECT 131.150 80.540 131.410 80.860 ;
        RECT 136.210 80.540 136.470 80.860 ;
        RECT 121.550 72.630 121.690 80.540 ;
        RECT 124.710 79.860 124.970 80.180 ;
        RECT 127.930 79.860 128.190 80.180 ;
        RECT 131.150 79.860 131.410 80.180 ;
        RECT 134.370 79.860 134.630 80.180 ;
        RECT 124.770 72.630 124.910 79.860 ;
        RECT 127.990 72.630 128.130 79.860 ;
        RECT 131.210 72.630 131.350 79.860 ;
        RECT 134.430 72.630 134.570 79.860 ;
        RECT 63.520 68.630 63.800 72.630 ;
        RECT 69.960 68.630 70.240 72.630 ;
        RECT 73.180 68.630 73.460 72.630 ;
        RECT 76.400 68.630 76.680 72.630 ;
        RECT 79.620 68.630 79.900 72.630 ;
        RECT 82.840 68.630 83.120 72.630 ;
        RECT 86.060 68.630 86.340 72.630 ;
        RECT 89.280 68.630 89.560 72.630 ;
        RECT 92.500 68.630 92.780 72.630 ;
        RECT 95.720 68.630 96.000 72.630 ;
        RECT 98.940 68.630 99.220 72.630 ;
        RECT 102.160 68.630 102.440 72.630 ;
        RECT 105.380 68.630 105.660 72.630 ;
        RECT 108.600 68.630 108.880 72.630 ;
        RECT 111.820 68.630 112.100 72.630 ;
        RECT 115.040 68.630 115.320 72.630 ;
        RECT 118.260 68.630 118.540 72.630 ;
        RECT 121.480 68.630 121.760 72.630 ;
        RECT 124.700 68.630 124.980 72.630 ;
        RECT 127.920 68.630 128.200 72.630 ;
        RECT 131.140 68.630 131.420 72.630 ;
        RECT 134.360 68.630 134.640 72.630 ;
        RECT 26.640 56.255 26.920 60.255 ;
        RECT 29.860 56.255 30.140 60.255 ;
        RECT 33.080 56.255 33.360 60.255 ;
        RECT 36.300 56.255 36.580 60.255 ;
        RECT 39.520 56.255 39.800 60.255 ;
        RECT 26.710 48.380 26.850 56.255 ;
        RECT 29.930 49.820 30.070 56.255 ;
        RECT 29.930 49.680 30.990 49.820 ;
        RECT 28.300 48.545 29.840 48.915 ;
        RECT 26.650 48.060 26.910 48.380 ;
        RECT 18.370 47.040 18.630 47.360 ;
        RECT 22.970 47.040 23.230 47.360 ;
        RECT 23.430 47.040 23.690 47.360 ;
        RECT 18.430 45.660 18.570 47.040 ;
        RECT 23.030 45.660 23.170 47.040 ;
        RECT 18.370 45.340 18.630 45.660 ;
        RECT 22.970 45.340 23.230 45.660 ;
        RECT 23.490 45.175 23.630 47.040 ;
        RECT 25.270 46.360 25.530 46.680 ;
        RECT 30.330 46.360 30.590 46.680 ;
        RECT 25.330 45.320 25.470 46.360 ;
        RECT 23.420 44.805 23.700 45.175 ;
        RECT 25.270 45.000 25.530 45.320 ;
        RECT 26.190 44.660 26.450 44.980 ;
        RECT 27.560 44.805 27.840 45.175 ;
        RECT 23.890 43.640 24.150 43.960 ;
        RECT 23.950 41.920 24.090 43.640 ;
        RECT 24.800 43.445 25.080 43.815 ;
        RECT 23.890 41.600 24.150 41.920 ;
        RECT 16.070 41.260 16.330 41.580 ;
        RECT 13.760 40.045 14.040 40.415 ;
        RECT 16.130 40.220 16.270 41.260 ;
        RECT 21.130 40.920 21.390 41.240 ;
        RECT 21.590 40.920 21.850 41.240 ;
        RECT 13.770 39.900 14.030 40.045 ;
        RECT 16.070 39.900 16.330 40.220 ;
        RECT 21.190 39.540 21.330 40.920 ;
        RECT 21.650 40.220 21.790 40.920 ;
        RECT 23.950 40.220 24.090 41.600 ;
        RECT 21.590 39.900 21.850 40.220 ;
        RECT 23.890 39.900 24.150 40.220 ;
        RECT 21.130 39.220 21.390 39.540 ;
        RECT 19.750 38.880 20.010 39.200 ;
        RECT 16.530 38.540 16.790 38.860 ;
        RECT 16.590 36.820 16.730 38.540 ;
        RECT 16.530 36.500 16.790 36.820 ;
        RECT 19.810 36.140 19.950 38.880 ;
        RECT 23.950 36.480 24.090 39.900 ;
        RECT 21.130 36.160 21.390 36.480 ;
        RECT 23.890 36.160 24.150 36.480 ;
        RECT 19.750 35.820 20.010 36.140 ;
        RECT 14.230 35.480 14.490 35.800 ;
        RECT 18.830 35.480 19.090 35.800 ;
        RECT 14.290 34.440 14.430 35.480 ;
        RECT 14.230 34.120 14.490 34.440 ;
        RECT 13.760 33.245 14.040 33.615 ;
        RECT 13.830 29.340 13.970 33.245 ;
        RECT 14.230 32.760 14.490 33.080 ;
        RECT 14.290 31.380 14.430 32.760 ;
        RECT 18.890 32.060 19.030 35.480 ;
        RECT 18.830 31.740 19.090 32.060 ;
        RECT 14.230 31.060 14.490 31.380 ;
        RECT 13.770 29.020 14.030 29.340 ;
        RECT 14.290 28.660 14.430 31.060 ;
        RECT 19.290 30.040 19.550 30.360 ;
        RECT 19.350 29.340 19.490 30.040 ;
        RECT 19.290 29.020 19.550 29.340 ;
        RECT 14.230 28.340 14.490 28.660 ;
        RECT 19.810 28.320 19.950 35.820 ;
        RECT 21.190 34.100 21.330 36.160 ;
        RECT 24.870 34.440 25.010 43.445 ;
        RECT 26.250 42.940 26.390 44.660 ;
        RECT 26.190 42.620 26.450 42.940 ;
        RECT 26.190 39.900 26.450 40.220 ;
        RECT 27.110 39.900 27.370 40.220 ;
        RECT 26.250 36.820 26.390 39.900 ;
        RECT 27.170 37.500 27.310 39.900 ;
        RECT 27.110 37.180 27.370 37.500 ;
        RECT 26.190 36.500 26.450 36.820 ;
        RECT 24.810 34.120 25.070 34.440 ;
        RECT 21.130 33.780 21.390 34.100 ;
        RECT 27.170 32.060 27.310 37.180 ;
        RECT 27.630 32.060 27.770 44.805 ;
        RECT 28.300 43.105 29.840 43.475 ;
        RECT 30.390 41.920 30.530 46.360 ;
        RECT 30.850 44.300 30.990 49.680 ;
        RECT 33.150 48.380 33.290 56.255 ;
        RECT 33.090 48.060 33.350 48.380 ;
        RECT 31.250 47.720 31.510 48.040 ;
        RECT 30.790 43.980 31.050 44.300 ;
        RECT 31.310 42.940 31.450 47.720 ;
        RECT 36.370 47.360 36.510 56.255 ;
        RECT 39.590 48.380 39.730 56.255 ;
        RECT 46.880 53.645 47.160 54.015 ;
        RECT 44.120 50.245 44.400 50.615 ;
        RECT 39.530 48.060 39.790 48.380 ;
        RECT 38.150 47.720 38.410 48.040 ;
        RECT 33.550 47.040 33.810 47.360 ;
        RECT 36.310 47.040 36.570 47.360 ;
        RECT 31.600 45.825 33.140 46.195 ;
        RECT 33.610 45.660 33.750 47.040 ;
        RECT 34.010 46.360 34.270 46.680 ;
        RECT 33.550 45.340 33.810 45.660 ;
        RECT 34.070 45.320 34.210 46.360 ;
        RECT 34.010 45.000 34.270 45.320 ;
        RECT 38.210 44.980 38.350 47.720 ;
        RECT 44.190 47.360 44.330 50.245 ;
        RECT 46.950 47.360 47.090 53.645 ;
        RECT 41.370 47.040 41.630 47.360 ;
        RECT 44.130 47.040 44.390 47.360 ;
        RECT 45.510 47.215 45.770 47.360 ;
        RECT 39.990 46.360 40.250 46.680 ;
        RECT 34.930 44.660 35.190 44.980 ;
        RECT 36.310 44.660 36.570 44.980 ;
        RECT 38.150 44.660 38.410 44.980 ;
        RECT 31.710 44.320 31.970 44.640 ;
        RECT 31.250 42.620 31.510 42.940 ;
        RECT 31.770 41.920 31.910 44.320 ;
        RECT 34.470 43.640 34.730 43.960 ;
        RECT 34.530 42.260 34.670 43.640 ;
        RECT 34.470 41.940 34.730 42.260 ;
        RECT 34.990 41.920 35.130 44.660 ;
        RECT 35.850 44.320 36.110 44.640 ;
        RECT 30.330 41.600 30.590 41.920 ;
        RECT 30.790 41.600 31.050 41.920 ;
        RECT 31.710 41.600 31.970 41.920 ;
        RECT 33.550 41.600 33.810 41.920 ;
        RECT 34.010 41.600 34.270 41.920 ;
        RECT 34.930 41.600 35.190 41.920 ;
        RECT 30.330 40.920 30.590 41.240 ;
        RECT 28.300 37.665 29.840 38.035 ;
        RECT 28.300 32.225 29.840 32.595 ;
        RECT 27.110 31.740 27.370 32.060 ;
        RECT 27.570 31.740 27.830 32.060 ;
        RECT 22.050 30.720 22.310 31.040 ;
        RECT 19.290 28.000 19.550 28.320 ;
        RECT 19.750 28.000 20.010 28.320 ;
        RECT 14.230 27.660 14.490 27.980 ;
        RECT 13.760 26.445 14.040 26.815 ;
        RECT 13.830 22.540 13.970 26.445 ;
        RECT 14.290 25.940 14.430 27.660 ;
        RECT 16.530 27.320 16.790 27.640 ;
        RECT 14.230 25.620 14.490 25.940 ;
        RECT 16.590 25.260 16.730 27.320 ;
        RECT 16.530 24.940 16.790 25.260 ;
        RECT 14.230 22.560 14.490 22.880 ;
        RECT 13.770 22.220 14.030 22.540 ;
        RECT 14.290 21.180 14.430 22.560 ;
        RECT 19.350 22.540 19.490 28.000 ;
        RECT 22.110 26.620 22.250 30.720 ;
        RECT 27.170 29.000 27.310 31.740 ;
        RECT 30.390 31.040 30.530 40.920 ;
        RECT 30.850 40.220 30.990 41.600 ;
        RECT 31.600 40.385 33.140 40.755 ;
        RECT 30.790 39.900 31.050 40.220 ;
        RECT 30.790 39.220 31.050 39.540 ;
        RECT 30.850 33.080 30.990 39.220 ;
        RECT 31.250 38.200 31.510 38.520 ;
        RECT 31.310 34.180 31.450 38.200 ;
        RECT 33.610 37.500 33.750 41.600 ;
        RECT 33.550 37.180 33.810 37.500 ;
        RECT 34.070 36.900 34.210 41.600 ;
        RECT 35.910 39.880 36.050 44.320 ;
        RECT 36.370 42.940 36.510 44.660 ;
        RECT 37.230 43.640 37.490 43.960 ;
        RECT 36.310 42.620 36.570 42.940 ;
        RECT 36.370 42.340 36.510 42.620 ;
        RECT 36.370 42.200 36.970 42.340 ;
        RECT 36.310 41.260 36.570 41.580 ;
        RECT 35.850 39.560 36.110 39.880 ;
        RECT 34.470 38.880 34.730 39.200 ;
        RECT 33.610 36.760 34.210 36.900 ;
        RECT 33.610 35.800 33.750 36.760 ;
        RECT 34.530 36.480 34.670 38.880 ;
        RECT 34.930 36.840 35.190 37.160 ;
        RECT 34.470 36.160 34.730 36.480 ;
        RECT 34.010 35.820 34.270 36.140 ;
        RECT 33.550 35.480 33.810 35.800 ;
        RECT 31.600 34.945 33.140 35.315 ;
        RECT 31.310 34.040 31.910 34.180 ;
        RECT 31.250 33.440 31.510 33.760 ;
        RECT 30.790 32.760 31.050 33.080 ;
        RECT 27.570 30.720 27.830 31.040 ;
        RECT 30.330 30.720 30.590 31.040 ;
        RECT 27.630 29.340 27.770 30.720 ;
        RECT 27.570 29.020 27.830 29.340 ;
        RECT 25.730 28.680 25.990 29.000 ;
        RECT 27.110 28.680 27.370 29.000 ;
        RECT 22.050 26.300 22.310 26.620 ;
        RECT 21.130 25.280 21.390 25.600 ;
        RECT 19.290 22.220 19.550 22.540 ;
        RECT 18.830 21.880 19.090 22.200 ;
        RECT 14.230 20.860 14.490 21.180 ;
        RECT 14.290 17.780 14.430 20.860 ;
        RECT 16.990 19.500 17.250 19.820 ;
        RECT 17.050 18.460 17.190 19.500 ;
        RECT 18.890 18.460 19.030 21.880 ;
        RECT 19.350 18.460 19.490 22.220 ;
        RECT 21.190 20.500 21.330 25.280 ;
        RECT 22.110 23.220 22.250 26.300 ;
        RECT 22.050 22.900 22.310 23.220 ;
        RECT 25.790 22.880 25.930 28.680 ;
        RECT 27.110 27.660 27.370 27.980 ;
        RECT 27.170 25.260 27.310 27.660 ;
        RECT 28.300 26.785 29.840 27.155 ;
        RECT 27.110 24.940 27.370 25.260 ;
        RECT 21.590 22.560 21.850 22.880 ;
        RECT 25.730 22.560 25.990 22.880 ;
        RECT 21.130 20.180 21.390 20.500 ;
        RECT 21.650 18.460 21.790 22.560 ;
        RECT 16.990 18.140 17.250 18.460 ;
        RECT 18.830 18.140 19.090 18.460 ;
        RECT 19.290 18.140 19.550 18.460 ;
        RECT 21.590 18.140 21.850 18.460 ;
        RECT 23.890 18.140 24.150 18.460 ;
        RECT 14.230 17.460 14.490 17.780 ;
        RECT 11.460 16.925 11.740 17.295 ;
        RECT 11.470 16.780 11.730 16.925 ;
        RECT 23.950 14.720 24.090 18.140 ;
        RECT 25.790 17.440 25.930 22.560 ;
        RECT 30.330 21.880 30.590 22.200 ;
        RECT 28.300 21.345 29.840 21.715 ;
        RECT 30.390 18.460 30.530 21.880 ;
        RECT 30.850 20.160 30.990 32.760 ;
        RECT 31.310 31.040 31.450 33.440 ;
        RECT 31.770 31.720 31.910 34.040 ;
        RECT 31.710 31.400 31.970 31.720 ;
        RECT 31.250 30.720 31.510 31.040 ;
        RECT 31.600 29.505 33.140 29.875 ;
        RECT 33.610 28.320 33.750 35.480 ;
        RECT 34.070 34.780 34.210 35.820 ;
        RECT 34.010 34.460 34.270 34.780 ;
        RECT 34.990 31.380 35.130 36.840 ;
        RECT 35.390 35.820 35.650 36.140 ;
        RECT 34.930 31.060 35.190 31.380 ;
        RECT 34.470 29.250 34.730 29.340 ;
        RECT 34.990 29.250 35.130 31.060 ;
        RECT 34.470 29.110 35.130 29.250 ;
        RECT 34.470 29.020 34.730 29.110 ;
        RECT 33.550 28.000 33.810 28.320 ;
        RECT 34.010 28.000 34.270 28.320 ;
        RECT 34.070 24.920 34.210 28.000 ;
        RECT 34.990 26.020 35.130 29.110 ;
        RECT 35.450 26.280 35.590 35.820 ;
        RECT 35.910 33.080 36.050 39.560 ;
        RECT 36.370 38.860 36.510 41.260 ;
        RECT 36.310 38.540 36.570 38.860 ;
        RECT 36.370 34.780 36.510 38.540 ;
        RECT 36.310 34.460 36.570 34.780 ;
        RECT 35.850 32.760 36.110 33.080 ;
        RECT 35.910 31.720 36.050 32.760 ;
        RECT 35.850 31.400 36.110 31.720 ;
        RECT 35.850 27.660 36.110 27.980 ;
        RECT 34.530 25.940 35.130 26.020 ;
        RECT 35.390 25.960 35.650 26.280 ;
        RECT 34.470 25.880 35.130 25.940 ;
        RECT 34.470 25.620 34.730 25.880 ;
        RECT 31.250 24.600 31.510 24.920 ;
        RECT 34.010 24.600 34.270 24.920 ;
        RECT 31.310 23.220 31.450 24.600 ;
        RECT 31.600 24.065 33.140 24.435 ;
        RECT 31.250 22.900 31.510 23.220 ;
        RECT 31.310 21.180 31.450 22.900 ;
        RECT 31.250 20.860 31.510 21.180 ;
        RECT 30.790 19.840 31.050 20.160 ;
        RECT 30.330 18.140 30.590 18.460 ;
        RECT 31.310 18.120 31.450 20.860 ;
        RECT 31.600 18.625 33.140 18.995 ;
        RECT 31.250 17.860 31.510 18.120 ;
        RECT 30.390 17.800 31.510 17.860 ;
        RECT 30.390 17.720 31.450 17.800 ;
        RECT 25.730 17.120 25.990 17.440 ;
        RECT 28.300 15.905 29.840 16.275 ;
        RECT 23.890 14.400 24.150 14.720 ;
        RECT 28.950 14.630 29.210 14.720 ;
        RECT 30.390 14.630 30.530 17.720 ;
        RECT 31.250 16.440 31.510 16.760 ;
        RECT 28.950 14.490 30.530 14.630 ;
        RECT 28.950 14.400 29.210 14.490 ;
        RECT 31.310 14.380 31.450 16.440 ;
        RECT 34.070 15.740 34.210 24.600 ;
        RECT 35.910 23.560 36.050 27.660 ;
        RECT 36.830 26.620 36.970 42.200 ;
        RECT 37.290 41.920 37.430 43.640 ;
        RECT 37.230 41.600 37.490 41.920 ;
        RECT 40.050 39.540 40.190 46.360 ;
        RECT 40.900 44.890 41.180 45.175 ;
        RECT 40.510 44.805 41.180 44.890 ;
        RECT 40.510 44.750 41.170 44.805 ;
        RECT 40.510 39.880 40.650 44.750 ;
        RECT 40.910 44.660 41.170 44.750 ;
        RECT 41.430 44.300 41.570 47.040 ;
        RECT 45.500 46.845 45.780 47.215 ;
        RECT 46.890 47.040 47.150 47.360 ;
        RECT 43.670 46.360 43.930 46.680 ;
        RECT 46.430 46.360 46.690 46.680 ;
        RECT 41.370 43.980 41.630 44.300 ;
        RECT 41.430 42.940 41.570 43.980 ;
        RECT 43.210 43.640 43.470 43.960 ;
        RECT 41.370 42.620 41.630 42.940 ;
        RECT 43.270 41.920 43.410 43.640 ;
        RECT 43.210 41.600 43.470 41.920 ;
        RECT 43.730 40.220 43.870 46.360 ;
        RECT 44.130 44.660 44.390 44.980 ;
        RECT 44.190 42.940 44.330 44.660 ;
        RECT 44.590 43.980 44.850 44.300 ;
        RECT 44.130 42.620 44.390 42.940 ;
        RECT 44.650 42.340 44.790 43.980 ;
        RECT 44.190 42.200 44.790 42.340 ;
        RECT 43.670 39.900 43.930 40.220 ;
        RECT 40.450 39.560 40.710 39.880 ;
        RECT 40.910 39.560 41.170 39.880 ;
        RECT 39.990 39.220 40.250 39.540 ;
        RECT 38.150 38.200 38.410 38.520 ;
        RECT 38.210 32.060 38.350 38.200 ;
        RECT 39.070 35.480 39.330 35.800 ;
        RECT 39.130 34.100 39.270 35.480 ;
        RECT 40.050 34.100 40.190 39.220 ;
        RECT 40.970 38.860 41.110 39.560 ;
        RECT 43.730 39.540 43.870 39.900 ;
        RECT 43.670 39.220 43.930 39.540 ;
        RECT 40.910 38.540 41.170 38.860 ;
        RECT 40.970 36.480 41.110 38.540 ;
        RECT 41.830 36.840 42.090 37.160 ;
        RECT 40.910 36.160 41.170 36.480 ;
        RECT 39.070 33.780 39.330 34.100 ;
        RECT 39.990 33.780 40.250 34.100 ;
        RECT 38.150 31.740 38.410 32.060 ;
        RECT 37.690 30.040 37.950 30.360 ;
        RECT 36.770 26.300 37.030 26.620 ;
        RECT 35.850 23.240 36.110 23.560 ;
        RECT 35.910 18.460 36.050 23.240 ;
        RECT 36.830 23.220 36.970 26.300 ;
        RECT 36.770 22.900 37.030 23.220 ;
        RECT 35.850 18.140 36.110 18.460 ;
        RECT 36.830 17.440 36.970 22.900 ;
        RECT 37.750 22.880 37.890 30.040 ;
        RECT 38.210 28.660 38.350 31.740 ;
        RECT 41.890 31.460 42.030 36.840 ;
        RECT 42.750 36.500 43.010 36.820 ;
        RECT 42.290 32.760 42.550 33.080 ;
        RECT 40.970 31.320 42.030 31.460 ;
        RECT 40.970 31.040 41.110 31.320 ;
        RECT 40.910 30.720 41.170 31.040 ;
        RECT 41.830 30.720 42.090 31.040 ;
        RECT 40.450 30.040 40.710 30.360 ;
        RECT 41.890 30.215 42.030 30.720 ;
        RECT 42.350 30.700 42.490 32.760 ;
        RECT 42.290 30.380 42.550 30.700 ;
        RECT 40.510 28.660 40.650 30.040 ;
        RECT 41.820 29.845 42.100 30.215 ;
        RECT 42.350 29.000 42.490 30.380 ;
        RECT 42.290 28.680 42.550 29.000 ;
        RECT 38.150 28.340 38.410 28.660 ;
        RECT 40.450 28.340 40.710 28.660 ;
        RECT 39.520 26.445 39.800 26.815 ;
        RECT 37.690 22.560 37.950 22.880 ;
        RECT 37.750 22.200 37.890 22.560 ;
        RECT 37.690 21.880 37.950 22.200 ;
        RECT 39.590 20.160 39.730 26.445 ;
        RECT 42.350 25.940 42.490 28.680 ;
        RECT 42.810 26.620 42.950 36.500 ;
        RECT 43.730 36.480 43.870 39.220 ;
        RECT 44.190 36.480 44.330 42.200 ;
        RECT 44.590 41.600 44.850 41.920 ;
        RECT 44.650 37.015 44.790 41.600 ;
        RECT 45.510 40.920 45.770 41.240 ;
        RECT 45.970 40.920 46.230 41.240 ;
        RECT 45.050 39.220 45.310 39.540 ;
        RECT 45.110 37.500 45.250 39.220 ;
        RECT 45.050 37.180 45.310 37.500 ;
        RECT 44.580 36.645 44.860 37.015 ;
        RECT 45.570 36.900 45.710 40.920 ;
        RECT 46.030 40.220 46.170 40.920 ;
        RECT 45.970 39.900 46.230 40.220 ;
        RECT 46.490 39.540 46.630 46.360 ;
        RECT 46.890 44.660 47.150 44.980 ;
        RECT 46.950 43.815 47.090 44.660 ;
        RECT 46.880 43.445 47.160 43.815 ;
        RECT 46.890 41.600 47.150 41.920 ;
        RECT 46.950 40.415 47.090 41.600 ;
        RECT 46.880 40.045 47.160 40.415 ;
        RECT 46.430 39.220 46.690 39.540 ;
        RECT 46.490 37.160 46.630 39.220 ;
        RECT 45.570 36.760 46.170 36.900 ;
        RECT 46.430 36.840 46.690 37.160 ;
        RECT 46.030 36.480 46.170 36.760 ;
        RECT 43.670 36.160 43.930 36.480 ;
        RECT 44.130 36.160 44.390 36.480 ;
        RECT 45.510 36.160 45.770 36.480 ;
        RECT 45.970 36.160 46.230 36.480 ;
        RECT 44.190 31.720 44.330 36.160 ;
        RECT 44.590 33.780 44.850 34.100 ;
        RECT 44.130 31.400 44.390 31.720 ;
        RECT 44.650 31.040 44.790 33.780 ;
        RECT 45.570 32.060 45.710 36.160 ;
        RECT 46.030 34.100 46.170 36.160 ;
        RECT 45.970 33.780 46.230 34.100 ;
        RECT 46.890 33.780 47.150 34.100 ;
        RECT 46.950 33.615 47.090 33.780 ;
        RECT 46.880 33.245 47.160 33.615 ;
        RECT 45.510 31.740 45.770 32.060 ;
        RECT 44.130 30.720 44.390 31.040 ;
        RECT 44.590 30.720 44.850 31.040 ;
        RECT 44.190 29.340 44.330 30.720 ;
        RECT 45.050 30.380 45.310 30.700 ;
        RECT 44.130 29.020 44.390 29.340 ;
        RECT 43.670 28.340 43.930 28.660 ;
        RECT 44.130 28.340 44.390 28.660 ;
        RECT 42.750 26.300 43.010 26.620 ;
        RECT 42.290 25.620 42.550 25.940 ;
        RECT 39.990 25.280 40.250 25.600 ;
        RECT 42.750 25.280 43.010 25.600 ;
        RECT 40.050 22.200 40.190 25.280 ;
        RECT 40.910 24.600 41.170 24.920 ;
        RECT 40.970 23.900 41.110 24.600 ;
        RECT 40.910 23.580 41.170 23.900 ;
        RECT 42.810 22.880 42.950 25.280 ;
        RECT 43.200 23.045 43.480 23.415 ;
        RECT 43.210 22.900 43.470 23.045 ;
        RECT 42.750 22.560 43.010 22.880 ;
        RECT 39.990 21.880 40.250 22.200 ;
        RECT 38.150 19.840 38.410 20.160 ;
        RECT 39.530 19.840 39.790 20.160 ;
        RECT 36.770 17.120 37.030 17.440 ;
        RECT 37.230 17.120 37.490 17.440 ;
        RECT 34.010 15.420 34.270 15.740 ;
        RECT 37.290 15.400 37.430 17.120 ;
        RECT 38.210 16.615 38.350 19.840 ;
        RECT 38.140 16.245 38.420 16.615 ;
        RECT 37.230 15.080 37.490 15.400 ;
        RECT 37.290 14.720 37.430 15.080 ;
        RECT 40.050 14.720 40.190 21.880 ;
        RECT 42.810 21.180 42.950 22.560 ;
        RECT 43.730 22.200 43.870 28.340 ;
        RECT 43.670 21.880 43.930 22.200 ;
        RECT 42.750 20.860 43.010 21.180 ;
        RECT 43.210 20.520 43.470 20.840 ;
        RECT 40.910 20.015 41.170 20.160 ;
        RECT 40.900 19.645 41.180 20.015 ;
        RECT 42.290 19.160 42.550 19.480 ;
        RECT 42.750 19.160 43.010 19.480 ;
        RECT 42.350 17.440 42.490 19.160 ;
        RECT 42.810 17.780 42.950 19.160 ;
        RECT 42.750 17.460 43.010 17.780 ;
        RECT 42.290 17.120 42.550 17.440 ;
        RECT 42.350 15.060 42.490 17.120 ;
        RECT 43.270 15.400 43.410 20.520 ;
        RECT 43.730 20.160 43.870 21.880 ;
        RECT 44.190 21.180 44.330 28.340 ;
        RECT 44.590 28.000 44.850 28.320 ;
        RECT 44.650 23.900 44.790 28.000 ;
        RECT 45.110 25.600 45.250 30.380 ;
        RECT 45.970 28.340 46.230 28.660 ;
        RECT 45.050 25.280 45.310 25.600 ;
        RECT 45.510 25.280 45.770 25.600 ;
        RECT 44.590 23.580 44.850 23.900 ;
        RECT 45.110 23.560 45.250 25.280 ;
        RECT 45.050 23.240 45.310 23.560 ;
        RECT 44.590 22.900 44.850 23.220 ;
        RECT 44.130 20.860 44.390 21.180 ;
        RECT 44.650 20.160 44.790 22.900 ;
        RECT 43.670 19.840 43.930 20.160 ;
        RECT 44.590 19.840 44.850 20.160 ;
        RECT 43.730 15.740 43.870 19.840 ;
        RECT 45.570 18.460 45.710 25.280 ;
        RECT 46.030 22.880 46.170 28.340 ;
        RECT 45.970 22.560 46.230 22.880 ;
        RECT 46.890 22.220 47.150 22.540 ;
        RECT 46.430 20.180 46.690 20.500 ;
        RECT 45.970 19.840 46.230 20.160 ;
        RECT 45.510 18.140 45.770 18.460 ;
        RECT 46.030 15.740 46.170 19.840 ;
        RECT 43.670 15.420 43.930 15.740 ;
        RECT 45.970 15.420 46.230 15.740 ;
        RECT 43.210 15.080 43.470 15.400 ;
        RECT 42.290 14.740 42.550 15.060 ;
        RECT 37.230 14.400 37.490 14.720 ;
        RECT 39.990 14.400 40.250 14.720 ;
        RECT 42.750 14.400 43.010 14.720 ;
        RECT 31.250 14.060 31.510 14.380 ;
        RECT 26.650 13.720 26.910 14.040 ;
        RECT 29.410 13.720 29.670 14.040 ;
        RECT 33.550 13.720 33.810 14.040 ;
        RECT 39.530 13.720 39.790 14.040 ;
        RECT 26.710 6.490 26.850 13.720 ;
        RECT 29.470 8.340 29.610 13.720 ;
        RECT 31.600 13.185 33.140 13.555 ;
        RECT 33.610 8.340 33.750 13.720 ;
        RECT 29.470 8.200 30.070 8.340 ;
        RECT 29.930 6.490 30.070 8.200 ;
        RECT 33.150 8.200 33.750 8.340 ;
        RECT 33.150 6.490 33.290 8.200 ;
        RECT 39.590 6.490 39.730 13.720 ;
        RECT 42.810 13.215 42.950 14.400 ;
        RECT 42.740 12.845 43.020 13.215 ;
        RECT 46.490 9.815 46.630 20.180 ;
        RECT 46.950 20.160 47.090 22.220 ;
        RECT 46.890 19.840 47.150 20.160 ;
        RECT 46.950 17.440 47.090 19.840 ;
        RECT 46.890 17.120 47.150 17.440 ;
        RECT 46.420 9.445 46.700 9.815 ;
        RECT 26.640 2.490 26.920 6.490 ;
        RECT 29.860 2.490 30.140 6.490 ;
        RECT 33.080 2.490 33.360 6.490 ;
        RECT 39.520 2.490 39.800 6.490 ;
      LAYER met3 ;
        RECT 36.260 204.465 37.840 204.795 ;
        RECT 32.960 201.745 34.540 202.075 ;
        RECT 36.260 199.025 37.840 199.355 ;
        RECT 11.910 198.320 15.910 198.470 ;
        RECT 11.910 198.020 17.120 198.320 ;
        RECT 11.910 197.870 15.910 198.020 ;
        RECT 12.435 196.960 12.765 196.975 ;
        RECT 16.820 196.960 17.120 198.020 ;
        RECT 12.435 196.660 17.120 196.960 ;
        RECT 12.435 196.645 12.765 196.660 ;
        RECT 32.960 196.305 34.540 196.635 ;
        RECT 36.260 193.585 37.840 193.915 ;
        RECT 32.960 190.865 34.540 191.195 ;
        RECT 36.260 188.145 37.840 188.475 ;
        RECT 79.595 186.090 79.925 186.095 ;
        RECT 79.340 186.080 79.925 186.090 ;
        RECT 79.140 185.780 79.925 186.080 ;
        RECT 79.340 185.770 79.925 185.780 ;
        RECT 79.595 185.765 79.925 185.770 ;
        RECT 32.960 185.425 34.540 185.755 ;
        RECT 67.635 184.040 67.965 184.055 ;
        RECT 75.455 184.040 75.785 184.055 ;
        RECT 83.275 184.040 83.605 184.055 ;
        RECT 67.635 183.740 83.605 184.040 ;
        RECT 67.635 183.725 67.965 183.740 ;
        RECT 75.455 183.725 75.785 183.740 ;
        RECT 83.275 183.725 83.605 183.740 ;
        RECT 117.775 184.050 118.105 184.055 ;
        RECT 117.775 184.040 118.360 184.050 ;
        RECT 117.775 183.740 118.560 184.040 ;
        RECT 117.775 183.730 118.360 183.740 ;
        RECT 117.775 183.725 118.105 183.730 ;
        RECT 115.015 183.360 115.345 183.375 ;
        RECT 120.535 183.360 120.865 183.375 ;
        RECT 115.015 183.060 120.865 183.360 ;
        RECT 115.015 183.045 115.345 183.060 ;
        RECT 120.535 183.045 120.865 183.060 ;
        RECT 36.260 182.705 37.840 183.035 ;
        RECT 141.235 181.320 141.565 181.335 ;
        RECT 144.570 181.320 148.570 181.470 ;
        RECT 141.235 181.020 148.570 181.320 ;
        RECT 141.235 181.005 141.565 181.020 ;
        RECT 144.570 180.870 148.570 181.020 ;
        RECT 32.960 179.985 34.540 180.315 ;
        RECT 34.515 179.280 34.845 179.295 ;
        RECT 37.275 179.280 37.605 179.295 ;
        RECT 34.515 178.980 37.605 179.280 ;
        RECT 34.515 178.965 34.845 178.980 ;
        RECT 37.275 178.965 37.605 178.980 ;
        RECT 140.775 177.920 141.105 177.935 ;
        RECT 144.570 177.920 148.570 178.070 ;
        RECT 140.775 177.620 148.570 177.920 ;
        RECT 140.775 177.605 141.105 177.620 ;
        RECT 36.260 177.265 37.840 177.595 ;
        RECT 144.570 177.470 148.570 177.620 ;
        RECT 110.875 177.240 111.205 177.255 ;
        RECT 116.855 177.240 117.185 177.255 ;
        RECT 110.875 176.940 117.185 177.240 ;
        RECT 110.875 176.925 111.205 176.940 ;
        RECT 116.855 176.925 117.185 176.940 ;
        RECT 115.015 175.880 115.345 175.895 ;
        RECT 123.755 175.880 124.085 175.895 ;
        RECT 115.015 175.580 124.085 175.880 ;
        RECT 115.015 175.565 115.345 175.580 ;
        RECT 123.755 175.565 124.085 175.580 ;
        RECT 16.115 175.200 16.445 175.215 ;
        RECT 15.900 174.885 16.445 175.200 ;
        RECT 15.900 174.670 16.200 174.885 ;
        RECT 11.910 174.220 16.200 174.670 ;
        RECT 32.960 174.545 34.540 174.875 ;
        RECT 138.935 174.520 139.265 174.535 ;
        RECT 144.570 174.520 148.570 174.670 ;
        RECT 138.935 174.220 148.570 174.520 ;
        RECT 11.910 174.070 15.910 174.220 ;
        RECT 138.935 174.205 139.265 174.220 ;
        RECT 144.570 174.070 148.570 174.220 ;
        RECT 75.455 173.840 75.785 173.855 ;
        RECT 77.295 173.840 77.625 173.855 ;
        RECT 80.515 173.840 80.845 173.855 ;
        RECT 75.455 173.540 80.845 173.840 ;
        RECT 75.455 173.525 75.785 173.540 ;
        RECT 77.295 173.525 77.625 173.540 ;
        RECT 80.515 173.525 80.845 173.540 ;
        RECT 113.635 173.160 113.965 173.175 ;
        RECT 120.535 173.160 120.865 173.175 ;
        RECT 113.635 172.860 120.865 173.160 ;
        RECT 113.635 172.845 113.965 172.860 ;
        RECT 120.535 172.845 120.865 172.860 ;
        RECT 118.695 172.480 119.025 172.495 ;
        RECT 121.915 172.490 122.245 172.495 ;
        RECT 121.660 172.480 122.245 172.490 ;
        RECT 118.695 172.180 121.080 172.480 ;
        RECT 121.460 172.180 122.245 172.480 ;
        RECT 118.695 172.165 119.025 172.180 ;
        RECT 36.260 171.825 37.840 172.155 ;
        RECT 120.780 171.815 121.080 172.180 ;
        RECT 121.660 172.170 122.245 172.180 ;
        RECT 121.915 172.165 122.245 172.170 ;
        RECT 75.915 171.800 76.245 171.815 ;
        RECT 81.895 171.800 82.225 171.815 ;
        RECT 75.915 171.500 82.225 171.800 ;
        RECT 75.915 171.485 76.245 171.500 ;
        RECT 81.895 171.485 82.225 171.500 ;
        RECT 111.335 171.800 111.665 171.815 ;
        RECT 117.980 171.800 118.360 171.810 ;
        RECT 118.695 171.800 119.025 171.815 ;
        RECT 120.780 171.800 121.325 171.815 ;
        RECT 121.915 171.800 122.245 171.815 ;
        RECT 111.335 171.500 119.025 171.800 ;
        RECT 120.540 171.500 122.245 171.800 ;
        RECT 111.335 171.485 111.665 171.500 ;
        RECT 117.980 171.490 118.360 171.500 ;
        RECT 118.695 171.485 119.025 171.500 ;
        RECT 120.995 171.485 121.325 171.500 ;
        RECT 121.915 171.485 122.245 171.500 ;
        RECT 69.475 171.120 69.805 171.135 ;
        RECT 79.135 171.120 79.465 171.135 ;
        RECT 69.475 170.820 79.465 171.120 ;
        RECT 69.475 170.805 69.805 170.820 ;
        RECT 79.135 170.805 79.465 170.820 ;
        RECT 141.695 171.120 142.025 171.135 ;
        RECT 144.570 171.120 148.570 171.270 ;
        RECT 141.695 170.820 148.570 171.120 ;
        RECT 141.695 170.805 142.025 170.820 ;
        RECT 144.570 170.670 148.570 170.820 ;
        RECT 32.960 169.105 34.540 169.435 ;
        RECT 132.495 167.720 132.825 167.735 ;
        RECT 144.570 167.720 148.570 167.870 ;
        RECT 132.495 167.420 148.570 167.720 ;
        RECT 132.495 167.405 132.825 167.420 ;
        RECT 144.570 167.270 148.570 167.420 ;
        RECT 36.260 166.385 37.840 166.715 ;
        RECT 35.180 165.000 35.560 165.010 ;
        RECT 35.895 165.000 36.225 165.015 ;
        RECT 35.180 164.700 36.225 165.000 ;
        RECT 35.180 164.690 35.560 164.700 ;
        RECT 35.895 164.685 36.225 164.700 ;
        RECT 138.935 164.320 139.265 164.335 ;
        RECT 144.570 164.320 148.570 164.470 ;
        RECT 138.935 164.020 148.570 164.320 ;
        RECT 138.935 164.005 139.265 164.020 ;
        RECT 32.960 163.665 34.540 163.995 ;
        RECT 144.570 163.870 148.570 164.020 ;
        RECT 116.855 162.960 117.185 162.975 ;
        RECT 123.295 162.960 123.625 162.975 ;
        RECT 116.855 162.660 123.625 162.960 ;
        RECT 116.855 162.645 117.185 162.660 ;
        RECT 123.295 162.645 123.625 162.660 ;
        RECT 119.155 162.280 119.485 162.295 ;
        RECT 120.535 162.280 120.865 162.295 ;
        RECT 121.915 162.280 122.245 162.295 ;
        RECT 119.155 161.980 122.245 162.280 ;
        RECT 119.155 161.965 119.485 161.980 ;
        RECT 120.535 161.965 120.865 161.980 ;
        RECT 121.915 161.965 122.245 161.980 ;
        RECT 16.115 161.600 16.445 161.615 ;
        RECT 15.900 161.285 16.445 161.600 ;
        RECT 117.775 161.600 118.105 161.615 ;
        RECT 121.455 161.600 121.785 161.615 ;
        RECT 117.775 161.300 121.785 161.600 ;
        RECT 117.775 161.285 118.105 161.300 ;
        RECT 121.455 161.285 121.785 161.300 ;
        RECT 15.900 161.070 16.200 161.285 ;
        RECT 11.910 160.620 16.200 161.070 ;
        RECT 36.260 160.945 37.840 161.275 ;
        RECT 52.915 160.920 53.245 160.935 ;
        RECT 56.135 160.920 56.465 160.935 ;
        RECT 79.595 160.930 79.925 160.935 ;
        RECT 52.915 160.620 56.465 160.920 ;
        RECT 11.910 160.470 15.910 160.620 ;
        RECT 52.915 160.605 53.245 160.620 ;
        RECT 56.135 160.605 56.465 160.620 ;
        RECT 79.340 160.920 79.925 160.930 ;
        RECT 140.775 160.920 141.105 160.935 ;
        RECT 144.570 160.920 148.570 161.070 ;
        RECT 79.340 160.620 80.150 160.920 ;
        RECT 140.775 160.620 148.570 160.920 ;
        RECT 79.340 160.610 79.925 160.620 ;
        RECT 79.595 160.605 79.925 160.610 ;
        RECT 140.775 160.605 141.105 160.620 ;
        RECT 144.570 160.470 148.570 160.620 ;
        RECT 111.335 160.240 111.665 160.255 ;
        RECT 115.475 160.240 115.805 160.255 ;
        RECT 111.335 159.940 115.805 160.240 ;
        RECT 111.335 159.925 111.665 159.940 ;
        RECT 115.475 159.925 115.805 159.940 ;
        RECT 32.960 158.225 34.540 158.555 ;
        RECT 140.775 157.520 141.105 157.535 ;
        RECT 144.570 157.520 148.570 157.670 ;
        RECT 140.775 157.220 148.570 157.520 ;
        RECT 140.775 157.205 141.105 157.220 ;
        RECT 144.570 157.070 148.570 157.220 ;
        RECT 36.260 155.505 37.840 155.835 ;
        RECT 140.775 154.120 141.105 154.135 ;
        RECT 144.570 154.120 148.570 154.270 ;
        RECT 140.775 153.820 148.570 154.120 ;
        RECT 140.775 153.805 141.105 153.820 ;
        RECT 144.570 153.670 148.570 153.820 ;
        RECT 32.960 152.785 34.540 153.115 ;
        RECT 142.155 150.720 142.485 150.735 ;
        RECT 144.570 150.720 148.570 150.870 ;
        RECT 142.155 150.420 148.570 150.720 ;
        RECT 142.155 150.405 142.485 150.420 ;
        RECT 36.260 150.065 37.840 150.395 ;
        RECT 144.570 150.270 148.570 150.420 ;
        RECT 16.115 148.000 16.445 148.015 ;
        RECT 15.900 147.685 16.445 148.000 ;
        RECT 15.900 147.470 16.200 147.685 ;
        RECT 11.910 147.020 16.200 147.470 ;
        RECT 32.960 147.345 34.540 147.675 ;
        RECT 140.775 147.320 141.105 147.335 ;
        RECT 144.570 147.320 148.570 147.470 ;
        RECT 140.775 147.020 148.570 147.320 ;
        RECT 11.910 146.870 15.910 147.020 ;
        RECT 140.775 147.005 141.105 147.020 ;
        RECT 144.570 146.870 148.570 147.020 ;
        RECT 121.455 146.650 121.785 146.655 ;
        RECT 121.455 146.640 122.040 146.650 ;
        RECT 121.230 146.340 122.040 146.640 ;
        RECT 121.455 146.330 122.040 146.340 ;
        RECT 121.455 146.325 121.785 146.330 ;
        RECT 36.260 144.625 37.840 144.955 ;
        RECT 11.910 143.920 15.910 144.070 ;
        RECT 19.335 143.920 19.665 143.935 ;
        RECT 11.910 143.620 19.665 143.920 ;
        RECT 11.910 143.470 15.910 143.620 ;
        RECT 19.335 143.605 19.665 143.620 ;
        RECT 138.935 143.920 139.265 143.935 ;
        RECT 144.570 143.920 148.570 144.070 ;
        RECT 138.935 143.620 148.570 143.920 ;
        RECT 138.935 143.605 139.265 143.620 ;
        RECT 144.570 143.470 148.570 143.620 ;
        RECT 32.960 141.905 34.540 142.235 ;
        RECT 32.215 140.520 32.545 140.535 ;
        RECT 41.415 140.520 41.745 140.535 ;
        RECT 32.215 140.220 41.745 140.520 ;
        RECT 32.215 140.205 32.545 140.220 ;
        RECT 41.415 140.205 41.745 140.220 ;
        RECT 140.775 140.520 141.105 140.535 ;
        RECT 144.570 140.520 148.570 140.670 ;
        RECT 140.775 140.220 148.570 140.520 ;
        RECT 140.775 140.205 141.105 140.220 ;
        RECT 144.570 140.070 148.570 140.220 ;
        RECT 36.260 139.185 37.840 139.515 ;
        RECT 87.415 138.480 87.745 138.495 ;
        RECT 90.175 138.480 90.505 138.495 ;
        RECT 87.415 138.180 90.505 138.480 ;
        RECT 87.415 138.165 87.745 138.180 ;
        RECT 90.175 138.165 90.505 138.180 ;
        RECT 120.075 138.480 120.405 138.495 ;
        RECT 125.595 138.480 125.925 138.495 ;
        RECT 133.875 138.480 134.205 138.495 ;
        RECT 120.075 138.180 134.205 138.480 ;
        RECT 120.075 138.165 120.405 138.180 ;
        RECT 125.595 138.165 125.925 138.180 ;
        RECT 133.875 138.165 134.205 138.180 ;
        RECT 138.935 137.120 139.265 137.135 ;
        RECT 144.570 137.120 148.570 137.270 ;
        RECT 138.935 136.820 148.570 137.120 ;
        RECT 138.935 136.805 139.265 136.820 ;
        RECT 32.960 136.465 34.540 136.795 ;
        RECT 144.570 136.670 148.570 136.820 ;
        RECT 36.260 133.745 37.840 134.075 ;
        RECT 140.775 133.720 141.105 133.735 ;
        RECT 144.570 133.720 148.570 133.870 ;
        RECT 140.775 133.420 148.570 133.720 ;
        RECT 140.775 133.405 141.105 133.420 ;
        RECT 144.570 133.270 148.570 133.420 ;
        RECT 32.960 131.025 34.540 131.355 ;
        RECT 118.695 130.320 119.025 130.335 ;
        RECT 138.015 130.320 138.345 130.335 ;
        RECT 118.695 130.020 138.345 130.320 ;
        RECT 118.695 130.005 119.025 130.020 ;
        RECT 138.015 130.005 138.345 130.020 ;
        RECT 140.775 130.320 141.105 130.335 ;
        RECT 144.570 130.320 148.570 130.470 ;
        RECT 140.775 130.020 148.570 130.320 ;
        RECT 140.775 130.005 141.105 130.020 ;
        RECT 144.570 129.870 148.570 130.020 ;
        RECT 120.075 129.640 120.405 129.655 ;
        RECT 124.675 129.640 125.005 129.655 ;
        RECT 120.075 129.340 125.005 129.640 ;
        RECT 120.075 129.325 120.405 129.340 ;
        RECT 124.675 129.325 125.005 129.340 ;
        RECT 36.260 128.305 37.840 128.635 ;
        RECT 35.180 127.600 35.560 127.610 ;
        RECT 35.895 127.600 36.225 127.615 ;
        RECT 37.735 127.600 38.065 127.615 ;
        RECT 35.180 127.300 38.065 127.600 ;
        RECT 35.180 127.290 35.560 127.300 ;
        RECT 35.895 127.285 36.225 127.300 ;
        RECT 37.735 127.285 38.065 127.300 ;
        RECT 140.775 126.920 141.105 126.935 ;
        RECT 144.570 126.920 148.570 127.070 ;
        RECT 140.775 126.620 148.570 126.920 ;
        RECT 140.775 126.605 141.105 126.620 ;
        RECT 144.570 126.470 148.570 126.620 ;
        RECT 32.960 125.585 34.540 125.915 ;
        RECT 48.775 124.200 49.105 124.215 ;
        RECT 52.915 124.200 53.245 124.215 ;
        RECT 48.775 123.900 53.245 124.200 ;
        RECT 48.775 123.885 49.105 123.900 ;
        RECT 52.915 123.885 53.245 123.900 ;
        RECT 140.775 123.520 141.105 123.535 ;
        RECT 144.570 123.520 148.570 123.670 ;
        RECT 140.775 123.220 148.570 123.520 ;
        RECT 140.775 123.205 141.105 123.220 ;
        RECT 36.260 122.865 37.840 123.195 ;
        RECT 144.570 123.070 148.570 123.220 ;
        RECT 32.960 120.145 34.540 120.475 ;
        RECT 140.775 120.120 141.105 120.135 ;
        RECT 144.570 120.120 148.570 120.270 ;
        RECT 140.775 119.820 148.570 120.120 ;
        RECT 140.775 119.805 141.105 119.820 ;
        RECT 144.570 119.670 148.570 119.820 ;
        RECT 36.260 117.425 37.840 117.755 ;
        RECT 138.935 116.720 139.265 116.735 ;
        RECT 144.570 116.720 148.570 116.870 ;
        RECT 138.935 116.420 148.570 116.720 ;
        RECT 138.935 116.405 139.265 116.420 ;
        RECT 144.570 116.270 148.570 116.420 ;
        RECT 32.960 114.705 34.540 115.035 ;
        RECT 34.515 113.320 34.845 113.335 ;
        RECT 40.035 113.320 40.365 113.335 ;
        RECT 42.795 113.320 43.125 113.335 ;
        RECT 34.515 113.020 43.125 113.320 ;
        RECT 34.515 113.005 34.845 113.020 ;
        RECT 40.035 113.005 40.365 113.020 ;
        RECT 42.795 113.005 43.125 113.020 ;
        RECT 140.775 113.320 141.105 113.335 ;
        RECT 144.570 113.320 148.570 113.470 ;
        RECT 140.775 113.020 148.570 113.320 ;
        RECT 140.775 113.005 141.105 113.020 ;
        RECT 144.570 112.870 148.570 113.020 ;
        RECT 36.260 111.985 37.840 112.315 ;
        RECT 66.715 109.920 67.045 109.935 ;
        RECT 72.695 109.920 73.025 109.935 ;
        RECT 66.715 109.620 73.025 109.920 ;
        RECT 66.715 109.605 67.045 109.620 ;
        RECT 72.695 109.605 73.025 109.620 ;
        RECT 142.615 109.920 142.945 109.935 ;
        RECT 144.570 109.920 148.570 110.070 ;
        RECT 142.615 109.620 148.570 109.920 ;
        RECT 142.615 109.605 142.945 109.620 ;
        RECT 32.960 109.265 34.540 109.595 ;
        RECT 144.570 109.470 148.570 109.620 ;
        RECT 36.260 106.545 37.840 106.875 ;
        RECT 140.775 106.520 141.105 106.535 ;
        RECT 144.570 106.520 148.570 106.670 ;
        RECT 140.775 106.220 148.570 106.520 ;
        RECT 140.775 106.205 141.105 106.220 ;
        RECT 144.570 106.070 148.570 106.220 ;
        RECT 95.235 105.840 95.565 105.855 ;
        RECT 120.995 105.840 121.325 105.855 ;
        RECT 95.235 105.540 121.325 105.840 ;
        RECT 95.235 105.525 95.565 105.540 ;
        RECT 120.995 105.525 121.325 105.540 ;
        RECT 69.935 105.160 70.265 105.175 ;
        RECT 74.075 105.160 74.405 105.175 ;
        RECT 69.935 104.860 74.405 105.160 ;
        RECT 69.935 104.845 70.265 104.860 ;
        RECT 74.075 104.845 74.405 104.860 ;
        RECT 107.655 105.160 107.985 105.175 ;
        RECT 128.355 105.160 128.685 105.175 ;
        RECT 107.655 104.860 128.685 105.160 ;
        RECT 107.655 104.845 107.985 104.860 ;
        RECT 128.355 104.845 128.685 104.860 ;
        RECT 32.960 103.825 34.540 104.155 ;
        RECT 138.935 103.120 139.265 103.135 ;
        RECT 144.570 103.120 148.570 103.270 ;
        RECT 138.935 102.820 148.570 103.120 ;
        RECT 138.935 102.805 139.265 102.820 ;
        RECT 144.570 102.670 148.570 102.820 ;
        RECT 36.260 101.105 37.840 101.435 ;
        RECT 140.775 99.720 141.105 99.735 ;
        RECT 144.570 99.720 148.570 99.870 ;
        RECT 140.775 99.420 148.570 99.720 ;
        RECT 140.775 99.405 141.105 99.420 ;
        RECT 144.570 99.270 148.570 99.420 ;
        RECT 32.960 98.385 34.540 98.715 ;
        RECT 124.675 98.360 125.005 98.375 ;
        RECT 135.715 98.360 136.045 98.375 ;
        RECT 124.675 98.060 136.045 98.360 ;
        RECT 124.675 98.045 125.005 98.060 ;
        RECT 135.715 98.045 136.045 98.060 ;
        RECT 88.795 97.680 89.125 97.695 ;
        RECT 137.555 97.680 137.885 97.695 ;
        RECT 88.795 97.380 137.885 97.680 ;
        RECT 88.795 97.365 89.125 97.380 ;
        RECT 137.555 97.365 137.885 97.380 ;
        RECT 88.795 96.320 89.125 96.335 ;
        RECT 119.155 96.320 119.485 96.335 ;
        RECT 88.795 96.020 119.485 96.320 ;
        RECT 88.795 96.005 89.125 96.020 ;
        RECT 119.155 96.005 119.485 96.020 ;
        RECT 140.775 96.320 141.105 96.335 ;
        RECT 144.570 96.320 148.570 96.470 ;
        RECT 140.775 96.020 148.570 96.320 ;
        RECT 140.775 96.005 141.105 96.020 ;
        RECT 36.260 95.665 37.840 95.995 ;
        RECT 144.570 95.870 148.570 96.020 ;
        RECT 32.960 92.945 34.540 93.275 ;
        RECT 140.775 92.920 141.105 92.935 ;
        RECT 144.570 92.920 148.570 93.070 ;
        RECT 140.775 92.620 148.570 92.920 ;
        RECT 140.775 92.605 141.105 92.620 ;
        RECT 144.570 92.470 148.570 92.620 ;
        RECT 36.260 90.225 37.840 90.555 ;
        RECT 112.715 89.520 113.045 89.535 ;
        RECT 114.555 89.520 114.885 89.535 ;
        RECT 112.715 89.220 114.885 89.520 ;
        RECT 112.715 89.205 113.045 89.220 ;
        RECT 114.555 89.205 114.885 89.220 ;
        RECT 138.935 89.520 139.265 89.535 ;
        RECT 144.570 89.520 148.570 89.670 ;
        RECT 138.935 89.220 148.570 89.520 ;
        RECT 138.935 89.205 139.265 89.220 ;
        RECT 144.570 89.070 148.570 89.220 ;
        RECT 99.375 88.840 99.705 88.855 ;
        RECT 129.275 88.840 129.605 88.855 ;
        RECT 99.375 88.540 129.605 88.840 ;
        RECT 99.375 88.525 99.705 88.540 ;
        RECT 129.275 88.525 129.605 88.540 ;
        RECT 32.960 87.505 34.540 87.835 ;
        RECT 110.415 86.810 110.745 86.815 ;
        RECT 110.415 86.800 111.000 86.810 ;
        RECT 114.555 86.800 114.885 86.815 ;
        RECT 131.115 86.800 131.445 86.815 ;
        RECT 110.415 86.500 111.200 86.800 ;
        RECT 114.555 86.500 131.445 86.800 ;
        RECT 110.415 86.490 111.000 86.500 ;
        RECT 110.415 86.485 110.745 86.490 ;
        RECT 114.555 86.485 114.885 86.500 ;
        RECT 131.115 86.485 131.445 86.500 ;
        RECT 140.775 86.120 141.105 86.135 ;
        RECT 144.570 86.120 148.570 86.270 ;
        RECT 140.775 85.820 148.570 86.120 ;
        RECT 140.775 85.805 141.105 85.820 ;
        RECT 144.570 85.670 148.570 85.820 ;
        RECT 109.035 85.440 109.365 85.455 ;
        RECT 116.395 85.440 116.725 85.455 ;
        RECT 109.035 85.140 116.725 85.440 ;
        RECT 109.035 85.125 109.365 85.140 ;
        RECT 116.395 85.125 116.725 85.140 ;
        RECT 36.260 84.785 37.840 85.115 ;
        RECT 110.415 84.770 110.745 84.775 ;
        RECT 110.415 84.760 111.000 84.770 ;
        RECT 110.190 84.460 111.000 84.760 ;
        RECT 110.415 84.450 111.000 84.460 ;
        RECT 112.715 84.760 113.045 84.775 ;
        RECT 119.155 84.760 119.485 84.775 ;
        RECT 112.715 84.460 119.485 84.760 ;
        RECT 110.415 84.445 110.745 84.450 ;
        RECT 112.715 84.445 113.045 84.460 ;
        RECT 119.155 84.445 119.485 84.460 ;
        RECT 96.615 84.080 96.945 84.095 ;
        RECT 97.535 84.080 97.865 84.095 ;
        RECT 122.375 84.080 122.705 84.095 ;
        RECT 96.615 83.780 122.705 84.080 ;
        RECT 96.615 83.765 96.945 83.780 ;
        RECT 97.535 83.765 97.865 83.780 ;
        RECT 122.375 83.765 122.705 83.780 ;
        RECT 115.015 83.400 115.345 83.415 ;
        RECT 117.315 83.400 117.645 83.415 ;
        RECT 115.015 83.100 117.645 83.400 ;
        RECT 115.015 83.085 115.345 83.100 ;
        RECT 117.315 83.085 117.645 83.100 ;
        RECT 140.775 82.720 141.105 82.735 ;
        RECT 144.570 82.720 148.570 82.870 ;
        RECT 140.775 82.420 148.570 82.720 ;
        RECT 140.775 82.405 141.105 82.420 ;
        RECT 32.960 82.065 34.540 82.395 ;
        RECT 144.570 82.270 148.570 82.420 ;
        RECT 36.260 79.345 37.840 79.675 ;
        RECT 46.855 53.980 47.185 53.995 ;
        RECT 50.275 53.980 54.275 54.130 ;
        RECT 46.855 53.680 54.275 53.980 ;
        RECT 46.855 53.665 47.185 53.680 ;
        RECT 50.275 53.530 54.275 53.680 ;
        RECT 44.095 50.580 44.425 50.595 ;
        RECT 50.275 50.580 54.275 50.730 ;
        RECT 44.095 50.280 54.275 50.580 ;
        RECT 44.095 50.265 44.425 50.280 ;
        RECT 50.275 50.130 54.275 50.280 ;
        RECT 28.280 48.565 29.860 48.895 ;
        RECT 45.475 47.180 45.805 47.195 ;
        RECT 50.275 47.180 54.275 47.330 ;
        RECT 45.475 46.880 54.275 47.180 ;
        RECT 45.475 46.865 45.805 46.880 ;
        RECT 50.275 46.730 54.275 46.880 ;
        RECT 31.580 45.845 33.160 46.175 ;
        RECT 23.395 45.140 23.725 45.155 ;
        RECT 27.535 45.140 27.865 45.155 ;
        RECT 40.875 45.140 41.205 45.155 ;
        RECT 23.395 44.840 41.205 45.140 ;
        RECT 23.395 44.825 23.725 44.840 ;
        RECT 27.535 44.825 27.865 44.840 ;
        RECT 40.875 44.825 41.205 44.840 ;
        RECT 7.230 43.780 11.230 43.930 ;
        RECT 24.775 43.780 25.105 43.795 ;
        RECT 7.230 43.480 25.105 43.780 ;
        RECT 7.230 43.330 11.230 43.480 ;
        RECT 24.775 43.465 25.105 43.480 ;
        RECT 46.855 43.780 47.185 43.795 ;
        RECT 50.275 43.780 54.275 43.930 ;
        RECT 46.855 43.480 54.275 43.780 ;
        RECT 46.855 43.465 47.185 43.480 ;
        RECT 28.280 43.125 29.860 43.455 ;
        RECT 50.275 43.330 54.275 43.480 ;
        RECT 7.230 40.380 11.230 40.530 ;
        RECT 31.580 40.405 33.160 40.735 ;
        RECT 13.735 40.380 14.065 40.395 ;
        RECT 7.230 40.080 14.065 40.380 ;
        RECT 7.230 39.930 11.230 40.080 ;
        RECT 13.735 40.065 14.065 40.080 ;
        RECT 46.855 40.380 47.185 40.395 ;
        RECT 50.275 40.380 54.275 40.530 ;
        RECT 46.855 40.080 54.275 40.380 ;
        RECT 46.855 40.065 47.185 40.080 ;
        RECT 50.275 39.930 54.275 40.080 ;
        RECT 28.280 37.685 29.860 38.015 ;
        RECT 44.555 36.980 44.885 36.995 ;
        RECT 50.275 36.980 54.275 37.130 ;
        RECT 44.555 36.680 54.275 36.980 ;
        RECT 44.555 36.665 44.885 36.680 ;
        RECT 50.275 36.530 54.275 36.680 ;
        RECT 31.580 34.965 33.160 35.295 ;
        RECT 7.230 33.580 11.230 33.730 ;
        RECT 13.735 33.580 14.065 33.595 ;
        RECT 7.230 33.280 14.065 33.580 ;
        RECT 7.230 33.130 11.230 33.280 ;
        RECT 13.735 33.265 14.065 33.280 ;
        RECT 46.855 33.580 47.185 33.595 ;
        RECT 50.275 33.580 54.275 33.730 ;
        RECT 46.855 33.280 54.275 33.580 ;
        RECT 46.855 33.265 47.185 33.280 ;
        RECT 50.275 33.130 54.275 33.280 ;
        RECT 28.280 32.245 29.860 32.575 ;
        RECT 41.795 30.180 42.125 30.195 ;
        RECT 50.275 30.180 54.275 30.330 ;
        RECT 41.795 29.880 54.275 30.180 ;
        RECT 41.795 29.865 42.125 29.880 ;
        RECT 31.580 29.525 33.160 29.855 ;
        RECT 50.275 29.730 54.275 29.880 ;
        RECT 7.230 26.780 11.230 26.930 ;
        RECT 28.280 26.805 29.860 27.135 ;
        RECT 13.735 26.780 14.065 26.795 ;
        RECT 7.230 26.480 14.065 26.780 ;
        RECT 7.230 26.330 11.230 26.480 ;
        RECT 13.735 26.465 14.065 26.480 ;
        RECT 39.495 26.780 39.825 26.795 ;
        RECT 50.275 26.780 54.275 26.930 ;
        RECT 39.495 26.480 54.275 26.780 ;
        RECT 39.495 26.465 39.825 26.480 ;
        RECT 50.275 26.330 54.275 26.480 ;
        RECT 31.580 24.085 33.160 24.415 ;
        RECT 43.175 23.380 43.505 23.395 ;
        RECT 50.275 23.380 54.275 23.530 ;
        RECT 43.175 23.080 54.275 23.380 ;
        RECT 43.175 23.065 43.505 23.080 ;
        RECT 50.275 22.930 54.275 23.080 ;
        RECT 28.280 21.365 29.860 21.695 ;
        RECT 40.875 19.980 41.205 19.995 ;
        RECT 50.275 19.980 54.275 20.130 ;
        RECT 40.875 19.680 54.275 19.980 ;
        RECT 40.875 19.665 41.205 19.680 ;
        RECT 50.275 19.530 54.275 19.680 ;
        RECT 31.580 18.645 33.160 18.975 ;
        RECT 11.435 17.260 11.765 17.275 ;
        RECT 11.220 16.945 11.765 17.260 ;
        RECT 11.220 16.730 11.520 16.945 ;
        RECT 7.230 16.280 11.520 16.730 ;
        RECT 38.115 16.580 38.445 16.595 ;
        RECT 50.275 16.580 54.275 16.730 ;
        RECT 38.115 16.280 54.275 16.580 ;
        RECT 7.230 16.130 11.230 16.280 ;
        RECT 38.115 16.265 38.445 16.280 ;
        RECT 28.280 15.925 29.860 16.255 ;
        RECT 50.275 16.130 54.275 16.280 ;
        RECT 31.580 13.205 33.160 13.535 ;
        RECT 42.715 13.180 43.045 13.195 ;
        RECT 50.275 13.180 54.275 13.330 ;
        RECT 42.715 12.880 54.275 13.180 ;
        RECT 42.715 12.865 43.045 12.880 ;
        RECT 50.275 12.730 54.275 12.880 ;
        RECT 46.395 9.780 46.725 9.795 ;
        RECT 50.275 9.780 54.275 9.930 ;
        RECT 46.395 9.480 54.275 9.780 ;
        RECT 46.395 9.465 46.725 9.480 ;
        RECT 50.275 9.330 54.275 9.480 ;
      LAYER met4 ;
        RECT 64.090 225.055 64.145 225.385 ;
        RECT 66.455 224.965 66.550 225.295 ;
        RECT 69.305 225.135 69.310 225.465 ;
        RECT 69.610 225.135 69.635 225.465 ;
        RECT 71.995 224.895 72.070 225.225 ;
        RECT 74.785 224.945 74.830 225.275 ;
        RECT 77.515 224.760 77.590 225.085 ;
        RECT 80.295 224.925 80.350 225.255 ;
        RECT 83.025 224.760 83.110 225.085 ;
        RECT 85.795 224.915 85.870 225.245 ;
        RECT 88.535 224.915 88.630 225.245 ;
        RECT 91.350 224.835 91.390 225.165 ;
        RECT 94.125 224.815 94.150 225.145 ;
        RECT 94.450 224.815 94.455 225.145 ;
        RECT 77.515 224.755 77.845 224.760 ;
        RECT 83.025 224.755 83.355 224.760 ;
        RECT 6.000 197.560 6.140 199.160 ;
        RECT 32.950 79.270 34.550 204.870 ;
        RECT 35.205 164.685 35.535 165.015 ;
        RECT 35.220 127.615 35.520 164.685 ;
        RECT 35.205 127.285 35.535 127.615 ;
        RECT 36.250 79.270 37.850 204.870 ;
        RECT 79.365 185.765 79.695 186.095 ;
        RECT 79.380 160.935 79.680 185.765 ;
        RECT 118.005 183.725 118.335 184.055 ;
        RECT 118.020 171.815 118.320 183.725 ;
        RECT 121.685 172.165 122.015 172.495 ;
        RECT 118.005 171.485 118.335 171.815 ;
        RECT 79.365 160.605 79.695 160.935 ;
        RECT 121.700 146.655 122.000 172.165 ;
        RECT 121.685 146.325 122.015 146.655 ;
        RECT 110.645 86.485 110.975 86.815 ;
        RECT 110.660 84.775 110.960 86.485 ;
        RECT 110.645 84.445 110.975 84.775 ;
        RECT 28.270 13.130 29.870 48.970 ;
        RECT 31.570 13.130 33.170 48.970 ;
  END
END tt_um_tim2305_adc_dac
END LIBRARY

