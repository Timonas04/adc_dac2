MACRO bit4_encoder
  CLASS BLOCK ;
  FOREIGN bit4_encoder ;
  ORIGIN 0.000 0.000 ;
  SIZE 47.045 BY 57.765 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 46.480 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 46.480 ;
    END
  END VPWR
  PIN bus0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 53.765 22.910 57.765 ;
    END
  END bus0[0]
  PIN bus0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END bus0[1]
  PIN bus0[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END bus0[2]
  PIN bus0[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END bus0[3]
  PIN bus1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 53.765 26.130 57.765 ;
    END
  END bus1[0]
  PIN bus1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END bus1[1]
  PIN bus1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END bus1[2]
  PIN bus1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END bus1[3]
  PIN bus2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 53.765 32.570 57.765 ;
    END
  END bus2[0]
  PIN bus2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 19.410 53.765 19.690 57.765 ;
    END
  END bus2[1]
  PIN bus2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END bus2[2]
  PIN bus2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END bus2[3]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END clk
  PIN compr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 6.840 47.045 7.440 ;
    END
  END compr[0]
  PIN compr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 51.040 47.045 51.640 ;
    END
  END compr[10]
  PIN compr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 44.240 47.045 44.840 ;
    END
  END compr[11]
  PIN compr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 37.440 47.045 38.040 ;
    END
  END compr[12]
  PIN compr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 47.640 47.045 48.240 ;
    END
  END compr[13]
  PIN compr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 29.070 53.765 29.350 57.765 ;
    END
  END compr[14]
  PIN compr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 17.040 47.045 17.640 ;
    END
  END compr[1]
  PIN compr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 20.440 47.045 21.040 ;
    END
  END compr[2]
  PIN compr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 13.640 47.045 14.240 ;
    END
  END compr[3]
  PIN compr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 10.240 47.045 10.840 ;
    END
  END compr[4]
  PIN compr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 23.840 47.045 24.440 ;
    END
  END compr[5]
  PIN compr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 27.240 47.045 27.840 ;
    END
  END compr[6]
  PIN compr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 30.640 47.045 31.240 ;
    END
  END compr[7]
  PIN compr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 34.040 47.045 34.640 ;
    END
  END compr[8]
  PIN compr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 43.045 40.840 47.045 41.440 ;
    END
  END compr[9]
  OBS
      LAYER nwell ;
        RECT 5.330 44.825 41.590 46.430 ;
      LAYER pwell ;
        RECT 5.525 43.625 6.895 44.435 ;
        RECT 6.905 43.625 12.415 44.435 ;
        RECT 13.830 44.305 15.175 44.535 ;
        RECT 13.345 43.625 15.175 44.305 ;
        RECT 15.315 43.625 18.315 44.535 ;
        RECT 18.415 43.710 18.845 44.495 ;
        RECT 22.440 44.305 23.360 44.535 ;
        RECT 19.895 43.625 23.360 44.305 ;
        RECT 24.385 44.305 25.730 44.535 ;
        RECT 28.880 44.305 29.800 44.535 ;
        RECT 24.385 43.625 26.215 44.305 ;
        RECT 26.335 43.625 29.800 44.305 ;
        RECT 29.905 43.625 31.275 44.405 ;
        RECT 31.295 43.710 31.725 44.495 ;
        RECT 32.665 44.305 34.010 44.535 ;
        RECT 32.665 43.625 34.495 44.305 ;
        RECT 34.505 43.625 35.875 44.435 ;
        RECT 35.885 43.625 37.255 44.405 ;
        RECT 37.265 43.625 38.635 44.405 ;
        RECT 38.645 43.625 40.015 44.405 ;
        RECT 40.025 43.625 41.395 44.435 ;
        RECT 5.665 43.415 5.835 43.625 ;
        RECT 7.045 43.415 7.215 43.625 ;
        RECT 10.720 43.465 10.840 43.575 ;
        RECT 12.575 43.470 12.735 43.580 ;
        RECT 13.485 43.435 13.655 43.625 ;
        RECT 18.085 43.415 18.255 43.625 ;
        RECT 18.545 43.415 18.715 43.605 ;
        RECT 19.015 43.470 19.175 43.580 ;
        RECT 19.925 43.435 20.095 43.625 ;
        RECT 23.615 43.470 23.775 43.580 ;
        RECT 25.905 43.435 26.075 43.625 ;
        RECT 26.365 43.435 26.535 43.625 ;
        RECT 30.055 43.605 30.225 43.625 ;
        RECT 27.745 43.435 27.915 43.605 ;
        RECT 27.745 43.415 27.910 43.435 ;
        RECT 28.205 43.415 28.375 43.605 ;
        RECT 30.045 43.435 30.225 43.605 ;
        RECT 30.045 43.415 30.215 43.435 ;
        RECT 31.885 43.415 32.055 43.605 ;
        RECT 34.185 43.435 34.355 43.625 ;
        RECT 34.645 43.435 34.815 43.625 ;
        RECT 35.105 43.415 35.275 43.605 ;
        RECT 36.945 43.435 37.115 43.625 ;
        RECT 38.325 43.435 38.495 43.625 ;
        RECT 39.695 43.415 39.865 43.625 ;
        RECT 41.085 43.415 41.255 43.625 ;
        RECT 5.525 42.605 6.895 43.415 ;
        RECT 6.905 42.605 10.575 43.415 ;
        RECT 11.085 42.735 18.395 43.415 ;
        RECT 18.405 42.735 25.715 43.415 ;
        RECT 11.085 42.505 12.435 42.735 ;
        RECT 13.970 42.515 14.880 42.735 ;
        RECT 21.920 42.515 22.830 42.735 ;
        RECT 24.365 42.505 25.715 42.735 ;
        RECT 26.075 42.735 27.910 43.415 ;
        RECT 28.065 42.735 29.895 43.415 ;
        RECT 26.075 42.505 27.005 42.735 ;
        RECT 28.550 42.505 29.895 42.735 ;
        RECT 29.915 42.505 31.265 43.415 ;
        RECT 31.295 42.545 31.725 43.330 ;
        RECT 31.825 42.505 34.825 43.415 ;
        RECT 35.075 42.735 38.540 43.415 ;
        RECT 37.620 42.505 38.540 42.735 ;
        RECT 38.645 42.635 40.015 43.415 ;
        RECT 40.025 42.605 41.395 43.415 ;
      LAYER nwell ;
        RECT 5.330 39.385 41.590 42.215 ;
      LAYER pwell ;
        RECT 5.525 38.185 6.895 38.995 ;
        RECT 10.420 38.865 11.330 39.085 ;
        RECT 12.865 38.865 14.215 39.095 ;
        RECT 6.905 38.185 14.215 38.865 ;
        RECT 14.360 38.865 15.280 39.095 ;
        RECT 14.360 38.185 17.825 38.865 ;
        RECT 18.415 38.270 18.845 39.055 ;
        RECT 18.865 38.865 19.795 39.095 ;
        RECT 24.515 38.865 25.445 39.095 ;
        RECT 18.865 38.185 22.765 38.865 ;
        RECT 23.610 38.185 25.445 38.865 ;
        RECT 25.775 38.185 27.125 39.095 ;
        RECT 30.660 38.865 31.570 39.085 ;
        RECT 33.105 38.865 34.455 39.095 ;
        RECT 36.015 38.865 36.945 39.095 ;
        RECT 27.145 38.185 34.455 38.865 ;
        RECT 35.110 38.185 36.945 38.865 ;
        RECT 37.265 38.185 38.635 38.965 ;
        RECT 38.645 38.185 40.015 38.965 ;
        RECT 40.025 38.185 41.395 38.995 ;
        RECT 5.665 37.975 5.835 38.185 ;
        RECT 7.045 37.995 7.215 38.185 ;
        RECT 8.425 37.975 8.595 38.165 ;
        RECT 9.160 37.975 9.330 38.165 ;
        RECT 13.025 37.975 13.195 38.165 ;
        RECT 17.625 37.995 17.795 38.185 ;
        RECT 18.080 38.025 18.200 38.135 ;
        RECT 19.280 37.995 19.450 38.185 ;
        RECT 23.610 38.165 23.775 38.185 ;
        RECT 23.145 38.135 23.315 38.165 ;
        RECT 23.140 38.025 23.315 38.135 ;
        RECT 23.145 37.975 23.315 38.025 ;
        RECT 23.605 37.995 23.775 38.165 ;
        RECT 26.825 37.975 26.995 38.185 ;
        RECT 27.285 37.975 27.455 38.185 ;
        RECT 35.110 38.165 35.275 38.185 ;
        RECT 5.525 37.165 6.895 37.975 ;
        RECT 6.905 37.295 8.735 37.975 ;
        RECT 8.745 37.295 12.645 37.975 ;
        RECT 6.905 37.065 8.250 37.295 ;
        RECT 8.745 37.065 9.675 37.295 ;
        RECT 12.885 37.165 14.255 37.975 ;
        RECT 14.350 37.295 23.455 37.975 ;
        RECT 23.560 37.295 27.025 37.975 ;
        RECT 23.560 37.065 24.480 37.295 ;
        RECT 27.145 37.165 28.515 37.975 ;
        RECT 28.670 37.945 28.840 38.165 ;
        RECT 31.885 37.975 32.055 38.165 ;
        RECT 34.640 38.025 34.760 38.135 ;
        RECT 35.105 37.995 35.275 38.165 ;
        RECT 35.565 37.975 35.735 38.165 ;
        RECT 37.405 37.995 37.575 38.185 ;
        RECT 39.255 38.020 39.415 38.130 ;
        RECT 39.695 37.995 39.865 38.185 ;
        RECT 41.085 37.975 41.255 38.185 ;
        RECT 30.330 37.945 31.275 37.975 ;
        RECT 28.525 37.265 31.275 37.945 ;
        RECT 30.330 37.065 31.275 37.265 ;
        RECT 31.295 37.105 31.725 37.890 ;
        RECT 31.825 37.065 35.275 37.975 ;
        RECT 35.505 37.065 38.955 37.975 ;
        RECT 40.025 37.165 41.395 37.975 ;
      LAYER nwell ;
        RECT 5.330 33.945 41.590 36.775 ;
      LAYER pwell ;
        RECT 5.525 32.745 6.895 33.555 ;
        RECT 6.905 33.425 7.835 33.655 ;
        RECT 14.560 33.425 15.470 33.645 ;
        RECT 17.005 33.425 18.355 33.655 ;
        RECT 6.905 32.745 10.805 33.425 ;
        RECT 11.045 32.745 18.355 33.425 ;
        RECT 18.415 32.830 18.845 33.615 ;
        RECT 22.380 33.425 23.290 33.645 ;
        RECT 24.825 33.425 26.175 33.655 ;
        RECT 18.865 32.745 26.175 33.425 ;
        RECT 26.685 33.425 28.050 33.655 ;
        RECT 26.685 32.745 29.895 33.425 ;
        RECT 30.905 32.745 33.905 33.655 ;
        RECT 34.045 32.745 35.395 33.655 ;
        RECT 35.965 32.745 39.415 33.655 ;
        RECT 40.025 32.745 41.395 33.555 ;
        RECT 5.665 32.535 5.835 32.745 ;
        RECT 7.320 32.555 7.490 32.745 ;
        RECT 11.185 32.555 11.355 32.745 ;
        RECT 13.945 32.535 14.115 32.725 ;
        RECT 14.405 32.535 14.575 32.725 ;
        RECT 17.160 32.585 17.280 32.695 ;
        RECT 17.625 32.535 17.795 32.725 ;
        RECT 19.005 32.555 19.175 32.745 ;
        RECT 26.360 32.585 26.480 32.695 ;
        RECT 29.580 32.555 29.750 32.745 ;
        RECT 30.045 32.535 30.215 32.725 ;
        RECT 30.515 32.580 30.675 32.690 ;
        RECT 30.965 32.555 31.135 32.745 ;
        RECT 34.190 32.725 34.360 32.745 ;
        RECT 5.525 31.725 6.895 32.535 ;
        RECT 6.945 31.855 14.255 32.535 ;
        RECT 6.945 31.625 8.295 31.855 ;
        RECT 9.830 31.635 10.740 31.855 ;
        RECT 14.265 31.725 17.015 32.535 ;
        RECT 17.485 31.855 26.590 32.535 ;
        RECT 26.780 31.855 30.245 32.535 ;
        RECT 31.880 32.505 32.050 32.725 ;
        RECT 34.185 32.555 34.360 32.725 ;
        RECT 35.560 32.585 35.680 32.695 ;
        RECT 36.025 32.555 36.195 32.745 ;
        RECT 36.940 32.585 37.060 32.695 ;
        RECT 34.185 32.535 34.355 32.555 ;
        RECT 38.320 32.535 38.490 32.725 ;
        RECT 39.705 32.695 39.875 32.725 ;
        RECT 39.700 32.585 39.875 32.695 ;
        RECT 39.705 32.535 39.875 32.585 ;
        RECT 41.085 32.535 41.255 32.745 ;
        RECT 33.080 32.505 34.035 32.535 ;
        RECT 26.780 31.625 27.700 31.855 ;
        RECT 31.295 31.665 31.725 32.450 ;
        RECT 31.755 31.825 34.035 32.505 ;
        RECT 33.080 31.625 34.035 31.825 ;
        RECT 34.045 31.725 36.795 32.535 ;
        RECT 37.285 31.625 38.635 32.535 ;
        RECT 38.645 31.755 40.015 32.535 ;
        RECT 40.025 31.725 41.395 32.535 ;
      LAYER nwell ;
        RECT 5.330 28.505 41.590 31.335 ;
      LAYER pwell ;
        RECT 5.525 27.305 6.895 28.115 ;
        RECT 6.905 27.305 8.275 28.115 ;
        RECT 10.940 27.985 11.860 28.215 ;
        RECT 8.395 27.305 11.860 27.985 ;
        RECT 12.060 27.985 12.980 28.215 ;
        RECT 12.060 27.305 15.525 27.985 ;
        RECT 15.645 27.305 18.395 28.115 ;
        RECT 18.415 27.390 18.845 28.175 ;
        RECT 18.885 27.305 20.235 28.215 ;
        RECT 20.315 27.305 24.375 28.215 ;
        RECT 24.480 27.985 25.400 28.215 ;
        RECT 24.480 27.305 27.945 27.985 ;
        RECT 28.065 27.305 29.435 28.115 ;
        RECT 29.445 28.015 30.395 28.215 ;
        RECT 29.445 27.335 33.115 28.015 ;
        RECT 29.445 27.305 30.395 27.335 ;
        RECT 5.665 27.095 5.835 27.305 ;
        RECT 7.045 27.115 7.215 27.305 ;
        RECT 8.425 27.095 8.595 27.305 ;
        RECT 8.880 27.145 9.000 27.255 ;
        RECT 9.620 27.095 9.790 27.285 ;
        RECT 13.485 27.095 13.655 27.285 ;
        RECT 15.325 27.115 15.495 27.305 ;
        RECT 15.785 27.115 15.955 27.305 ;
        RECT 19.920 27.115 20.090 27.305 ;
        RECT 21.120 27.095 21.290 27.285 ;
        RECT 24.065 27.115 24.235 27.305 ;
        RECT 27.745 27.115 27.915 27.305 ;
        RECT 28.205 27.095 28.375 27.305 ;
        RECT 28.665 27.095 28.835 27.285 ;
        RECT 32.800 27.115 32.970 27.335 ;
        RECT 33.125 27.305 34.475 28.215 ;
        RECT 34.505 27.305 35.875 28.085 ;
        RECT 36.025 27.305 39.475 28.215 ;
        RECT 40.025 27.305 41.395 28.115 ;
        RECT 33.270 27.115 33.440 27.305 ;
        RECT 34.655 27.285 34.825 27.305 ;
        RECT 34.640 27.115 34.825 27.285 ;
        RECT 35.115 27.140 35.275 27.250 ;
        RECT 34.640 27.095 34.810 27.115 ;
        RECT 39.245 27.095 39.415 27.305 ;
        RECT 39.700 27.145 39.820 27.255 ;
        RECT 41.085 27.095 41.255 27.305 ;
        RECT 5.525 26.285 6.895 27.095 ;
        RECT 6.905 26.415 8.735 27.095 ;
        RECT 9.205 26.415 13.105 27.095 ;
        RECT 13.345 26.415 20.655 27.095 ;
        RECT 6.905 26.185 8.250 26.415 ;
        RECT 9.205 26.185 10.135 26.415 ;
        RECT 16.860 26.195 17.770 26.415 ;
        RECT 19.305 26.185 20.655 26.415 ;
        RECT 20.705 26.415 24.605 27.095 ;
        RECT 24.940 26.415 28.405 27.095 ;
        RECT 20.705 26.185 21.635 26.415 ;
        RECT 24.940 26.185 25.860 26.415 ;
        RECT 28.525 26.285 31.275 27.095 ;
        RECT 31.295 26.225 31.725 27.010 ;
        RECT 32.035 26.185 34.955 27.095 ;
        RECT 36.025 26.185 39.475 27.095 ;
        RECT 40.025 26.285 41.395 27.095 ;
      LAYER nwell ;
        RECT 5.330 23.065 41.590 25.895 ;
      LAYER pwell ;
        RECT 5.525 21.865 6.895 22.675 ;
        RECT 10.420 22.545 11.330 22.765 ;
        RECT 12.865 22.545 14.215 22.775 ;
        RECT 6.905 21.865 14.215 22.545 ;
        RECT 14.265 21.865 17.935 22.675 ;
        RECT 18.415 21.950 18.845 22.735 ;
        RECT 22.380 22.545 23.290 22.765 ;
        RECT 24.825 22.545 26.175 22.775 ;
        RECT 28.070 22.545 29.435 22.775 ;
        RECT 18.865 21.865 26.175 22.545 ;
        RECT 26.225 21.865 29.435 22.545 ;
        RECT 29.445 21.865 32.195 22.675 ;
        RECT 35.320 22.545 36.240 22.775 ;
        RECT 32.775 21.865 36.240 22.545 ;
        RECT 36.425 21.865 39.425 22.775 ;
        RECT 40.025 21.865 41.395 22.675 ;
        RECT 5.665 21.655 5.835 21.865 ;
        RECT 7.045 21.675 7.215 21.865 ;
        RECT 8.425 21.655 8.595 21.845 ;
        RECT 8.895 21.700 9.055 21.810 ;
        RECT 9.805 21.655 9.975 21.845 ;
        RECT 13.495 21.700 13.655 21.810 ;
        RECT 14.405 21.655 14.575 21.865 ;
        RECT 18.080 21.705 18.200 21.815 ;
        RECT 19.005 21.675 19.175 21.865 ;
        RECT 21.490 21.655 21.660 21.845 ;
        RECT 22.225 21.655 22.395 21.845 ;
        RECT 24.065 21.655 24.235 21.845 ;
        RECT 26.370 21.675 26.540 21.865 ;
        RECT 29.585 21.675 29.755 21.865 ;
        RECT 32.160 21.655 32.330 21.845 ;
        RECT 32.340 21.705 32.460 21.815 ;
        RECT 32.805 21.675 32.975 21.865 ;
        RECT 36.025 21.655 36.195 21.845 ;
        RECT 36.485 21.675 36.655 21.865 ;
        RECT 5.525 20.845 6.895 21.655 ;
        RECT 6.905 20.975 8.735 21.655 ;
        RECT 9.775 20.975 13.240 21.655 ;
        RECT 14.375 20.975 17.840 21.655 ;
        RECT 18.175 20.975 22.075 21.655 ;
        RECT 6.905 20.745 8.250 20.975 ;
        RECT 12.320 20.745 13.240 20.975 ;
        RECT 16.920 20.745 17.840 20.975 ;
        RECT 21.145 20.745 22.075 20.975 ;
        RECT 22.085 20.845 23.915 21.655 ;
        RECT 23.925 20.975 31.235 21.655 ;
        RECT 27.440 20.755 28.350 20.975 ;
        RECT 29.885 20.745 31.235 20.975 ;
        RECT 31.295 20.785 31.725 21.570 ;
        RECT 31.745 20.975 35.645 21.655 ;
        RECT 31.745 20.745 32.675 20.975 ;
        RECT 35.885 20.875 37.255 21.655 ;
        RECT 37.265 21.625 38.210 21.655 ;
        RECT 39.700 21.625 39.870 21.845 ;
        RECT 41.085 21.655 41.255 21.865 ;
        RECT 37.265 20.945 40.015 21.625 ;
        RECT 37.265 20.745 38.210 20.945 ;
        RECT 40.025 20.845 41.395 21.655 ;
      LAYER nwell ;
        RECT 5.330 17.625 41.590 20.455 ;
      LAYER pwell ;
        RECT 5.525 16.425 6.895 17.235 ;
        RECT 6.945 17.105 8.295 17.335 ;
        RECT 9.830 17.105 10.740 17.325 ;
        RECT 6.945 16.425 14.255 17.105 ;
        RECT 14.265 16.425 17.935 17.235 ;
        RECT 18.415 16.510 18.845 17.295 ;
        RECT 18.865 16.425 27.970 17.105 ;
        RECT 28.065 16.425 29.435 17.235 ;
        RECT 29.445 16.425 30.815 17.205 ;
        RECT 30.825 16.425 32.195 17.205 ;
        RECT 32.205 16.425 33.575 17.205 ;
        RECT 33.585 16.425 34.955 17.205 ;
        RECT 34.985 16.425 36.335 17.335 ;
        RECT 36.425 16.425 39.875 17.335 ;
        RECT 40.025 16.425 41.395 17.235 ;
        RECT 5.665 16.215 5.835 16.425 ;
        RECT 8.425 16.215 8.595 16.405 ;
        RECT 8.895 16.260 9.055 16.370 ;
        RECT 10.080 16.215 10.250 16.405 ;
        RECT 13.945 16.215 14.115 16.425 ;
        RECT 14.405 16.235 14.575 16.425 ;
        RECT 17.625 16.215 17.795 16.405 ;
        RECT 18.080 16.265 18.200 16.375 ;
        RECT 19.005 16.235 19.175 16.425 ;
        RECT 25.905 16.215 26.075 16.405 ;
        RECT 26.640 16.215 26.810 16.405 ;
        RECT 28.205 16.235 28.375 16.425 ;
        RECT 29.585 16.235 29.755 16.425 ;
        RECT 30.515 16.260 30.675 16.370 ;
        RECT 30.965 16.235 31.135 16.425 ;
        RECT 32.345 16.235 32.515 16.425 ;
        RECT 33.725 16.235 33.895 16.425 ;
        RECT 35.105 16.215 35.275 16.405 ;
        RECT 35.575 16.260 35.735 16.370 ;
        RECT 36.020 16.235 36.190 16.425 ;
        RECT 36.485 16.235 36.655 16.425 ;
        RECT 38.785 16.215 38.955 16.405 ;
        RECT 39.255 16.260 39.415 16.370 ;
        RECT 41.085 16.215 41.255 16.425 ;
        RECT 5.525 15.405 6.895 16.215 ;
        RECT 6.905 15.535 8.735 16.215 ;
        RECT 9.665 15.535 13.565 16.215 ;
        RECT 6.905 15.305 8.250 15.535 ;
        RECT 9.665 15.305 10.595 15.535 ;
        RECT 13.805 15.405 17.475 16.215 ;
        RECT 17.485 15.405 18.855 16.215 ;
        RECT 18.905 15.535 26.215 16.215 ;
        RECT 26.225 15.535 30.125 16.215 ;
        RECT 18.905 15.305 20.255 15.535 ;
        RECT 21.790 15.315 22.700 15.535 ;
        RECT 26.225 15.305 27.155 15.535 ;
        RECT 31.295 15.345 31.725 16.130 ;
        RECT 31.840 15.535 35.305 16.215 ;
        RECT 31.840 15.305 32.760 15.535 ;
        RECT 36.345 15.305 39.095 16.215 ;
        RECT 40.025 15.405 41.395 16.215 ;
      LAYER nwell ;
        RECT 5.330 12.185 41.590 15.015 ;
      LAYER pwell ;
        RECT 5.525 10.985 6.895 11.795 ;
        RECT 6.905 10.985 12.415 11.795 ;
        RECT 12.425 10.985 16.095 11.795 ;
        RECT 17.050 11.665 18.395 11.895 ;
        RECT 16.565 10.985 18.395 11.665 ;
        RECT 18.415 11.070 18.845 11.855 ;
        RECT 19.325 11.665 20.670 11.895 ;
        RECT 24.680 11.665 25.590 11.885 ;
        RECT 27.125 11.665 28.475 11.895 ;
        RECT 19.325 10.985 21.155 11.665 ;
        RECT 21.165 10.985 28.475 11.665 ;
        RECT 28.525 11.665 29.870 11.895 ;
        RECT 28.525 10.985 30.355 11.665 ;
        RECT 31.295 11.070 31.725 11.855 ;
        RECT 33.150 11.665 34.495 11.895 ;
        RECT 32.665 10.985 34.495 11.665 ;
        RECT 34.505 10.985 35.875 11.765 ;
        RECT 38.625 11.665 39.555 11.895 ;
        RECT 36.805 10.985 39.555 11.665 ;
        RECT 40.025 10.985 41.395 11.795 ;
        RECT 5.665 10.795 5.835 10.985 ;
        RECT 7.045 10.795 7.215 10.985 ;
        RECT 12.565 10.795 12.735 10.985 ;
        RECT 16.240 10.825 16.360 10.935 ;
        RECT 16.705 10.795 16.875 10.985 ;
        RECT 19.000 10.825 19.120 10.935 ;
        RECT 20.845 10.795 21.015 10.985 ;
        RECT 21.305 10.795 21.475 10.985 ;
        RECT 30.045 10.795 30.215 10.985 ;
        RECT 30.515 10.830 30.675 10.940 ;
        RECT 31.895 10.830 32.055 10.940 ;
        RECT 32.805 10.795 32.975 10.985 ;
        RECT 35.555 10.795 35.725 10.985 ;
        RECT 36.035 10.830 36.195 10.940 ;
        RECT 36.945 10.795 37.115 10.985 ;
        RECT 39.700 10.825 39.820 10.935 ;
        RECT 41.085 10.795 41.255 10.985 ;
      LAYER li1 ;
        RECT 5.520 46.155 41.400 46.325 ;
        RECT 5.605 45.065 6.815 46.155 ;
        RECT 6.985 45.720 12.330 46.155 ;
        RECT 5.605 44.355 6.125 44.895 ;
        RECT 6.295 44.525 6.815 45.065 ;
        RECT 5.605 43.605 6.815 44.355 ;
        RECT 8.570 44.150 8.910 44.980 ;
        RECT 10.390 44.470 10.740 45.720 ;
        RECT 13.515 45.225 13.685 45.985 ;
        RECT 13.900 45.395 14.230 46.155 ;
        RECT 13.515 45.055 14.230 45.225 ;
        RECT 14.400 45.080 14.655 45.985 ;
        RECT 13.425 44.505 13.780 44.875 ;
        RECT 14.060 44.845 14.230 45.055 ;
        RECT 14.060 44.515 14.315 44.845 ;
        RECT 14.060 44.325 14.230 44.515 ;
        RECT 14.485 44.350 14.655 45.080 ;
        RECT 14.830 45.005 15.090 46.155 ;
        RECT 15.275 45.355 15.605 46.155 ;
        RECT 15.785 45.815 17.215 45.985 ;
        RECT 15.785 45.185 16.035 45.815 ;
        RECT 15.265 45.015 16.035 45.185 ;
        RECT 13.515 44.155 14.230 44.325 ;
        RECT 6.985 43.605 12.330 44.150 ;
        RECT 13.515 43.775 13.685 44.155 ;
        RECT 13.900 43.605 14.230 43.985 ;
        RECT 14.400 43.775 14.655 44.350 ;
        RECT 14.830 43.605 15.090 44.445 ;
        RECT 15.265 44.345 15.435 45.015 ;
        RECT 15.605 44.515 16.010 44.845 ;
        RECT 16.225 44.515 16.475 45.645 ;
        RECT 16.675 44.845 16.875 45.645 ;
        RECT 17.045 45.135 17.215 45.815 ;
        RECT 17.385 45.305 17.700 46.155 ;
        RECT 17.875 45.355 18.315 45.985 ;
        RECT 17.045 44.965 17.835 45.135 ;
        RECT 16.675 44.515 16.920 44.845 ;
        RECT 17.105 44.515 17.495 44.795 ;
        RECT 17.665 44.515 17.835 44.965 ;
        RECT 18.005 44.345 18.315 45.355 ;
        RECT 18.485 44.990 18.775 46.155 ;
        RECT 19.980 45.525 20.265 45.985 ;
        RECT 20.435 45.695 20.705 46.155 ;
        RECT 19.980 45.305 20.935 45.525 ;
        RECT 19.865 44.575 20.555 45.135 ;
        RECT 20.725 44.405 20.935 45.305 ;
        RECT 15.265 43.775 15.755 44.345 ;
        RECT 15.925 44.175 17.085 44.345 ;
        RECT 15.925 43.775 16.155 44.175 ;
        RECT 16.325 43.605 16.745 44.005 ;
        RECT 16.915 43.775 17.085 44.175 ;
        RECT 17.255 43.605 17.705 44.345 ;
        RECT 17.875 43.785 18.315 44.345 ;
        RECT 18.485 43.605 18.775 44.330 ;
        RECT 19.980 44.235 20.935 44.405 ;
        RECT 21.105 45.135 21.505 45.985 ;
        RECT 21.695 45.525 21.975 45.985 ;
        RECT 22.495 45.695 22.820 46.155 ;
        RECT 21.695 45.305 22.820 45.525 ;
        RECT 21.105 44.575 22.200 45.135 ;
        RECT 22.370 44.845 22.820 45.305 ;
        RECT 22.990 45.015 23.375 45.985 ;
        RECT 19.980 43.775 20.265 44.235 ;
        RECT 20.435 43.605 20.705 44.065 ;
        RECT 21.105 43.775 21.505 44.575 ;
        RECT 22.370 44.515 22.925 44.845 ;
        RECT 22.370 44.405 22.820 44.515 ;
        RECT 21.695 44.235 22.820 44.405 ;
        RECT 23.095 44.345 23.375 45.015 ;
        RECT 24.470 45.005 24.730 46.155 ;
        RECT 24.905 45.080 25.160 45.985 ;
        RECT 25.330 45.395 25.660 46.155 ;
        RECT 25.875 45.225 26.045 45.985 ;
        RECT 26.420 45.525 26.705 45.985 ;
        RECT 26.875 45.695 27.145 46.155 ;
        RECT 26.420 45.305 27.375 45.525 ;
        RECT 21.695 43.775 21.975 44.235 ;
        RECT 22.495 43.605 22.820 44.065 ;
        RECT 22.990 43.775 23.375 44.345 ;
        RECT 24.470 43.605 24.730 44.445 ;
        RECT 24.905 44.350 25.075 45.080 ;
        RECT 25.330 45.055 26.045 45.225 ;
        RECT 25.330 44.845 25.500 45.055 ;
        RECT 25.245 44.515 25.500 44.845 ;
        RECT 24.905 43.775 25.160 44.350 ;
        RECT 25.330 44.325 25.500 44.515 ;
        RECT 25.780 44.505 26.135 44.875 ;
        RECT 26.305 44.575 26.995 45.135 ;
        RECT 27.165 44.405 27.375 45.305 ;
        RECT 25.330 44.155 26.045 44.325 ;
        RECT 25.330 43.605 25.660 43.985 ;
        RECT 25.875 43.775 26.045 44.155 ;
        RECT 26.420 44.235 27.375 44.405 ;
        RECT 27.545 45.135 27.945 45.985 ;
        RECT 28.135 45.525 28.415 45.985 ;
        RECT 28.935 45.695 29.260 46.155 ;
        RECT 28.135 45.305 29.260 45.525 ;
        RECT 27.545 44.575 28.640 45.135 ;
        RECT 28.810 44.845 29.260 45.305 ;
        RECT 29.430 45.015 29.815 45.985 ;
        RECT 30.065 45.225 30.245 45.985 ;
        RECT 30.425 45.395 30.755 46.155 ;
        RECT 30.065 45.055 30.740 45.225 ;
        RECT 30.925 45.080 31.195 45.985 ;
        RECT 26.420 43.775 26.705 44.235 ;
        RECT 26.875 43.605 27.145 44.065 ;
        RECT 27.545 43.775 27.945 44.575 ;
        RECT 28.810 44.515 29.365 44.845 ;
        RECT 28.810 44.405 29.260 44.515 ;
        RECT 28.135 44.235 29.260 44.405 ;
        RECT 29.535 44.345 29.815 45.015 ;
        RECT 30.570 44.910 30.740 45.055 ;
        RECT 30.005 44.505 30.345 44.875 ;
        RECT 30.570 44.580 30.845 44.910 ;
        RECT 28.135 43.775 28.415 44.235 ;
        RECT 28.935 43.605 29.260 44.065 ;
        RECT 29.430 43.775 29.815 44.345 ;
        RECT 30.570 44.325 30.740 44.580 ;
        RECT 30.075 44.155 30.740 44.325 ;
        RECT 31.015 44.280 31.195 45.080 ;
        RECT 31.365 44.990 31.655 46.155 ;
        RECT 32.750 45.005 33.010 46.155 ;
        RECT 33.185 45.080 33.440 45.985 ;
        RECT 33.610 45.395 33.940 46.155 ;
        RECT 34.155 45.225 34.325 45.985 ;
        RECT 30.075 43.775 30.245 44.155 ;
        RECT 30.425 43.605 30.755 43.985 ;
        RECT 30.935 43.775 31.195 44.280 ;
        RECT 31.365 43.605 31.655 44.330 ;
        RECT 32.750 43.605 33.010 44.445 ;
        RECT 33.185 44.350 33.355 45.080 ;
        RECT 33.610 45.055 34.325 45.225 ;
        RECT 34.585 45.065 35.795 46.155 ;
        RECT 33.610 44.845 33.780 45.055 ;
        RECT 33.525 44.515 33.780 44.845 ;
        RECT 33.185 43.775 33.440 44.350 ;
        RECT 33.610 44.325 33.780 44.515 ;
        RECT 34.060 44.505 34.415 44.875 ;
        RECT 34.585 44.355 35.105 44.895 ;
        RECT 35.275 44.525 35.795 45.065 ;
        RECT 35.965 45.080 36.235 45.985 ;
        RECT 36.405 45.395 36.735 46.155 ;
        RECT 36.915 45.225 37.085 45.985 ;
        RECT 33.610 44.155 34.325 44.325 ;
        RECT 33.610 43.605 33.940 43.985 ;
        RECT 34.155 43.775 34.325 44.155 ;
        RECT 34.585 43.605 35.795 44.355 ;
        RECT 35.965 44.280 36.135 45.080 ;
        RECT 36.420 45.055 37.085 45.225 ;
        RECT 37.345 45.080 37.615 45.985 ;
        RECT 37.785 45.395 38.115 46.155 ;
        RECT 38.295 45.225 38.465 45.985 ;
        RECT 36.420 44.910 36.590 45.055 ;
        RECT 36.305 44.580 36.590 44.910 ;
        RECT 36.420 44.325 36.590 44.580 ;
        RECT 36.825 44.505 37.155 44.875 ;
        RECT 35.965 43.775 36.225 44.280 ;
        RECT 36.420 44.155 37.085 44.325 ;
        RECT 36.405 43.605 36.735 43.985 ;
        RECT 36.915 43.775 37.085 44.155 ;
        RECT 37.345 44.280 37.515 45.080 ;
        RECT 37.800 45.055 38.465 45.225 ;
        RECT 38.725 45.080 38.995 45.985 ;
        RECT 39.165 45.395 39.495 46.155 ;
        RECT 39.675 45.225 39.855 45.985 ;
        RECT 37.800 44.910 37.970 45.055 ;
        RECT 37.685 44.580 37.970 44.910 ;
        RECT 37.800 44.325 37.970 44.580 ;
        RECT 38.205 44.505 38.535 44.875 ;
        RECT 37.345 43.775 37.605 44.280 ;
        RECT 37.800 44.155 38.465 44.325 ;
        RECT 37.785 43.605 38.115 43.985 ;
        RECT 38.295 43.775 38.465 44.155 ;
        RECT 38.725 44.280 38.905 45.080 ;
        RECT 39.180 45.055 39.855 45.225 ;
        RECT 40.105 45.065 41.315 46.155 ;
        RECT 39.180 44.910 39.350 45.055 ;
        RECT 39.075 44.580 39.350 44.910 ;
        RECT 39.180 44.325 39.350 44.580 ;
        RECT 39.575 44.505 39.915 44.875 ;
        RECT 40.105 44.525 40.625 45.065 ;
        RECT 40.795 44.355 41.315 44.895 ;
        RECT 38.725 43.775 38.985 44.280 ;
        RECT 39.180 44.155 39.845 44.325 ;
        RECT 39.165 43.605 39.495 43.985 ;
        RECT 39.675 43.775 39.845 44.155 ;
        RECT 40.105 43.605 41.315 44.355 ;
        RECT 5.520 43.435 41.400 43.605 ;
        RECT 5.605 42.685 6.815 43.435 ;
        RECT 5.605 42.145 6.125 42.685 ;
        RECT 6.985 42.665 10.495 43.435 ;
        RECT 11.175 42.780 11.505 43.215 ;
        RECT 11.675 42.825 11.845 43.435 ;
        RECT 11.125 42.695 11.505 42.780 ;
        RECT 12.015 42.695 12.345 43.220 ;
        RECT 12.605 42.905 12.815 43.435 ;
        RECT 13.090 42.985 13.875 43.155 ;
        RECT 14.045 42.985 14.450 43.155 ;
        RECT 6.295 41.975 6.815 42.515 ;
        RECT 6.985 42.145 8.635 42.665 ;
        RECT 11.125 42.655 11.350 42.695 ;
        RECT 8.805 41.975 10.495 42.495 ;
        RECT 5.605 40.885 6.815 41.975 ;
        RECT 6.985 40.885 10.495 41.975 ;
        RECT 11.125 42.075 11.295 42.655 ;
        RECT 12.015 42.525 12.215 42.695 ;
        RECT 13.090 42.525 13.260 42.985 ;
        RECT 11.465 42.195 12.215 42.525 ;
        RECT 12.385 42.195 13.260 42.525 ;
        RECT 11.125 42.025 11.340 42.075 ;
        RECT 11.125 41.945 11.515 42.025 ;
        RECT 11.185 41.100 11.515 41.945 ;
        RECT 12.025 41.990 12.215 42.195 ;
        RECT 11.685 40.885 11.855 41.895 ;
        RECT 12.025 41.615 12.920 41.990 ;
        RECT 12.025 41.055 12.365 41.615 ;
        RECT 12.595 40.885 12.910 41.385 ;
        RECT 13.090 41.355 13.260 42.195 ;
        RECT 13.430 42.485 13.895 42.815 ;
        RECT 14.280 42.755 14.450 42.985 ;
        RECT 14.630 42.935 15.000 43.435 ;
        RECT 15.320 42.985 15.995 43.155 ;
        RECT 16.190 42.985 16.525 43.155 ;
        RECT 13.430 41.525 13.750 42.485 ;
        RECT 14.280 42.455 15.110 42.755 ;
        RECT 13.920 41.555 14.110 42.275 ;
        RECT 14.280 41.385 14.450 42.455 ;
        RECT 14.910 42.425 15.110 42.455 ;
        RECT 14.620 42.205 14.790 42.275 ;
        RECT 15.320 42.205 15.490 42.985 ;
        RECT 16.355 42.845 16.525 42.985 ;
        RECT 16.695 42.975 16.945 43.435 ;
        RECT 14.620 42.035 15.490 42.205 ;
        RECT 15.660 42.565 16.185 42.785 ;
        RECT 16.355 42.715 16.580 42.845 ;
        RECT 14.620 41.945 15.130 42.035 ;
        RECT 13.090 41.185 13.975 41.355 ;
        RECT 14.200 41.055 14.450 41.385 ;
        RECT 14.620 40.885 14.790 41.685 ;
        RECT 14.960 41.330 15.130 41.945 ;
        RECT 15.660 41.865 15.830 42.565 ;
        RECT 15.300 41.500 15.830 41.865 ;
        RECT 16.000 41.800 16.240 42.395 ;
        RECT 16.410 41.610 16.580 42.715 ;
        RECT 16.750 41.855 17.030 42.805 ;
        RECT 16.275 41.480 16.580 41.610 ;
        RECT 14.960 41.160 16.065 41.330 ;
        RECT 16.275 41.055 16.525 41.480 ;
        RECT 16.695 40.885 16.960 41.345 ;
        RECT 17.200 41.055 17.385 43.175 ;
        RECT 17.555 43.055 17.885 43.435 ;
        RECT 18.055 42.885 18.225 43.175 ;
        RECT 17.560 42.715 18.225 42.885 ;
        RECT 18.575 42.885 18.745 43.175 ;
        RECT 18.915 43.055 19.245 43.435 ;
        RECT 18.575 42.715 19.240 42.885 ;
        RECT 17.560 41.725 17.790 42.715 ;
        RECT 17.960 41.895 18.310 42.545 ;
        RECT 18.490 41.895 18.840 42.545 ;
        RECT 19.010 41.725 19.240 42.715 ;
        RECT 17.560 41.555 18.225 41.725 ;
        RECT 17.555 40.885 17.885 41.385 ;
        RECT 18.055 41.055 18.225 41.555 ;
        RECT 18.575 41.555 19.240 41.725 ;
        RECT 18.575 41.055 18.745 41.555 ;
        RECT 18.915 40.885 19.245 41.385 ;
        RECT 19.415 41.055 19.600 43.175 ;
        RECT 19.855 42.975 20.105 43.435 ;
        RECT 20.275 42.985 20.610 43.155 ;
        RECT 20.805 42.985 21.480 43.155 ;
        RECT 20.275 42.845 20.445 42.985 ;
        RECT 19.770 41.855 20.050 42.805 ;
        RECT 20.220 42.715 20.445 42.845 ;
        RECT 20.220 41.610 20.390 42.715 ;
        RECT 20.615 42.565 21.140 42.785 ;
        RECT 20.560 41.800 20.800 42.395 ;
        RECT 20.970 41.865 21.140 42.565 ;
        RECT 21.310 42.205 21.480 42.985 ;
        RECT 21.800 42.935 22.170 43.435 ;
        RECT 22.350 42.985 22.755 43.155 ;
        RECT 22.925 42.985 23.710 43.155 ;
        RECT 22.350 42.755 22.520 42.985 ;
        RECT 21.690 42.455 22.520 42.755 ;
        RECT 22.905 42.485 23.370 42.815 ;
        RECT 21.690 42.425 21.890 42.455 ;
        RECT 22.010 42.205 22.180 42.275 ;
        RECT 21.310 42.035 22.180 42.205 ;
        RECT 21.670 41.945 22.180 42.035 ;
        RECT 20.220 41.480 20.525 41.610 ;
        RECT 20.970 41.500 21.500 41.865 ;
        RECT 19.840 40.885 20.105 41.345 ;
        RECT 20.275 41.055 20.525 41.480 ;
        RECT 21.670 41.330 21.840 41.945 ;
        RECT 20.735 41.160 21.840 41.330 ;
        RECT 22.010 40.885 22.180 41.685 ;
        RECT 22.350 41.385 22.520 42.455 ;
        RECT 22.690 41.555 22.880 42.275 ;
        RECT 23.050 41.525 23.370 42.485 ;
        RECT 23.540 42.525 23.710 42.985 ;
        RECT 23.985 42.905 24.195 43.435 ;
        RECT 24.455 42.695 24.785 43.220 ;
        RECT 24.955 42.825 25.125 43.435 ;
        RECT 25.295 42.780 25.625 43.215 ;
        RECT 25.295 42.695 25.675 42.780 ;
        RECT 24.585 42.525 24.785 42.695 ;
        RECT 25.450 42.655 25.675 42.695 ;
        RECT 23.540 42.195 24.415 42.525 ;
        RECT 24.585 42.195 25.335 42.525 ;
        RECT 22.350 41.055 22.600 41.385 ;
        RECT 23.540 41.355 23.710 42.195 ;
        RECT 24.585 41.990 24.775 42.195 ;
        RECT 25.505 42.075 25.675 42.655 ;
        RECT 25.460 42.025 25.675 42.075 ;
        RECT 23.880 41.615 24.775 41.990 ;
        RECT 25.285 41.945 25.675 42.025 ;
        RECT 25.880 42.695 26.495 43.265 ;
        RECT 26.665 42.925 26.880 43.435 ;
        RECT 27.110 42.925 27.390 43.255 ;
        RECT 27.570 42.925 27.810 43.435 ;
        RECT 22.825 41.185 23.710 41.355 ;
        RECT 23.890 40.885 24.205 41.385 ;
        RECT 24.435 41.055 24.775 41.615 ;
        RECT 24.945 40.885 25.115 41.895 ;
        RECT 25.285 41.100 25.615 41.945 ;
        RECT 25.880 41.675 26.195 42.695 ;
        RECT 26.365 42.025 26.535 42.525 ;
        RECT 26.785 42.195 27.050 42.755 ;
        RECT 27.220 42.025 27.390 42.925 ;
        RECT 28.235 42.885 28.405 43.265 ;
        RECT 28.620 43.055 28.950 43.435 ;
        RECT 27.560 42.195 27.915 42.755 ;
        RECT 28.235 42.715 28.950 42.885 ;
        RECT 28.145 42.165 28.500 42.535 ;
        RECT 28.780 42.525 28.950 42.715 ;
        RECT 29.120 42.690 29.375 43.265 ;
        RECT 28.780 42.195 29.035 42.525 ;
        RECT 26.365 41.855 27.790 42.025 ;
        RECT 28.780 41.985 28.950 42.195 ;
        RECT 25.880 41.055 26.415 41.675 ;
        RECT 26.585 40.885 26.915 41.685 ;
        RECT 27.400 41.680 27.790 41.855 ;
        RECT 28.235 41.815 28.950 41.985 ;
        RECT 29.205 41.960 29.375 42.690 ;
        RECT 29.550 42.595 29.810 43.435 ;
        RECT 30.025 42.615 30.255 43.435 ;
        RECT 30.425 42.635 30.755 43.265 ;
        RECT 30.005 42.195 30.335 42.445 ;
        RECT 30.505 42.035 30.755 42.635 ;
        RECT 30.925 42.615 31.135 43.435 ;
        RECT 31.365 42.710 31.655 43.435 ;
        RECT 31.825 42.695 32.265 43.255 ;
        RECT 32.435 42.695 32.885 43.435 ;
        RECT 33.055 42.865 33.225 43.265 ;
        RECT 33.395 43.035 33.815 43.435 ;
        RECT 33.985 42.865 34.215 43.265 ;
        RECT 33.055 42.695 34.215 42.865 ;
        RECT 34.385 42.695 34.875 43.265 ;
        RECT 28.235 41.055 28.405 41.815 ;
        RECT 28.620 40.885 28.950 41.645 ;
        RECT 29.120 41.055 29.375 41.960 ;
        RECT 29.550 40.885 29.810 42.035 ;
        RECT 30.025 40.885 30.255 42.025 ;
        RECT 30.425 41.055 30.755 42.035 ;
        RECT 30.925 40.885 31.135 42.025 ;
        RECT 31.365 40.885 31.655 42.050 ;
        RECT 31.825 41.685 32.135 42.695 ;
        RECT 32.305 42.075 32.475 42.525 ;
        RECT 32.645 42.245 33.035 42.525 ;
        RECT 33.220 42.195 33.465 42.525 ;
        RECT 32.305 41.905 33.095 42.075 ;
        RECT 31.825 41.055 32.265 41.685 ;
        RECT 32.440 40.885 32.755 41.735 ;
        RECT 32.925 41.225 33.095 41.905 ;
        RECT 33.265 41.395 33.465 42.195 ;
        RECT 33.665 41.395 33.915 42.525 ;
        RECT 34.130 42.195 34.535 42.525 ;
        RECT 34.705 42.025 34.875 42.695 ;
        RECT 35.160 42.805 35.445 43.265 ;
        RECT 35.615 42.975 35.885 43.435 ;
        RECT 35.160 42.635 36.115 42.805 ;
        RECT 34.105 41.855 34.875 42.025 ;
        RECT 35.045 41.905 35.735 42.465 ;
        RECT 34.105 41.225 34.355 41.855 ;
        RECT 35.905 41.735 36.115 42.635 ;
        RECT 32.925 41.055 34.355 41.225 ;
        RECT 34.535 40.885 34.865 41.685 ;
        RECT 35.160 41.515 36.115 41.735 ;
        RECT 36.285 42.465 36.685 43.265 ;
        RECT 36.875 42.805 37.155 43.265 ;
        RECT 37.675 42.975 38.000 43.435 ;
        RECT 36.875 42.635 38.000 42.805 ;
        RECT 38.170 42.695 38.555 43.265 ;
        RECT 37.550 42.525 38.000 42.635 ;
        RECT 36.285 41.905 37.380 42.465 ;
        RECT 37.550 42.195 38.105 42.525 ;
        RECT 35.160 41.055 35.445 41.515 ;
        RECT 35.615 40.885 35.885 41.345 ;
        RECT 36.285 41.055 36.685 41.905 ;
        RECT 37.550 41.735 38.000 42.195 ;
        RECT 38.275 42.025 38.555 42.695 ;
        RECT 36.875 41.515 38.000 41.735 ;
        RECT 36.875 41.055 37.155 41.515 ;
        RECT 37.675 40.885 38.000 41.345 ;
        RECT 38.170 41.055 38.555 42.025 ;
        RECT 38.725 42.760 38.985 43.265 ;
        RECT 39.165 43.055 39.495 43.435 ;
        RECT 39.675 42.885 39.845 43.265 ;
        RECT 38.725 41.960 38.905 42.760 ;
        RECT 39.180 42.715 39.845 42.885 ;
        RECT 39.180 42.460 39.350 42.715 ;
        RECT 40.105 42.685 41.315 43.435 ;
        RECT 39.075 42.130 39.350 42.460 ;
        RECT 39.575 42.165 39.915 42.535 ;
        RECT 39.180 41.985 39.350 42.130 ;
        RECT 38.725 41.055 38.995 41.960 ;
        RECT 39.180 41.815 39.855 41.985 ;
        RECT 39.165 40.885 39.495 41.645 ;
        RECT 39.675 41.055 39.855 41.815 ;
        RECT 40.105 41.975 40.625 42.515 ;
        RECT 40.795 42.145 41.315 42.685 ;
        RECT 40.105 40.885 41.315 41.975 ;
        RECT 5.520 40.715 41.400 40.885 ;
        RECT 5.605 39.625 6.815 40.715 ;
        RECT 7.075 40.045 7.245 40.545 ;
        RECT 7.415 40.215 7.745 40.715 ;
        RECT 7.075 39.875 7.740 40.045 ;
        RECT 5.605 38.915 6.125 39.455 ;
        RECT 6.295 39.085 6.815 39.625 ;
        RECT 6.990 39.055 7.340 39.705 ;
        RECT 5.605 38.165 6.815 38.915 ;
        RECT 7.510 38.885 7.740 39.875 ;
        RECT 7.075 38.715 7.740 38.885 ;
        RECT 7.075 38.425 7.245 38.715 ;
        RECT 7.415 38.165 7.745 38.545 ;
        RECT 7.915 38.425 8.100 40.545 ;
        RECT 8.340 40.255 8.605 40.715 ;
        RECT 8.775 40.120 9.025 40.545 ;
        RECT 9.235 40.270 10.340 40.440 ;
        RECT 8.720 39.990 9.025 40.120 ;
        RECT 8.270 38.795 8.550 39.745 ;
        RECT 8.720 38.885 8.890 39.990 ;
        RECT 9.060 39.205 9.300 39.800 ;
        RECT 9.470 39.735 10.000 40.100 ;
        RECT 9.470 39.035 9.640 39.735 ;
        RECT 10.170 39.655 10.340 40.270 ;
        RECT 10.510 39.915 10.680 40.715 ;
        RECT 10.850 40.215 11.100 40.545 ;
        RECT 11.325 40.245 12.210 40.415 ;
        RECT 10.170 39.565 10.680 39.655 ;
        RECT 8.720 38.755 8.945 38.885 ;
        RECT 9.115 38.815 9.640 39.035 ;
        RECT 9.810 39.395 10.680 39.565 ;
        RECT 8.355 38.165 8.605 38.625 ;
        RECT 8.775 38.615 8.945 38.755 ;
        RECT 9.810 38.615 9.980 39.395 ;
        RECT 10.510 39.325 10.680 39.395 ;
        RECT 10.190 39.145 10.390 39.175 ;
        RECT 10.850 39.145 11.020 40.215 ;
        RECT 11.190 39.325 11.380 40.045 ;
        RECT 10.190 38.845 11.020 39.145 ;
        RECT 11.550 39.115 11.870 40.075 ;
        RECT 8.775 38.445 9.110 38.615 ;
        RECT 9.305 38.445 9.980 38.615 ;
        RECT 10.300 38.165 10.670 38.665 ;
        RECT 10.850 38.615 11.020 38.845 ;
        RECT 11.405 38.785 11.870 39.115 ;
        RECT 12.040 39.405 12.210 40.245 ;
        RECT 12.390 40.215 12.705 40.715 ;
        RECT 12.935 39.985 13.275 40.545 ;
        RECT 12.380 39.610 13.275 39.985 ;
        RECT 13.445 39.705 13.615 40.715 ;
        RECT 13.085 39.405 13.275 39.610 ;
        RECT 13.785 39.655 14.115 40.500 ;
        RECT 13.785 39.575 14.175 39.655 ;
        RECT 13.960 39.525 14.175 39.575 ;
        RECT 12.040 39.075 12.915 39.405 ;
        RECT 13.085 39.075 13.835 39.405 ;
        RECT 12.040 38.615 12.210 39.075 ;
        RECT 13.085 38.905 13.285 39.075 ;
        RECT 14.005 38.945 14.175 39.525 ;
        RECT 13.950 38.905 14.175 38.945 ;
        RECT 10.850 38.445 11.255 38.615 ;
        RECT 11.425 38.445 12.210 38.615 ;
        RECT 12.485 38.165 12.695 38.695 ;
        RECT 12.955 38.380 13.285 38.905 ;
        RECT 13.795 38.820 14.175 38.905 ;
        RECT 14.345 39.575 14.730 40.545 ;
        RECT 14.900 40.255 15.225 40.715 ;
        RECT 15.745 40.085 16.025 40.545 ;
        RECT 14.900 39.865 16.025 40.085 ;
        RECT 14.345 38.905 14.625 39.575 ;
        RECT 14.900 39.405 15.350 39.865 ;
        RECT 16.215 39.695 16.615 40.545 ;
        RECT 17.015 40.255 17.285 40.715 ;
        RECT 17.455 40.085 17.740 40.545 ;
        RECT 14.795 39.075 15.350 39.405 ;
        RECT 15.520 39.135 16.615 39.695 ;
        RECT 14.900 38.965 15.350 39.075 ;
        RECT 13.455 38.165 13.625 38.775 ;
        RECT 13.795 38.385 14.125 38.820 ;
        RECT 14.345 38.335 14.730 38.905 ;
        RECT 14.900 38.795 16.025 38.965 ;
        RECT 14.900 38.165 15.225 38.625 ;
        RECT 15.745 38.335 16.025 38.795 ;
        RECT 16.215 38.335 16.615 39.135 ;
        RECT 16.785 39.865 17.740 40.085 ;
        RECT 16.785 38.965 16.995 39.865 ;
        RECT 17.165 39.135 17.855 39.695 ;
        RECT 18.485 39.550 18.775 40.715 ;
        RECT 18.950 39.575 19.285 40.545 ;
        RECT 19.455 39.575 19.625 40.715 ;
        RECT 19.795 40.375 21.825 40.545 ;
        RECT 16.785 38.795 17.740 38.965 ;
        RECT 18.950 38.905 19.120 39.575 ;
        RECT 19.795 39.405 19.965 40.375 ;
        RECT 19.290 39.075 19.545 39.405 ;
        RECT 19.770 39.075 19.965 39.405 ;
        RECT 20.135 40.035 21.260 40.205 ;
        RECT 19.375 38.905 19.545 39.075 ;
        RECT 20.135 38.905 20.305 40.035 ;
        RECT 17.015 38.165 17.285 38.625 ;
        RECT 17.455 38.335 17.740 38.795 ;
        RECT 18.485 38.165 18.775 38.890 ;
        RECT 18.950 38.335 19.205 38.905 ;
        RECT 19.375 38.735 20.305 38.905 ;
        RECT 20.475 39.695 21.485 39.865 ;
        RECT 20.475 38.895 20.645 39.695 ;
        RECT 20.850 39.355 21.125 39.495 ;
        RECT 20.845 39.185 21.125 39.355 ;
        RECT 20.130 38.700 20.305 38.735 ;
        RECT 19.375 38.165 19.705 38.565 ;
        RECT 20.130 38.335 20.660 38.700 ;
        RECT 20.850 38.335 21.125 39.185 ;
        RECT 21.295 38.335 21.485 39.695 ;
        RECT 21.655 39.710 21.825 40.375 ;
        RECT 21.995 39.955 22.165 40.715 ;
        RECT 22.400 39.955 22.915 40.365 ;
        RECT 21.655 39.520 22.405 39.710 ;
        RECT 22.575 39.145 22.915 39.955 ;
        RECT 23.730 39.745 24.120 39.920 ;
        RECT 24.605 39.915 24.935 40.715 ;
        RECT 25.105 39.925 25.640 40.545 ;
        RECT 23.730 39.575 25.155 39.745 ;
        RECT 21.685 38.975 22.915 39.145 ;
        RECT 21.665 38.165 22.175 38.700 ;
        RECT 22.395 38.370 22.640 38.975 ;
        RECT 23.605 38.845 23.960 39.405 ;
        RECT 24.130 38.675 24.300 39.575 ;
        RECT 24.470 38.845 24.735 39.405 ;
        RECT 24.985 39.075 25.155 39.575 ;
        RECT 25.325 38.905 25.640 39.925 ;
        RECT 25.905 39.575 26.115 40.715 ;
        RECT 26.285 39.565 26.615 40.545 ;
        RECT 26.785 39.575 27.015 40.715 ;
        RECT 27.315 40.045 27.485 40.545 ;
        RECT 27.655 40.215 27.985 40.715 ;
        RECT 27.315 39.875 27.980 40.045 ;
        RECT 23.710 38.165 23.950 38.675 ;
        RECT 24.130 38.345 24.410 38.675 ;
        RECT 24.640 38.165 24.855 38.675 ;
        RECT 25.025 38.335 25.640 38.905 ;
        RECT 25.905 38.165 26.115 38.985 ;
        RECT 26.285 38.965 26.535 39.565 ;
        RECT 26.705 39.155 27.035 39.405 ;
        RECT 27.230 39.055 27.580 39.705 ;
        RECT 26.285 38.335 26.615 38.965 ;
        RECT 26.785 38.165 27.015 38.985 ;
        RECT 27.750 38.885 27.980 39.875 ;
        RECT 27.315 38.715 27.980 38.885 ;
        RECT 27.315 38.425 27.485 38.715 ;
        RECT 27.655 38.165 27.985 38.545 ;
        RECT 28.155 38.425 28.340 40.545 ;
        RECT 28.580 40.255 28.845 40.715 ;
        RECT 29.015 40.120 29.265 40.545 ;
        RECT 29.475 40.270 30.580 40.440 ;
        RECT 28.960 39.990 29.265 40.120 ;
        RECT 28.510 38.795 28.790 39.745 ;
        RECT 28.960 38.885 29.130 39.990 ;
        RECT 29.300 39.205 29.540 39.800 ;
        RECT 29.710 39.735 30.240 40.100 ;
        RECT 29.710 39.035 29.880 39.735 ;
        RECT 30.410 39.655 30.580 40.270 ;
        RECT 30.750 39.915 30.920 40.715 ;
        RECT 31.090 40.215 31.340 40.545 ;
        RECT 31.565 40.245 32.450 40.415 ;
        RECT 30.410 39.565 30.920 39.655 ;
        RECT 28.960 38.755 29.185 38.885 ;
        RECT 29.355 38.815 29.880 39.035 ;
        RECT 30.050 39.395 30.920 39.565 ;
        RECT 28.595 38.165 28.845 38.625 ;
        RECT 29.015 38.615 29.185 38.755 ;
        RECT 30.050 38.615 30.220 39.395 ;
        RECT 30.750 39.325 30.920 39.395 ;
        RECT 30.430 39.145 30.630 39.175 ;
        RECT 31.090 39.145 31.260 40.215 ;
        RECT 31.430 39.325 31.620 40.045 ;
        RECT 30.430 38.845 31.260 39.145 ;
        RECT 31.790 39.115 32.110 40.075 ;
        RECT 29.015 38.445 29.350 38.615 ;
        RECT 29.545 38.445 30.220 38.615 ;
        RECT 30.540 38.165 30.910 38.665 ;
        RECT 31.090 38.615 31.260 38.845 ;
        RECT 31.645 38.785 32.110 39.115 ;
        RECT 32.280 39.405 32.450 40.245 ;
        RECT 32.630 40.215 32.945 40.715 ;
        RECT 33.175 39.985 33.515 40.545 ;
        RECT 32.620 39.610 33.515 39.985 ;
        RECT 33.685 39.705 33.855 40.715 ;
        RECT 33.325 39.405 33.515 39.610 ;
        RECT 34.025 39.655 34.355 40.500 ;
        RECT 35.230 39.745 35.620 39.920 ;
        RECT 36.105 39.915 36.435 40.715 ;
        RECT 36.605 39.925 37.140 40.545 ;
        RECT 34.025 39.575 34.415 39.655 ;
        RECT 35.230 39.575 36.655 39.745 ;
        RECT 34.200 39.525 34.415 39.575 ;
        RECT 32.280 39.075 33.155 39.405 ;
        RECT 33.325 39.075 34.075 39.405 ;
        RECT 32.280 38.615 32.450 39.075 ;
        RECT 33.325 38.905 33.525 39.075 ;
        RECT 34.245 38.945 34.415 39.525 ;
        RECT 34.190 38.905 34.415 38.945 ;
        RECT 31.090 38.445 31.495 38.615 ;
        RECT 31.665 38.445 32.450 38.615 ;
        RECT 32.725 38.165 32.935 38.695 ;
        RECT 33.195 38.380 33.525 38.905 ;
        RECT 34.035 38.820 34.415 38.905 ;
        RECT 35.105 38.845 35.460 39.405 ;
        RECT 33.695 38.165 33.865 38.775 ;
        RECT 34.035 38.385 34.365 38.820 ;
        RECT 35.630 38.675 35.800 39.575 ;
        RECT 35.970 38.845 36.235 39.405 ;
        RECT 36.485 39.075 36.655 39.575 ;
        RECT 36.825 38.905 37.140 39.925 ;
        RECT 37.435 39.785 37.605 40.545 ;
        RECT 37.785 39.955 38.115 40.715 ;
        RECT 37.435 39.615 38.100 39.785 ;
        RECT 38.285 39.640 38.555 40.545 ;
        RECT 37.930 39.470 38.100 39.615 ;
        RECT 37.365 39.065 37.695 39.435 ;
        RECT 37.930 39.140 38.215 39.470 ;
        RECT 35.210 38.165 35.450 38.675 ;
        RECT 35.630 38.345 35.910 38.675 ;
        RECT 36.140 38.165 36.355 38.675 ;
        RECT 36.525 38.335 37.140 38.905 ;
        RECT 37.930 38.885 38.100 39.140 ;
        RECT 37.435 38.715 38.100 38.885 ;
        RECT 38.385 38.840 38.555 39.640 ;
        RECT 37.435 38.335 37.605 38.715 ;
        RECT 37.785 38.165 38.115 38.545 ;
        RECT 38.295 38.335 38.555 38.840 ;
        RECT 38.725 39.640 38.995 40.545 ;
        RECT 39.165 39.955 39.495 40.715 ;
        RECT 39.675 39.785 39.855 40.545 ;
        RECT 38.725 38.840 38.905 39.640 ;
        RECT 39.180 39.615 39.855 39.785 ;
        RECT 40.105 39.625 41.315 40.715 ;
        RECT 39.180 39.470 39.350 39.615 ;
        RECT 39.075 39.140 39.350 39.470 ;
        RECT 39.180 38.885 39.350 39.140 ;
        RECT 39.575 39.065 39.915 39.435 ;
        RECT 40.105 39.085 40.625 39.625 ;
        RECT 40.795 38.915 41.315 39.455 ;
        RECT 38.725 38.335 38.985 38.840 ;
        RECT 39.180 38.715 39.845 38.885 ;
        RECT 39.165 38.165 39.495 38.545 ;
        RECT 39.675 38.335 39.845 38.715 ;
        RECT 40.105 38.165 41.315 38.915 ;
        RECT 5.520 37.995 41.400 38.165 ;
        RECT 5.605 37.245 6.815 37.995 ;
        RECT 5.605 36.705 6.125 37.245 ;
        RECT 6.990 37.155 7.250 37.995 ;
        RECT 7.425 37.250 7.680 37.825 ;
        RECT 7.850 37.615 8.180 37.995 ;
        RECT 8.395 37.445 8.565 37.825 ;
        RECT 7.850 37.275 8.565 37.445 ;
        RECT 6.295 36.535 6.815 37.075 ;
        RECT 5.605 35.445 6.815 36.535 ;
        RECT 6.990 35.445 7.250 36.595 ;
        RECT 7.425 36.520 7.595 37.250 ;
        RECT 7.850 37.085 8.020 37.275 ;
        RECT 8.830 37.255 9.085 37.825 ;
        RECT 9.255 37.595 9.585 37.995 ;
        RECT 10.010 37.460 10.540 37.825 ;
        RECT 10.730 37.655 11.005 37.825 ;
        RECT 10.725 37.485 11.005 37.655 ;
        RECT 10.010 37.425 10.185 37.460 ;
        RECT 9.255 37.255 10.185 37.425 ;
        RECT 7.765 36.755 8.020 37.085 ;
        RECT 7.850 36.545 8.020 36.755 ;
        RECT 8.300 36.725 8.655 37.095 ;
        RECT 8.830 36.585 9.000 37.255 ;
        RECT 9.255 37.085 9.425 37.255 ;
        RECT 9.170 36.755 9.425 37.085 ;
        RECT 9.650 36.755 9.845 37.085 ;
        RECT 7.425 35.615 7.680 36.520 ;
        RECT 7.850 36.375 8.565 36.545 ;
        RECT 7.850 35.445 8.180 36.205 ;
        RECT 8.395 35.615 8.565 36.375 ;
        RECT 8.830 35.615 9.165 36.585 ;
        RECT 9.335 35.445 9.505 36.585 ;
        RECT 9.675 35.785 9.845 36.755 ;
        RECT 10.015 36.125 10.185 37.255 ;
        RECT 10.355 36.465 10.525 37.265 ;
        RECT 10.730 36.665 11.005 37.485 ;
        RECT 11.175 36.465 11.365 37.825 ;
        RECT 11.545 37.460 12.055 37.995 ;
        RECT 12.275 37.185 12.520 37.790 ;
        RECT 12.965 37.245 14.175 37.995 ;
        RECT 14.435 37.515 14.735 37.995 ;
        RECT 14.905 37.345 15.165 37.800 ;
        RECT 15.335 37.515 15.595 37.995 ;
        RECT 15.775 37.345 16.035 37.800 ;
        RECT 16.205 37.515 16.455 37.995 ;
        RECT 16.635 37.345 16.895 37.800 ;
        RECT 17.065 37.515 17.315 37.995 ;
        RECT 17.495 37.345 17.755 37.800 ;
        RECT 17.925 37.515 18.170 37.995 ;
        RECT 18.340 37.345 18.615 37.800 ;
        RECT 18.785 37.515 19.030 37.995 ;
        RECT 19.200 37.345 19.460 37.800 ;
        RECT 19.630 37.515 19.890 37.995 ;
        RECT 20.060 37.345 20.320 37.800 ;
        RECT 20.490 37.515 20.750 37.995 ;
        RECT 20.920 37.345 21.180 37.800 ;
        RECT 21.350 37.435 21.610 37.995 ;
        RECT 11.565 37.015 12.795 37.185 ;
        RECT 10.355 36.295 11.365 36.465 ;
        RECT 11.535 36.450 12.285 36.640 ;
        RECT 10.015 35.955 11.140 36.125 ;
        RECT 11.535 35.785 11.705 36.450 ;
        RECT 12.455 36.205 12.795 37.015 ;
        RECT 12.965 36.705 13.485 37.245 ;
        RECT 14.435 37.175 21.180 37.345 ;
        RECT 13.655 36.535 14.175 37.075 ;
        RECT 9.675 35.615 11.705 35.785 ;
        RECT 11.875 35.445 12.045 36.205 ;
        RECT 12.280 35.795 12.795 36.205 ;
        RECT 12.965 35.445 14.175 36.535 ;
        RECT 14.435 36.585 15.600 37.175 ;
        RECT 21.780 37.005 22.030 37.815 ;
        RECT 22.210 37.470 22.470 37.995 ;
        RECT 22.640 37.005 22.890 37.815 ;
        RECT 23.070 37.485 23.375 37.995 ;
        RECT 15.770 36.755 22.890 37.005 ;
        RECT 23.060 36.755 23.375 37.315 ;
        RECT 23.545 37.255 23.930 37.825 ;
        RECT 24.100 37.535 24.425 37.995 ;
        RECT 24.945 37.365 25.225 37.825 ;
        RECT 14.435 36.360 21.180 36.585 ;
        RECT 14.435 35.445 14.705 36.190 ;
        RECT 14.875 35.620 15.165 36.360 ;
        RECT 15.775 36.345 21.180 36.360 ;
        RECT 15.335 35.450 15.590 36.175 ;
        RECT 15.775 35.620 16.035 36.345 ;
        RECT 16.205 35.450 16.450 36.175 ;
        RECT 16.635 35.620 16.895 36.345 ;
        RECT 17.065 35.450 17.310 36.175 ;
        RECT 17.495 35.620 17.755 36.345 ;
        RECT 17.925 35.450 18.170 36.175 ;
        RECT 18.340 35.620 18.600 36.345 ;
        RECT 18.770 35.450 19.030 36.175 ;
        RECT 19.200 35.620 19.460 36.345 ;
        RECT 19.630 35.450 19.890 36.175 ;
        RECT 20.060 35.620 20.320 36.345 ;
        RECT 20.490 35.450 20.750 36.175 ;
        RECT 20.920 35.620 21.180 36.345 ;
        RECT 21.350 35.450 21.610 36.245 ;
        RECT 21.780 35.620 22.030 36.755 ;
        RECT 15.335 35.445 21.610 35.450 ;
        RECT 22.210 35.445 22.470 36.255 ;
        RECT 22.645 35.615 22.890 36.755 ;
        RECT 23.545 36.585 23.825 37.255 ;
        RECT 24.100 37.195 25.225 37.365 ;
        RECT 24.100 37.085 24.550 37.195 ;
        RECT 23.995 36.755 24.550 37.085 ;
        RECT 25.415 37.025 25.815 37.825 ;
        RECT 26.215 37.535 26.485 37.995 ;
        RECT 26.655 37.365 26.940 37.825 ;
        RECT 23.070 35.445 23.365 36.255 ;
        RECT 23.545 35.615 23.930 36.585 ;
        RECT 24.100 36.295 24.550 36.755 ;
        RECT 24.720 36.465 25.815 37.025 ;
        RECT 24.100 36.075 25.225 36.295 ;
        RECT 24.100 35.445 24.425 35.905 ;
        RECT 24.945 35.615 25.225 36.075 ;
        RECT 25.415 35.615 25.815 36.465 ;
        RECT 25.985 37.195 26.940 37.365 ;
        RECT 27.225 37.245 28.435 37.995 ;
        RECT 28.615 37.495 28.945 37.995 ;
        RECT 29.145 37.425 29.315 37.775 ;
        RECT 29.515 37.595 29.845 37.995 ;
        RECT 30.015 37.425 30.185 37.775 ;
        RECT 30.355 37.595 30.735 37.995 ;
        RECT 25.985 36.295 26.195 37.195 ;
        RECT 26.365 36.465 27.055 37.025 ;
        RECT 27.225 36.705 27.745 37.245 ;
        RECT 27.915 36.535 28.435 37.075 ;
        RECT 28.610 36.755 28.960 37.325 ;
        RECT 29.145 37.255 30.755 37.425 ;
        RECT 30.925 37.320 31.195 37.665 ;
        RECT 30.585 37.085 30.755 37.255 ;
        RECT 25.985 36.075 26.940 36.295 ;
        RECT 26.215 35.445 26.485 35.905 ;
        RECT 26.655 35.615 26.940 36.075 ;
        RECT 27.225 35.445 28.435 36.535 ;
        RECT 28.610 36.295 28.930 36.585 ;
        RECT 29.130 36.465 29.840 37.085 ;
        RECT 30.010 36.755 30.415 37.085 ;
        RECT 30.585 36.755 30.855 37.085 ;
        RECT 30.585 36.585 30.755 36.755 ;
        RECT 31.025 36.585 31.195 37.320 ;
        RECT 31.365 37.270 31.655 37.995 ;
        RECT 31.825 37.255 32.185 37.630 ;
        RECT 32.450 37.255 32.620 37.995 ;
        RECT 32.900 37.425 33.070 37.630 ;
        RECT 32.900 37.255 33.440 37.425 ;
        RECT 30.030 36.415 30.755 36.585 ;
        RECT 30.030 36.295 30.200 36.415 ;
        RECT 28.610 36.125 30.200 36.295 ;
        RECT 28.610 35.665 30.265 35.955 ;
        RECT 30.435 35.445 30.715 36.245 ;
        RECT 30.925 35.615 31.195 36.585 ;
        RECT 31.365 35.445 31.655 36.610 ;
        RECT 31.825 36.600 32.080 37.255 ;
        RECT 32.250 36.755 32.600 37.085 ;
        RECT 32.770 36.755 33.100 37.085 ;
        RECT 31.825 35.615 32.165 36.600 ;
        RECT 32.335 36.215 32.600 36.755 ;
        RECT 33.270 36.555 33.440 37.255 ;
        RECT 32.815 36.385 33.440 36.555 ;
        RECT 33.610 36.625 33.780 37.825 ;
        RECT 34.010 37.345 34.340 37.825 ;
        RECT 34.510 37.525 34.680 37.995 ;
        RECT 34.850 37.345 35.180 37.810 ;
        RECT 34.010 37.175 35.180 37.345 ;
        RECT 35.505 37.255 35.865 37.630 ;
        RECT 36.130 37.255 36.300 37.995 ;
        RECT 36.580 37.425 36.750 37.630 ;
        RECT 36.580 37.255 37.120 37.425 ;
        RECT 33.950 36.795 34.520 37.005 ;
        RECT 34.690 36.795 35.335 37.005 ;
        RECT 33.610 36.215 34.315 36.625 ;
        RECT 35.505 36.600 35.760 37.255 ;
        RECT 35.930 36.755 36.280 37.085 ;
        RECT 36.450 36.755 36.780 37.085 ;
        RECT 32.335 36.045 34.315 36.215 ;
        RECT 32.335 35.445 32.745 35.875 ;
        RECT 33.490 35.445 33.820 35.865 ;
        RECT 33.990 35.615 34.315 36.045 ;
        RECT 34.790 35.445 35.120 36.545 ;
        RECT 35.505 35.615 35.845 36.600 ;
        RECT 36.015 36.215 36.280 36.755 ;
        RECT 36.950 36.555 37.120 37.255 ;
        RECT 36.495 36.385 37.120 36.555 ;
        RECT 37.290 36.625 37.460 37.825 ;
        RECT 37.690 37.345 38.020 37.825 ;
        RECT 38.190 37.525 38.360 37.995 ;
        RECT 38.530 37.345 38.860 37.810 ;
        RECT 37.690 37.175 38.860 37.345 ;
        RECT 40.105 37.245 41.315 37.995 ;
        RECT 37.630 36.795 38.200 37.005 ;
        RECT 38.370 36.795 39.015 37.005 ;
        RECT 37.290 36.215 37.995 36.625 ;
        RECT 36.015 36.045 37.995 36.215 ;
        RECT 36.015 35.445 36.425 35.875 ;
        RECT 37.170 35.445 37.500 35.865 ;
        RECT 37.670 35.615 37.995 36.045 ;
        RECT 38.470 35.445 38.800 36.545 ;
        RECT 40.105 36.535 40.625 37.075 ;
        RECT 40.795 36.705 41.315 37.245 ;
        RECT 40.105 35.445 41.315 36.535 ;
        RECT 5.520 35.275 41.400 35.445 ;
        RECT 5.605 34.185 6.815 35.275 ;
        RECT 5.605 33.475 6.125 34.015 ;
        RECT 6.295 33.645 6.815 34.185 ;
        RECT 6.990 34.135 7.325 35.105 ;
        RECT 7.495 34.135 7.665 35.275 ;
        RECT 7.835 34.935 9.865 35.105 ;
        RECT 5.605 32.725 6.815 33.475 ;
        RECT 6.990 33.465 7.160 34.135 ;
        RECT 7.835 33.965 8.005 34.935 ;
        RECT 7.330 33.635 7.585 33.965 ;
        RECT 7.810 33.635 8.005 33.965 ;
        RECT 8.175 34.595 9.300 34.765 ;
        RECT 7.415 33.465 7.585 33.635 ;
        RECT 8.175 33.465 8.345 34.595 ;
        RECT 6.990 32.895 7.245 33.465 ;
        RECT 7.415 33.295 8.345 33.465 ;
        RECT 8.515 34.255 9.525 34.425 ;
        RECT 8.515 33.455 8.685 34.255 ;
        RECT 8.170 33.260 8.345 33.295 ;
        RECT 7.415 32.725 7.745 33.125 ;
        RECT 8.170 32.895 8.700 33.260 ;
        RECT 8.890 33.235 9.165 34.055 ;
        RECT 8.885 33.065 9.165 33.235 ;
        RECT 8.890 32.895 9.165 33.065 ;
        RECT 9.335 32.895 9.525 34.255 ;
        RECT 9.695 34.270 9.865 34.935 ;
        RECT 10.035 34.515 10.205 35.275 ;
        RECT 10.440 34.515 10.955 34.925 ;
        RECT 9.695 34.080 10.445 34.270 ;
        RECT 10.615 33.705 10.955 34.515 ;
        RECT 11.215 34.605 11.385 35.105 ;
        RECT 11.555 34.775 11.885 35.275 ;
        RECT 11.215 34.435 11.880 34.605 ;
        RECT 9.725 33.535 10.955 33.705 ;
        RECT 11.130 33.615 11.480 34.265 ;
        RECT 9.705 32.725 10.215 33.260 ;
        RECT 10.435 32.930 10.680 33.535 ;
        RECT 11.650 33.445 11.880 34.435 ;
        RECT 11.215 33.275 11.880 33.445 ;
        RECT 11.215 32.985 11.385 33.275 ;
        RECT 11.555 32.725 11.885 33.105 ;
        RECT 12.055 32.985 12.240 35.105 ;
        RECT 12.480 34.815 12.745 35.275 ;
        RECT 12.915 34.680 13.165 35.105 ;
        RECT 13.375 34.830 14.480 35.000 ;
        RECT 12.860 34.550 13.165 34.680 ;
        RECT 12.410 33.355 12.690 34.305 ;
        RECT 12.860 33.445 13.030 34.550 ;
        RECT 13.200 33.765 13.440 34.360 ;
        RECT 13.610 34.295 14.140 34.660 ;
        RECT 13.610 33.595 13.780 34.295 ;
        RECT 14.310 34.215 14.480 34.830 ;
        RECT 14.650 34.475 14.820 35.275 ;
        RECT 14.990 34.775 15.240 35.105 ;
        RECT 15.465 34.805 16.350 34.975 ;
        RECT 14.310 34.125 14.820 34.215 ;
        RECT 12.860 33.315 13.085 33.445 ;
        RECT 13.255 33.375 13.780 33.595 ;
        RECT 13.950 33.955 14.820 34.125 ;
        RECT 12.495 32.725 12.745 33.185 ;
        RECT 12.915 33.175 13.085 33.315 ;
        RECT 13.950 33.175 14.120 33.955 ;
        RECT 14.650 33.885 14.820 33.955 ;
        RECT 14.330 33.705 14.530 33.735 ;
        RECT 14.990 33.705 15.160 34.775 ;
        RECT 15.330 33.885 15.520 34.605 ;
        RECT 14.330 33.405 15.160 33.705 ;
        RECT 15.690 33.675 16.010 34.635 ;
        RECT 12.915 33.005 13.250 33.175 ;
        RECT 13.445 33.005 14.120 33.175 ;
        RECT 14.440 32.725 14.810 33.225 ;
        RECT 14.990 33.175 15.160 33.405 ;
        RECT 15.545 33.345 16.010 33.675 ;
        RECT 16.180 33.965 16.350 34.805 ;
        RECT 16.530 34.775 16.845 35.275 ;
        RECT 17.075 34.545 17.415 35.105 ;
        RECT 16.520 34.170 17.415 34.545 ;
        RECT 17.585 34.265 17.755 35.275 ;
        RECT 17.225 33.965 17.415 34.170 ;
        RECT 17.925 34.215 18.255 35.060 ;
        RECT 17.925 34.135 18.315 34.215 ;
        RECT 18.100 34.085 18.315 34.135 ;
        RECT 18.485 34.110 18.775 35.275 ;
        RECT 19.035 34.605 19.205 35.105 ;
        RECT 19.375 34.775 19.705 35.275 ;
        RECT 19.035 34.435 19.700 34.605 ;
        RECT 16.180 33.635 17.055 33.965 ;
        RECT 17.225 33.635 17.975 33.965 ;
        RECT 16.180 33.175 16.350 33.635 ;
        RECT 17.225 33.465 17.425 33.635 ;
        RECT 18.145 33.505 18.315 34.085 ;
        RECT 18.950 33.615 19.300 34.265 ;
        RECT 18.090 33.465 18.315 33.505 ;
        RECT 14.990 33.005 15.395 33.175 ;
        RECT 15.565 33.005 16.350 33.175 ;
        RECT 16.625 32.725 16.835 33.255 ;
        RECT 17.095 32.940 17.425 33.465 ;
        RECT 17.935 33.380 18.315 33.465 ;
        RECT 17.595 32.725 17.765 33.335 ;
        RECT 17.935 32.945 18.265 33.380 ;
        RECT 18.485 32.725 18.775 33.450 ;
        RECT 19.470 33.445 19.700 34.435 ;
        RECT 19.035 33.275 19.700 33.445 ;
        RECT 19.035 32.985 19.205 33.275 ;
        RECT 19.375 32.725 19.705 33.105 ;
        RECT 19.875 32.985 20.060 35.105 ;
        RECT 20.300 34.815 20.565 35.275 ;
        RECT 20.735 34.680 20.985 35.105 ;
        RECT 21.195 34.830 22.300 35.000 ;
        RECT 20.680 34.550 20.985 34.680 ;
        RECT 20.230 33.355 20.510 34.305 ;
        RECT 20.680 33.445 20.850 34.550 ;
        RECT 21.020 33.765 21.260 34.360 ;
        RECT 21.430 34.295 21.960 34.660 ;
        RECT 21.430 33.595 21.600 34.295 ;
        RECT 22.130 34.215 22.300 34.830 ;
        RECT 22.470 34.475 22.640 35.275 ;
        RECT 22.810 34.775 23.060 35.105 ;
        RECT 23.285 34.805 24.170 34.975 ;
        RECT 22.130 34.125 22.640 34.215 ;
        RECT 20.680 33.315 20.905 33.445 ;
        RECT 21.075 33.375 21.600 33.595 ;
        RECT 21.770 33.955 22.640 34.125 ;
        RECT 20.315 32.725 20.565 33.185 ;
        RECT 20.735 33.175 20.905 33.315 ;
        RECT 21.770 33.175 21.940 33.955 ;
        RECT 22.470 33.885 22.640 33.955 ;
        RECT 22.150 33.705 22.350 33.735 ;
        RECT 22.810 33.705 22.980 34.775 ;
        RECT 23.150 33.885 23.340 34.605 ;
        RECT 22.150 33.405 22.980 33.705 ;
        RECT 23.510 33.675 23.830 34.635 ;
        RECT 20.735 33.005 21.070 33.175 ;
        RECT 21.265 33.005 21.940 33.175 ;
        RECT 22.260 32.725 22.630 33.225 ;
        RECT 22.810 33.175 22.980 33.405 ;
        RECT 23.365 33.345 23.830 33.675 ;
        RECT 24.000 33.965 24.170 34.805 ;
        RECT 24.350 34.775 24.665 35.275 ;
        RECT 24.895 34.545 25.235 35.105 ;
        RECT 24.340 34.170 25.235 34.545 ;
        RECT 25.405 34.265 25.575 35.275 ;
        RECT 25.045 33.965 25.235 34.170 ;
        RECT 25.745 34.215 26.075 35.060 ;
        RECT 26.765 34.320 27.035 35.275 ;
        RECT 27.220 34.220 27.525 35.005 ;
        RECT 27.705 34.805 28.390 35.275 ;
        RECT 27.700 34.285 28.395 34.595 ;
        RECT 25.745 34.135 26.135 34.215 ;
        RECT 25.920 34.085 26.135 34.135 ;
        RECT 24.000 33.635 24.875 33.965 ;
        RECT 25.045 33.635 25.795 33.965 ;
        RECT 24.000 33.175 24.170 33.635 ;
        RECT 25.045 33.465 25.245 33.635 ;
        RECT 25.965 33.505 26.135 34.085 ;
        RECT 25.910 33.465 26.135 33.505 ;
        RECT 22.810 33.005 23.215 33.175 ;
        RECT 23.385 33.005 24.170 33.175 ;
        RECT 24.445 32.725 24.655 33.255 ;
        RECT 24.915 32.940 25.245 33.465 ;
        RECT 25.755 33.380 26.135 33.465 ;
        RECT 27.220 33.415 27.395 34.220 ;
        RECT 28.570 34.115 28.855 35.060 ;
        RECT 29.055 34.825 29.385 35.275 ;
        RECT 29.555 34.655 29.725 35.085 ;
        RECT 27.995 33.965 28.855 34.115 ;
        RECT 27.565 33.945 28.855 33.965 ;
        RECT 29.045 34.425 29.725 34.655 ;
        RECT 30.905 34.475 31.345 35.105 ;
        RECT 27.565 33.585 28.555 33.945 ;
        RECT 29.045 33.775 29.280 34.425 ;
        RECT 25.415 32.725 25.585 33.335 ;
        RECT 25.755 32.945 26.085 33.380 ;
        RECT 26.765 32.725 27.035 33.360 ;
        RECT 27.220 32.895 27.455 33.415 ;
        RECT 28.385 33.250 28.555 33.585 ;
        RECT 28.725 33.445 29.280 33.775 ;
        RECT 29.065 33.295 29.280 33.445 ;
        RECT 29.450 33.575 29.750 34.255 ;
        RECT 29.450 33.405 29.755 33.575 ;
        RECT 30.905 33.465 31.215 34.475 ;
        RECT 31.520 34.425 31.835 35.275 ;
        RECT 32.005 34.935 33.435 35.105 ;
        RECT 32.005 34.255 32.175 34.935 ;
        RECT 31.385 34.085 32.175 34.255 ;
        RECT 31.385 33.635 31.555 34.085 ;
        RECT 32.345 33.965 32.545 34.765 ;
        RECT 31.725 33.635 32.115 33.915 ;
        RECT 32.300 33.635 32.545 33.965 ;
        RECT 32.745 33.635 32.995 34.765 ;
        RECT 33.185 34.305 33.435 34.935 ;
        RECT 33.615 34.475 33.945 35.275 ;
        RECT 34.135 34.305 34.465 35.090 ;
        RECT 33.185 34.135 33.955 34.305 ;
        RECT 34.135 34.135 34.815 34.305 ;
        RECT 34.995 34.135 35.325 35.275 ;
        RECT 33.210 33.635 33.615 33.965 ;
        RECT 33.785 33.465 33.955 34.135 ;
        RECT 34.125 33.715 34.475 33.965 ;
        RECT 34.645 33.535 34.815 34.135 ;
        RECT 35.965 34.120 36.305 35.105 ;
        RECT 36.475 34.845 36.885 35.275 ;
        RECT 37.630 34.855 37.960 35.275 ;
        RECT 38.130 34.675 38.455 35.105 ;
        RECT 36.475 34.505 38.455 34.675 ;
        RECT 34.985 33.715 35.335 33.965 ;
        RECT 27.625 32.725 28.025 33.220 ;
        RECT 28.385 33.055 28.785 33.250 ;
        RECT 28.615 32.910 28.785 33.055 ;
        RECT 29.065 32.920 29.305 33.295 ;
        RECT 29.475 32.725 29.805 33.230 ;
        RECT 30.905 32.905 31.345 33.465 ;
        RECT 31.515 32.725 31.965 33.465 ;
        RECT 32.135 33.295 33.295 33.465 ;
        RECT 32.135 32.895 32.305 33.295 ;
        RECT 32.475 32.725 32.895 33.125 ;
        RECT 33.065 32.895 33.295 33.295 ;
        RECT 33.465 32.895 33.955 33.465 ;
        RECT 34.145 32.725 34.385 33.535 ;
        RECT 34.555 32.895 34.885 33.535 ;
        RECT 35.055 32.725 35.325 33.535 ;
        RECT 35.965 33.465 36.220 34.120 ;
        RECT 36.475 33.965 36.740 34.505 ;
        RECT 36.955 34.165 37.580 34.335 ;
        RECT 36.390 33.635 36.740 33.965 ;
        RECT 36.910 33.635 37.240 33.965 ;
        RECT 37.410 33.465 37.580 34.165 ;
        RECT 35.965 33.090 36.325 33.465 ;
        RECT 36.590 32.725 36.760 33.465 ;
        RECT 37.040 33.295 37.580 33.465 ;
        RECT 37.750 34.095 38.455 34.505 ;
        RECT 38.930 34.175 39.260 35.275 ;
        RECT 40.105 34.185 41.315 35.275 ;
        RECT 37.040 33.090 37.210 33.295 ;
        RECT 37.750 32.895 37.920 34.095 ;
        RECT 38.090 33.715 38.660 33.925 ;
        RECT 38.830 33.715 39.475 33.925 ;
        RECT 40.105 33.645 40.625 34.185 ;
        RECT 38.150 33.375 39.320 33.545 ;
        RECT 40.795 33.475 41.315 34.015 ;
        RECT 38.150 32.895 38.480 33.375 ;
        RECT 38.650 32.725 38.820 33.195 ;
        RECT 38.990 32.910 39.320 33.375 ;
        RECT 40.105 32.725 41.315 33.475 ;
        RECT 5.520 32.555 41.400 32.725 ;
        RECT 5.605 31.805 6.815 32.555 ;
        RECT 7.035 31.900 7.365 32.335 ;
        RECT 7.535 31.945 7.705 32.555 ;
        RECT 6.985 31.815 7.365 31.900 ;
        RECT 7.875 31.815 8.205 32.340 ;
        RECT 8.465 32.025 8.675 32.555 ;
        RECT 8.950 32.105 9.735 32.275 ;
        RECT 9.905 32.105 10.310 32.275 ;
        RECT 5.605 31.265 6.125 31.805 ;
        RECT 6.985 31.775 7.210 31.815 ;
        RECT 6.295 31.095 6.815 31.635 ;
        RECT 5.605 30.005 6.815 31.095 ;
        RECT 6.985 31.195 7.155 31.775 ;
        RECT 7.875 31.645 8.075 31.815 ;
        RECT 8.950 31.645 9.120 32.105 ;
        RECT 7.325 31.315 8.075 31.645 ;
        RECT 8.245 31.315 9.120 31.645 ;
        RECT 6.985 31.145 7.200 31.195 ;
        RECT 6.985 31.065 7.375 31.145 ;
        RECT 7.045 30.220 7.375 31.065 ;
        RECT 7.885 31.110 8.075 31.315 ;
        RECT 7.545 30.005 7.715 31.015 ;
        RECT 7.885 30.735 8.780 31.110 ;
        RECT 7.885 30.175 8.225 30.735 ;
        RECT 8.455 30.005 8.770 30.505 ;
        RECT 8.950 30.475 9.120 31.315 ;
        RECT 9.290 31.605 9.755 31.935 ;
        RECT 10.140 31.875 10.310 32.105 ;
        RECT 10.490 32.055 10.860 32.555 ;
        RECT 11.180 32.105 11.855 32.275 ;
        RECT 12.050 32.105 12.385 32.275 ;
        RECT 9.290 30.645 9.610 31.605 ;
        RECT 10.140 31.575 10.970 31.875 ;
        RECT 9.780 30.675 9.970 31.395 ;
        RECT 10.140 30.505 10.310 31.575 ;
        RECT 10.770 31.545 10.970 31.575 ;
        RECT 10.480 31.325 10.650 31.395 ;
        RECT 11.180 31.325 11.350 32.105 ;
        RECT 12.215 31.965 12.385 32.105 ;
        RECT 12.555 32.095 12.805 32.555 ;
        RECT 10.480 31.155 11.350 31.325 ;
        RECT 11.520 31.685 12.045 31.905 ;
        RECT 12.215 31.835 12.440 31.965 ;
        RECT 10.480 31.065 10.990 31.155 ;
        RECT 8.950 30.305 9.835 30.475 ;
        RECT 10.060 30.175 10.310 30.505 ;
        RECT 10.480 30.005 10.650 30.805 ;
        RECT 10.820 30.450 10.990 31.065 ;
        RECT 11.520 30.985 11.690 31.685 ;
        RECT 11.160 30.620 11.690 30.985 ;
        RECT 11.860 30.920 12.100 31.515 ;
        RECT 12.270 30.730 12.440 31.835 ;
        RECT 12.610 30.975 12.890 31.925 ;
        RECT 12.135 30.600 12.440 30.730 ;
        RECT 10.820 30.280 11.925 30.450 ;
        RECT 12.135 30.175 12.385 30.600 ;
        RECT 12.555 30.005 12.820 30.465 ;
        RECT 13.060 30.175 13.245 32.295 ;
        RECT 13.415 32.175 13.745 32.555 ;
        RECT 13.915 32.005 14.085 32.295 ;
        RECT 13.420 31.835 14.085 32.005 ;
        RECT 13.420 30.845 13.650 31.835 ;
        RECT 14.345 31.785 16.935 32.555 ;
        RECT 17.565 32.045 17.870 32.555 ;
        RECT 13.820 31.015 14.170 31.665 ;
        RECT 14.345 31.265 15.555 31.785 ;
        RECT 15.725 31.095 16.935 31.615 ;
        RECT 17.565 31.315 17.880 31.875 ;
        RECT 18.050 31.565 18.300 32.375 ;
        RECT 18.470 32.030 18.730 32.555 ;
        RECT 18.910 31.565 19.160 32.375 ;
        RECT 19.330 31.995 19.590 32.555 ;
        RECT 19.760 31.905 20.020 32.360 ;
        RECT 20.190 32.075 20.450 32.555 ;
        RECT 20.620 31.905 20.880 32.360 ;
        RECT 21.050 32.075 21.310 32.555 ;
        RECT 21.480 31.905 21.740 32.360 ;
        RECT 21.910 32.075 22.155 32.555 ;
        RECT 22.325 31.905 22.600 32.360 ;
        RECT 22.770 32.075 23.015 32.555 ;
        RECT 23.185 31.905 23.445 32.360 ;
        RECT 23.625 32.075 23.875 32.555 ;
        RECT 24.045 31.905 24.305 32.360 ;
        RECT 24.485 32.075 24.735 32.555 ;
        RECT 24.905 31.905 25.165 32.360 ;
        RECT 25.345 32.075 25.605 32.555 ;
        RECT 25.775 31.905 26.035 32.360 ;
        RECT 26.205 32.075 26.505 32.555 ;
        RECT 19.760 31.735 26.505 31.905 ;
        RECT 18.050 31.315 25.170 31.565 ;
        RECT 13.420 30.675 14.085 30.845 ;
        RECT 13.415 30.005 13.745 30.505 ;
        RECT 13.915 30.175 14.085 30.675 ;
        RECT 14.345 30.005 16.935 31.095 ;
        RECT 17.575 30.005 17.870 30.815 ;
        RECT 18.050 30.175 18.295 31.315 ;
        RECT 18.470 30.005 18.730 30.815 ;
        RECT 18.910 30.180 19.160 31.315 ;
        RECT 25.340 31.145 26.505 31.735 ;
        RECT 19.760 30.920 26.505 31.145 ;
        RECT 26.765 31.815 27.150 32.385 ;
        RECT 27.320 32.095 27.645 32.555 ;
        RECT 28.165 31.925 28.445 32.385 ;
        RECT 26.765 31.145 27.045 31.815 ;
        RECT 27.320 31.755 28.445 31.925 ;
        RECT 27.320 31.645 27.770 31.755 ;
        RECT 27.215 31.315 27.770 31.645 ;
        RECT 28.635 31.585 29.035 32.385 ;
        RECT 29.435 32.095 29.705 32.555 ;
        RECT 29.875 31.925 30.160 32.385 ;
        RECT 19.760 30.905 25.165 30.920 ;
        RECT 19.330 30.010 19.590 30.805 ;
        RECT 19.760 30.180 20.020 30.905 ;
        RECT 20.190 30.010 20.450 30.735 ;
        RECT 20.620 30.180 20.880 30.905 ;
        RECT 21.050 30.010 21.310 30.735 ;
        RECT 21.480 30.180 21.740 30.905 ;
        RECT 21.910 30.010 22.170 30.735 ;
        RECT 22.340 30.180 22.600 30.905 ;
        RECT 22.770 30.010 23.015 30.735 ;
        RECT 23.185 30.180 23.445 30.905 ;
        RECT 23.630 30.010 23.875 30.735 ;
        RECT 24.045 30.180 24.305 30.905 ;
        RECT 24.490 30.010 24.735 30.735 ;
        RECT 24.905 30.180 25.165 30.905 ;
        RECT 25.350 30.010 25.605 30.735 ;
        RECT 25.775 30.180 26.065 30.920 ;
        RECT 19.330 30.005 25.605 30.010 ;
        RECT 26.235 30.005 26.505 30.750 ;
        RECT 26.765 30.175 27.150 31.145 ;
        RECT 27.320 30.855 27.770 31.315 ;
        RECT 27.940 31.025 29.035 31.585 ;
        RECT 27.320 30.635 28.445 30.855 ;
        RECT 27.320 30.005 27.645 30.465 ;
        RECT 28.165 30.175 28.445 30.635 ;
        RECT 28.635 30.175 29.035 31.025 ;
        RECT 29.205 31.755 30.160 31.925 ;
        RECT 31.365 31.830 31.655 32.555 ;
        RECT 31.840 31.985 32.095 32.335 ;
        RECT 32.265 32.155 32.595 32.555 ;
        RECT 32.765 31.985 32.935 32.335 ;
        RECT 33.105 32.155 33.485 32.555 ;
        RECT 31.840 31.815 33.505 31.985 ;
        RECT 33.675 31.880 33.950 32.225 ;
        RECT 29.205 30.855 29.415 31.755 ;
        RECT 33.335 31.645 33.505 31.815 ;
        RECT 29.585 31.025 30.275 31.585 ;
        RECT 31.825 31.315 32.170 31.645 ;
        RECT 32.340 31.315 33.165 31.645 ;
        RECT 33.335 31.315 33.610 31.645 ;
        RECT 29.205 30.635 30.160 30.855 ;
        RECT 29.435 30.005 29.705 30.465 ;
        RECT 29.875 30.175 30.160 30.635 ;
        RECT 31.365 30.005 31.655 31.170 ;
        RECT 31.845 30.855 32.170 31.145 ;
        RECT 32.340 31.025 32.535 31.315 ;
        RECT 33.335 31.145 33.505 31.315 ;
        RECT 33.780 31.145 33.950 31.880 ;
        RECT 34.125 31.785 36.715 32.555 ;
        RECT 34.125 31.265 35.335 31.785 ;
        RECT 37.355 31.745 37.625 32.555 ;
        RECT 37.795 31.745 38.125 32.385 ;
        RECT 38.295 31.745 38.535 32.555 ;
        RECT 38.725 31.880 38.985 32.385 ;
        RECT 39.165 32.175 39.495 32.555 ;
        RECT 39.675 32.005 39.845 32.385 ;
        RECT 32.845 30.975 33.505 31.145 ;
        RECT 32.845 30.855 33.015 30.975 ;
        RECT 31.845 30.685 33.015 30.855 ;
        RECT 31.825 30.225 33.015 30.515 ;
        RECT 33.185 30.005 33.465 30.805 ;
        RECT 33.675 30.175 33.950 31.145 ;
        RECT 35.505 31.095 36.715 31.615 ;
        RECT 37.345 31.315 37.695 31.565 ;
        RECT 37.865 31.145 38.035 31.745 ;
        RECT 38.205 31.315 38.555 31.565 ;
        RECT 34.125 30.005 36.715 31.095 ;
        RECT 37.355 30.005 37.685 31.145 ;
        RECT 37.865 30.975 38.545 31.145 ;
        RECT 38.215 30.190 38.545 30.975 ;
        RECT 38.725 31.080 38.895 31.880 ;
        RECT 39.180 31.835 39.845 32.005 ;
        RECT 39.180 31.580 39.350 31.835 ;
        RECT 40.105 31.805 41.315 32.555 ;
        RECT 39.065 31.250 39.350 31.580 ;
        RECT 39.585 31.285 39.915 31.655 ;
        RECT 39.180 31.105 39.350 31.250 ;
        RECT 38.725 30.175 38.995 31.080 ;
        RECT 39.180 30.935 39.845 31.105 ;
        RECT 39.165 30.005 39.495 30.765 ;
        RECT 39.675 30.175 39.845 30.935 ;
        RECT 40.105 31.095 40.625 31.635 ;
        RECT 40.795 31.265 41.315 31.805 ;
        RECT 40.105 30.005 41.315 31.095 ;
        RECT 5.520 29.835 41.400 30.005 ;
        RECT 5.605 28.745 6.815 29.835 ;
        RECT 6.985 28.745 8.195 29.835 ;
        RECT 8.480 29.205 8.765 29.665 ;
        RECT 8.935 29.375 9.205 29.835 ;
        RECT 8.480 28.985 9.435 29.205 ;
        RECT 5.605 28.035 6.125 28.575 ;
        RECT 6.295 28.205 6.815 28.745 ;
        RECT 6.985 28.035 7.505 28.575 ;
        RECT 7.675 28.205 8.195 28.745 ;
        RECT 8.365 28.255 9.055 28.815 ;
        RECT 9.225 28.085 9.435 28.985 ;
        RECT 5.605 27.285 6.815 28.035 ;
        RECT 6.985 27.285 8.195 28.035 ;
        RECT 8.480 27.915 9.435 28.085 ;
        RECT 9.605 28.815 10.005 29.665 ;
        RECT 10.195 29.205 10.475 29.665 ;
        RECT 10.995 29.375 11.320 29.835 ;
        RECT 10.195 28.985 11.320 29.205 ;
        RECT 9.605 28.255 10.700 28.815 ;
        RECT 10.870 28.525 11.320 28.985 ;
        RECT 11.490 28.695 11.875 29.665 ;
        RECT 8.480 27.455 8.765 27.915 ;
        RECT 8.935 27.285 9.205 27.745 ;
        RECT 9.605 27.455 10.005 28.255 ;
        RECT 10.870 28.195 11.425 28.525 ;
        RECT 10.870 28.085 11.320 28.195 ;
        RECT 10.195 27.915 11.320 28.085 ;
        RECT 11.595 28.025 11.875 28.695 ;
        RECT 10.195 27.455 10.475 27.915 ;
        RECT 10.995 27.285 11.320 27.745 ;
        RECT 11.490 27.455 11.875 28.025 ;
        RECT 12.045 28.695 12.430 29.665 ;
        RECT 12.600 29.375 12.925 29.835 ;
        RECT 13.445 29.205 13.725 29.665 ;
        RECT 12.600 28.985 13.725 29.205 ;
        RECT 12.045 28.025 12.325 28.695 ;
        RECT 12.600 28.525 13.050 28.985 ;
        RECT 13.915 28.815 14.315 29.665 ;
        RECT 14.715 29.375 14.985 29.835 ;
        RECT 15.155 29.205 15.440 29.665 ;
        RECT 12.495 28.195 13.050 28.525 ;
        RECT 13.220 28.255 14.315 28.815 ;
        RECT 12.600 28.085 13.050 28.195 ;
        RECT 12.045 27.455 12.430 28.025 ;
        RECT 12.600 27.915 13.725 28.085 ;
        RECT 12.600 27.285 12.925 27.745 ;
        RECT 13.445 27.455 13.725 27.915 ;
        RECT 13.915 27.455 14.315 28.255 ;
        RECT 14.485 28.985 15.440 29.205 ;
        RECT 14.485 28.085 14.695 28.985 ;
        RECT 14.865 28.255 15.555 28.815 ;
        RECT 15.725 28.745 18.315 29.835 ;
        RECT 14.485 27.915 15.440 28.085 ;
        RECT 14.715 27.285 14.985 27.745 ;
        RECT 15.155 27.455 15.440 27.915 ;
        RECT 15.725 28.055 16.935 28.575 ;
        RECT 17.105 28.225 18.315 28.745 ;
        RECT 18.485 28.670 18.775 29.835 ;
        RECT 18.955 28.695 19.285 29.835 ;
        RECT 19.815 28.865 20.145 29.650 ;
        RECT 19.465 28.695 20.145 28.865 ;
        RECT 20.445 28.715 20.775 29.835 ;
        RECT 18.945 28.275 19.295 28.525 ;
        RECT 19.465 28.095 19.635 28.695 ;
        RECT 19.805 28.275 20.155 28.525 ;
        RECT 20.385 28.275 20.895 28.525 ;
        RECT 21.105 28.275 21.475 29.590 ;
        RECT 21.645 28.275 21.975 29.590 ;
        RECT 22.185 28.275 22.515 29.590 ;
        RECT 22.785 28.945 23.035 29.665 ;
        RECT 23.205 29.115 23.535 29.835 ;
        RECT 22.785 28.655 23.535 28.945 ;
        RECT 23.770 28.655 24.295 29.665 ;
        RECT 23.275 28.485 23.535 28.655 ;
        RECT 22.685 28.275 23.105 28.485 ;
        RECT 23.275 28.275 23.855 28.485 ;
        RECT 23.275 28.105 23.645 28.275 ;
        RECT 15.725 27.285 18.315 28.055 ;
        RECT 18.485 27.285 18.775 28.010 ;
        RECT 18.955 27.285 19.225 28.095 ;
        RECT 19.395 27.455 19.725 28.095 ;
        RECT 19.895 27.285 20.135 28.095 ;
        RECT 20.425 27.935 22.725 28.105 ;
        RECT 20.425 27.455 20.755 27.935 ;
        RECT 20.925 27.285 21.255 27.745 ;
        RECT 21.470 27.455 21.800 27.935 ;
        RECT 22.000 27.285 22.330 27.745 ;
        RECT 22.555 27.615 22.725 27.935 ;
        RECT 22.895 27.915 23.645 28.105 ;
        RECT 24.025 28.085 24.295 28.655 ;
        RECT 22.895 27.470 23.225 27.915 ;
        RECT 23.495 27.285 23.665 27.745 ;
        RECT 23.955 27.455 24.295 28.085 ;
        RECT 24.465 28.695 24.850 29.665 ;
        RECT 25.020 29.375 25.345 29.835 ;
        RECT 25.865 29.205 26.145 29.665 ;
        RECT 25.020 28.985 26.145 29.205 ;
        RECT 24.465 28.025 24.745 28.695 ;
        RECT 25.020 28.525 25.470 28.985 ;
        RECT 26.335 28.815 26.735 29.665 ;
        RECT 27.135 29.375 27.405 29.835 ;
        RECT 27.575 29.205 27.860 29.665 ;
        RECT 24.915 28.195 25.470 28.525 ;
        RECT 25.640 28.255 26.735 28.815 ;
        RECT 25.020 28.085 25.470 28.195 ;
        RECT 24.465 27.455 24.850 28.025 ;
        RECT 25.020 27.915 26.145 28.085 ;
        RECT 25.020 27.285 25.345 27.745 ;
        RECT 25.865 27.455 26.145 27.915 ;
        RECT 26.335 27.455 26.735 28.255 ;
        RECT 26.905 28.985 27.860 29.205 ;
        RECT 26.905 28.085 27.115 28.985 ;
        RECT 27.285 28.255 27.975 28.815 ;
        RECT 28.145 28.745 29.355 29.835 ;
        RECT 26.905 27.915 27.860 28.085 ;
        RECT 27.135 27.285 27.405 27.745 ;
        RECT 27.575 27.455 27.860 27.915 ;
        RECT 28.145 28.035 28.665 28.575 ;
        RECT 28.835 28.205 29.355 28.745 ;
        RECT 29.525 28.695 29.800 29.665 ;
        RECT 30.010 29.035 30.290 29.835 ;
        RECT 30.460 29.325 32.510 29.615 ;
        RECT 30.460 28.985 32.090 29.155 ;
        RECT 30.460 28.865 30.630 28.985 ;
        RECT 29.970 28.695 30.630 28.865 ;
        RECT 28.145 27.285 29.355 28.035 ;
        RECT 29.525 27.960 29.695 28.695 ;
        RECT 29.970 28.525 30.140 28.695 ;
        RECT 29.865 28.195 30.140 28.525 ;
        RECT 30.310 28.195 30.690 28.525 ;
        RECT 30.860 28.195 31.600 28.815 ;
        RECT 31.770 28.695 32.090 28.985 ;
        RECT 32.285 28.525 32.525 29.120 ;
        RECT 32.695 28.760 33.035 29.835 ;
        RECT 33.215 28.865 33.545 29.650 ;
        RECT 33.215 28.695 33.895 28.865 ;
        RECT 34.075 28.695 34.405 29.835 ;
        RECT 34.665 28.905 34.845 29.665 ;
        RECT 35.025 29.075 35.355 29.835 ;
        RECT 34.665 28.735 35.340 28.905 ;
        RECT 35.525 28.760 35.795 29.665 ;
        RECT 31.870 28.195 32.525 28.525 ;
        RECT 29.970 28.025 30.140 28.195 ;
        RECT 29.525 27.615 29.800 27.960 ;
        RECT 29.970 27.855 31.555 28.025 ;
        RECT 29.990 27.285 30.370 27.685 ;
        RECT 30.540 27.505 30.710 27.855 ;
        RECT 30.880 27.285 31.210 27.685 ;
        RECT 31.385 27.505 31.555 27.855 ;
        RECT 31.755 27.285 32.085 27.785 ;
        RECT 32.280 27.505 32.525 28.195 ;
        RECT 32.695 27.955 33.035 28.525 ;
        RECT 33.205 28.275 33.555 28.525 ;
        RECT 33.725 28.095 33.895 28.695 ;
        RECT 35.170 28.590 35.340 28.735 ;
        RECT 34.065 28.275 34.415 28.525 ;
        RECT 34.605 28.185 34.945 28.555 ;
        RECT 35.170 28.260 35.445 28.590 ;
        RECT 32.695 27.285 33.035 27.785 ;
        RECT 33.225 27.285 33.465 28.095 ;
        RECT 33.635 27.455 33.965 28.095 ;
        RECT 34.135 27.285 34.405 28.095 ;
        RECT 35.170 28.005 35.340 28.260 ;
        RECT 34.675 27.835 35.340 28.005 ;
        RECT 35.615 27.960 35.795 28.760 ;
        RECT 36.180 28.735 36.510 29.835 ;
        RECT 36.985 29.235 37.310 29.665 ;
        RECT 37.480 29.415 37.810 29.835 ;
        RECT 38.555 29.405 38.965 29.835 ;
        RECT 36.985 29.065 38.965 29.235 ;
        RECT 36.985 28.655 37.690 29.065 ;
        RECT 35.965 28.275 36.610 28.485 ;
        RECT 36.780 28.275 37.350 28.485 ;
        RECT 34.675 27.455 34.845 27.835 ;
        RECT 35.025 27.285 35.355 27.665 ;
        RECT 35.535 27.455 35.795 27.960 ;
        RECT 36.120 27.935 37.290 28.105 ;
        RECT 36.120 27.470 36.450 27.935 ;
        RECT 36.620 27.285 36.790 27.755 ;
        RECT 36.960 27.455 37.290 27.935 ;
        RECT 37.520 27.455 37.690 28.655 ;
        RECT 37.860 28.725 38.485 28.895 ;
        RECT 37.860 28.025 38.030 28.725 ;
        RECT 38.700 28.525 38.965 29.065 ;
        RECT 39.135 28.680 39.475 29.665 ;
        RECT 38.200 28.195 38.530 28.525 ;
        RECT 38.700 28.195 39.050 28.525 ;
        RECT 39.220 28.025 39.475 28.680 ;
        RECT 40.105 28.745 41.315 29.835 ;
        RECT 40.105 28.205 40.625 28.745 ;
        RECT 40.795 28.035 41.315 28.575 ;
        RECT 37.860 27.855 38.400 28.025 ;
        RECT 38.230 27.650 38.400 27.855 ;
        RECT 38.680 27.285 38.850 28.025 ;
        RECT 39.115 27.650 39.475 28.025 ;
        RECT 40.105 27.285 41.315 28.035 ;
        RECT 5.520 27.115 41.400 27.285 ;
        RECT 5.605 26.365 6.815 27.115 ;
        RECT 5.605 25.825 6.125 26.365 ;
        RECT 6.990 26.275 7.250 27.115 ;
        RECT 7.425 26.370 7.680 26.945 ;
        RECT 7.850 26.735 8.180 27.115 ;
        RECT 8.395 26.565 8.565 26.945 ;
        RECT 7.850 26.395 8.565 26.565 ;
        RECT 6.295 25.655 6.815 26.195 ;
        RECT 5.605 24.565 6.815 25.655 ;
        RECT 6.990 24.565 7.250 25.715 ;
        RECT 7.425 25.640 7.595 26.370 ;
        RECT 7.850 26.205 8.020 26.395 ;
        RECT 9.290 26.375 9.545 26.945 ;
        RECT 9.715 26.715 10.045 27.115 ;
        RECT 10.470 26.580 11.000 26.945 ;
        RECT 11.190 26.775 11.465 26.945 ;
        RECT 11.185 26.605 11.465 26.775 ;
        RECT 10.470 26.545 10.645 26.580 ;
        RECT 9.715 26.375 10.645 26.545 ;
        RECT 7.765 25.875 8.020 26.205 ;
        RECT 7.850 25.665 8.020 25.875 ;
        RECT 8.300 25.845 8.655 26.215 ;
        RECT 9.290 25.705 9.460 26.375 ;
        RECT 9.715 26.205 9.885 26.375 ;
        RECT 9.630 25.875 9.885 26.205 ;
        RECT 10.110 25.875 10.305 26.205 ;
        RECT 7.425 24.735 7.680 25.640 ;
        RECT 7.850 25.495 8.565 25.665 ;
        RECT 7.850 24.565 8.180 25.325 ;
        RECT 8.395 24.735 8.565 25.495 ;
        RECT 9.290 24.735 9.625 25.705 ;
        RECT 9.795 24.565 9.965 25.705 ;
        RECT 10.135 24.905 10.305 25.875 ;
        RECT 10.475 25.245 10.645 26.375 ;
        RECT 10.815 25.585 10.985 26.385 ;
        RECT 11.190 25.785 11.465 26.605 ;
        RECT 11.635 25.585 11.825 26.945 ;
        RECT 12.005 26.580 12.515 27.115 ;
        RECT 12.735 26.305 12.980 26.910 ;
        RECT 13.515 26.565 13.685 26.855 ;
        RECT 13.855 26.735 14.185 27.115 ;
        RECT 13.515 26.395 14.180 26.565 ;
        RECT 12.025 26.135 13.255 26.305 ;
        RECT 10.815 25.415 11.825 25.585 ;
        RECT 11.995 25.570 12.745 25.760 ;
        RECT 10.475 25.075 11.600 25.245 ;
        RECT 11.995 24.905 12.165 25.570 ;
        RECT 12.915 25.325 13.255 26.135 ;
        RECT 13.430 25.575 13.780 26.225 ;
        RECT 13.950 25.405 14.180 26.395 ;
        RECT 10.135 24.735 12.165 24.905 ;
        RECT 12.335 24.565 12.505 25.325 ;
        RECT 12.740 24.915 13.255 25.325 ;
        RECT 13.515 25.235 14.180 25.405 ;
        RECT 13.515 24.735 13.685 25.235 ;
        RECT 13.855 24.565 14.185 25.065 ;
        RECT 14.355 24.735 14.540 26.855 ;
        RECT 14.795 26.655 15.045 27.115 ;
        RECT 15.215 26.665 15.550 26.835 ;
        RECT 15.745 26.665 16.420 26.835 ;
        RECT 15.215 26.525 15.385 26.665 ;
        RECT 14.710 25.535 14.990 26.485 ;
        RECT 15.160 26.395 15.385 26.525 ;
        RECT 15.160 25.290 15.330 26.395 ;
        RECT 15.555 26.245 16.080 26.465 ;
        RECT 15.500 25.480 15.740 26.075 ;
        RECT 15.910 25.545 16.080 26.245 ;
        RECT 16.250 25.885 16.420 26.665 ;
        RECT 16.740 26.615 17.110 27.115 ;
        RECT 17.290 26.665 17.695 26.835 ;
        RECT 17.865 26.665 18.650 26.835 ;
        RECT 17.290 26.435 17.460 26.665 ;
        RECT 16.630 26.135 17.460 26.435 ;
        RECT 17.845 26.165 18.310 26.495 ;
        RECT 16.630 26.105 16.830 26.135 ;
        RECT 16.950 25.885 17.120 25.955 ;
        RECT 16.250 25.715 17.120 25.885 ;
        RECT 16.610 25.625 17.120 25.715 ;
        RECT 15.160 25.160 15.465 25.290 ;
        RECT 15.910 25.180 16.440 25.545 ;
        RECT 14.780 24.565 15.045 25.025 ;
        RECT 15.215 24.735 15.465 25.160 ;
        RECT 16.610 25.010 16.780 25.625 ;
        RECT 15.675 24.840 16.780 25.010 ;
        RECT 16.950 24.565 17.120 25.365 ;
        RECT 17.290 25.065 17.460 26.135 ;
        RECT 17.630 25.235 17.820 25.955 ;
        RECT 17.990 25.205 18.310 26.165 ;
        RECT 18.480 26.205 18.650 26.665 ;
        RECT 18.925 26.585 19.135 27.115 ;
        RECT 19.395 26.375 19.725 26.900 ;
        RECT 19.895 26.505 20.065 27.115 ;
        RECT 20.235 26.460 20.565 26.895 ;
        RECT 20.235 26.375 20.615 26.460 ;
        RECT 19.525 26.205 19.725 26.375 ;
        RECT 20.390 26.335 20.615 26.375 ;
        RECT 18.480 25.875 19.355 26.205 ;
        RECT 19.525 25.875 20.275 26.205 ;
        RECT 17.290 24.735 17.540 25.065 ;
        RECT 18.480 25.035 18.650 25.875 ;
        RECT 19.525 25.670 19.715 25.875 ;
        RECT 20.445 25.755 20.615 26.335 ;
        RECT 20.400 25.705 20.615 25.755 ;
        RECT 18.820 25.295 19.715 25.670 ;
        RECT 20.225 25.625 20.615 25.705 ;
        RECT 20.790 26.375 21.045 26.945 ;
        RECT 21.215 26.715 21.545 27.115 ;
        RECT 21.970 26.580 22.500 26.945 ;
        RECT 21.970 26.545 22.145 26.580 ;
        RECT 21.215 26.375 22.145 26.545 ;
        RECT 20.790 25.705 20.960 26.375 ;
        RECT 21.215 26.205 21.385 26.375 ;
        RECT 21.130 25.875 21.385 26.205 ;
        RECT 21.610 25.875 21.805 26.205 ;
        RECT 17.765 24.865 18.650 25.035 ;
        RECT 18.830 24.565 19.145 25.065 ;
        RECT 19.375 24.735 19.715 25.295 ;
        RECT 19.885 24.565 20.055 25.575 ;
        RECT 20.225 24.780 20.555 25.625 ;
        RECT 20.790 24.735 21.125 25.705 ;
        RECT 21.295 24.565 21.465 25.705 ;
        RECT 21.635 24.905 21.805 25.875 ;
        RECT 21.975 25.245 22.145 26.375 ;
        RECT 22.315 25.585 22.485 26.385 ;
        RECT 22.690 26.095 22.965 26.945 ;
        RECT 22.685 25.925 22.965 26.095 ;
        RECT 22.690 25.785 22.965 25.925 ;
        RECT 23.135 25.585 23.325 26.945 ;
        RECT 23.505 26.580 24.015 27.115 ;
        RECT 24.235 26.305 24.480 26.910 ;
        RECT 24.925 26.375 25.310 26.945 ;
        RECT 25.480 26.655 25.805 27.115 ;
        RECT 26.325 26.485 26.605 26.945 ;
        RECT 23.525 26.135 24.755 26.305 ;
        RECT 22.315 25.415 23.325 25.585 ;
        RECT 23.495 25.570 24.245 25.760 ;
        RECT 21.975 25.075 23.100 25.245 ;
        RECT 23.495 24.905 23.665 25.570 ;
        RECT 24.415 25.325 24.755 26.135 ;
        RECT 21.635 24.735 23.665 24.905 ;
        RECT 23.835 24.565 24.005 25.325 ;
        RECT 24.240 24.915 24.755 25.325 ;
        RECT 24.925 25.705 25.205 26.375 ;
        RECT 25.480 26.315 26.605 26.485 ;
        RECT 25.480 26.205 25.930 26.315 ;
        RECT 25.375 25.875 25.930 26.205 ;
        RECT 26.795 26.145 27.195 26.945 ;
        RECT 27.595 26.655 27.865 27.115 ;
        RECT 28.035 26.485 28.320 26.945 ;
        RECT 24.925 24.735 25.310 25.705 ;
        RECT 25.480 25.415 25.930 25.875 ;
        RECT 26.100 25.585 27.195 26.145 ;
        RECT 25.480 25.195 26.605 25.415 ;
        RECT 25.480 24.565 25.805 25.025 ;
        RECT 26.325 24.735 26.605 25.195 ;
        RECT 26.795 24.735 27.195 25.585 ;
        RECT 27.365 26.315 28.320 26.485 ;
        RECT 28.605 26.345 31.195 27.115 ;
        RECT 31.365 26.390 31.655 27.115 ;
        RECT 32.155 26.715 32.485 27.115 ;
        RECT 32.655 26.545 32.985 26.885 ;
        RECT 34.035 26.715 34.365 27.115 ;
        RECT 32.000 26.375 34.365 26.545 ;
        RECT 34.535 26.390 34.865 26.900 ;
        RECT 27.365 25.415 27.575 26.315 ;
        RECT 27.745 25.585 28.435 26.145 ;
        RECT 28.605 25.825 29.815 26.345 ;
        RECT 29.985 25.655 31.195 26.175 ;
        RECT 27.365 25.195 28.320 25.415 ;
        RECT 27.595 24.565 27.865 25.025 ;
        RECT 28.035 24.735 28.320 25.195 ;
        RECT 28.605 24.565 31.195 25.655 ;
        RECT 31.365 24.565 31.655 25.730 ;
        RECT 32.000 25.375 32.170 26.375 ;
        RECT 34.195 26.205 34.365 26.375 ;
        RECT 32.340 25.545 32.585 26.205 ;
        RECT 32.800 25.545 33.065 26.205 ;
        RECT 33.260 25.545 33.545 26.205 ;
        RECT 33.720 25.875 34.025 26.205 ;
        RECT 34.195 25.875 34.505 26.205 ;
        RECT 33.720 25.545 33.935 25.875 ;
        RECT 32.000 25.205 32.455 25.375 ;
        RECT 32.125 24.775 32.455 25.205 ;
        RECT 32.635 25.205 33.925 25.375 ;
        RECT 32.635 24.785 32.885 25.205 ;
        RECT 33.115 24.565 33.445 25.035 ;
        RECT 33.675 24.785 33.925 25.205 ;
        RECT 34.115 24.565 34.365 25.705 ;
        RECT 34.675 25.625 34.865 26.390 ;
        RECT 36.120 26.465 36.450 26.930 ;
        RECT 36.620 26.645 36.790 27.115 ;
        RECT 36.960 26.465 37.290 26.945 ;
        RECT 36.120 26.295 37.290 26.465 ;
        RECT 35.965 25.915 36.610 26.125 ;
        RECT 36.780 25.915 37.350 26.125 ;
        RECT 37.520 25.745 37.690 26.945 ;
        RECT 38.230 26.545 38.400 26.750 ;
        RECT 34.535 24.775 34.865 25.625 ;
        RECT 36.180 24.565 36.510 25.665 ;
        RECT 36.985 25.335 37.690 25.745 ;
        RECT 37.860 26.375 38.400 26.545 ;
        RECT 38.680 26.375 38.850 27.115 ;
        RECT 39.245 26.750 39.415 26.775 ;
        RECT 39.115 26.375 39.475 26.750 ;
        RECT 37.860 25.675 38.030 26.375 ;
        RECT 38.200 25.875 38.530 26.205 ;
        RECT 38.700 25.875 39.050 26.205 ;
        RECT 37.860 25.505 38.485 25.675 ;
        RECT 38.700 25.335 38.965 25.875 ;
        RECT 39.220 25.720 39.475 26.375 ;
        RECT 40.105 26.365 41.315 27.115 ;
        RECT 36.985 25.165 38.965 25.335 ;
        RECT 36.985 24.735 37.310 25.165 ;
        RECT 37.480 24.565 37.810 24.985 ;
        RECT 38.555 24.565 38.965 24.995 ;
        RECT 39.135 24.735 39.475 25.720 ;
        RECT 40.105 25.655 40.625 26.195 ;
        RECT 40.795 25.825 41.315 26.365 ;
        RECT 40.105 24.565 41.315 25.655 ;
        RECT 5.520 24.395 41.400 24.565 ;
        RECT 5.605 23.305 6.815 24.395 ;
        RECT 7.075 23.725 7.245 24.225 ;
        RECT 7.415 23.895 7.745 24.395 ;
        RECT 7.075 23.555 7.740 23.725 ;
        RECT 5.605 22.595 6.125 23.135 ;
        RECT 6.295 22.765 6.815 23.305 ;
        RECT 6.990 22.735 7.340 23.385 ;
        RECT 5.605 21.845 6.815 22.595 ;
        RECT 7.510 22.565 7.740 23.555 ;
        RECT 7.075 22.395 7.740 22.565 ;
        RECT 7.075 22.105 7.245 22.395 ;
        RECT 7.415 21.845 7.745 22.225 ;
        RECT 7.915 22.105 8.100 24.225 ;
        RECT 8.340 23.935 8.605 24.395 ;
        RECT 8.775 23.800 9.025 24.225 ;
        RECT 9.235 23.950 10.340 24.120 ;
        RECT 8.720 23.670 9.025 23.800 ;
        RECT 8.270 22.475 8.550 23.425 ;
        RECT 8.720 22.565 8.890 23.670 ;
        RECT 9.060 22.885 9.300 23.480 ;
        RECT 9.470 23.415 10.000 23.780 ;
        RECT 9.470 22.715 9.640 23.415 ;
        RECT 10.170 23.335 10.340 23.950 ;
        RECT 10.510 23.595 10.680 24.395 ;
        RECT 10.850 23.895 11.100 24.225 ;
        RECT 11.325 23.925 12.210 24.095 ;
        RECT 10.170 23.245 10.680 23.335 ;
        RECT 8.720 22.435 8.945 22.565 ;
        RECT 9.115 22.495 9.640 22.715 ;
        RECT 9.810 23.075 10.680 23.245 ;
        RECT 8.355 21.845 8.605 22.305 ;
        RECT 8.775 22.295 8.945 22.435 ;
        RECT 9.810 22.295 9.980 23.075 ;
        RECT 10.510 23.005 10.680 23.075 ;
        RECT 10.190 22.825 10.390 22.855 ;
        RECT 10.850 22.825 11.020 23.895 ;
        RECT 11.190 23.005 11.380 23.725 ;
        RECT 10.190 22.525 11.020 22.825 ;
        RECT 11.550 22.795 11.870 23.755 ;
        RECT 8.775 22.125 9.110 22.295 ;
        RECT 9.305 22.125 9.980 22.295 ;
        RECT 10.300 21.845 10.670 22.345 ;
        RECT 10.850 22.295 11.020 22.525 ;
        RECT 11.405 22.465 11.870 22.795 ;
        RECT 12.040 23.085 12.210 23.925 ;
        RECT 12.390 23.895 12.705 24.395 ;
        RECT 12.935 23.665 13.275 24.225 ;
        RECT 12.380 23.290 13.275 23.665 ;
        RECT 13.445 23.385 13.615 24.395 ;
        RECT 13.085 23.085 13.275 23.290 ;
        RECT 13.785 23.335 14.115 24.180 ;
        RECT 13.785 23.255 14.175 23.335 ;
        RECT 14.345 23.305 17.855 24.395 ;
        RECT 13.960 23.205 14.175 23.255 ;
        RECT 12.040 22.755 12.915 23.085 ;
        RECT 13.085 22.755 13.835 23.085 ;
        RECT 12.040 22.295 12.210 22.755 ;
        RECT 13.085 22.585 13.285 22.755 ;
        RECT 14.005 22.625 14.175 23.205 ;
        RECT 13.950 22.585 14.175 22.625 ;
        RECT 10.850 22.125 11.255 22.295 ;
        RECT 11.425 22.125 12.210 22.295 ;
        RECT 12.485 21.845 12.695 22.375 ;
        RECT 12.955 22.060 13.285 22.585 ;
        RECT 13.795 22.500 14.175 22.585 ;
        RECT 14.345 22.615 15.995 23.135 ;
        RECT 16.165 22.785 17.855 23.305 ;
        RECT 18.485 23.230 18.775 24.395 ;
        RECT 19.035 23.725 19.205 24.225 ;
        RECT 19.375 23.895 19.705 24.395 ;
        RECT 19.035 23.555 19.700 23.725 ;
        RECT 18.950 22.735 19.300 23.385 ;
        RECT 13.455 21.845 13.625 22.455 ;
        RECT 13.795 22.065 14.125 22.500 ;
        RECT 14.345 21.845 17.855 22.615 ;
        RECT 18.485 21.845 18.775 22.570 ;
        RECT 19.470 22.565 19.700 23.555 ;
        RECT 19.035 22.395 19.700 22.565 ;
        RECT 19.035 22.105 19.205 22.395 ;
        RECT 19.375 21.845 19.705 22.225 ;
        RECT 19.875 22.105 20.060 24.225 ;
        RECT 20.300 23.935 20.565 24.395 ;
        RECT 20.735 23.800 20.985 24.225 ;
        RECT 21.195 23.950 22.300 24.120 ;
        RECT 20.680 23.670 20.985 23.800 ;
        RECT 20.230 22.475 20.510 23.425 ;
        RECT 20.680 22.565 20.850 23.670 ;
        RECT 21.020 22.885 21.260 23.480 ;
        RECT 21.430 23.415 21.960 23.780 ;
        RECT 21.430 22.715 21.600 23.415 ;
        RECT 22.130 23.335 22.300 23.950 ;
        RECT 22.470 23.595 22.640 24.395 ;
        RECT 22.810 23.895 23.060 24.225 ;
        RECT 23.285 23.925 24.170 24.095 ;
        RECT 22.130 23.245 22.640 23.335 ;
        RECT 20.680 22.435 20.905 22.565 ;
        RECT 21.075 22.495 21.600 22.715 ;
        RECT 21.770 23.075 22.640 23.245 ;
        RECT 20.315 21.845 20.565 22.305 ;
        RECT 20.735 22.295 20.905 22.435 ;
        RECT 21.770 22.295 21.940 23.075 ;
        RECT 22.470 23.005 22.640 23.075 ;
        RECT 22.150 22.825 22.350 22.855 ;
        RECT 22.810 22.825 22.980 23.895 ;
        RECT 23.150 23.005 23.340 23.725 ;
        RECT 22.150 22.525 22.980 22.825 ;
        RECT 23.510 22.795 23.830 23.755 ;
        RECT 20.735 22.125 21.070 22.295 ;
        RECT 21.265 22.125 21.940 22.295 ;
        RECT 22.260 21.845 22.630 22.345 ;
        RECT 22.810 22.295 22.980 22.525 ;
        RECT 23.365 22.465 23.830 22.795 ;
        RECT 24.000 23.085 24.170 23.925 ;
        RECT 24.350 23.895 24.665 24.395 ;
        RECT 24.895 23.665 25.235 24.225 ;
        RECT 24.340 23.290 25.235 23.665 ;
        RECT 25.405 23.385 25.575 24.395 ;
        RECT 25.045 23.085 25.235 23.290 ;
        RECT 25.745 23.335 26.075 24.180 ;
        RECT 26.395 23.775 26.565 24.205 ;
        RECT 26.735 23.945 27.065 24.395 ;
        RECT 26.395 23.545 27.075 23.775 ;
        RECT 25.745 23.255 26.135 23.335 ;
        RECT 25.920 23.205 26.135 23.255 ;
        RECT 26.365 23.205 26.670 23.375 ;
        RECT 24.000 22.755 24.875 23.085 ;
        RECT 25.045 22.755 25.795 23.085 ;
        RECT 24.000 22.295 24.170 22.755 ;
        RECT 25.045 22.585 25.245 22.755 ;
        RECT 25.965 22.625 26.135 23.205 ;
        RECT 25.910 22.585 26.135 22.625 ;
        RECT 22.810 22.125 23.215 22.295 ;
        RECT 23.385 22.125 24.170 22.295 ;
        RECT 24.445 21.845 24.655 22.375 ;
        RECT 24.915 22.060 25.245 22.585 ;
        RECT 25.755 22.500 26.135 22.585 ;
        RECT 26.370 22.525 26.670 23.205 ;
        RECT 26.840 22.895 27.075 23.545 ;
        RECT 27.265 23.235 27.550 24.180 ;
        RECT 27.730 23.925 28.415 24.395 ;
        RECT 27.725 23.405 28.420 23.715 ;
        RECT 28.595 23.340 28.900 24.125 ;
        RECT 29.085 23.440 29.355 24.395 ;
        RECT 27.265 23.085 28.125 23.235 ;
        RECT 27.265 23.065 28.555 23.085 ;
        RECT 26.840 22.565 27.395 22.895 ;
        RECT 27.565 22.705 28.555 23.065 ;
        RECT 25.415 21.845 25.585 22.455 ;
        RECT 25.755 22.065 26.085 22.500 ;
        RECT 26.840 22.415 27.055 22.565 ;
        RECT 26.315 21.845 26.645 22.350 ;
        RECT 26.815 22.040 27.055 22.415 ;
        RECT 27.565 22.370 27.735 22.705 ;
        RECT 28.725 22.535 28.900 23.340 ;
        RECT 29.525 23.305 32.115 24.395 ;
        RECT 32.860 23.765 33.145 24.225 ;
        RECT 33.315 23.935 33.585 24.395 ;
        RECT 32.860 23.545 33.815 23.765 ;
        RECT 27.335 22.175 27.735 22.370 ;
        RECT 27.335 22.030 27.505 22.175 ;
        RECT 28.095 21.845 28.495 22.340 ;
        RECT 28.665 22.015 28.900 22.535 ;
        RECT 29.525 22.615 30.735 23.135 ;
        RECT 30.905 22.785 32.115 23.305 ;
        RECT 32.745 22.815 33.435 23.375 ;
        RECT 33.605 22.645 33.815 23.545 ;
        RECT 29.085 21.845 29.355 22.480 ;
        RECT 29.525 21.845 32.115 22.615 ;
        RECT 32.860 22.475 33.815 22.645 ;
        RECT 33.985 23.375 34.385 24.225 ;
        RECT 34.575 23.765 34.855 24.225 ;
        RECT 35.375 23.935 35.700 24.395 ;
        RECT 34.575 23.545 35.700 23.765 ;
        RECT 33.985 22.815 35.080 23.375 ;
        RECT 35.250 23.085 35.700 23.545 ;
        RECT 35.870 23.255 36.255 24.225 ;
        RECT 32.860 22.015 33.145 22.475 ;
        RECT 33.315 21.845 33.585 22.305 ;
        RECT 33.985 22.015 34.385 22.815 ;
        RECT 35.250 22.755 35.805 23.085 ;
        RECT 35.250 22.645 35.700 22.755 ;
        RECT 34.575 22.475 35.700 22.645 ;
        RECT 35.975 22.585 36.255 23.255 ;
        RECT 34.575 22.015 34.855 22.475 ;
        RECT 35.375 21.845 35.700 22.305 ;
        RECT 35.870 22.015 36.255 22.585 ;
        RECT 36.425 23.595 36.865 24.225 ;
        RECT 36.425 22.585 36.735 23.595 ;
        RECT 37.040 23.545 37.355 24.395 ;
        RECT 37.525 24.055 38.955 24.225 ;
        RECT 37.525 23.375 37.695 24.055 ;
        RECT 36.905 23.205 37.695 23.375 ;
        RECT 36.905 22.755 37.075 23.205 ;
        RECT 37.865 23.085 38.065 23.885 ;
        RECT 37.245 22.755 37.635 23.035 ;
        RECT 37.820 22.755 38.065 23.085 ;
        RECT 38.265 22.755 38.515 23.885 ;
        RECT 38.705 23.425 38.955 24.055 ;
        RECT 39.135 23.595 39.465 24.395 ;
        RECT 38.705 23.255 39.475 23.425 ;
        RECT 38.730 22.755 39.135 23.085 ;
        RECT 39.305 22.585 39.475 23.255 ;
        RECT 40.105 23.305 41.315 24.395 ;
        RECT 40.105 22.765 40.625 23.305 ;
        RECT 40.795 22.595 41.315 23.135 ;
        RECT 36.425 22.025 36.865 22.585 ;
        RECT 37.035 21.845 37.485 22.585 ;
        RECT 37.655 22.415 38.815 22.585 ;
        RECT 37.655 22.015 37.825 22.415 ;
        RECT 37.995 21.845 38.415 22.245 ;
        RECT 38.585 22.015 38.815 22.415 ;
        RECT 38.985 22.015 39.475 22.585 ;
        RECT 40.105 21.845 41.315 22.595 ;
        RECT 5.520 21.675 41.400 21.845 ;
        RECT 5.605 20.925 6.815 21.675 ;
        RECT 5.605 20.385 6.125 20.925 ;
        RECT 6.990 20.835 7.250 21.675 ;
        RECT 7.425 20.930 7.680 21.505 ;
        RECT 7.850 21.295 8.180 21.675 ;
        RECT 8.395 21.125 8.565 21.505 ;
        RECT 7.850 20.955 8.565 21.125 ;
        RECT 9.860 21.045 10.145 21.505 ;
        RECT 10.315 21.215 10.585 21.675 ;
        RECT 6.295 20.215 6.815 20.755 ;
        RECT 5.605 19.125 6.815 20.215 ;
        RECT 6.990 19.125 7.250 20.275 ;
        RECT 7.425 20.200 7.595 20.930 ;
        RECT 7.850 20.765 8.020 20.955 ;
        RECT 9.860 20.875 10.815 21.045 ;
        RECT 7.765 20.435 8.020 20.765 ;
        RECT 7.850 20.225 8.020 20.435 ;
        RECT 8.300 20.405 8.655 20.775 ;
        RECT 7.425 19.295 7.680 20.200 ;
        RECT 7.850 20.055 8.565 20.225 ;
        RECT 9.745 20.145 10.435 20.705 ;
        RECT 7.850 19.125 8.180 19.885 ;
        RECT 8.395 19.295 8.565 20.055 ;
        RECT 10.605 19.975 10.815 20.875 ;
        RECT 9.860 19.755 10.815 19.975 ;
        RECT 10.985 20.705 11.385 21.505 ;
        RECT 11.575 21.045 11.855 21.505 ;
        RECT 12.375 21.215 12.700 21.675 ;
        RECT 11.575 20.875 12.700 21.045 ;
        RECT 12.870 20.935 13.255 21.505 ;
        RECT 12.250 20.765 12.700 20.875 ;
        RECT 10.985 20.145 12.080 20.705 ;
        RECT 12.250 20.435 12.805 20.765 ;
        RECT 9.860 19.295 10.145 19.755 ;
        RECT 10.315 19.125 10.585 19.585 ;
        RECT 10.985 19.295 11.385 20.145 ;
        RECT 12.250 19.975 12.700 20.435 ;
        RECT 12.975 20.265 13.255 20.935 ;
        RECT 14.460 21.045 14.745 21.505 ;
        RECT 14.915 21.215 15.185 21.675 ;
        RECT 14.460 20.875 15.415 21.045 ;
        RECT 11.575 19.755 12.700 19.975 ;
        RECT 11.575 19.295 11.855 19.755 ;
        RECT 12.375 19.125 12.700 19.585 ;
        RECT 12.870 19.295 13.255 20.265 ;
        RECT 14.345 20.145 15.035 20.705 ;
        RECT 15.205 19.975 15.415 20.875 ;
        RECT 14.460 19.755 15.415 19.975 ;
        RECT 15.585 20.705 15.985 21.505 ;
        RECT 16.175 21.045 16.455 21.505 ;
        RECT 16.975 21.215 17.300 21.675 ;
        RECT 16.175 20.875 17.300 21.045 ;
        RECT 17.470 20.935 17.855 21.505 ;
        RECT 16.850 20.765 17.300 20.875 ;
        RECT 15.585 20.145 16.680 20.705 ;
        RECT 16.850 20.435 17.405 20.765 ;
        RECT 14.460 19.295 14.745 19.755 ;
        RECT 14.915 19.125 15.185 19.585 ;
        RECT 15.585 19.295 15.985 20.145 ;
        RECT 16.850 19.975 17.300 20.435 ;
        RECT 17.575 20.265 17.855 20.935 ;
        RECT 18.300 20.865 18.545 21.470 ;
        RECT 18.765 21.140 19.275 21.675 ;
        RECT 16.175 19.755 17.300 19.975 ;
        RECT 16.175 19.295 16.455 19.755 ;
        RECT 16.975 19.125 17.300 19.585 ;
        RECT 17.470 19.295 17.855 20.265 ;
        RECT 18.025 20.695 19.255 20.865 ;
        RECT 18.025 19.885 18.365 20.695 ;
        RECT 18.535 20.130 19.285 20.320 ;
        RECT 18.025 19.475 18.540 19.885 ;
        RECT 18.775 19.125 18.945 19.885 ;
        RECT 19.115 19.465 19.285 20.130 ;
        RECT 19.455 20.145 19.645 21.505 ;
        RECT 19.815 20.655 20.090 21.505 ;
        RECT 20.280 21.140 20.810 21.505 ;
        RECT 21.235 21.275 21.565 21.675 ;
        RECT 20.635 21.105 20.810 21.140 ;
        RECT 19.815 20.485 20.095 20.655 ;
        RECT 19.815 20.345 20.090 20.485 ;
        RECT 20.295 20.145 20.465 20.945 ;
        RECT 19.455 19.975 20.465 20.145 ;
        RECT 20.635 20.935 21.565 21.105 ;
        RECT 21.735 20.935 21.990 21.505 ;
        RECT 20.635 19.805 20.805 20.935 ;
        RECT 21.395 20.765 21.565 20.935 ;
        RECT 19.680 19.635 20.805 19.805 ;
        RECT 20.975 20.435 21.170 20.765 ;
        RECT 21.395 20.435 21.650 20.765 ;
        RECT 20.975 19.465 21.145 20.435 ;
        RECT 21.820 20.265 21.990 20.935 ;
        RECT 22.165 20.905 23.835 21.675 ;
        RECT 24.095 21.125 24.265 21.415 ;
        RECT 24.435 21.295 24.765 21.675 ;
        RECT 24.095 20.955 24.760 21.125 ;
        RECT 22.165 20.385 22.915 20.905 ;
        RECT 19.115 19.295 21.145 19.465 ;
        RECT 21.315 19.125 21.485 20.265 ;
        RECT 21.655 19.295 21.990 20.265 ;
        RECT 23.085 20.215 23.835 20.735 ;
        RECT 22.165 19.125 23.835 20.215 ;
        RECT 24.010 20.135 24.360 20.785 ;
        RECT 24.530 19.965 24.760 20.955 ;
        RECT 24.095 19.795 24.760 19.965 ;
        RECT 24.095 19.295 24.265 19.795 ;
        RECT 24.435 19.125 24.765 19.625 ;
        RECT 24.935 19.295 25.120 21.415 ;
        RECT 25.375 21.215 25.625 21.675 ;
        RECT 25.795 21.225 26.130 21.395 ;
        RECT 26.325 21.225 27.000 21.395 ;
        RECT 25.795 21.085 25.965 21.225 ;
        RECT 25.290 20.095 25.570 21.045 ;
        RECT 25.740 20.955 25.965 21.085 ;
        RECT 25.740 19.850 25.910 20.955 ;
        RECT 26.135 20.805 26.660 21.025 ;
        RECT 26.080 20.040 26.320 20.635 ;
        RECT 26.490 20.105 26.660 20.805 ;
        RECT 26.830 20.445 27.000 21.225 ;
        RECT 27.320 21.175 27.690 21.675 ;
        RECT 27.870 21.225 28.275 21.395 ;
        RECT 28.445 21.225 29.230 21.395 ;
        RECT 27.870 20.995 28.040 21.225 ;
        RECT 27.210 20.695 28.040 20.995 ;
        RECT 28.425 20.725 28.890 21.055 ;
        RECT 27.210 20.665 27.410 20.695 ;
        RECT 27.530 20.445 27.700 20.515 ;
        RECT 26.830 20.275 27.700 20.445 ;
        RECT 27.190 20.185 27.700 20.275 ;
        RECT 25.740 19.720 26.045 19.850 ;
        RECT 26.490 19.740 27.020 20.105 ;
        RECT 25.360 19.125 25.625 19.585 ;
        RECT 25.795 19.295 26.045 19.720 ;
        RECT 27.190 19.570 27.360 20.185 ;
        RECT 26.255 19.400 27.360 19.570 ;
        RECT 27.530 19.125 27.700 19.925 ;
        RECT 27.870 19.625 28.040 20.695 ;
        RECT 28.210 19.795 28.400 20.515 ;
        RECT 28.570 19.765 28.890 20.725 ;
        RECT 29.060 20.765 29.230 21.225 ;
        RECT 29.505 21.145 29.715 21.675 ;
        RECT 29.975 20.935 30.305 21.460 ;
        RECT 30.475 21.065 30.645 21.675 ;
        RECT 30.815 21.020 31.145 21.455 ;
        RECT 30.815 20.935 31.195 21.020 ;
        RECT 31.365 20.950 31.655 21.675 ;
        RECT 30.105 20.765 30.305 20.935 ;
        RECT 30.970 20.895 31.195 20.935 ;
        RECT 29.060 20.435 29.935 20.765 ;
        RECT 30.105 20.435 30.855 20.765 ;
        RECT 27.870 19.295 28.120 19.625 ;
        RECT 29.060 19.595 29.230 20.435 ;
        RECT 30.105 20.230 30.295 20.435 ;
        RECT 31.025 20.315 31.195 20.895 ;
        RECT 30.980 20.265 31.195 20.315 ;
        RECT 31.830 20.935 32.085 21.505 ;
        RECT 32.255 21.275 32.585 21.675 ;
        RECT 33.010 21.140 33.540 21.505 ;
        RECT 33.730 21.335 34.005 21.505 ;
        RECT 33.725 21.165 34.005 21.335 ;
        RECT 33.010 21.105 33.185 21.140 ;
        RECT 32.255 20.935 33.185 21.105 ;
        RECT 29.400 19.855 30.295 20.230 ;
        RECT 30.805 20.185 31.195 20.265 ;
        RECT 28.345 19.425 29.230 19.595 ;
        RECT 29.410 19.125 29.725 19.625 ;
        RECT 29.955 19.295 30.295 19.855 ;
        RECT 30.465 19.125 30.635 20.135 ;
        RECT 30.805 19.340 31.135 20.185 ;
        RECT 31.365 19.125 31.655 20.290 ;
        RECT 31.830 20.265 32.000 20.935 ;
        RECT 32.255 20.765 32.425 20.935 ;
        RECT 32.170 20.435 32.425 20.765 ;
        RECT 32.650 20.435 32.845 20.765 ;
        RECT 31.830 19.295 32.165 20.265 ;
        RECT 32.335 19.125 32.505 20.265 ;
        RECT 32.675 19.465 32.845 20.435 ;
        RECT 33.015 19.805 33.185 20.935 ;
        RECT 33.355 20.145 33.525 20.945 ;
        RECT 33.730 20.345 34.005 21.165 ;
        RECT 34.175 20.145 34.365 21.505 ;
        RECT 34.545 21.140 35.055 21.675 ;
        RECT 35.275 20.865 35.520 21.470 ;
        RECT 36.055 21.125 36.225 21.505 ;
        RECT 36.405 21.295 36.735 21.675 ;
        RECT 36.055 20.955 36.720 21.125 ;
        RECT 36.915 21.000 37.175 21.505 ;
        RECT 34.565 20.695 35.795 20.865 ;
        RECT 33.355 19.975 34.365 20.145 ;
        RECT 34.535 20.130 35.285 20.320 ;
        RECT 33.015 19.635 34.140 19.805 ;
        RECT 34.535 19.465 34.705 20.130 ;
        RECT 35.455 19.885 35.795 20.695 ;
        RECT 35.985 20.405 36.315 20.775 ;
        RECT 36.550 20.700 36.720 20.955 ;
        RECT 36.550 20.370 36.835 20.700 ;
        RECT 36.550 20.225 36.720 20.370 ;
        RECT 32.675 19.295 34.705 19.465 ;
        RECT 34.875 19.125 35.045 19.885 ;
        RECT 35.280 19.475 35.795 19.885 ;
        RECT 36.055 20.055 36.720 20.225 ;
        RECT 37.005 20.200 37.175 21.000 ;
        RECT 36.055 19.295 36.225 20.055 ;
        RECT 36.405 19.125 36.735 19.885 ;
        RECT 36.905 19.295 37.175 20.200 ;
        RECT 37.345 21.000 37.615 21.345 ;
        RECT 37.805 21.275 38.185 21.675 ;
        RECT 38.355 21.105 38.525 21.455 ;
        RECT 38.695 21.275 39.025 21.675 ;
        RECT 39.225 21.105 39.395 21.455 ;
        RECT 39.595 21.175 39.925 21.675 ;
        RECT 37.345 20.265 37.515 21.000 ;
        RECT 37.785 20.935 39.395 21.105 ;
        RECT 37.785 20.765 37.955 20.935 ;
        RECT 37.685 20.435 37.955 20.765 ;
        RECT 38.125 20.435 38.530 20.765 ;
        RECT 37.785 20.265 37.955 20.435 ;
        RECT 37.345 19.295 37.615 20.265 ;
        RECT 37.785 20.095 38.510 20.265 ;
        RECT 38.700 20.145 39.410 20.765 ;
        RECT 39.580 20.435 39.930 21.005 ;
        RECT 40.105 20.925 41.315 21.675 ;
        RECT 38.340 19.975 38.510 20.095 ;
        RECT 39.610 19.975 39.930 20.265 ;
        RECT 37.825 19.125 38.105 19.925 ;
        RECT 38.340 19.805 39.930 19.975 ;
        RECT 40.105 20.215 40.625 20.755 ;
        RECT 40.795 20.385 41.315 20.925 ;
        RECT 38.275 19.345 39.930 19.635 ;
        RECT 40.105 19.125 41.315 20.215 ;
        RECT 5.520 18.955 41.400 19.125 ;
        RECT 5.605 17.865 6.815 18.955 ;
        RECT 7.045 17.895 7.375 18.740 ;
        RECT 7.545 17.945 7.715 18.955 ;
        RECT 7.885 18.225 8.225 18.785 ;
        RECT 8.455 18.455 8.770 18.955 ;
        RECT 8.950 18.485 9.835 18.655 ;
        RECT 5.605 17.155 6.125 17.695 ;
        RECT 6.295 17.325 6.815 17.865 ;
        RECT 6.985 17.815 7.375 17.895 ;
        RECT 7.885 17.850 8.780 18.225 ;
        RECT 6.985 17.765 7.200 17.815 ;
        RECT 6.985 17.185 7.155 17.765 ;
        RECT 7.885 17.645 8.075 17.850 ;
        RECT 8.950 17.645 9.120 18.485 ;
        RECT 10.060 18.455 10.310 18.785 ;
        RECT 7.325 17.315 8.075 17.645 ;
        RECT 8.245 17.315 9.120 17.645 ;
        RECT 5.605 16.405 6.815 17.155 ;
        RECT 6.985 17.145 7.210 17.185 ;
        RECT 7.875 17.145 8.075 17.315 ;
        RECT 6.985 17.060 7.365 17.145 ;
        RECT 7.035 16.625 7.365 17.060 ;
        RECT 7.535 16.405 7.705 17.015 ;
        RECT 7.875 16.620 8.205 17.145 ;
        RECT 8.465 16.405 8.675 16.935 ;
        RECT 8.950 16.855 9.120 17.315 ;
        RECT 9.290 17.355 9.610 18.315 ;
        RECT 9.780 17.565 9.970 18.285 ;
        RECT 10.140 17.385 10.310 18.455 ;
        RECT 10.480 18.155 10.650 18.955 ;
        RECT 10.820 18.510 11.925 18.680 ;
        RECT 10.820 17.895 10.990 18.510 ;
        RECT 12.135 18.360 12.385 18.785 ;
        RECT 12.555 18.495 12.820 18.955 ;
        RECT 11.160 17.975 11.690 18.340 ;
        RECT 12.135 18.230 12.440 18.360 ;
        RECT 10.480 17.805 10.990 17.895 ;
        RECT 10.480 17.635 11.350 17.805 ;
        RECT 10.480 17.565 10.650 17.635 ;
        RECT 10.770 17.385 10.970 17.415 ;
        RECT 9.290 17.025 9.755 17.355 ;
        RECT 10.140 17.085 10.970 17.385 ;
        RECT 10.140 16.855 10.310 17.085 ;
        RECT 8.950 16.685 9.735 16.855 ;
        RECT 9.905 16.685 10.310 16.855 ;
        RECT 10.490 16.405 10.860 16.905 ;
        RECT 11.180 16.855 11.350 17.635 ;
        RECT 11.520 17.275 11.690 17.975 ;
        RECT 11.860 17.445 12.100 18.040 ;
        RECT 11.520 17.055 12.045 17.275 ;
        RECT 12.270 17.125 12.440 18.230 ;
        RECT 12.215 16.995 12.440 17.125 ;
        RECT 12.610 17.035 12.890 17.985 ;
        RECT 12.215 16.855 12.385 16.995 ;
        RECT 11.180 16.685 11.855 16.855 ;
        RECT 12.050 16.685 12.385 16.855 ;
        RECT 12.555 16.405 12.805 16.865 ;
        RECT 13.060 16.665 13.245 18.785 ;
        RECT 13.415 18.455 13.745 18.955 ;
        RECT 13.915 18.285 14.085 18.785 ;
        RECT 13.420 18.115 14.085 18.285 ;
        RECT 13.420 17.125 13.650 18.115 ;
        RECT 13.820 17.295 14.170 17.945 ;
        RECT 14.345 17.865 17.855 18.955 ;
        RECT 14.345 17.175 15.995 17.695 ;
        RECT 16.165 17.345 17.855 17.865 ;
        RECT 18.485 17.790 18.775 18.955 ;
        RECT 18.955 18.145 19.250 18.955 ;
        RECT 19.430 17.645 19.675 18.785 ;
        RECT 19.850 18.145 20.110 18.955 ;
        RECT 20.710 18.950 26.985 18.955 ;
        RECT 20.290 17.645 20.540 18.780 ;
        RECT 20.710 18.155 20.970 18.950 ;
        RECT 21.140 18.055 21.400 18.780 ;
        RECT 21.570 18.225 21.830 18.950 ;
        RECT 22.000 18.055 22.260 18.780 ;
        RECT 22.430 18.225 22.690 18.950 ;
        RECT 22.860 18.055 23.120 18.780 ;
        RECT 23.290 18.225 23.550 18.950 ;
        RECT 23.720 18.055 23.980 18.780 ;
        RECT 24.150 18.225 24.395 18.950 ;
        RECT 24.565 18.055 24.825 18.780 ;
        RECT 25.010 18.225 25.255 18.950 ;
        RECT 25.425 18.055 25.685 18.780 ;
        RECT 25.870 18.225 26.115 18.950 ;
        RECT 26.285 18.055 26.545 18.780 ;
        RECT 26.730 18.225 26.985 18.950 ;
        RECT 21.140 18.040 26.545 18.055 ;
        RECT 27.155 18.040 27.445 18.780 ;
        RECT 27.615 18.210 27.885 18.955 ;
        RECT 21.140 17.815 27.885 18.040 ;
        RECT 28.145 17.865 29.355 18.955 ;
        RECT 13.420 16.955 14.085 17.125 ;
        RECT 13.415 16.405 13.745 16.785 ;
        RECT 13.915 16.665 14.085 16.955 ;
        RECT 14.345 16.405 17.855 17.175 ;
        RECT 18.485 16.405 18.775 17.130 ;
        RECT 18.945 17.085 19.260 17.645 ;
        RECT 19.430 17.395 26.550 17.645 ;
        RECT 18.945 16.405 19.250 16.915 ;
        RECT 19.430 16.585 19.680 17.395 ;
        RECT 19.850 16.405 20.110 16.930 ;
        RECT 20.290 16.585 20.540 17.395 ;
        RECT 26.720 17.225 27.885 17.815 ;
        RECT 21.140 17.055 27.885 17.225 ;
        RECT 28.145 17.155 28.665 17.695 ;
        RECT 28.835 17.325 29.355 17.865 ;
        RECT 29.615 18.025 29.785 18.785 ;
        RECT 29.965 18.195 30.295 18.955 ;
        RECT 29.615 17.855 30.280 18.025 ;
        RECT 30.465 17.880 30.735 18.785 ;
        RECT 30.110 17.710 30.280 17.855 ;
        RECT 29.545 17.305 29.875 17.675 ;
        RECT 30.110 17.380 30.395 17.710 ;
        RECT 20.710 16.405 20.970 16.965 ;
        RECT 21.140 16.600 21.400 17.055 ;
        RECT 21.570 16.405 21.830 16.885 ;
        RECT 22.000 16.600 22.260 17.055 ;
        RECT 22.430 16.405 22.690 16.885 ;
        RECT 22.860 16.600 23.120 17.055 ;
        RECT 23.290 16.405 23.535 16.885 ;
        RECT 23.705 16.600 23.980 17.055 ;
        RECT 24.150 16.405 24.395 16.885 ;
        RECT 24.565 16.600 24.825 17.055 ;
        RECT 25.005 16.405 25.255 16.885 ;
        RECT 25.425 16.600 25.685 17.055 ;
        RECT 25.865 16.405 26.115 16.885 ;
        RECT 26.285 16.600 26.545 17.055 ;
        RECT 26.725 16.405 26.985 16.885 ;
        RECT 27.155 16.600 27.415 17.055 ;
        RECT 27.585 16.405 27.885 16.885 ;
        RECT 28.145 16.405 29.355 17.155 ;
        RECT 30.110 17.125 30.280 17.380 ;
        RECT 29.615 16.955 30.280 17.125 ;
        RECT 30.565 17.080 30.735 17.880 ;
        RECT 30.995 18.025 31.165 18.785 ;
        RECT 31.345 18.195 31.675 18.955 ;
        RECT 30.995 17.855 31.660 18.025 ;
        RECT 31.845 17.880 32.115 18.785 ;
        RECT 31.490 17.710 31.660 17.855 ;
        RECT 30.925 17.305 31.255 17.675 ;
        RECT 31.490 17.380 31.775 17.710 ;
        RECT 31.490 17.125 31.660 17.380 ;
        RECT 29.615 16.575 29.785 16.955 ;
        RECT 29.965 16.405 30.295 16.785 ;
        RECT 30.475 16.575 30.735 17.080 ;
        RECT 30.995 16.955 31.660 17.125 ;
        RECT 31.945 17.080 32.115 17.880 ;
        RECT 32.375 18.025 32.545 18.785 ;
        RECT 32.725 18.195 33.055 18.955 ;
        RECT 32.375 17.855 33.040 18.025 ;
        RECT 33.225 17.880 33.495 18.785 ;
        RECT 32.870 17.710 33.040 17.855 ;
        RECT 32.305 17.305 32.635 17.675 ;
        RECT 32.870 17.380 33.155 17.710 ;
        RECT 32.870 17.125 33.040 17.380 ;
        RECT 30.995 16.575 31.165 16.955 ;
        RECT 31.345 16.405 31.675 16.785 ;
        RECT 31.855 16.575 32.115 17.080 ;
        RECT 32.375 16.955 33.040 17.125 ;
        RECT 33.325 17.080 33.495 17.880 ;
        RECT 33.755 18.025 33.925 18.785 ;
        RECT 34.105 18.195 34.435 18.955 ;
        RECT 33.755 17.855 34.420 18.025 ;
        RECT 34.605 17.880 34.875 18.785 ;
        RECT 34.250 17.710 34.420 17.855 ;
        RECT 33.685 17.305 34.015 17.675 ;
        RECT 34.250 17.380 34.535 17.710 ;
        RECT 34.250 17.125 34.420 17.380 ;
        RECT 32.375 16.575 32.545 16.955 ;
        RECT 32.725 16.405 33.055 16.785 ;
        RECT 33.235 16.575 33.495 17.080 ;
        RECT 33.755 16.955 34.420 17.125 ;
        RECT 34.705 17.080 34.875 17.880 ;
        RECT 35.055 17.815 35.385 18.955 ;
        RECT 35.915 17.985 36.245 18.770 ;
        RECT 35.565 17.815 36.245 17.985 ;
        RECT 35.045 17.395 35.395 17.645 ;
        RECT 35.565 17.215 35.735 17.815 ;
        RECT 36.425 17.800 36.765 18.785 ;
        RECT 36.935 18.525 37.345 18.955 ;
        RECT 38.090 18.535 38.420 18.955 ;
        RECT 38.590 18.355 38.915 18.785 ;
        RECT 36.935 18.185 38.915 18.355 ;
        RECT 35.905 17.395 36.255 17.645 ;
        RECT 33.755 16.575 33.925 16.955 ;
        RECT 34.105 16.405 34.435 16.785 ;
        RECT 34.615 16.575 34.875 17.080 ;
        RECT 35.055 16.405 35.325 17.215 ;
        RECT 35.495 16.575 35.825 17.215 ;
        RECT 35.995 16.405 36.235 17.215 ;
        RECT 36.425 17.145 36.680 17.800 ;
        RECT 36.935 17.645 37.200 18.185 ;
        RECT 37.415 17.845 38.040 18.015 ;
        RECT 36.850 17.315 37.200 17.645 ;
        RECT 37.370 17.315 37.700 17.645 ;
        RECT 37.870 17.145 38.040 17.845 ;
        RECT 36.425 16.770 36.785 17.145 ;
        RECT 37.050 16.405 37.220 17.145 ;
        RECT 37.500 16.975 38.040 17.145 ;
        RECT 38.210 17.775 38.915 18.185 ;
        RECT 39.390 17.855 39.720 18.955 ;
        RECT 40.105 17.865 41.315 18.955 ;
        RECT 37.500 16.770 37.670 16.975 ;
        RECT 38.210 16.575 38.380 17.775 ;
        RECT 38.550 17.395 39.120 17.605 ;
        RECT 39.290 17.395 39.935 17.605 ;
        RECT 40.105 17.325 40.625 17.865 ;
        RECT 38.610 17.055 39.780 17.225 ;
        RECT 40.795 17.155 41.315 17.695 ;
        RECT 38.610 16.575 38.940 17.055 ;
        RECT 39.110 16.405 39.280 16.875 ;
        RECT 39.450 16.590 39.780 17.055 ;
        RECT 40.105 16.405 41.315 17.155 ;
        RECT 5.520 16.235 41.400 16.405 ;
        RECT 5.605 15.485 6.815 16.235 ;
        RECT 5.605 14.945 6.125 15.485 ;
        RECT 6.990 15.395 7.250 16.235 ;
        RECT 7.425 15.490 7.680 16.065 ;
        RECT 7.850 15.855 8.180 16.235 ;
        RECT 8.395 15.685 8.565 16.065 ;
        RECT 7.850 15.515 8.565 15.685 ;
        RECT 6.295 14.775 6.815 15.315 ;
        RECT 5.605 13.685 6.815 14.775 ;
        RECT 6.990 13.685 7.250 14.835 ;
        RECT 7.425 14.760 7.595 15.490 ;
        RECT 7.850 15.325 8.020 15.515 ;
        RECT 9.750 15.495 10.005 16.065 ;
        RECT 10.175 15.835 10.505 16.235 ;
        RECT 10.930 15.700 11.460 16.065 ;
        RECT 11.650 15.895 11.925 16.065 ;
        RECT 11.645 15.725 11.925 15.895 ;
        RECT 10.930 15.665 11.105 15.700 ;
        RECT 10.175 15.495 11.105 15.665 ;
        RECT 7.765 14.995 8.020 15.325 ;
        RECT 7.850 14.785 8.020 14.995 ;
        RECT 8.300 14.965 8.655 15.335 ;
        RECT 9.750 14.825 9.920 15.495 ;
        RECT 10.175 15.325 10.345 15.495 ;
        RECT 10.090 14.995 10.345 15.325 ;
        RECT 10.570 14.995 10.765 15.325 ;
        RECT 7.425 13.855 7.680 14.760 ;
        RECT 7.850 14.615 8.565 14.785 ;
        RECT 7.850 13.685 8.180 14.445 ;
        RECT 8.395 13.855 8.565 14.615 ;
        RECT 9.750 13.855 10.085 14.825 ;
        RECT 10.255 13.685 10.425 14.825 ;
        RECT 10.595 14.025 10.765 14.995 ;
        RECT 10.935 14.365 11.105 15.495 ;
        RECT 11.275 14.705 11.445 15.505 ;
        RECT 11.650 14.905 11.925 15.725 ;
        RECT 12.095 14.705 12.285 16.065 ;
        RECT 12.465 15.700 12.975 16.235 ;
        RECT 13.195 15.425 13.440 16.030 ;
        RECT 13.885 15.465 17.395 16.235 ;
        RECT 17.565 15.485 18.775 16.235 ;
        RECT 18.995 15.580 19.325 16.015 ;
        RECT 19.495 15.625 19.665 16.235 ;
        RECT 18.945 15.495 19.325 15.580 ;
        RECT 19.835 15.495 20.165 16.020 ;
        RECT 20.425 15.705 20.635 16.235 ;
        RECT 20.910 15.785 21.695 15.955 ;
        RECT 21.865 15.785 22.270 15.955 ;
        RECT 12.485 15.255 13.715 15.425 ;
        RECT 11.275 14.535 12.285 14.705 ;
        RECT 12.455 14.690 13.205 14.880 ;
        RECT 10.935 14.195 12.060 14.365 ;
        RECT 12.455 14.025 12.625 14.690 ;
        RECT 13.375 14.445 13.715 15.255 ;
        RECT 13.885 14.945 15.535 15.465 ;
        RECT 15.705 14.775 17.395 15.295 ;
        RECT 17.565 14.945 18.085 15.485 ;
        RECT 18.945 15.455 19.170 15.495 ;
        RECT 18.255 14.775 18.775 15.315 ;
        RECT 10.595 13.855 12.625 14.025 ;
        RECT 12.795 13.685 12.965 14.445 ;
        RECT 13.200 14.035 13.715 14.445 ;
        RECT 13.885 13.685 17.395 14.775 ;
        RECT 17.565 13.685 18.775 14.775 ;
        RECT 18.945 14.875 19.115 15.455 ;
        RECT 19.835 15.325 20.035 15.495 ;
        RECT 20.910 15.325 21.080 15.785 ;
        RECT 19.285 14.995 20.035 15.325 ;
        RECT 20.205 14.995 21.080 15.325 ;
        RECT 18.945 14.825 19.160 14.875 ;
        RECT 18.945 14.745 19.335 14.825 ;
        RECT 19.005 13.900 19.335 14.745 ;
        RECT 19.845 14.790 20.035 14.995 ;
        RECT 19.505 13.685 19.675 14.695 ;
        RECT 19.845 14.415 20.740 14.790 ;
        RECT 19.845 13.855 20.185 14.415 ;
        RECT 20.415 13.685 20.730 14.185 ;
        RECT 20.910 14.155 21.080 14.995 ;
        RECT 21.250 15.285 21.715 15.615 ;
        RECT 22.100 15.555 22.270 15.785 ;
        RECT 22.450 15.735 22.820 16.235 ;
        RECT 23.140 15.785 23.815 15.955 ;
        RECT 24.010 15.785 24.345 15.955 ;
        RECT 21.250 14.325 21.570 15.285 ;
        RECT 22.100 15.255 22.930 15.555 ;
        RECT 21.740 14.355 21.930 15.075 ;
        RECT 22.100 14.185 22.270 15.255 ;
        RECT 22.730 15.225 22.930 15.255 ;
        RECT 22.440 15.005 22.610 15.075 ;
        RECT 23.140 15.005 23.310 15.785 ;
        RECT 24.175 15.645 24.345 15.785 ;
        RECT 24.515 15.775 24.765 16.235 ;
        RECT 22.440 14.835 23.310 15.005 ;
        RECT 23.480 15.365 24.005 15.585 ;
        RECT 24.175 15.515 24.400 15.645 ;
        RECT 22.440 14.745 22.950 14.835 ;
        RECT 20.910 13.985 21.795 14.155 ;
        RECT 22.020 13.855 22.270 14.185 ;
        RECT 22.440 13.685 22.610 14.485 ;
        RECT 22.780 14.130 22.950 14.745 ;
        RECT 23.480 14.665 23.650 15.365 ;
        RECT 23.120 14.300 23.650 14.665 ;
        RECT 23.820 14.600 24.060 15.195 ;
        RECT 24.230 14.410 24.400 15.515 ;
        RECT 24.570 14.655 24.850 15.605 ;
        RECT 24.095 14.280 24.400 14.410 ;
        RECT 22.780 13.960 23.885 14.130 ;
        RECT 24.095 13.855 24.345 14.280 ;
        RECT 24.515 13.685 24.780 14.145 ;
        RECT 25.020 13.855 25.205 15.975 ;
        RECT 25.375 15.855 25.705 16.235 ;
        RECT 25.875 15.685 26.045 15.975 ;
        RECT 25.380 15.515 26.045 15.685 ;
        RECT 25.380 14.525 25.610 15.515 ;
        RECT 26.310 15.495 26.565 16.065 ;
        RECT 26.735 15.835 27.065 16.235 ;
        RECT 27.490 15.700 28.020 16.065 ;
        RECT 27.490 15.665 27.665 15.700 ;
        RECT 26.735 15.495 27.665 15.665 ;
        RECT 25.780 14.695 26.130 15.345 ;
        RECT 26.310 14.825 26.480 15.495 ;
        RECT 26.735 15.325 26.905 15.495 ;
        RECT 26.650 14.995 26.905 15.325 ;
        RECT 27.130 14.995 27.325 15.325 ;
        RECT 25.380 14.355 26.045 14.525 ;
        RECT 25.375 13.685 25.705 14.185 ;
        RECT 25.875 13.855 26.045 14.355 ;
        RECT 26.310 13.855 26.645 14.825 ;
        RECT 26.815 13.685 26.985 14.825 ;
        RECT 27.155 14.025 27.325 14.995 ;
        RECT 27.495 14.365 27.665 15.495 ;
        RECT 27.835 14.705 28.005 15.505 ;
        RECT 28.210 15.215 28.485 16.065 ;
        RECT 28.205 15.045 28.485 15.215 ;
        RECT 28.210 14.905 28.485 15.045 ;
        RECT 28.655 14.705 28.845 16.065 ;
        RECT 29.025 15.700 29.535 16.235 ;
        RECT 29.755 15.425 30.000 16.030 ;
        RECT 31.365 15.510 31.655 16.235 ;
        RECT 31.825 15.495 32.210 16.065 ;
        RECT 32.380 15.775 32.705 16.235 ;
        RECT 33.225 15.605 33.505 16.065 ;
        RECT 29.045 15.255 30.275 15.425 ;
        RECT 27.835 14.535 28.845 14.705 ;
        RECT 29.015 14.690 29.765 14.880 ;
        RECT 27.495 14.195 28.620 14.365 ;
        RECT 29.015 14.025 29.185 14.690 ;
        RECT 29.935 14.445 30.275 15.255 ;
        RECT 27.155 13.855 29.185 14.025 ;
        RECT 29.355 13.685 29.525 14.445 ;
        RECT 29.760 14.035 30.275 14.445 ;
        RECT 31.365 13.685 31.655 14.850 ;
        RECT 31.825 14.825 32.105 15.495 ;
        RECT 32.380 15.435 33.505 15.605 ;
        RECT 32.380 15.325 32.830 15.435 ;
        RECT 32.275 14.995 32.830 15.325 ;
        RECT 33.695 15.265 34.095 16.065 ;
        RECT 34.495 15.775 34.765 16.235 ;
        RECT 34.935 15.605 35.220 16.065 ;
        RECT 31.825 13.855 32.210 14.825 ;
        RECT 32.380 14.535 32.830 14.995 ;
        RECT 33.000 14.705 34.095 15.265 ;
        RECT 32.380 14.315 33.505 14.535 ;
        RECT 32.380 13.685 32.705 14.145 ;
        RECT 33.225 13.855 33.505 14.315 ;
        RECT 33.695 13.855 34.095 14.705 ;
        RECT 34.265 15.435 35.220 15.605 ;
        RECT 36.425 15.605 36.765 16.065 ;
        RECT 36.935 15.775 37.105 16.235 ;
        RECT 37.735 15.800 38.095 16.065 ;
        RECT 37.740 15.795 38.095 15.800 ;
        RECT 37.745 15.785 38.095 15.795 ;
        RECT 37.750 15.780 38.095 15.785 ;
        RECT 37.755 15.770 38.095 15.780 ;
        RECT 38.335 15.775 38.505 16.235 ;
        RECT 37.760 15.765 38.095 15.770 ;
        RECT 37.770 15.755 38.095 15.765 ;
        RECT 37.780 15.745 38.095 15.755 ;
        RECT 37.275 15.605 37.605 15.685 ;
        RECT 34.265 14.535 34.475 15.435 ;
        RECT 36.425 15.415 37.605 15.605 ;
        RECT 37.795 15.605 38.095 15.745 ;
        RECT 37.795 15.415 38.505 15.605 ;
        RECT 34.645 14.705 35.335 15.265 ;
        RECT 36.425 15.045 36.755 15.245 ;
        RECT 37.065 15.225 37.395 15.245 ;
        RECT 36.945 15.045 37.395 15.225 ;
        RECT 36.425 14.705 36.655 15.045 ;
        RECT 34.265 14.315 35.220 14.535 ;
        RECT 34.495 13.685 34.765 14.145 ;
        RECT 34.935 13.855 35.220 14.315 ;
        RECT 36.435 13.685 36.765 14.405 ;
        RECT 36.945 13.930 37.160 15.045 ;
        RECT 37.565 15.015 38.035 15.245 ;
        RECT 38.220 14.845 38.505 15.415 ;
        RECT 38.675 15.290 39.015 16.065 ;
        RECT 40.105 15.485 41.315 16.235 ;
        RECT 37.355 14.630 38.505 14.845 ;
        RECT 37.355 13.855 37.685 14.630 ;
        RECT 37.855 13.685 38.565 14.460 ;
        RECT 38.735 13.855 39.015 15.290 ;
        RECT 40.105 14.775 40.625 15.315 ;
        RECT 40.795 14.945 41.315 15.485 ;
        RECT 40.105 13.685 41.315 14.775 ;
        RECT 5.520 13.515 41.400 13.685 ;
        RECT 5.605 12.425 6.815 13.515 ;
        RECT 6.985 13.080 12.330 13.515 ;
        RECT 5.605 11.715 6.125 12.255 ;
        RECT 6.295 11.885 6.815 12.425 ;
        RECT 5.605 10.965 6.815 11.715 ;
        RECT 8.570 11.510 8.910 12.340 ;
        RECT 10.390 11.830 10.740 13.080 ;
        RECT 12.505 12.425 16.015 13.515 ;
        RECT 12.505 11.735 14.155 12.255 ;
        RECT 14.325 11.905 16.015 12.425 ;
        RECT 16.735 12.585 16.905 13.345 ;
        RECT 17.120 12.755 17.450 13.515 ;
        RECT 16.735 12.415 17.450 12.585 ;
        RECT 17.620 12.440 17.875 13.345 ;
        RECT 16.645 11.865 17.000 12.235 ;
        RECT 17.280 12.205 17.450 12.415 ;
        RECT 17.280 11.875 17.535 12.205 ;
        RECT 6.985 10.965 12.330 11.510 ;
        RECT 12.505 10.965 16.015 11.735 ;
        RECT 17.280 11.685 17.450 11.875 ;
        RECT 17.705 11.710 17.875 12.440 ;
        RECT 18.050 12.365 18.310 13.515 ;
        RECT 18.485 12.350 18.775 13.515 ;
        RECT 19.410 12.365 19.670 13.515 ;
        RECT 19.845 12.440 20.100 13.345 ;
        RECT 20.270 12.755 20.600 13.515 ;
        RECT 20.815 12.585 20.985 13.345 ;
        RECT 21.335 12.845 21.505 13.345 ;
        RECT 21.675 13.015 22.005 13.515 ;
        RECT 21.335 12.675 22.000 12.845 ;
        RECT 16.735 11.515 17.450 11.685 ;
        RECT 16.735 11.135 16.905 11.515 ;
        RECT 17.120 10.965 17.450 11.345 ;
        RECT 17.620 11.135 17.875 11.710 ;
        RECT 18.050 10.965 18.310 11.805 ;
        RECT 18.485 10.965 18.775 11.690 ;
        RECT 19.410 10.965 19.670 11.805 ;
        RECT 19.845 11.710 20.015 12.440 ;
        RECT 20.270 12.415 20.985 12.585 ;
        RECT 20.270 12.205 20.440 12.415 ;
        RECT 20.185 11.875 20.440 12.205 ;
        RECT 19.845 11.135 20.100 11.710 ;
        RECT 20.270 11.685 20.440 11.875 ;
        RECT 20.720 11.865 21.075 12.235 ;
        RECT 21.250 11.855 21.600 12.505 ;
        RECT 21.770 11.685 22.000 12.675 ;
        RECT 20.270 11.515 20.985 11.685 ;
        RECT 20.270 10.965 20.600 11.345 ;
        RECT 20.815 11.135 20.985 11.515 ;
        RECT 21.335 11.515 22.000 11.685 ;
        RECT 21.335 11.225 21.505 11.515 ;
        RECT 21.675 10.965 22.005 11.345 ;
        RECT 22.175 11.225 22.360 13.345 ;
        RECT 22.600 13.055 22.865 13.515 ;
        RECT 23.035 12.920 23.285 13.345 ;
        RECT 23.495 13.070 24.600 13.240 ;
        RECT 22.980 12.790 23.285 12.920 ;
        RECT 22.530 11.595 22.810 12.545 ;
        RECT 22.980 11.685 23.150 12.790 ;
        RECT 23.320 12.005 23.560 12.600 ;
        RECT 23.730 12.535 24.260 12.900 ;
        RECT 23.730 11.835 23.900 12.535 ;
        RECT 24.430 12.455 24.600 13.070 ;
        RECT 24.770 12.715 24.940 13.515 ;
        RECT 25.110 13.015 25.360 13.345 ;
        RECT 25.585 13.045 26.470 13.215 ;
        RECT 24.430 12.365 24.940 12.455 ;
        RECT 22.980 11.555 23.205 11.685 ;
        RECT 23.375 11.615 23.900 11.835 ;
        RECT 24.070 12.195 24.940 12.365 ;
        RECT 22.615 10.965 22.865 11.425 ;
        RECT 23.035 11.415 23.205 11.555 ;
        RECT 24.070 11.415 24.240 12.195 ;
        RECT 24.770 12.125 24.940 12.195 ;
        RECT 24.450 11.945 24.650 11.975 ;
        RECT 25.110 11.945 25.280 13.015 ;
        RECT 25.450 12.125 25.640 12.845 ;
        RECT 24.450 11.645 25.280 11.945 ;
        RECT 25.810 11.915 26.130 12.875 ;
        RECT 23.035 11.245 23.370 11.415 ;
        RECT 23.565 11.245 24.240 11.415 ;
        RECT 24.560 10.965 24.930 11.465 ;
        RECT 25.110 11.415 25.280 11.645 ;
        RECT 25.665 11.585 26.130 11.915 ;
        RECT 26.300 12.205 26.470 13.045 ;
        RECT 26.650 13.015 26.965 13.515 ;
        RECT 27.195 12.785 27.535 13.345 ;
        RECT 26.640 12.410 27.535 12.785 ;
        RECT 27.705 12.505 27.875 13.515 ;
        RECT 27.345 12.205 27.535 12.410 ;
        RECT 28.045 12.455 28.375 13.300 ;
        RECT 28.045 12.375 28.435 12.455 ;
        RECT 28.220 12.325 28.435 12.375 ;
        RECT 28.610 12.365 28.870 13.515 ;
        RECT 29.045 12.440 29.300 13.345 ;
        RECT 29.470 12.755 29.800 13.515 ;
        RECT 30.015 12.585 30.185 13.345 ;
        RECT 26.300 11.875 27.175 12.205 ;
        RECT 27.345 11.875 28.095 12.205 ;
        RECT 26.300 11.415 26.470 11.875 ;
        RECT 27.345 11.705 27.545 11.875 ;
        RECT 28.265 11.745 28.435 12.325 ;
        RECT 28.210 11.705 28.435 11.745 ;
        RECT 25.110 11.245 25.515 11.415 ;
        RECT 25.685 11.245 26.470 11.415 ;
        RECT 26.745 10.965 26.955 11.495 ;
        RECT 27.215 11.180 27.545 11.705 ;
        RECT 28.055 11.620 28.435 11.705 ;
        RECT 27.715 10.965 27.885 11.575 ;
        RECT 28.055 11.185 28.385 11.620 ;
        RECT 28.610 10.965 28.870 11.805 ;
        RECT 29.045 11.710 29.215 12.440 ;
        RECT 29.470 12.415 30.185 12.585 ;
        RECT 29.470 12.205 29.640 12.415 ;
        RECT 31.365 12.350 31.655 13.515 ;
        RECT 32.835 12.585 33.005 13.345 ;
        RECT 33.220 12.755 33.550 13.515 ;
        RECT 32.835 12.415 33.550 12.585 ;
        RECT 33.720 12.440 33.975 13.345 ;
        RECT 29.385 11.875 29.640 12.205 ;
        RECT 29.045 11.135 29.300 11.710 ;
        RECT 29.470 11.685 29.640 11.875 ;
        RECT 29.920 11.865 30.275 12.235 ;
        RECT 32.745 11.865 33.100 12.235 ;
        RECT 33.380 12.205 33.550 12.415 ;
        RECT 33.380 11.875 33.635 12.205 ;
        RECT 29.470 11.515 30.185 11.685 ;
        RECT 29.470 10.965 29.800 11.345 ;
        RECT 30.015 11.135 30.185 11.515 ;
        RECT 31.365 10.965 31.655 11.690 ;
        RECT 33.380 11.685 33.550 11.875 ;
        RECT 33.805 11.710 33.975 12.440 ;
        RECT 34.150 12.365 34.410 13.515 ;
        RECT 34.585 12.440 34.855 13.345 ;
        RECT 35.025 12.755 35.355 13.515 ;
        RECT 35.535 12.585 35.715 13.345 ;
        RECT 36.975 12.895 37.145 13.325 ;
        RECT 37.315 13.065 37.645 13.515 ;
        RECT 36.975 12.665 37.650 12.895 ;
        RECT 32.835 11.515 33.550 11.685 ;
        RECT 32.835 11.135 33.005 11.515 ;
        RECT 33.220 10.965 33.550 11.345 ;
        RECT 33.720 11.135 33.975 11.710 ;
        RECT 34.150 10.965 34.410 11.805 ;
        RECT 34.585 11.640 34.765 12.440 ;
        RECT 35.040 12.415 35.715 12.585 ;
        RECT 35.040 12.270 35.210 12.415 ;
        RECT 34.935 11.940 35.210 12.270 ;
        RECT 35.040 11.685 35.210 11.940 ;
        RECT 35.435 11.865 35.775 12.235 ;
        RECT 34.585 11.135 34.845 11.640 ;
        RECT 35.040 11.515 35.705 11.685 ;
        RECT 36.945 11.645 37.245 12.495 ;
        RECT 37.415 12.015 37.650 12.665 ;
        RECT 37.820 12.355 38.105 13.300 ;
        RECT 38.285 13.045 38.970 13.515 ;
        RECT 38.280 12.525 38.975 12.835 ;
        RECT 39.150 12.460 39.455 13.245 ;
        RECT 37.820 12.205 38.680 12.355 ;
        RECT 37.820 12.185 39.105 12.205 ;
        RECT 37.415 11.685 37.950 12.015 ;
        RECT 38.120 11.825 39.105 12.185 ;
        RECT 37.415 11.535 37.635 11.685 ;
        RECT 35.025 10.965 35.355 11.345 ;
        RECT 35.535 11.135 35.705 11.515 ;
        RECT 36.890 10.965 37.225 11.470 ;
        RECT 37.395 11.160 37.635 11.535 ;
        RECT 38.120 11.490 38.290 11.825 ;
        RECT 39.280 11.655 39.455 12.460 ;
        RECT 40.105 12.425 41.315 13.515 ;
        RECT 40.105 11.885 40.625 12.425 ;
        RECT 40.795 11.715 41.315 12.255 ;
        RECT 37.915 11.295 38.290 11.490 ;
        RECT 37.915 11.150 38.085 11.295 ;
        RECT 38.650 10.965 39.045 11.460 ;
        RECT 39.215 11.135 39.455 11.655 ;
        RECT 40.105 10.965 41.315 11.715 ;
        RECT 5.520 10.795 41.400 10.965 ;
      LAYER met1 ;
        RECT 5.520 46.000 41.400 46.480 ;
        RECT 14.345 45.800 14.635 45.845 ;
        RECT 19.390 45.800 19.710 45.860 ;
        RECT 14.345 45.660 19.710 45.800 ;
        RECT 14.345 45.615 14.635 45.660 ;
        RECT 19.390 45.600 19.710 45.660 ;
        RECT 24.925 45.800 25.215 45.845 ;
        RECT 25.830 45.800 26.150 45.860 ;
        RECT 24.925 45.660 26.150 45.800 ;
        RECT 24.925 45.615 25.215 45.660 ;
        RECT 25.830 45.600 26.150 45.660 ;
        RECT 32.270 45.800 32.590 45.860 ;
        RECT 33.205 45.800 33.495 45.845 ;
        RECT 32.270 45.660 33.495 45.800 ;
        RECT 32.270 45.600 32.590 45.660 ;
        RECT 33.205 45.615 33.495 45.660 ;
        RECT 16.645 45.460 16.935 45.505 ;
        RECT 23.990 45.460 24.310 45.520 ;
        RECT 30.890 45.460 31.210 45.520 ;
        RECT 16.645 45.320 24.310 45.460 ;
        RECT 16.645 45.275 16.935 45.320 ;
        RECT 23.990 45.260 24.310 45.320 ;
        RECT 25.460 45.320 31.210 45.460 ;
        RECT 19.865 45.120 20.155 45.165 ;
        RECT 13.500 44.980 20.155 45.120 ;
        RECT 11.110 44.780 11.430 44.840 ;
        RECT 13.500 44.825 13.640 44.980 ;
        RECT 19.865 44.935 20.155 44.980 ;
        RECT 13.425 44.780 13.715 44.825 ;
        RECT 11.110 44.640 13.715 44.780 ;
        RECT 11.110 44.580 11.430 44.640 ;
        RECT 13.425 44.595 13.715 44.640 ;
        RECT 15.710 44.580 16.030 44.840 ;
        RECT 16.170 44.580 16.490 44.840 ;
        RECT 17.105 44.780 17.395 44.825 ;
        RECT 25.460 44.780 25.600 45.320 ;
        RECT 30.890 45.260 31.210 45.320 ;
        RECT 17.105 44.640 25.600 44.780 ;
        RECT 25.845 44.780 26.135 44.825 ;
        RECT 26.290 44.780 26.610 44.840 ;
        RECT 25.845 44.640 26.610 44.780 ;
        RECT 17.105 44.595 17.395 44.640 ;
        RECT 25.845 44.595 26.135 44.640 ;
        RECT 26.290 44.580 26.610 44.640 ;
        RECT 29.050 44.780 29.370 44.840 ;
        RECT 29.985 44.780 30.275 44.825 ;
        RECT 29.050 44.640 30.275 44.780 ;
        RECT 29.050 44.580 29.370 44.640 ;
        RECT 29.985 44.595 30.275 44.640 ;
        RECT 34.110 44.580 34.430 44.840 ;
        RECT 36.870 44.580 37.190 44.840 ;
        RECT 38.250 44.580 38.570 44.840 ;
        RECT 39.630 44.580 39.950 44.840 ;
        RECT 18.010 43.900 18.330 44.160 ;
        RECT 23.070 43.900 23.390 44.160 ;
        RECT 26.750 44.100 27.070 44.160 ;
        RECT 29.525 44.100 29.815 44.145 ;
        RECT 26.750 43.960 29.815 44.100 ;
        RECT 26.750 43.900 27.070 43.960 ;
        RECT 29.525 43.915 29.815 43.960 ;
        RECT 32.730 44.100 33.050 44.160 ;
        RECT 35.965 44.100 36.255 44.145 ;
        RECT 32.730 43.960 36.255 44.100 ;
        RECT 32.730 43.900 33.050 43.960 ;
        RECT 35.965 43.915 36.255 43.960 ;
        RECT 36.410 44.100 36.730 44.160 ;
        RECT 37.345 44.100 37.635 44.145 ;
        RECT 36.410 43.960 37.635 44.100 ;
        RECT 36.410 43.900 36.730 43.960 ;
        RECT 37.345 43.915 37.635 43.960 ;
        RECT 38.725 44.100 39.015 44.145 ;
        RECT 39.170 44.100 39.490 44.160 ;
        RECT 38.725 43.960 39.490 44.100 ;
        RECT 38.725 43.915 39.015 43.960 ;
        RECT 39.170 43.900 39.490 43.960 ;
        RECT 5.520 43.280 41.400 43.760 ;
        RECT 11.110 42.880 11.430 43.140 ;
        RECT 15.710 43.080 16.030 43.140 ;
        RECT 25.385 43.080 25.675 43.125 ;
        RECT 26.290 43.080 26.610 43.140 ;
        RECT 15.710 42.940 21.000 43.080 ;
        RECT 15.710 42.880 16.030 42.940 ;
        RECT 18.010 42.740 18.330 42.800 ;
        RECT 19.710 42.740 20.000 42.785 ;
        RECT 18.010 42.600 20.000 42.740 ;
        RECT 20.860 42.740 21.000 42.940 ;
        RECT 25.385 42.940 26.610 43.080 ;
        RECT 25.385 42.895 25.675 42.940 ;
        RECT 26.290 42.880 26.610 42.940 ;
        RECT 25.845 42.740 26.135 42.785 ;
        RECT 20.860 42.600 26.135 42.740 ;
        RECT 18.010 42.540 18.330 42.600 ;
        RECT 19.710 42.555 20.000 42.600 ;
        RECT 25.845 42.555 26.135 42.600 ;
        RECT 26.750 42.540 27.070 42.800 ;
        RECT 16.745 42.400 17.035 42.445 ;
        RECT 18.930 42.400 19.250 42.460 ;
        RECT 16.745 42.260 19.250 42.400 ;
        RECT 16.745 42.215 17.035 42.260 ;
        RECT 18.930 42.200 19.250 42.260 ;
        RECT 27.670 42.200 27.990 42.460 ;
        RECT 28.145 42.215 28.435 42.445 ;
        RECT 29.050 42.400 29.370 42.460 ;
        RECT 29.985 42.400 30.275 42.445 ;
        RECT 29.050 42.260 30.275 42.400 ;
        RECT 13.435 42.060 13.725 42.105 ;
        RECT 15.955 42.060 16.245 42.105 ;
        RECT 17.145 42.060 17.435 42.105 ;
        RECT 13.435 41.920 17.435 42.060 ;
        RECT 13.435 41.875 13.725 41.920 ;
        RECT 15.955 41.875 16.245 41.920 ;
        RECT 17.145 41.875 17.435 41.920 ;
        RECT 18.025 42.060 18.315 42.105 ;
        RECT 18.485 42.060 18.775 42.105 ;
        RECT 18.025 41.920 18.775 42.060 ;
        RECT 18.025 41.875 18.315 41.920 ;
        RECT 18.485 41.875 18.775 41.920 ;
        RECT 19.365 42.060 19.655 42.105 ;
        RECT 20.555 42.060 20.845 42.105 ;
        RECT 23.075 42.060 23.365 42.105 ;
        RECT 19.365 41.920 23.365 42.060 ;
        RECT 19.365 41.875 19.655 41.920 ;
        RECT 20.555 41.875 20.845 41.920 ;
        RECT 23.075 41.875 23.365 41.920 ;
        RECT 24.450 42.060 24.770 42.120 ;
        RECT 28.220 42.060 28.360 42.215 ;
        RECT 29.050 42.200 29.370 42.260 ;
        RECT 29.985 42.215 30.275 42.260 ;
        RECT 30.890 42.400 31.210 42.460 ;
        RECT 32.745 42.400 33.035 42.445 ;
        RECT 30.890 42.260 33.035 42.400 ;
        RECT 30.890 42.200 31.210 42.260 ;
        RECT 32.745 42.215 33.035 42.260 ;
        RECT 33.650 42.200 33.970 42.460 ;
        RECT 34.125 42.400 34.415 42.445 ;
        RECT 36.870 42.400 37.190 42.460 ;
        RECT 34.125 42.260 37.190 42.400 ;
        RECT 34.125 42.215 34.415 42.260 ;
        RECT 36.870 42.200 37.190 42.260 ;
        RECT 39.630 42.200 39.950 42.460 ;
        RECT 24.450 41.920 28.360 42.060 ;
        RECT 28.590 42.060 28.910 42.120 ;
        RECT 30.980 42.060 31.120 42.200 ;
        RECT 28.590 41.920 31.120 42.060 ;
        RECT 13.870 41.720 14.160 41.765 ;
        RECT 15.440 41.720 15.730 41.765 ;
        RECT 17.540 41.720 17.830 41.765 ;
        RECT 13.870 41.580 17.830 41.720 ;
        RECT 13.870 41.535 14.160 41.580 ;
        RECT 15.440 41.535 15.730 41.580 ;
        RECT 17.540 41.535 17.830 41.580 ;
        RECT 16.630 41.380 16.950 41.440 ;
        RECT 18.560 41.380 18.700 41.875 ;
        RECT 24.450 41.860 24.770 41.920 ;
        RECT 28.590 41.860 28.910 41.920 ;
        RECT 35.045 41.875 35.335 42.105 ;
        RECT 18.970 41.720 19.260 41.765 ;
        RECT 21.070 41.720 21.360 41.765 ;
        RECT 22.640 41.720 22.930 41.765 ;
        RECT 18.970 41.580 22.930 41.720 ;
        RECT 18.970 41.535 19.260 41.580 ;
        RECT 21.070 41.535 21.360 41.580 ;
        RECT 22.640 41.535 22.930 41.580 ;
        RECT 23.530 41.720 23.850 41.780 ;
        RECT 29.065 41.720 29.355 41.765 ;
        RECT 23.530 41.580 29.355 41.720 ;
        RECT 23.530 41.520 23.850 41.580 ;
        RECT 29.065 41.535 29.355 41.580 ;
        RECT 30.445 41.720 30.735 41.765 ;
        RECT 33.205 41.720 33.495 41.765 ;
        RECT 30.445 41.580 33.495 41.720 ;
        RECT 30.445 41.535 30.735 41.580 ;
        RECT 33.205 41.535 33.495 41.580 ;
        RECT 34.110 41.720 34.430 41.780 ;
        RECT 35.120 41.720 35.260 41.875 ;
        RECT 34.110 41.580 35.260 41.720 ;
        RECT 37.330 41.720 37.650 41.780 ;
        RECT 38.725 41.720 39.015 41.765 ;
        RECT 37.330 41.580 39.015 41.720 ;
        RECT 34.110 41.520 34.430 41.580 ;
        RECT 37.330 41.520 37.650 41.580 ;
        RECT 38.725 41.535 39.015 41.580 ;
        RECT 27.210 41.380 27.530 41.440 ;
        RECT 16.630 41.240 27.530 41.380 ;
        RECT 16.630 41.180 16.950 41.240 ;
        RECT 27.210 41.180 27.530 41.240 ;
        RECT 29.970 41.380 30.290 41.440 ;
        RECT 31.825 41.380 32.115 41.425 ;
        RECT 29.970 41.240 32.115 41.380 ;
        RECT 29.970 41.180 30.290 41.240 ;
        RECT 31.825 41.195 32.115 41.240 ;
        RECT 35.950 41.380 36.270 41.440 ;
        RECT 38.265 41.380 38.555 41.425 ;
        RECT 35.950 41.240 38.555 41.380 ;
        RECT 35.950 41.180 36.270 41.240 ;
        RECT 38.265 41.195 38.555 41.240 ;
        RECT 5.520 40.560 41.400 41.040 ;
        RECT 18.930 40.160 19.250 40.420 ;
        RECT 23.990 40.360 24.310 40.420 ;
        RECT 26.305 40.360 26.595 40.405 ;
        RECT 29.050 40.360 29.370 40.420 ;
        RECT 23.990 40.220 26.595 40.360 ;
        RECT 23.990 40.160 24.310 40.220 ;
        RECT 26.305 40.175 26.595 40.220 ;
        RECT 27.300 40.220 32.500 40.360 ;
        RECT 7.470 40.020 7.760 40.065 ;
        RECT 9.570 40.020 9.860 40.065 ;
        RECT 11.140 40.020 11.430 40.065 ;
        RECT 27.300 40.020 27.440 40.220 ;
        RECT 29.050 40.160 29.370 40.220 ;
        RECT 7.470 39.880 11.430 40.020 ;
        RECT 7.470 39.835 7.760 39.880 ;
        RECT 9.570 39.835 9.860 39.880 ;
        RECT 11.140 39.835 11.430 39.880 ;
        RECT 22.240 39.880 27.440 40.020 ;
        RECT 27.710 40.020 28.000 40.065 ;
        RECT 29.810 40.020 30.100 40.065 ;
        RECT 31.380 40.020 31.670 40.065 ;
        RECT 27.710 39.880 31.670 40.020 ;
        RECT 22.240 39.725 22.380 39.880 ;
        RECT 27.710 39.835 28.000 39.880 ;
        RECT 29.810 39.835 30.100 39.880 ;
        RECT 31.380 39.835 31.670 39.880 ;
        RECT 7.865 39.680 8.155 39.725 ;
        RECT 9.055 39.680 9.345 39.725 ;
        RECT 11.575 39.680 11.865 39.725 ;
        RECT 7.865 39.540 11.865 39.680 ;
        RECT 7.865 39.495 8.155 39.540 ;
        RECT 9.055 39.495 9.345 39.540 ;
        RECT 11.575 39.495 11.865 39.540 ;
        RECT 22.165 39.495 22.455 39.725 ;
        RECT 27.210 39.480 27.530 39.740 ;
        RECT 28.105 39.680 28.395 39.725 ;
        RECT 29.295 39.680 29.585 39.725 ;
        RECT 31.815 39.680 32.105 39.725 ;
        RECT 28.105 39.540 32.105 39.680 ;
        RECT 28.105 39.495 28.395 39.540 ;
        RECT 29.295 39.495 29.585 39.540 ;
        RECT 31.815 39.495 32.105 39.540 ;
        RECT 6.985 39.340 7.275 39.385 ;
        RECT 16.630 39.340 16.950 39.400 ;
        RECT 6.985 39.200 16.950 39.340 ;
        RECT 6.985 39.155 7.275 39.200 ;
        RECT 16.630 39.140 16.950 39.200 ;
        RECT 17.105 39.155 17.395 39.385 ;
        RECT 20.785 39.340 21.075 39.385 ;
        RECT 23.070 39.340 23.390 39.400 ;
        RECT 20.785 39.200 23.390 39.340 ;
        RECT 20.785 39.155 21.075 39.200 ;
        RECT 8.320 39.000 8.610 39.045 ;
        RECT 8.810 39.000 9.130 39.060 ;
        RECT 17.180 39.000 17.320 39.155 ;
        RECT 23.070 39.140 23.390 39.200 ;
        RECT 23.530 39.140 23.850 39.400 ;
        RECT 24.450 39.340 24.770 39.400 ;
        RECT 26.290 39.340 26.610 39.400 ;
        RECT 24.450 39.200 26.610 39.340 ;
        RECT 24.450 39.140 24.770 39.200 ;
        RECT 26.290 39.140 26.610 39.200 ;
        RECT 26.750 39.340 27.070 39.400 ;
        RECT 27.670 39.340 27.990 39.400 ;
        RECT 26.750 39.200 27.990 39.340 ;
        RECT 26.750 39.140 27.070 39.200 ;
        RECT 27.670 39.140 27.990 39.200 ;
        RECT 28.560 39.340 28.850 39.385 ;
        RECT 29.970 39.340 30.290 39.400 ;
        RECT 28.560 39.200 30.290 39.340 ;
        RECT 32.360 39.340 32.500 40.220 ;
        RECT 34.110 40.160 34.430 40.420 ;
        RECT 36.870 40.160 37.190 40.420 ;
        RECT 35.045 39.340 35.335 39.385 ;
        RECT 32.360 39.200 35.335 39.340 ;
        RECT 28.560 39.155 28.850 39.200 ;
        RECT 29.970 39.140 30.290 39.200 ;
        RECT 35.045 39.155 35.335 39.200 ;
        RECT 35.950 39.140 36.270 39.400 ;
        RECT 37.330 39.140 37.650 39.400 ;
        RECT 39.630 39.140 39.950 39.400 ;
        RECT 8.320 38.860 9.130 39.000 ;
        RECT 8.320 38.815 8.610 38.860 ;
        RECT 8.810 38.800 9.130 38.860 ;
        RECT 13.960 38.860 17.320 39.000 ;
        RECT 21.245 39.000 21.535 39.045 ;
        RECT 29.050 39.000 29.370 39.060 ;
        RECT 21.245 38.860 29.370 39.000 ;
        RECT 13.960 38.720 14.100 38.860 ;
        RECT 21.245 38.815 21.535 38.860 ;
        RECT 29.050 38.800 29.370 38.860 ;
        RECT 13.870 38.460 14.190 38.720 ;
        RECT 14.330 38.460 14.650 38.720 ;
        RECT 23.070 38.660 23.390 38.720 ;
        RECT 25.385 38.660 25.675 38.705 ;
        RECT 23.070 38.520 25.675 38.660 ;
        RECT 23.070 38.460 23.390 38.520 ;
        RECT 25.385 38.475 25.675 38.520 ;
        RECT 38.250 38.460 38.570 38.720 ;
        RECT 38.710 38.460 39.030 38.720 ;
        RECT 5.520 37.840 41.400 38.320 ;
        RECT 6.510 37.640 6.830 37.700 ;
        RECT 7.445 37.640 7.735 37.685 ;
        RECT 6.510 37.500 7.735 37.640 ;
        RECT 6.510 37.440 6.830 37.500 ;
        RECT 7.445 37.455 7.735 37.500 ;
        RECT 8.810 37.440 9.130 37.700 ;
        RECT 10.665 37.640 10.955 37.685 ;
        RECT 14.330 37.640 14.650 37.700 ;
        RECT 10.665 37.500 14.650 37.640 ;
        RECT 10.665 37.455 10.955 37.500 ;
        RECT 14.330 37.440 14.650 37.500 ;
        RECT 16.630 37.640 16.950 37.700 ;
        RECT 18.930 37.640 19.250 37.700 ;
        RECT 16.630 37.500 19.250 37.640 ;
        RECT 16.630 37.440 16.950 37.500 ;
        RECT 18.930 37.440 19.250 37.500 ;
        RECT 19.850 37.640 20.170 37.700 ;
        RECT 23.530 37.640 23.850 37.700 ;
        RECT 36.410 37.640 36.730 37.700 ;
        RECT 19.850 37.500 23.850 37.640 ;
        RECT 19.850 37.440 20.170 37.500 ;
        RECT 23.530 37.440 23.850 37.500 ;
        RECT 30.060 37.500 36.730 37.640 ;
        RECT 28.590 37.100 28.910 37.360 ;
        RECT 8.365 36.960 8.655 37.005 ;
        RECT 13.870 36.960 14.190 37.020 ;
        RECT 8.365 36.820 14.190 36.960 ;
        RECT 8.365 36.775 8.655 36.820 ;
        RECT 13.870 36.760 14.190 36.820 ;
        RECT 23.085 36.960 23.375 37.005 ;
        RECT 23.530 36.960 23.850 37.020 ;
        RECT 30.060 37.005 30.200 37.500 ;
        RECT 36.410 37.440 36.730 37.500 ;
        RECT 38.710 37.440 39.030 37.700 ;
        RECT 31.825 37.300 32.115 37.345 ;
        RECT 33.190 37.300 33.510 37.360 ;
        RECT 31.825 37.160 33.510 37.300 ;
        RECT 31.825 37.115 32.115 37.160 ;
        RECT 33.190 37.100 33.510 37.160 ;
        RECT 33.650 37.300 33.970 37.360 ;
        RECT 38.800 37.300 38.940 37.440 ;
        RECT 33.650 37.160 38.940 37.300 ;
        RECT 33.650 37.100 33.970 37.160 ;
        RECT 23.085 36.820 23.850 36.960 ;
        RECT 23.085 36.775 23.375 36.820 ;
        RECT 23.530 36.760 23.850 36.820 ;
        RECT 29.985 36.775 30.275 37.005 ;
        RECT 32.730 36.760 33.050 37.020 ;
        RECT 35.120 37.005 35.260 37.160 ;
        RECT 34.125 36.775 34.415 37.005 ;
        RECT 35.045 36.775 35.335 37.005 ;
        RECT 11.125 36.435 11.415 36.665 ;
        RECT 12.045 36.620 12.335 36.665 ;
        RECT 12.490 36.620 12.810 36.680 ;
        RECT 12.045 36.480 12.810 36.620 ;
        RECT 12.045 36.435 12.335 36.480 ;
        RECT 9.270 36.280 9.590 36.340 ;
        RECT 11.200 36.280 11.340 36.435 ;
        RECT 12.490 36.420 12.810 36.480 ;
        RECT 26.765 36.620 27.055 36.665 ;
        RECT 27.210 36.620 27.530 36.680 ;
        RECT 26.765 36.480 27.530 36.620 ;
        RECT 26.765 36.435 27.055 36.480 ;
        RECT 27.210 36.420 27.530 36.480 ;
        RECT 29.525 36.620 29.815 36.665 ;
        RECT 32.820 36.620 32.960 36.760 ;
        RECT 29.525 36.480 32.960 36.620 ;
        RECT 34.200 36.620 34.340 36.775 ;
        RECT 36.410 36.760 36.730 37.020 ;
        RECT 37.790 36.760 38.110 37.020 ;
        RECT 38.725 36.960 39.015 37.005 ;
        RECT 39.170 36.960 39.490 37.020 ;
        RECT 38.725 36.820 39.490 36.960 ;
        RECT 38.725 36.775 39.015 36.820 ;
        RECT 39.170 36.760 39.490 36.820 ;
        RECT 35.505 36.620 35.795 36.665 ;
        RECT 34.200 36.480 35.795 36.620 ;
        RECT 29.525 36.435 29.815 36.480 ;
        RECT 35.505 36.435 35.795 36.480 ;
        RECT 29.050 36.280 29.370 36.340 ;
        RECT 33.650 36.280 33.970 36.340 ;
        RECT 9.270 36.140 29.370 36.280 ;
        RECT 9.270 36.080 9.590 36.140 ;
        RECT 29.050 36.080 29.370 36.140 ;
        RECT 30.060 36.140 33.970 36.280 ;
        RECT 23.545 35.940 23.835 35.985 ;
        RECT 23.990 35.940 24.310 36.000 ;
        RECT 30.060 35.985 30.200 36.140 ;
        RECT 33.650 36.080 33.970 36.140 ;
        RECT 23.545 35.800 24.310 35.940 ;
        RECT 23.545 35.755 23.835 35.800 ;
        RECT 23.990 35.740 24.310 35.800 ;
        RECT 29.985 35.755 30.275 35.985 ;
        RECT 30.890 35.740 31.210 36.000 ;
        RECT 5.520 35.120 41.400 35.600 ;
        RECT 19.850 34.920 20.170 34.980 ;
        RECT 11.200 34.780 20.170 34.920 ;
        RECT 9.270 34.040 9.590 34.300 ;
        RECT 10.205 34.240 10.495 34.285 ;
        RECT 11.200 34.240 11.340 34.780 ;
        RECT 19.850 34.720 20.170 34.780 ;
        RECT 25.845 34.920 26.135 34.965 ;
        RECT 26.290 34.920 26.610 34.980 ;
        RECT 25.845 34.780 26.610 34.920 ;
        RECT 25.845 34.735 26.135 34.780 ;
        RECT 26.290 34.720 26.610 34.780 ;
        RECT 35.965 34.920 36.255 34.965 ;
        RECT 37.790 34.920 38.110 34.980 ;
        RECT 35.965 34.780 38.110 34.920 ;
        RECT 35.965 34.735 36.255 34.780 ;
        RECT 37.790 34.720 38.110 34.780 ;
        RECT 11.610 34.580 11.900 34.625 ;
        RECT 13.710 34.580 14.000 34.625 ;
        RECT 15.280 34.580 15.570 34.625 ;
        RECT 11.610 34.440 15.570 34.580 ;
        RECT 11.610 34.395 11.900 34.440 ;
        RECT 13.710 34.395 14.000 34.440 ;
        RECT 15.280 34.395 15.570 34.440 ;
        RECT 18.025 34.395 18.315 34.625 ;
        RECT 19.430 34.580 19.720 34.625 ;
        RECT 21.530 34.580 21.820 34.625 ;
        RECT 23.100 34.580 23.390 34.625 ;
        RECT 19.430 34.440 23.390 34.580 ;
        RECT 19.430 34.395 19.720 34.440 ;
        RECT 21.530 34.395 21.820 34.440 ;
        RECT 23.100 34.395 23.390 34.440 ;
        RECT 10.205 34.100 11.340 34.240 ;
        RECT 12.005 34.240 12.295 34.285 ;
        RECT 13.195 34.240 13.485 34.285 ;
        RECT 15.715 34.240 16.005 34.285 ;
        RECT 12.005 34.100 16.005 34.240 ;
        RECT 10.205 34.055 10.495 34.100 ;
        RECT 12.005 34.055 12.295 34.100 ;
        RECT 13.195 34.055 13.485 34.100 ;
        RECT 15.715 34.055 16.005 34.100 ;
        RECT 11.125 33.900 11.415 33.945 ;
        RECT 13.870 33.900 14.190 33.960 ;
        RECT 16.630 33.900 16.950 33.960 ;
        RECT 11.125 33.760 16.950 33.900 ;
        RECT 18.100 33.900 18.240 34.395 ;
        RECT 27.670 34.380 27.990 34.640 ;
        RECT 34.570 34.580 34.890 34.640 ;
        RECT 39.170 34.580 39.490 34.640 ;
        RECT 32.360 34.440 39.490 34.580 ;
        RECT 18.930 34.040 19.250 34.300 ;
        RECT 32.360 34.285 32.500 34.440 ;
        RECT 34.570 34.380 34.890 34.440 ;
        RECT 39.170 34.380 39.490 34.440 ;
        RECT 19.825 34.240 20.115 34.285 ;
        RECT 21.015 34.240 21.305 34.285 ;
        RECT 23.535 34.240 23.825 34.285 ;
        RECT 19.825 34.100 23.825 34.240 ;
        RECT 19.825 34.055 20.115 34.100 ;
        RECT 21.015 34.055 21.305 34.100 ;
        RECT 23.535 34.055 23.825 34.100 ;
        RECT 32.285 34.055 32.575 34.285 ;
        RECT 32.745 34.240 33.035 34.285 ;
        RECT 35.490 34.240 35.810 34.300 ;
        RECT 32.745 34.100 35.810 34.240 ;
        RECT 32.745 34.055 33.035 34.100 ;
        RECT 35.490 34.040 35.810 34.100 ;
        RECT 27.210 33.900 27.530 33.960 ;
        RECT 18.100 33.760 28.360 33.900 ;
        RECT 11.125 33.715 11.415 33.760 ;
        RECT 13.870 33.700 14.190 33.760 ;
        RECT 16.630 33.700 16.950 33.760 ;
        RECT 27.210 33.700 27.530 33.760 ;
        RECT 28.220 33.620 28.360 33.760 ;
        RECT 31.825 33.715 32.115 33.945 ;
        RECT 33.205 33.715 33.495 33.945 ;
        RECT 33.650 33.900 33.970 33.960 ;
        RECT 34.125 33.900 34.415 33.945 ;
        RECT 33.650 33.760 34.415 33.900 ;
        RECT 12.490 33.605 12.810 33.620 ;
        RECT 12.460 33.560 12.810 33.605 ;
        RECT 20.280 33.560 20.570 33.605 ;
        RECT 26.750 33.560 27.070 33.620 ;
        RECT 12.055 33.420 20.080 33.560 ;
        RECT 12.460 33.375 12.810 33.420 ;
        RECT 12.490 33.360 12.810 33.375 ;
        RECT 6.970 33.020 7.290 33.280 ;
        RECT 8.825 33.220 9.115 33.265 ;
        RECT 11.570 33.220 11.890 33.280 ;
        RECT 8.825 33.080 11.890 33.220 ;
        RECT 19.940 33.220 20.080 33.420 ;
        RECT 20.280 33.420 27.070 33.560 ;
        RECT 20.280 33.375 20.570 33.420 ;
        RECT 26.750 33.360 27.070 33.420 ;
        RECT 28.130 33.560 28.450 33.620 ;
        RECT 29.525 33.560 29.815 33.605 ;
        RECT 28.130 33.420 29.815 33.560 ;
        RECT 31.900 33.560 32.040 33.715 ;
        RECT 33.280 33.560 33.420 33.715 ;
        RECT 33.650 33.700 33.970 33.760 ;
        RECT 34.125 33.715 34.415 33.760 ;
        RECT 35.045 33.900 35.335 33.945 ;
        RECT 36.410 33.900 36.730 33.960 ;
        RECT 35.045 33.760 36.730 33.900 ;
        RECT 35.045 33.715 35.335 33.760 ;
        RECT 36.410 33.700 36.730 33.760 ;
        RECT 36.870 33.700 37.190 33.960 ;
        RECT 38.250 33.700 38.570 33.960 ;
        RECT 38.710 33.900 39.030 33.960 ;
        RECT 39.185 33.900 39.475 33.945 ;
        RECT 38.710 33.760 39.475 33.900 ;
        RECT 38.710 33.700 39.030 33.760 ;
        RECT 39.185 33.715 39.475 33.760 ;
        RECT 34.585 33.560 34.875 33.605 ;
        RECT 31.900 33.420 32.500 33.560 ;
        RECT 33.280 33.420 34.875 33.560 ;
        RECT 28.130 33.360 28.450 33.420 ;
        RECT 29.525 33.375 29.815 33.420 ;
        RECT 26.290 33.220 26.610 33.280 ;
        RECT 27.225 33.220 27.515 33.265 ;
        RECT 19.940 33.080 27.515 33.220 ;
        RECT 8.825 33.035 9.115 33.080 ;
        RECT 11.570 33.020 11.890 33.080 ;
        RECT 26.290 33.020 26.610 33.080 ;
        RECT 27.225 33.035 27.515 33.080 ;
        RECT 30.905 33.220 31.195 33.265 ;
        RECT 31.810 33.220 32.130 33.280 ;
        RECT 30.905 33.080 32.130 33.220 ;
        RECT 32.360 33.220 32.500 33.420 ;
        RECT 34.585 33.375 34.875 33.420 ;
        RECT 36.960 33.220 37.100 33.700 ;
        RECT 32.360 33.080 37.100 33.220 ;
        RECT 30.905 33.035 31.195 33.080 ;
        RECT 31.810 33.020 32.130 33.080 ;
        RECT 5.520 32.400 41.400 32.880 ;
        RECT 26.750 32.000 27.070 32.260 ;
        RECT 29.050 32.200 29.370 32.260 ;
        RECT 33.665 32.200 33.955 32.245 ;
        RECT 29.050 32.060 33.955 32.200 ;
        RECT 29.050 32.000 29.370 32.060 ;
        RECT 33.665 32.015 33.955 32.060 ;
        RECT 38.725 32.015 39.015 32.245 ;
        RECT 6.970 31.860 7.290 31.920 ;
        RECT 12.550 31.860 12.840 31.905 ;
        RECT 6.970 31.720 12.840 31.860 ;
        RECT 6.970 31.660 7.290 31.720 ;
        RECT 12.550 31.675 12.840 31.720 ;
        RECT 17.550 31.660 17.870 31.920 ;
        RECT 38.800 31.860 38.940 32.015 ;
        RECT 37.420 31.720 38.940 31.860 ;
        RECT 37.420 31.580 37.560 31.720 ;
        RECT 13.870 31.320 14.190 31.580 ;
        RECT 31.810 31.320 32.130 31.580 ;
        RECT 32.730 31.320 33.050 31.580 ;
        RECT 37.330 31.320 37.650 31.580 ;
        RECT 38.265 31.520 38.555 31.565 ;
        RECT 38.710 31.520 39.030 31.580 ;
        RECT 38.265 31.380 39.030 31.520 ;
        RECT 38.265 31.335 38.555 31.380 ;
        RECT 38.710 31.320 39.030 31.380 ;
        RECT 39.630 31.320 39.950 31.580 ;
        RECT 9.295 31.180 9.585 31.225 ;
        RECT 11.815 31.180 12.105 31.225 ;
        RECT 13.005 31.180 13.295 31.225 ;
        RECT 9.295 31.040 13.295 31.180 ;
        RECT 9.295 30.995 9.585 31.040 ;
        RECT 11.815 30.995 12.105 31.040 ;
        RECT 13.005 30.995 13.295 31.040 ;
        RECT 23.990 31.180 24.310 31.240 ;
        RECT 29.525 31.180 29.815 31.225 ;
        RECT 23.990 31.040 29.815 31.180 ;
        RECT 23.990 30.980 24.310 31.040 ;
        RECT 29.525 30.995 29.815 31.040 ;
        RECT 9.730 30.840 10.020 30.885 ;
        RECT 11.300 30.840 11.590 30.885 ;
        RECT 13.400 30.840 13.690 30.885 ;
        RECT 9.730 30.700 13.690 30.840 ;
        RECT 9.730 30.655 10.020 30.700 ;
        RECT 11.300 30.655 11.590 30.700 ;
        RECT 13.400 30.655 13.690 30.700 ;
        RECT 6.970 30.300 7.290 30.560 ;
        RECT 23.530 30.500 23.850 30.560 ;
        RECT 24.005 30.500 24.295 30.545 ;
        RECT 23.530 30.360 24.295 30.500 ;
        RECT 23.530 30.300 23.850 30.360 ;
        RECT 24.005 30.315 24.295 30.360 ;
        RECT 28.590 30.500 28.910 30.560 ;
        RECT 31.825 30.500 32.115 30.545 ;
        RECT 28.590 30.360 32.115 30.500 ;
        RECT 28.590 30.300 28.910 30.360 ;
        RECT 31.825 30.315 32.115 30.360 ;
        RECT 35.030 30.500 35.350 30.560 ;
        RECT 38.265 30.500 38.555 30.545 ;
        RECT 35.030 30.360 38.555 30.500 ;
        RECT 35.030 30.300 35.350 30.360 ;
        RECT 38.265 30.315 38.555 30.360 ;
        RECT 5.520 29.680 41.400 30.160 ;
        RECT 11.570 29.280 11.890 29.540 ;
        RECT 19.850 29.280 20.170 29.540 ;
        RECT 20.310 29.480 20.630 29.540 ;
        RECT 22.165 29.480 22.455 29.525 ;
        RECT 20.310 29.340 22.455 29.480 ;
        RECT 20.310 29.280 20.630 29.340 ;
        RECT 22.165 29.295 22.455 29.340 ;
        RECT 30.890 29.280 31.210 29.540 ;
        RECT 38.250 29.480 38.570 29.540 ;
        RECT 39.185 29.480 39.475 29.525 ;
        RECT 38.250 29.340 39.475 29.480 ;
        RECT 38.250 29.280 38.570 29.340 ;
        RECT 39.185 29.295 39.475 29.340 ;
        RECT 21.245 29.140 21.535 29.185 ;
        RECT 24.450 29.140 24.770 29.200 ;
        RECT 28.590 29.140 28.910 29.200 ;
        RECT 21.245 29.000 24.770 29.140 ;
        RECT 21.245 28.955 21.535 29.000 ;
        RECT 6.970 28.800 7.290 28.860 ;
        RECT 8.365 28.800 8.655 28.845 ;
        RECT 21.320 28.800 21.460 28.955 ;
        RECT 24.450 28.940 24.770 29.000 ;
        RECT 27.300 29.000 28.910 29.140 ;
        RECT 6.970 28.660 8.655 28.800 ;
        RECT 6.970 28.600 7.290 28.660 ;
        RECT 8.365 28.615 8.655 28.660 ;
        RECT 19.940 28.660 21.460 28.800 ;
        RECT 21.705 28.800 21.995 28.845 ;
        RECT 27.300 28.800 27.440 29.000 ;
        RECT 28.590 28.940 28.910 29.000 ;
        RECT 36.870 28.940 37.190 29.200 ;
        RECT 21.705 28.660 27.440 28.800 ;
        RECT 14.790 28.260 15.110 28.520 ;
        RECT 19.940 28.505 20.080 28.660 ;
        RECT 21.705 28.615 21.995 28.660 ;
        RECT 27.670 28.600 27.990 28.860 ;
        RECT 36.960 28.800 37.100 28.940 ;
        RECT 30.520 28.660 37.100 28.800 ;
        RECT 18.945 28.275 19.235 28.505 ;
        RECT 19.865 28.275 20.155 28.505 ;
        RECT 19.020 28.120 19.160 28.275 ;
        RECT 20.310 28.260 20.630 28.520 ;
        RECT 22.625 28.460 22.915 28.505 ;
        RECT 23.070 28.460 23.390 28.520 ;
        RECT 22.625 28.320 23.390 28.460 ;
        RECT 22.625 28.275 22.915 28.320 ;
        RECT 23.070 28.260 23.390 28.320 ;
        RECT 23.990 28.260 24.310 28.520 ;
        RECT 30.520 28.505 30.660 28.660 ;
        RECT 30.445 28.275 30.735 28.505 ;
        RECT 31.365 28.460 31.655 28.505 ;
        RECT 33.205 28.460 33.495 28.505 ;
        RECT 33.650 28.460 33.970 28.520 ;
        RECT 34.200 28.505 34.340 28.660 ;
        RECT 31.365 28.320 33.970 28.460 ;
        RECT 31.365 28.275 31.655 28.320 ;
        RECT 33.205 28.275 33.495 28.320 ;
        RECT 33.650 28.260 33.970 28.320 ;
        RECT 34.125 28.275 34.415 28.505 ;
        RECT 34.570 28.260 34.890 28.520 ;
        RECT 35.965 28.275 36.255 28.505 ;
        RECT 24.465 28.120 24.755 28.165 ;
        RECT 19.020 27.980 24.755 28.120 ;
        RECT 24.465 27.935 24.755 27.980 ;
        RECT 32.745 28.120 33.035 28.165 ;
        RECT 35.030 28.120 35.350 28.180 ;
        RECT 36.040 28.120 36.180 28.275 ;
        RECT 36.870 28.260 37.190 28.520 ;
        RECT 37.330 28.460 37.650 28.520 ;
        RECT 38.265 28.460 38.555 28.505 ;
        RECT 37.330 28.320 38.555 28.460 ;
        RECT 37.330 28.260 37.650 28.320 ;
        RECT 38.265 28.275 38.555 28.320 ;
        RECT 37.790 28.120 38.110 28.180 ;
        RECT 32.745 27.980 35.350 28.120 ;
        RECT 32.745 27.935 33.035 27.980 ;
        RECT 35.030 27.920 35.350 27.980 ;
        RECT 35.580 27.980 38.110 28.120 ;
        RECT 12.030 27.580 12.350 27.840 ;
        RECT 29.525 27.780 29.815 27.825 ;
        RECT 30.430 27.780 30.750 27.840 ;
        RECT 29.525 27.640 30.750 27.780 ;
        RECT 29.525 27.595 29.815 27.640 ;
        RECT 30.430 27.580 30.750 27.640 ;
        RECT 33.190 27.780 33.510 27.840 ;
        RECT 35.580 27.825 35.720 27.980 ;
        RECT 37.790 27.920 38.110 27.980 ;
        RECT 33.665 27.780 33.955 27.825 ;
        RECT 33.190 27.640 33.955 27.780 ;
        RECT 33.190 27.580 33.510 27.640 ;
        RECT 33.665 27.595 33.955 27.640 ;
        RECT 35.505 27.595 35.795 27.825 ;
        RECT 5.520 26.960 41.400 27.440 ;
        RECT 6.510 26.760 6.830 26.820 ;
        RECT 7.445 26.760 7.735 26.805 ;
        RECT 6.510 26.620 7.735 26.760 ;
        RECT 6.510 26.560 6.830 26.620 ;
        RECT 7.445 26.575 7.735 26.620 ;
        RECT 11.125 26.760 11.415 26.805 ;
        RECT 12.030 26.760 12.350 26.820 ;
        RECT 11.125 26.620 12.350 26.760 ;
        RECT 11.125 26.575 11.415 26.620 ;
        RECT 12.030 26.560 12.350 26.620 ;
        RECT 20.310 26.760 20.630 26.820 ;
        RECT 27.210 26.760 27.530 26.820 ;
        RECT 20.310 26.620 27.530 26.760 ;
        RECT 20.310 26.560 20.630 26.620 ;
        RECT 27.210 26.560 27.530 26.620 ;
        RECT 36.870 26.760 37.190 26.820 ;
        RECT 39.185 26.760 39.475 26.805 ;
        RECT 36.870 26.620 39.475 26.760 ;
        RECT 36.870 26.560 37.190 26.620 ;
        RECT 39.185 26.575 39.475 26.620 ;
        RECT 14.760 26.420 15.050 26.465 ;
        RECT 18.470 26.420 18.790 26.480 ;
        RECT 19.850 26.420 20.170 26.480 ;
        RECT 35.030 26.420 35.350 26.480 ;
        RECT 14.760 26.280 20.170 26.420 ;
        RECT 14.760 26.235 15.050 26.280 ;
        RECT 18.470 26.220 18.790 26.280 ;
        RECT 19.850 26.220 20.170 26.280 ;
        RECT 32.820 26.280 35.350 26.420 ;
        RECT 6.970 26.080 7.290 26.140 ;
        RECT 8.365 26.080 8.655 26.125 ;
        RECT 6.970 25.940 8.655 26.080 ;
        RECT 6.970 25.880 7.290 25.940 ;
        RECT 8.365 25.895 8.655 25.940 ;
        RECT 22.625 26.080 22.915 26.125 ;
        RECT 24.925 26.080 25.215 26.125 ;
        RECT 22.625 25.940 25.215 26.080 ;
        RECT 22.625 25.895 22.915 25.940 ;
        RECT 24.925 25.895 25.215 25.940 ;
        RECT 30.890 26.080 31.210 26.140 ;
        RECT 32.820 26.125 32.960 26.280 ;
        RECT 35.030 26.220 35.350 26.280 ;
        RECT 32.285 26.080 32.575 26.125 ;
        RECT 30.890 25.940 32.575 26.080 ;
        RECT 30.890 25.880 31.210 25.940 ;
        RECT 32.285 25.895 32.575 25.940 ;
        RECT 32.745 25.895 33.035 26.125 ;
        RECT 33.190 25.880 33.510 26.140 ;
        RECT 35.965 26.080 36.255 26.125 ;
        RECT 36.410 26.080 36.730 26.140 ;
        RECT 35.965 25.940 36.730 26.080 ;
        RECT 35.965 25.895 36.255 25.940 ;
        RECT 36.410 25.880 36.730 25.940 ;
        RECT 36.870 25.880 37.190 26.140 ;
        RECT 38.265 26.080 38.555 26.125 ;
        RECT 38.710 26.080 39.030 26.140 ;
        RECT 38.265 25.940 39.030 26.080 ;
        RECT 38.265 25.895 38.555 25.940 ;
        RECT 38.710 25.880 39.030 25.940 ;
        RECT 11.585 25.740 11.875 25.785 ;
        RECT 12.030 25.740 12.350 25.800 ;
        RECT 11.585 25.600 12.350 25.740 ;
        RECT 11.585 25.555 11.875 25.600 ;
        RECT 12.030 25.540 12.350 25.600 ;
        RECT 12.490 25.540 12.810 25.800 ;
        RECT 13.425 25.555 13.715 25.785 ;
        RECT 14.305 25.740 14.595 25.785 ;
        RECT 15.495 25.740 15.785 25.785 ;
        RECT 18.015 25.740 18.305 25.785 ;
        RECT 14.305 25.600 18.305 25.740 ;
        RECT 14.305 25.555 14.595 25.600 ;
        RECT 15.495 25.555 15.785 25.600 ;
        RECT 18.015 25.555 18.305 25.600 ;
        RECT 23.085 25.555 23.375 25.785 ;
        RECT 24.005 25.740 24.295 25.785 ;
        RECT 26.290 25.740 26.610 25.800 ;
        RECT 24.005 25.600 26.610 25.740 ;
        RECT 24.005 25.555 24.295 25.600 ;
        RECT 6.970 25.400 7.290 25.460 ;
        RECT 13.500 25.400 13.640 25.555 ;
        RECT 6.970 25.260 13.640 25.400 ;
        RECT 13.910 25.400 14.200 25.445 ;
        RECT 16.010 25.400 16.300 25.445 ;
        RECT 17.580 25.400 17.870 25.445 ;
        RECT 13.910 25.260 17.870 25.400 ;
        RECT 6.970 25.200 7.290 25.260 ;
        RECT 13.910 25.215 14.200 25.260 ;
        RECT 16.010 25.215 16.300 25.260 ;
        RECT 17.580 25.215 17.870 25.260 ;
        RECT 19.850 25.400 20.170 25.460 ;
        RECT 20.785 25.400 21.075 25.445 ;
        RECT 19.850 25.260 21.075 25.400 ;
        RECT 23.160 25.400 23.300 25.555 ;
        RECT 26.290 25.540 26.610 25.600 ;
        RECT 26.750 25.740 27.070 25.800 ;
        RECT 27.685 25.740 27.975 25.785 ;
        RECT 26.750 25.600 27.975 25.740 ;
        RECT 26.750 25.540 27.070 25.600 ;
        RECT 27.685 25.555 27.975 25.600 ;
        RECT 33.665 25.740 33.955 25.785 ;
        RECT 37.330 25.740 37.650 25.800 ;
        RECT 33.665 25.600 37.650 25.740 ;
        RECT 33.665 25.555 33.955 25.600 ;
        RECT 37.330 25.540 37.650 25.600 ;
        RECT 28.590 25.400 28.910 25.460 ;
        RECT 34.585 25.400 34.875 25.445 ;
        RECT 23.160 25.260 34.875 25.400 ;
        RECT 19.850 25.200 20.170 25.260 ;
        RECT 20.785 25.215 21.075 25.260 ;
        RECT 28.590 25.200 28.910 25.260 ;
        RECT 34.585 25.215 34.875 25.260 ;
        RECT 9.270 24.860 9.590 25.120 ;
        RECT 5.520 24.240 41.400 24.720 ;
        RECT 13.885 24.040 14.175 24.085 ;
        RECT 14.790 24.040 15.110 24.100 ;
        RECT 13.885 23.900 15.110 24.040 ;
        RECT 13.885 23.855 14.175 23.900 ;
        RECT 14.790 23.840 15.110 23.900 ;
        RECT 28.605 24.040 28.895 24.085 ;
        RECT 29.510 24.040 29.830 24.100 ;
        RECT 28.605 23.900 29.830 24.040 ;
        RECT 28.605 23.855 28.895 23.900 ;
        RECT 29.510 23.840 29.830 23.900 ;
        RECT 35.490 24.040 35.810 24.100 ;
        RECT 36.425 24.040 36.715 24.085 ;
        RECT 35.490 23.900 36.715 24.040 ;
        RECT 35.490 23.840 35.810 23.900 ;
        RECT 36.425 23.855 36.715 23.900 ;
        RECT 7.470 23.700 7.760 23.745 ;
        RECT 9.570 23.700 9.860 23.745 ;
        RECT 11.140 23.700 11.430 23.745 ;
        RECT 7.470 23.560 11.430 23.700 ;
        RECT 7.470 23.515 7.760 23.560 ;
        RECT 9.570 23.515 9.860 23.560 ;
        RECT 11.140 23.515 11.430 23.560 ;
        RECT 19.430 23.700 19.720 23.745 ;
        RECT 21.530 23.700 21.820 23.745 ;
        RECT 23.100 23.700 23.390 23.745 ;
        RECT 19.430 23.560 23.390 23.700 ;
        RECT 19.430 23.515 19.720 23.560 ;
        RECT 21.530 23.515 21.820 23.560 ;
        RECT 23.100 23.515 23.390 23.560 ;
        RECT 28.130 23.500 28.450 23.760 ;
        RECT 6.970 23.160 7.290 23.420 ;
        RECT 7.865 23.360 8.155 23.405 ;
        RECT 9.055 23.360 9.345 23.405 ;
        RECT 11.575 23.360 11.865 23.405 ;
        RECT 7.865 23.220 11.865 23.360 ;
        RECT 7.865 23.175 8.155 23.220 ;
        RECT 9.055 23.175 9.345 23.220 ;
        RECT 11.575 23.175 11.865 23.220 ;
        RECT 19.825 23.360 20.115 23.405 ;
        RECT 21.015 23.360 21.305 23.405 ;
        RECT 23.535 23.360 23.825 23.405 ;
        RECT 19.825 23.220 23.825 23.360 ;
        RECT 19.825 23.175 20.115 23.220 ;
        RECT 21.015 23.175 21.305 23.220 ;
        RECT 23.535 23.175 23.825 23.220 ;
        RECT 26.305 23.360 26.595 23.405 ;
        RECT 27.210 23.360 27.530 23.420 ;
        RECT 26.305 23.220 27.530 23.360 ;
        RECT 26.305 23.175 26.595 23.220 ;
        RECT 27.210 23.160 27.530 23.220 ;
        RECT 35.030 23.360 35.350 23.420 ;
        RECT 35.030 23.220 38.940 23.360 ;
        RECT 35.030 23.160 35.350 23.220 ;
        RECT 7.060 23.020 7.200 23.160 ;
        RECT 13.870 23.020 14.190 23.080 ;
        RECT 18.945 23.020 19.235 23.065 ;
        RECT 7.060 22.880 19.235 23.020 ;
        RECT 13.870 22.820 14.190 22.880 ;
        RECT 18.945 22.835 19.235 22.880 ;
        RECT 20.280 22.835 20.570 23.065 ;
        RECT 8.320 22.680 8.610 22.725 ;
        RECT 9.270 22.680 9.590 22.740 ;
        RECT 8.320 22.540 9.590 22.680 ;
        RECT 8.320 22.495 8.610 22.540 ;
        RECT 9.270 22.480 9.590 22.540 ;
        RECT 19.020 22.340 19.160 22.835 ;
        RECT 19.850 22.680 20.170 22.740 ;
        RECT 20.400 22.680 20.540 22.835 ;
        RECT 32.730 22.820 33.050 23.080 ;
        RECT 35.490 23.020 35.810 23.080 ;
        RECT 37.345 23.020 37.635 23.065 ;
        RECT 35.490 22.880 37.635 23.020 ;
        RECT 35.490 22.820 35.810 22.880 ;
        RECT 37.345 22.835 37.635 22.880 ;
        RECT 37.790 22.820 38.110 23.080 ;
        RECT 38.250 22.820 38.570 23.080 ;
        RECT 38.800 23.065 38.940 23.220 ;
        RECT 38.725 22.835 39.015 23.065 ;
        RECT 19.850 22.540 20.540 22.680 ;
        RECT 19.850 22.480 20.170 22.540 ;
        RECT 23.990 22.340 24.310 22.400 ;
        RECT 19.020 22.200 24.310 22.340 ;
        RECT 23.990 22.140 24.310 22.200 ;
        RECT 25.845 22.340 26.135 22.385 ;
        RECT 26.750 22.340 27.070 22.400 ;
        RECT 25.845 22.200 27.070 22.340 ;
        RECT 25.845 22.155 26.135 22.200 ;
        RECT 26.750 22.140 27.070 22.200 ;
        RECT 33.650 22.340 33.970 22.400 ;
        RECT 35.965 22.340 36.255 22.385 ;
        RECT 33.650 22.200 36.255 22.340 ;
        RECT 33.650 22.140 33.970 22.200 ;
        RECT 35.965 22.155 36.255 22.200 ;
        RECT 5.520 21.520 41.400 22.000 ;
        RECT 33.650 21.120 33.970 21.380 ;
        RECT 37.330 21.120 37.650 21.380 ;
        RECT 28.590 20.980 28.910 21.040 ;
        RECT 23.620 20.840 28.910 20.980 ;
        RECT 8.365 20.640 8.655 20.685 ;
        RECT 14.790 20.640 15.110 20.700 ;
        RECT 8.365 20.500 15.110 20.640 ;
        RECT 8.365 20.455 8.655 20.500 ;
        RECT 14.790 20.440 15.110 20.500 ;
        RECT 17.565 20.640 17.855 20.685 ;
        RECT 19.865 20.640 20.155 20.685 ;
        RECT 17.565 20.500 20.155 20.640 ;
        RECT 17.565 20.455 17.855 20.500 ;
        RECT 19.865 20.455 20.155 20.500 ;
        RECT 6.970 20.300 7.290 20.360 ;
        RECT 9.745 20.300 10.035 20.345 ;
        RECT 6.970 20.160 10.035 20.300 ;
        RECT 6.970 20.100 7.290 20.160 ;
        RECT 9.745 20.115 10.035 20.160 ;
        RECT 14.330 20.100 14.650 20.360 ;
        RECT 18.470 20.100 18.790 20.360 ;
        RECT 19.405 20.300 19.695 20.345 ;
        RECT 23.620 20.300 23.760 20.840 ;
        RECT 28.590 20.780 28.910 20.840 ;
        RECT 37.790 20.980 38.110 21.040 ;
        RECT 39.645 20.980 39.935 21.025 ;
        RECT 37.790 20.840 39.935 20.980 ;
        RECT 37.790 20.780 38.110 20.840 ;
        RECT 39.645 20.795 39.935 20.840 ;
        RECT 23.990 20.440 24.310 20.700 ;
        RECT 25.340 20.640 25.630 20.685 ;
        RECT 29.510 20.640 29.830 20.700 ;
        RECT 25.340 20.500 29.280 20.640 ;
        RECT 25.340 20.455 25.630 20.500 ;
        RECT 19.405 20.160 23.760 20.300 ;
        RECT 24.885 20.300 25.175 20.345 ;
        RECT 26.075 20.300 26.365 20.345 ;
        RECT 28.595 20.300 28.885 20.345 ;
        RECT 24.885 20.160 28.885 20.300 ;
        RECT 19.405 20.115 19.695 20.160 ;
        RECT 24.885 20.115 25.175 20.160 ;
        RECT 26.075 20.115 26.365 20.160 ;
        RECT 28.595 20.115 28.885 20.160 ;
        RECT 6.510 19.960 6.830 20.020 ;
        RECT 7.445 19.960 7.735 20.005 ;
        RECT 6.510 19.820 7.735 19.960 ;
        RECT 6.510 19.760 6.830 19.820 ;
        RECT 7.445 19.775 7.735 19.820 ;
        RECT 12.030 19.960 12.350 20.020 ;
        RECT 24.490 19.960 24.780 20.005 ;
        RECT 26.590 19.960 26.880 20.005 ;
        RECT 28.160 19.960 28.450 20.005 ;
        RECT 12.030 19.820 24.220 19.960 ;
        RECT 12.030 19.760 12.350 19.820 ;
        RECT 11.570 19.620 11.890 19.680 ;
        RECT 12.965 19.620 13.255 19.665 ;
        RECT 11.570 19.480 13.255 19.620 ;
        RECT 11.570 19.420 11.890 19.480 ;
        RECT 12.965 19.435 13.255 19.480 ;
        RECT 21.705 19.620 21.995 19.665 ;
        RECT 23.070 19.620 23.390 19.680 ;
        RECT 21.705 19.480 23.390 19.620 ;
        RECT 24.080 19.620 24.220 19.820 ;
        RECT 24.490 19.820 28.450 19.960 ;
        RECT 29.140 19.960 29.280 20.500 ;
        RECT 29.510 20.500 34.800 20.640 ;
        RECT 29.510 20.440 29.830 20.500 ;
        RECT 30.430 20.300 30.750 20.360 ;
        RECT 34.660 20.345 34.800 20.500 ;
        RECT 35.950 20.440 36.270 20.700 ;
        RECT 37.330 20.640 37.650 20.700 ;
        RECT 38.265 20.640 38.555 20.685 ;
        RECT 37.330 20.500 38.555 20.640 ;
        RECT 37.330 20.440 37.650 20.500 ;
        RECT 38.265 20.455 38.555 20.500 ;
        RECT 34.125 20.300 34.415 20.345 ;
        RECT 30.430 20.160 34.415 20.300 ;
        RECT 30.430 20.100 30.750 20.160 ;
        RECT 34.125 20.115 34.415 20.160 ;
        RECT 34.585 20.115 34.875 20.345 ;
        RECT 35.490 20.300 35.810 20.360 ;
        RECT 38.710 20.300 39.030 20.360 ;
        RECT 35.490 20.160 39.030 20.300 ;
        RECT 35.490 20.100 35.810 20.160 ;
        RECT 38.710 20.100 39.030 20.160 ;
        RECT 31.825 19.960 32.115 20.005 ;
        RECT 29.140 19.820 32.115 19.960 ;
        RECT 24.490 19.775 24.780 19.820 ;
        RECT 26.590 19.775 26.880 19.820 ;
        RECT 28.160 19.775 28.450 19.820 ;
        RECT 31.825 19.775 32.115 19.820 ;
        RECT 36.885 19.960 37.175 20.005 ;
        RECT 39.630 19.960 39.950 20.020 ;
        RECT 36.885 19.820 39.950 19.960 ;
        RECT 36.885 19.775 37.175 19.820 ;
        RECT 39.630 19.760 39.950 19.820 ;
        RECT 30.430 19.620 30.750 19.680 ;
        RECT 24.080 19.480 30.750 19.620 ;
        RECT 21.705 19.435 21.995 19.480 ;
        RECT 23.070 19.420 23.390 19.480 ;
        RECT 30.430 19.420 30.750 19.480 ;
        RECT 30.905 19.620 31.195 19.665 ;
        RECT 32.730 19.620 33.050 19.680 ;
        RECT 30.905 19.480 33.050 19.620 ;
        RECT 30.905 19.435 31.195 19.480 ;
        RECT 32.730 19.420 33.050 19.480 ;
        RECT 36.410 19.620 36.730 19.680 ;
        RECT 38.265 19.620 38.555 19.665 ;
        RECT 36.410 19.480 38.555 19.620 ;
        RECT 36.410 19.420 36.730 19.480 ;
        RECT 38.265 19.435 38.555 19.480 ;
        RECT 5.520 18.800 41.400 19.280 ;
        RECT 6.970 18.400 7.290 18.660 ;
        RECT 23.990 18.600 24.310 18.660 ;
        RECT 25.385 18.600 25.675 18.645 ;
        RECT 23.990 18.460 25.675 18.600 ;
        RECT 23.990 18.400 24.310 18.460 ;
        RECT 25.385 18.415 25.675 18.460 ;
        RECT 33.205 18.600 33.495 18.645 ;
        RECT 35.490 18.600 35.810 18.660 ;
        RECT 33.205 18.460 35.810 18.600 ;
        RECT 33.205 18.415 33.495 18.460 ;
        RECT 35.490 18.400 35.810 18.460 ;
        RECT 36.425 18.600 36.715 18.645 ;
        RECT 36.870 18.600 37.190 18.660 ;
        RECT 36.425 18.460 37.190 18.600 ;
        RECT 36.425 18.415 36.715 18.460 ;
        RECT 36.870 18.400 37.190 18.460 ;
        RECT 9.730 18.260 10.020 18.305 ;
        RECT 11.300 18.260 11.590 18.305 ;
        RECT 13.400 18.260 13.690 18.305 ;
        RECT 9.730 18.120 13.690 18.260 ;
        RECT 9.730 18.075 10.020 18.120 ;
        RECT 11.300 18.075 11.590 18.120 ;
        RECT 13.400 18.075 13.690 18.120 ;
        RECT 30.445 18.260 30.735 18.305 ;
        RECT 35.950 18.260 36.270 18.320 ;
        RECT 30.445 18.120 36.270 18.260 ;
        RECT 30.445 18.075 30.735 18.120 ;
        RECT 35.950 18.060 36.270 18.120 ;
        RECT 9.295 17.920 9.585 17.965 ;
        RECT 11.815 17.920 12.105 17.965 ;
        RECT 13.005 17.920 13.295 17.965 ;
        RECT 9.295 17.780 13.295 17.920 ;
        RECT 9.295 17.735 9.585 17.780 ;
        RECT 11.815 17.735 12.105 17.780 ;
        RECT 13.005 17.735 13.295 17.780 ;
        RECT 13.870 17.720 14.190 17.980 ;
        RECT 39.170 17.920 39.490 17.980 ;
        RECT 29.600 17.780 39.490 17.920 ;
        RECT 18.945 17.580 19.235 17.625 ;
        RECT 23.530 17.580 23.850 17.640 ;
        RECT 29.600 17.625 29.740 17.780 ;
        RECT 39.170 17.720 39.490 17.780 ;
        RECT 18.945 17.440 23.850 17.580 ;
        RECT 18.945 17.395 19.235 17.440 ;
        RECT 23.530 17.380 23.850 17.440 ;
        RECT 29.525 17.395 29.815 17.625 ;
        RECT 30.890 17.380 31.210 17.640 ;
        RECT 32.270 17.380 32.590 17.640 ;
        RECT 33.650 17.380 33.970 17.640 ;
        RECT 35.045 17.395 35.335 17.625 ;
        RECT 35.965 17.580 36.255 17.625 ;
        RECT 36.410 17.580 36.730 17.640 ;
        RECT 35.965 17.440 36.730 17.580 ;
        RECT 35.965 17.395 36.255 17.440 ;
        RECT 9.730 17.240 10.050 17.300 ;
        RECT 12.550 17.240 12.840 17.285 ;
        RECT 35.120 17.240 35.260 17.395 ;
        RECT 36.410 17.380 36.730 17.440 ;
        RECT 37.330 17.380 37.650 17.640 ;
        RECT 38.710 17.380 39.030 17.640 ;
        RECT 39.630 17.380 39.950 17.640 ;
        RECT 37.420 17.240 37.560 17.380 ;
        RECT 9.730 17.100 12.840 17.240 ;
        RECT 9.730 17.040 10.050 17.100 ;
        RECT 12.550 17.055 12.840 17.100 ;
        RECT 31.900 17.100 37.560 17.240 ;
        RECT 31.900 16.945 32.040 17.100 ;
        RECT 31.825 16.715 32.115 16.945 ;
        RECT 34.585 16.900 34.875 16.945 ;
        RECT 35.030 16.900 35.350 16.960 ;
        RECT 34.585 16.760 35.350 16.900 ;
        RECT 34.585 16.715 34.875 16.760 ;
        RECT 35.030 16.700 35.350 16.760 ;
        RECT 35.490 16.700 35.810 16.960 ;
        RECT 5.520 16.080 41.400 16.560 ;
        RECT 9.730 15.680 10.050 15.940 ;
        RECT 11.570 15.680 11.890 15.940 ;
        RECT 12.030 15.680 12.350 15.940 ;
        RECT 14.330 15.880 14.650 15.940 ;
        RECT 16.630 15.880 16.950 15.940 ;
        RECT 18.945 15.880 19.235 15.925 ;
        RECT 14.330 15.740 19.235 15.880 ;
        RECT 14.330 15.680 14.650 15.740 ;
        RECT 16.630 15.680 16.950 15.740 ;
        RECT 18.945 15.695 19.235 15.740 ;
        RECT 23.070 15.680 23.390 15.940 ;
        RECT 28.590 15.680 28.910 15.940 ;
        RECT 38.250 15.880 38.570 15.940 ;
        RECT 38.725 15.880 39.015 15.925 ;
        RECT 38.250 15.740 39.015 15.880 ;
        RECT 38.250 15.680 38.570 15.740 ;
        RECT 38.725 15.695 39.015 15.740 ;
        RECT 6.970 15.200 7.290 15.260 ;
        RECT 8.365 15.200 8.655 15.245 ;
        RECT 6.970 15.060 8.655 15.200 ;
        RECT 23.160 15.200 23.300 15.680 ;
        RECT 23.990 15.540 24.310 15.600 ;
        RECT 23.990 15.400 26.060 15.540 ;
        RECT 23.990 15.340 24.310 15.400 ;
        RECT 25.920 15.245 26.060 15.400 ;
        RECT 24.510 15.200 24.800 15.245 ;
        RECT 23.160 15.060 24.800 15.200 ;
        RECT 6.970 15.000 7.290 15.060 ;
        RECT 8.365 15.015 8.655 15.060 ;
        RECT 24.510 15.015 24.800 15.060 ;
        RECT 25.845 15.015 26.135 15.245 ;
        RECT 28.145 15.200 28.435 15.245 ;
        RECT 31.825 15.200 32.115 15.245 ;
        RECT 28.145 15.060 32.115 15.200 ;
        RECT 28.145 15.015 28.435 15.060 ;
        RECT 31.825 15.015 32.115 15.060 ;
        RECT 35.490 15.200 35.810 15.260 ;
        RECT 37.805 15.200 38.095 15.245 ;
        RECT 35.490 15.060 38.095 15.200 ;
        RECT 35.490 15.000 35.810 15.060 ;
        RECT 37.805 15.015 38.095 15.060 ;
        RECT 12.965 14.860 13.255 14.905 ;
        RECT 18.470 14.860 18.790 14.920 ;
        RECT 12.965 14.720 18.790 14.860 ;
        RECT 12.965 14.675 13.255 14.720 ;
        RECT 18.470 14.660 18.790 14.720 ;
        RECT 21.255 14.860 21.545 14.905 ;
        RECT 23.775 14.860 24.065 14.905 ;
        RECT 24.965 14.860 25.255 14.905 ;
        RECT 21.255 14.720 25.255 14.860 ;
        RECT 21.255 14.675 21.545 14.720 ;
        RECT 23.775 14.675 24.065 14.720 ;
        RECT 24.965 14.675 25.255 14.720 ;
        RECT 29.510 14.660 29.830 14.920 ;
        RECT 29.970 14.860 30.290 14.920 ;
        RECT 34.585 14.860 34.875 14.905 ;
        RECT 29.970 14.720 34.875 14.860 ;
        RECT 29.970 14.660 30.290 14.720 ;
        RECT 34.585 14.675 34.875 14.720 ;
        RECT 35.030 14.860 35.350 14.920 ;
        RECT 36.425 14.860 36.715 14.905 ;
        RECT 35.030 14.720 36.715 14.860 ;
        RECT 35.030 14.660 35.350 14.720 ;
        RECT 36.425 14.675 36.715 14.720 ;
        RECT 36.885 14.860 37.175 14.905 ;
        RECT 39.630 14.860 39.950 14.920 ;
        RECT 36.885 14.720 39.950 14.860 ;
        RECT 36.885 14.675 37.175 14.720 ;
        RECT 39.630 14.660 39.950 14.720 ;
        RECT 4.210 14.520 4.530 14.580 ;
        RECT 7.445 14.520 7.735 14.565 ;
        RECT 4.210 14.380 7.735 14.520 ;
        RECT 4.210 14.320 4.530 14.380 ;
        RECT 7.445 14.335 7.735 14.380 ;
        RECT 21.690 14.520 21.980 14.565 ;
        RECT 23.260 14.520 23.550 14.565 ;
        RECT 25.360 14.520 25.650 14.565 ;
        RECT 21.690 14.380 25.650 14.520 ;
        RECT 21.690 14.335 21.980 14.380 ;
        RECT 23.260 14.335 23.550 14.380 ;
        RECT 25.360 14.335 25.650 14.380 ;
        RECT 23.990 14.180 24.310 14.240 ;
        RECT 26.305 14.180 26.595 14.225 ;
        RECT 23.990 14.040 26.595 14.180 ;
        RECT 23.990 13.980 24.310 14.040 ;
        RECT 26.305 13.995 26.595 14.040 ;
        RECT 5.520 13.360 41.400 13.840 ;
        RECT 26.750 13.160 27.070 13.220 ;
        RECT 20.860 13.020 27.070 13.160 ;
        RECT 16.630 11.940 16.950 12.200 ;
        RECT 20.860 12.185 21.000 13.020 ;
        RECT 26.750 12.960 27.070 13.020 ;
        RECT 34.585 13.160 34.875 13.205 ;
        RECT 36.410 13.160 36.730 13.220 ;
        RECT 34.585 13.020 36.730 13.160 ;
        RECT 34.585 12.975 34.875 13.020 ;
        RECT 36.410 12.960 36.730 13.020 ;
        RECT 38.710 13.160 39.030 13.220 ;
        RECT 39.185 13.160 39.475 13.205 ;
        RECT 38.710 13.020 39.475 13.160 ;
        RECT 38.710 12.960 39.030 13.020 ;
        RECT 39.185 12.975 39.475 13.020 ;
        RECT 21.730 12.820 22.020 12.865 ;
        RECT 23.830 12.820 24.120 12.865 ;
        RECT 25.400 12.820 25.690 12.865 ;
        RECT 21.730 12.680 25.690 12.820 ;
        RECT 21.730 12.635 22.020 12.680 ;
        RECT 23.830 12.635 24.120 12.680 ;
        RECT 25.400 12.635 25.690 12.680 ;
        RECT 28.145 12.820 28.435 12.865 ;
        RECT 29.970 12.820 30.290 12.880 ;
        RECT 28.145 12.680 30.290 12.820 ;
        RECT 28.145 12.635 28.435 12.680 ;
        RECT 29.970 12.620 30.290 12.680 ;
        RECT 35.950 12.820 36.270 12.880 ;
        RECT 38.265 12.820 38.555 12.865 ;
        RECT 35.950 12.680 38.555 12.820 ;
        RECT 35.950 12.620 36.270 12.680 ;
        RECT 38.265 12.635 38.555 12.680 ;
        RECT 22.125 12.480 22.415 12.525 ;
        RECT 23.315 12.480 23.605 12.525 ;
        RECT 25.835 12.480 26.125 12.525 ;
        RECT 22.125 12.340 26.125 12.480 ;
        RECT 22.125 12.295 22.415 12.340 ;
        RECT 23.315 12.295 23.605 12.340 ;
        RECT 25.835 12.295 26.125 12.340 ;
        RECT 35.030 12.480 35.350 12.540 ;
        RECT 36.885 12.480 37.175 12.525 ;
        RECT 35.030 12.340 37.175 12.480 ;
        RECT 35.030 12.280 35.350 12.340 ;
        RECT 36.885 12.295 37.175 12.340 ;
        RECT 20.785 11.955 21.075 12.185 ;
        RECT 21.245 12.140 21.535 12.185 ;
        RECT 21.690 12.140 22.010 12.200 ;
        RECT 21.245 12.000 22.010 12.140 ;
        RECT 21.245 11.955 21.535 12.000 ;
        RECT 21.690 11.940 22.010 12.000 ;
        RECT 29.970 11.940 30.290 12.200 ;
        RECT 32.730 11.940 33.050 12.200 ;
        RECT 35.490 11.940 35.810 12.200 ;
        RECT 22.580 11.800 22.870 11.845 ;
        RECT 23.990 11.800 24.310 11.860 ;
        RECT 22.580 11.660 24.310 11.800 ;
        RECT 22.580 11.615 22.870 11.660 ;
        RECT 23.990 11.600 24.310 11.660 ;
        RECT 26.380 11.660 29.280 11.800 ;
        RECT 26.380 11.520 26.520 11.660 ;
        RECT 17.565 11.460 17.855 11.505 ;
        RECT 19.390 11.460 19.710 11.520 ;
        RECT 17.565 11.320 19.710 11.460 ;
        RECT 17.565 11.275 17.855 11.320 ;
        RECT 19.390 11.260 19.710 11.320 ;
        RECT 19.865 11.460 20.155 11.505 ;
        RECT 22.150 11.460 22.470 11.520 ;
        RECT 19.865 11.320 22.470 11.460 ;
        RECT 19.865 11.275 20.155 11.320 ;
        RECT 22.150 11.260 22.470 11.320 ;
        RECT 26.290 11.260 26.610 11.520 ;
        RECT 29.140 11.505 29.280 11.660 ;
        RECT 29.065 11.275 29.355 11.505 ;
        RECT 32.270 11.460 32.590 11.520 ;
        RECT 33.665 11.460 33.955 11.505 ;
        RECT 32.270 11.320 33.955 11.460 ;
        RECT 32.270 11.260 32.590 11.320 ;
        RECT 33.665 11.275 33.955 11.320 ;
        RECT 5.520 10.640 41.400 11.120 ;
      LAYER met2 ;
        RECT 19.480 45.890 19.620 53.765 ;
        RECT 22.700 47.330 22.840 53.765 ;
        RECT 22.700 47.190 23.760 47.330 ;
        RECT 21.070 46.055 22.610 46.425 ;
        RECT 19.420 45.570 19.680 45.890 ;
        RECT 11.140 44.550 11.400 44.870 ;
        RECT 15.740 44.550 16.000 44.870 ;
        RECT 16.200 44.550 16.460 44.870 ;
        RECT 11.200 43.170 11.340 44.550 ;
        RECT 15.800 43.170 15.940 44.550 ;
        RECT 11.140 42.850 11.400 43.170 ;
        RECT 15.740 42.850 16.000 43.170 ;
        RECT 16.260 42.685 16.400 44.550 ;
        RECT 18.040 43.870 18.300 44.190 ;
        RECT 23.100 43.870 23.360 44.190 ;
        RECT 18.100 42.830 18.240 43.870 ;
        RECT 16.190 42.315 16.470 42.685 ;
        RECT 18.040 42.510 18.300 42.830 ;
        RECT 18.960 42.170 19.220 42.490 ;
        RECT 20.330 42.315 20.610 42.685 ;
        RECT 16.660 41.150 16.920 41.470 ;
        RECT 16.720 39.430 16.860 41.150 ;
        RECT 17.570 40.955 17.850 41.325 ;
        RECT 16.660 39.110 16.920 39.430 ;
        RECT 8.840 38.770 9.100 39.090 ;
        RECT 6.530 37.555 6.810 37.925 ;
        RECT 8.900 37.730 9.040 38.770 ;
        RECT 13.900 38.430 14.160 38.750 ;
        RECT 14.360 38.430 14.620 38.750 ;
        RECT 6.540 37.410 6.800 37.555 ;
        RECT 8.840 37.410 9.100 37.730 ;
        RECT 13.960 37.050 14.100 38.430 ;
        RECT 14.420 37.730 14.560 38.430 ;
        RECT 16.720 37.730 16.860 39.110 ;
        RECT 14.360 37.410 14.620 37.730 ;
        RECT 16.660 37.410 16.920 37.730 ;
        RECT 13.900 36.730 14.160 37.050 ;
        RECT 12.520 36.390 12.780 36.710 ;
        RECT 9.300 36.050 9.560 36.370 ;
        RECT 9.360 34.330 9.500 36.050 ;
        RECT 9.300 34.010 9.560 34.330 ;
        RECT 12.580 33.650 12.720 36.390 ;
        RECT 16.720 33.990 16.860 37.410 ;
        RECT 13.900 33.670 14.160 33.990 ;
        RECT 16.660 33.670 16.920 33.990 ;
        RECT 12.520 33.330 12.780 33.650 ;
        RECT 7.000 32.990 7.260 33.310 ;
        RECT 11.600 32.990 11.860 33.310 ;
        RECT 7.060 31.950 7.200 32.990 ;
        RECT 7.000 31.630 7.260 31.950 ;
        RECT 6.530 30.755 6.810 31.125 ;
        RECT 6.600 26.850 6.740 30.755 ;
        RECT 7.000 30.270 7.260 30.590 ;
        RECT 7.060 28.890 7.200 30.270 ;
        RECT 11.660 29.570 11.800 32.990 ;
        RECT 11.600 29.250 11.860 29.570 ;
        RECT 7.000 28.570 7.260 28.890 ;
        RECT 6.540 26.530 6.800 26.850 ;
        RECT 7.060 26.170 7.200 28.570 ;
        RECT 12.060 27.550 12.320 27.870 ;
        RECT 12.120 26.850 12.260 27.550 ;
        RECT 12.060 26.530 12.320 26.850 ;
        RECT 7.000 25.850 7.260 26.170 ;
        RECT 12.580 25.830 12.720 33.330 ;
        RECT 13.960 31.610 14.100 33.670 ;
        RECT 17.640 31.950 17.780 40.955 ;
        RECT 19.020 40.450 19.160 42.170 ;
        RECT 18.960 40.130 19.220 40.450 ;
        RECT 18.960 37.410 19.220 37.730 ;
        RECT 19.880 37.410 20.140 37.730 ;
        RECT 19.020 34.330 19.160 37.410 ;
        RECT 19.940 35.010 20.080 37.410 ;
        RECT 19.880 34.690 20.140 35.010 ;
        RECT 18.960 34.010 19.220 34.330 ;
        RECT 17.580 31.630 17.840 31.950 ;
        RECT 13.900 31.290 14.160 31.610 ;
        RECT 19.940 29.570 20.080 34.690 ;
        RECT 20.400 29.570 20.540 42.315 ;
        RECT 21.070 40.615 22.610 40.985 ;
        RECT 23.160 39.430 23.300 43.870 ;
        RECT 23.620 41.810 23.760 47.190 ;
        RECT 25.920 45.890 26.060 53.765 ;
        RECT 25.860 45.570 26.120 45.890 ;
        RECT 24.020 45.230 24.280 45.550 ;
        RECT 23.560 41.490 23.820 41.810 ;
        RECT 24.080 40.450 24.220 45.230 ;
        RECT 29.140 44.870 29.280 53.765 ;
        RECT 32.360 45.890 32.500 53.765 ;
        RECT 39.650 51.155 39.930 51.525 ;
        RECT 36.890 47.755 37.170 48.125 ;
        RECT 32.300 45.570 32.560 45.890 ;
        RECT 30.920 45.230 31.180 45.550 ;
        RECT 26.320 44.550 26.580 44.870 ;
        RECT 29.080 44.550 29.340 44.870 ;
        RECT 24.370 43.335 25.910 43.705 ;
        RECT 26.380 43.170 26.520 44.550 ;
        RECT 26.780 43.870 27.040 44.190 ;
        RECT 26.320 42.850 26.580 43.170 ;
        RECT 26.840 42.830 26.980 43.870 ;
        RECT 26.780 42.510 27.040 42.830 ;
        RECT 30.980 42.490 31.120 45.230 ;
        RECT 36.960 44.870 37.100 47.755 ;
        RECT 39.720 44.870 39.860 51.155 ;
        RECT 34.140 44.550 34.400 44.870 ;
        RECT 36.900 44.550 37.160 44.870 ;
        RECT 38.280 44.725 38.540 44.870 ;
        RECT 32.760 43.870 33.020 44.190 ;
        RECT 27.700 42.170 27.960 42.490 ;
        RECT 29.080 42.170 29.340 42.490 ;
        RECT 30.920 42.170 31.180 42.490 ;
        RECT 24.480 41.830 24.740 42.150 ;
        RECT 24.020 40.130 24.280 40.450 ;
        RECT 24.540 39.430 24.680 41.830 ;
        RECT 27.240 41.150 27.500 41.470 ;
        RECT 27.300 39.770 27.440 41.150 ;
        RECT 27.240 39.450 27.500 39.770 ;
        RECT 27.760 39.430 27.900 42.170 ;
        RECT 28.620 41.830 28.880 42.150 ;
        RECT 23.100 39.110 23.360 39.430 ;
        RECT 23.560 39.110 23.820 39.430 ;
        RECT 24.480 39.110 24.740 39.430 ;
        RECT 26.320 39.110 26.580 39.430 ;
        RECT 26.780 39.110 27.040 39.430 ;
        RECT 27.700 39.110 27.960 39.430 ;
        RECT 23.100 38.430 23.360 38.750 ;
        RECT 21.070 35.175 22.610 35.545 ;
        RECT 21.070 29.735 22.610 30.105 ;
        RECT 19.880 29.250 20.140 29.570 ;
        RECT 20.340 29.250 20.600 29.570 ;
        RECT 14.820 28.230 15.080 28.550 ;
        RECT 12.060 25.510 12.320 25.830 ;
        RECT 12.520 25.510 12.780 25.830 ;
        RECT 7.000 25.170 7.260 25.490 ;
        RECT 6.530 23.955 6.810 24.325 ;
        RECT 6.600 20.050 6.740 23.955 ;
        RECT 7.060 23.450 7.200 25.170 ;
        RECT 9.300 24.830 9.560 25.150 ;
        RECT 7.000 23.130 7.260 23.450 ;
        RECT 9.360 22.770 9.500 24.830 ;
        RECT 9.300 22.450 9.560 22.770 ;
        RECT 7.000 20.070 7.260 20.390 ;
        RECT 6.540 19.730 6.800 20.050 ;
        RECT 7.060 18.690 7.200 20.070 ;
        RECT 12.120 20.050 12.260 25.510 ;
        RECT 14.880 24.130 15.020 28.230 ;
        RECT 19.940 26.510 20.080 29.250 ;
        RECT 23.160 28.550 23.300 38.430 ;
        RECT 23.620 37.730 23.760 39.110 ;
        RECT 24.370 37.895 25.910 38.265 ;
        RECT 23.560 37.410 23.820 37.730 ;
        RECT 23.560 36.730 23.820 37.050 ;
        RECT 23.620 30.590 23.760 36.730 ;
        RECT 24.020 35.710 24.280 36.030 ;
        RECT 24.080 31.690 24.220 35.710 ;
        RECT 26.380 35.010 26.520 39.110 ;
        RECT 26.320 34.690 26.580 35.010 ;
        RECT 26.840 34.410 26.980 39.110 ;
        RECT 28.680 37.390 28.820 41.830 ;
        RECT 29.140 40.450 29.280 42.170 ;
        RECT 30.000 41.150 30.260 41.470 ;
        RECT 29.080 40.130 29.340 40.450 ;
        RECT 29.140 39.850 29.280 40.130 ;
        RECT 29.140 39.710 29.740 39.850 ;
        RECT 29.080 38.770 29.340 39.090 ;
        RECT 28.620 37.070 28.880 37.390 ;
        RECT 27.240 36.390 27.500 36.710 ;
        RECT 26.380 34.270 26.980 34.410 ;
        RECT 26.380 33.310 26.520 34.270 ;
        RECT 27.300 33.990 27.440 36.390 ;
        RECT 27.700 34.350 27.960 34.670 ;
        RECT 27.240 33.670 27.500 33.990 ;
        RECT 26.780 33.330 27.040 33.650 ;
        RECT 26.320 32.990 26.580 33.310 ;
        RECT 24.370 32.455 25.910 32.825 ;
        RECT 24.080 31.550 24.680 31.690 ;
        RECT 24.020 30.950 24.280 31.270 ;
        RECT 23.560 30.270 23.820 30.590 ;
        RECT 20.340 28.230 20.600 28.550 ;
        RECT 23.100 28.230 23.360 28.550 ;
        RECT 20.400 26.850 20.540 28.230 ;
        RECT 20.340 26.530 20.600 26.850 ;
        RECT 18.500 26.190 18.760 26.510 ;
        RECT 19.880 26.190 20.140 26.510 ;
        RECT 14.820 23.810 15.080 24.130 ;
        RECT 13.900 22.790 14.160 23.110 ;
        RECT 12.060 19.730 12.320 20.050 ;
        RECT 11.600 19.390 11.860 19.710 ;
        RECT 7.000 18.370 7.260 18.690 ;
        RECT 7.060 15.290 7.200 18.370 ;
        RECT 9.760 17.010 10.020 17.330 ;
        RECT 9.820 15.970 9.960 17.010 ;
        RECT 11.660 15.970 11.800 19.390 ;
        RECT 12.120 15.970 12.260 19.730 ;
        RECT 13.960 18.010 14.100 22.790 ;
        RECT 14.880 20.730 15.020 23.810 ;
        RECT 14.820 20.410 15.080 20.730 ;
        RECT 18.560 20.390 18.700 26.190 ;
        RECT 19.880 25.170 20.140 25.490 ;
        RECT 19.940 22.770 20.080 25.170 ;
        RECT 21.070 24.295 22.610 24.665 ;
        RECT 19.880 22.450 20.140 22.770 ;
        RECT 14.360 20.070 14.620 20.390 ;
        RECT 18.500 20.070 18.760 20.390 ;
        RECT 13.900 17.690 14.160 18.010 ;
        RECT 14.420 15.970 14.560 20.070 ;
        RECT 9.760 15.650 10.020 15.970 ;
        RECT 11.600 15.650 11.860 15.970 ;
        RECT 12.060 15.650 12.320 15.970 ;
        RECT 14.360 15.650 14.620 15.970 ;
        RECT 16.660 15.650 16.920 15.970 ;
        RECT 7.000 14.970 7.260 15.290 ;
        RECT 4.230 14.435 4.510 14.805 ;
        RECT 4.240 14.290 4.500 14.435 ;
        RECT 16.720 12.230 16.860 15.650 ;
        RECT 18.560 14.950 18.700 20.070 ;
        RECT 23.100 19.390 23.360 19.710 ;
        RECT 21.070 18.855 22.610 19.225 ;
        RECT 23.160 15.970 23.300 19.390 ;
        RECT 23.620 17.670 23.760 30.270 ;
        RECT 24.080 28.550 24.220 30.950 ;
        RECT 24.540 29.230 24.680 31.550 ;
        RECT 24.480 28.910 24.740 29.230 ;
        RECT 24.020 28.230 24.280 28.550 ;
        RECT 24.370 27.015 25.910 27.385 ;
        RECT 26.380 25.830 26.520 32.990 ;
        RECT 26.840 32.290 26.980 33.330 ;
        RECT 26.780 31.970 27.040 32.290 ;
        RECT 27.760 28.890 27.900 34.350 ;
        RECT 28.160 33.330 28.420 33.650 ;
        RECT 27.700 28.570 27.960 28.890 ;
        RECT 27.240 26.760 27.500 26.850 ;
        RECT 27.760 26.760 27.900 28.570 ;
        RECT 27.240 26.620 27.900 26.760 ;
        RECT 27.240 26.530 27.500 26.620 ;
        RECT 26.320 25.510 26.580 25.830 ;
        RECT 26.780 25.510 27.040 25.830 ;
        RECT 26.840 22.430 26.980 25.510 ;
        RECT 27.760 23.530 27.900 26.620 ;
        RECT 28.220 23.790 28.360 33.330 ;
        RECT 28.680 30.590 28.820 37.070 ;
        RECT 29.140 36.370 29.280 38.770 ;
        RECT 29.080 36.050 29.340 36.370 ;
        RECT 29.140 32.290 29.280 36.050 ;
        RECT 29.080 31.970 29.340 32.290 ;
        RECT 28.620 30.270 28.880 30.590 ;
        RECT 28.680 29.230 28.820 30.270 ;
        RECT 28.620 28.910 28.880 29.230 ;
        RECT 28.620 25.170 28.880 25.490 ;
        RECT 27.300 23.450 27.900 23.530 ;
        RECT 28.160 23.470 28.420 23.790 ;
        RECT 27.240 23.390 27.900 23.450 ;
        RECT 27.240 23.130 27.500 23.390 ;
        RECT 24.020 22.110 24.280 22.430 ;
        RECT 26.780 22.110 27.040 22.430 ;
        RECT 24.080 20.730 24.220 22.110 ;
        RECT 24.370 21.575 25.910 21.945 ;
        RECT 24.020 20.410 24.280 20.730 ;
        RECT 24.080 18.690 24.220 20.410 ;
        RECT 24.020 18.370 24.280 18.690 ;
        RECT 23.560 17.350 23.820 17.670 ;
        RECT 23.100 15.650 23.360 15.970 ;
        RECT 24.080 15.630 24.220 18.370 ;
        RECT 24.370 16.135 25.910 16.505 ;
        RECT 24.020 15.370 24.280 15.630 ;
        RECT 23.160 15.310 24.280 15.370 ;
        RECT 23.160 15.230 24.220 15.310 ;
        RECT 18.500 14.630 18.760 14.950 ;
        RECT 21.070 13.415 22.610 13.785 ;
        RECT 16.660 11.910 16.920 12.230 ;
        RECT 21.720 12.140 21.980 12.230 ;
        RECT 23.160 12.140 23.300 15.230 ;
        RECT 24.020 13.950 24.280 14.270 ;
        RECT 21.720 12.000 23.300 12.140 ;
        RECT 21.720 11.910 21.980 12.000 ;
        RECT 24.080 11.890 24.220 13.950 ;
        RECT 26.840 13.250 26.980 22.110 ;
        RECT 28.680 21.070 28.820 25.170 ;
        RECT 29.600 24.130 29.740 39.710 ;
        RECT 30.060 39.430 30.200 41.150 ;
        RECT 30.000 39.110 30.260 39.430 ;
        RECT 32.820 37.050 32.960 43.870 ;
        RECT 33.670 42.400 33.950 42.685 ;
        RECT 33.280 42.315 33.950 42.400 ;
        RECT 33.280 42.260 33.940 42.315 ;
        RECT 33.280 37.390 33.420 42.260 ;
        RECT 33.680 42.170 33.940 42.260 ;
        RECT 34.200 41.810 34.340 44.550 ;
        RECT 38.270 44.355 38.550 44.725 ;
        RECT 39.660 44.550 39.920 44.870 ;
        RECT 36.440 43.870 36.700 44.190 ;
        RECT 39.200 43.870 39.460 44.190 ;
        RECT 34.140 41.490 34.400 41.810 ;
        RECT 34.200 40.450 34.340 41.490 ;
        RECT 35.980 41.150 36.240 41.470 ;
        RECT 34.140 40.130 34.400 40.450 ;
        RECT 36.040 39.430 36.180 41.150 ;
        RECT 35.980 39.110 36.240 39.430 ;
        RECT 36.500 37.730 36.640 43.870 ;
        RECT 36.900 42.170 37.160 42.490 ;
        RECT 36.960 40.450 37.100 42.170 ;
        RECT 37.360 41.490 37.620 41.810 ;
        RECT 36.900 40.130 37.160 40.450 ;
        RECT 37.420 39.850 37.560 41.490 ;
        RECT 36.960 39.710 37.560 39.850 ;
        RECT 36.440 37.410 36.700 37.730 ;
        RECT 33.220 37.070 33.480 37.390 ;
        RECT 33.680 37.070 33.940 37.390 ;
        RECT 32.760 36.730 33.020 37.050 ;
        RECT 30.920 35.710 31.180 36.030 ;
        RECT 30.980 29.570 31.120 35.710 ;
        RECT 31.840 32.990 32.100 33.310 ;
        RECT 31.900 31.610 32.040 32.990 ;
        RECT 32.820 31.610 32.960 36.730 ;
        RECT 33.740 36.370 33.880 37.070 ;
        RECT 36.500 37.050 36.640 37.410 ;
        RECT 36.440 36.730 36.700 37.050 ;
        RECT 33.680 36.050 33.940 36.370 ;
        RECT 33.740 33.990 33.880 36.050 ;
        RECT 34.600 34.350 34.860 34.670 ;
        RECT 33.680 33.670 33.940 33.990 ;
        RECT 31.840 31.290 32.100 31.610 ;
        RECT 32.760 31.290 33.020 31.610 ;
        RECT 30.920 29.250 31.180 29.570 ;
        RECT 30.460 27.550 30.720 27.870 ;
        RECT 29.540 23.810 29.800 24.130 ;
        RECT 28.620 20.750 28.880 21.070 ;
        RECT 28.680 15.970 28.820 20.750 ;
        RECT 29.600 20.730 29.740 23.810 ;
        RECT 29.540 20.410 29.800 20.730 ;
        RECT 28.620 15.650 28.880 15.970 ;
        RECT 29.600 14.950 29.740 20.410 ;
        RECT 30.520 20.390 30.660 27.550 ;
        RECT 30.980 26.170 31.120 29.250 ;
        RECT 34.660 28.970 34.800 34.350 ;
        RECT 35.520 34.010 35.780 34.330 ;
        RECT 35.060 30.270 35.320 30.590 ;
        RECT 33.740 28.830 34.800 28.970 ;
        RECT 33.740 28.550 33.880 28.830 ;
        RECT 33.680 28.230 33.940 28.550 ;
        RECT 34.600 28.230 34.860 28.550 ;
        RECT 33.220 27.550 33.480 27.870 ;
        RECT 34.660 27.725 34.800 28.230 ;
        RECT 35.120 28.210 35.260 30.270 ;
        RECT 35.060 27.890 35.320 28.210 ;
        RECT 33.280 26.170 33.420 27.550 ;
        RECT 34.590 27.355 34.870 27.725 ;
        RECT 35.120 26.510 35.260 27.890 ;
        RECT 35.060 26.190 35.320 26.510 ;
        RECT 30.920 25.850 31.180 26.170 ;
        RECT 33.220 25.850 33.480 26.170 ;
        RECT 32.290 23.955 32.570 24.325 ;
        RECT 30.460 20.070 30.720 20.390 ;
        RECT 30.520 19.710 30.660 20.070 ;
        RECT 30.460 19.390 30.720 19.710 ;
        RECT 32.360 17.670 32.500 23.955 ;
        RECT 35.120 23.450 35.260 26.190 ;
        RECT 35.580 24.130 35.720 34.010 ;
        RECT 36.500 33.990 36.640 36.730 ;
        RECT 36.960 33.990 37.100 39.710 ;
        RECT 37.360 39.110 37.620 39.430 ;
        RECT 37.420 34.525 37.560 39.110 ;
        RECT 38.280 38.430 38.540 38.750 ;
        RECT 38.740 38.430 39.000 38.750 ;
        RECT 37.820 36.730 38.080 37.050 ;
        RECT 37.880 35.010 38.020 36.730 ;
        RECT 37.820 34.690 38.080 35.010 ;
        RECT 37.350 34.155 37.630 34.525 ;
        RECT 38.340 34.410 38.480 38.430 ;
        RECT 38.800 37.730 38.940 38.430 ;
        RECT 38.740 37.410 39.000 37.730 ;
        RECT 39.260 37.050 39.400 43.870 ;
        RECT 39.660 42.170 39.920 42.490 ;
        RECT 39.720 41.325 39.860 42.170 ;
        RECT 39.650 40.955 39.930 41.325 ;
        RECT 39.660 39.110 39.920 39.430 ;
        RECT 39.720 37.925 39.860 39.110 ;
        RECT 39.650 37.555 39.930 37.925 ;
        RECT 39.200 36.730 39.460 37.050 ;
        RECT 39.260 34.670 39.400 36.730 ;
        RECT 38.340 34.270 38.940 34.410 ;
        RECT 39.200 34.350 39.460 34.670 ;
        RECT 38.800 33.990 38.940 34.270 ;
        RECT 36.440 33.670 36.700 33.990 ;
        RECT 36.900 33.670 37.160 33.990 ;
        RECT 38.280 33.670 38.540 33.990 ;
        RECT 38.740 33.670 39.000 33.990 ;
        RECT 36.960 29.230 37.100 33.670 ;
        RECT 37.360 31.290 37.620 31.610 ;
        RECT 36.900 28.910 37.160 29.230 ;
        RECT 37.420 28.550 37.560 31.290 ;
        RECT 38.340 29.570 38.480 33.670 ;
        RECT 38.800 31.610 38.940 33.670 ;
        RECT 38.740 31.290 39.000 31.610 ;
        RECT 39.660 31.290 39.920 31.610 ;
        RECT 39.720 31.125 39.860 31.290 ;
        RECT 39.650 30.755 39.930 31.125 ;
        RECT 38.280 29.250 38.540 29.570 ;
        RECT 36.900 28.230 37.160 28.550 ;
        RECT 37.360 28.230 37.620 28.550 ;
        RECT 36.960 26.850 37.100 28.230 ;
        RECT 37.820 27.890 38.080 28.210 ;
        RECT 36.900 26.530 37.160 26.850 ;
        RECT 36.440 25.850 36.700 26.170 ;
        RECT 36.900 25.850 37.160 26.170 ;
        RECT 35.520 23.810 35.780 24.130 ;
        RECT 35.060 23.130 35.320 23.450 ;
        RECT 32.760 22.790 33.020 23.110 ;
        RECT 35.520 22.790 35.780 23.110 ;
        RECT 32.820 19.710 32.960 22.790 ;
        RECT 33.680 22.110 33.940 22.430 ;
        RECT 33.740 21.410 33.880 22.110 ;
        RECT 33.680 21.090 33.940 21.410 ;
        RECT 35.580 20.390 35.720 22.790 ;
        RECT 35.970 20.555 36.250 20.925 ;
        RECT 35.980 20.410 36.240 20.555 ;
        RECT 35.520 20.070 35.780 20.390 ;
        RECT 32.760 19.390 33.020 19.710 ;
        RECT 30.920 17.350 31.180 17.670 ;
        RECT 32.300 17.350 32.560 17.670 ;
        RECT 29.540 14.630 29.800 14.950 ;
        RECT 30.000 14.630 30.260 14.950 ;
        RECT 26.780 12.930 27.040 13.250 ;
        RECT 30.060 12.910 30.200 14.630 ;
        RECT 30.980 14.125 31.120 17.350 ;
        RECT 30.910 13.755 31.190 14.125 ;
        RECT 30.000 12.590 30.260 12.910 ;
        RECT 30.060 12.230 30.200 12.590 ;
        RECT 32.820 12.230 32.960 19.390 ;
        RECT 35.580 18.690 35.720 20.070 ;
        RECT 36.500 19.710 36.640 25.850 ;
        RECT 36.440 19.390 36.700 19.710 ;
        RECT 35.520 18.370 35.780 18.690 ;
        RECT 35.980 18.030 36.240 18.350 ;
        RECT 33.680 17.525 33.940 17.670 ;
        RECT 33.670 17.155 33.950 17.525 ;
        RECT 35.060 16.670 35.320 16.990 ;
        RECT 35.520 16.670 35.780 16.990 ;
        RECT 35.120 14.950 35.260 16.670 ;
        RECT 35.580 15.290 35.720 16.670 ;
        RECT 35.520 14.970 35.780 15.290 ;
        RECT 35.060 14.630 35.320 14.950 ;
        RECT 35.120 12.570 35.260 14.630 ;
        RECT 36.040 12.910 36.180 18.030 ;
        RECT 36.500 17.670 36.640 19.390 ;
        RECT 36.960 18.690 37.100 25.850 ;
        RECT 37.360 25.510 37.620 25.830 ;
        RECT 37.420 21.410 37.560 25.510 ;
        RECT 37.880 23.110 38.020 27.890 ;
        RECT 38.740 25.850 39.000 26.170 ;
        RECT 37.820 22.790 38.080 23.110 ;
        RECT 38.280 22.790 38.540 23.110 ;
        RECT 37.360 21.090 37.620 21.410 ;
        RECT 37.880 21.070 38.020 22.790 ;
        RECT 37.820 20.750 38.080 21.070 ;
        RECT 37.360 20.410 37.620 20.730 ;
        RECT 36.900 18.370 37.160 18.690 ;
        RECT 37.420 17.670 37.560 20.410 ;
        RECT 36.440 17.350 36.700 17.670 ;
        RECT 37.360 17.350 37.620 17.670 ;
        RECT 36.500 13.250 36.640 17.350 ;
        RECT 38.340 15.970 38.480 22.790 ;
        RECT 38.800 20.390 38.940 25.850 ;
        RECT 38.740 20.070 39.000 20.390 ;
        RECT 39.660 19.730 39.920 20.050 ;
        RECT 39.200 17.690 39.460 18.010 ;
        RECT 38.740 17.350 39.000 17.670 ;
        RECT 38.280 15.650 38.540 15.970 ;
        RECT 38.800 13.250 38.940 17.350 ;
        RECT 36.440 12.930 36.700 13.250 ;
        RECT 38.740 12.930 39.000 13.250 ;
        RECT 35.980 12.590 36.240 12.910 ;
        RECT 35.060 12.250 35.320 12.570 ;
        RECT 30.000 11.910 30.260 12.230 ;
        RECT 32.760 11.910 33.020 12.230 ;
        RECT 35.520 11.910 35.780 12.230 ;
        RECT 24.020 11.570 24.280 11.890 ;
        RECT 19.420 11.230 19.680 11.550 ;
        RECT 22.180 11.230 22.440 11.550 ;
        RECT 26.320 11.230 26.580 11.550 ;
        RECT 32.300 11.230 32.560 11.550 ;
        RECT 19.480 4.000 19.620 11.230 ;
        RECT 22.240 5.850 22.380 11.230 ;
        RECT 24.370 10.695 25.910 11.065 ;
        RECT 26.380 5.850 26.520 11.230 ;
        RECT 22.240 5.710 22.840 5.850 ;
        RECT 22.700 4.000 22.840 5.710 ;
        RECT 25.920 5.710 26.520 5.850 ;
        RECT 25.920 4.000 26.060 5.710 ;
        RECT 32.360 4.000 32.500 11.230 ;
        RECT 35.580 10.725 35.720 11.910 ;
        RECT 35.510 10.355 35.790 10.725 ;
        RECT 39.260 7.325 39.400 17.690 ;
        RECT 39.720 17.670 39.860 19.730 ;
        RECT 39.660 17.350 39.920 17.670 ;
        RECT 39.720 14.950 39.860 17.350 ;
        RECT 39.660 14.630 39.920 14.950 ;
        RECT 39.190 6.955 39.470 7.325 ;
      LAYER met3 ;
        RECT 39.625 51.490 39.955 51.505 ;
        RECT 39.625 51.190 43.045 51.490 ;
        RECT 39.625 51.175 39.955 51.190 ;
        RECT 36.865 48.090 37.195 48.105 ;
        RECT 36.865 47.790 43.045 48.090 ;
        RECT 36.865 47.775 37.195 47.790 ;
        RECT 21.050 46.075 22.630 46.405 ;
        RECT 38.245 44.690 38.575 44.705 ;
        RECT 38.245 44.390 43.045 44.690 ;
        RECT 38.245 44.375 38.575 44.390 ;
        RECT 24.350 43.355 25.930 43.685 ;
        RECT 16.165 42.650 16.495 42.665 ;
        RECT 20.305 42.650 20.635 42.665 ;
        RECT 33.645 42.650 33.975 42.665 ;
        RECT 16.165 42.350 33.975 42.650 ;
        RECT 16.165 42.335 16.495 42.350 ;
        RECT 20.305 42.335 20.635 42.350 ;
        RECT 33.645 42.335 33.975 42.350 ;
        RECT 17.545 41.290 17.875 41.305 ;
        RECT 4.000 40.990 17.875 41.290 ;
        RECT 17.545 40.975 17.875 40.990 ;
        RECT 39.625 41.290 39.955 41.305 ;
        RECT 39.625 40.990 43.045 41.290 ;
        RECT 39.625 40.975 39.955 40.990 ;
        RECT 21.050 40.635 22.630 40.965 ;
        RECT 24.350 37.915 25.930 38.245 ;
        RECT 6.505 37.890 6.835 37.905 ;
        RECT 4.000 37.590 6.835 37.890 ;
        RECT 6.505 37.575 6.835 37.590 ;
        RECT 39.625 37.890 39.955 37.905 ;
        RECT 39.625 37.590 43.045 37.890 ;
        RECT 39.625 37.575 39.955 37.590 ;
        RECT 21.050 35.195 22.630 35.525 ;
        RECT 37.325 34.490 37.655 34.505 ;
        RECT 37.325 34.190 43.045 34.490 ;
        RECT 37.325 34.175 37.655 34.190 ;
        RECT 24.350 32.475 25.930 32.805 ;
        RECT 6.505 31.090 6.835 31.105 ;
        RECT 4.000 30.790 6.835 31.090 ;
        RECT 6.505 30.775 6.835 30.790 ;
        RECT 39.625 31.090 39.955 31.105 ;
        RECT 39.625 30.790 43.045 31.090 ;
        RECT 39.625 30.775 39.955 30.790 ;
        RECT 21.050 29.755 22.630 30.085 ;
        RECT 34.565 27.690 34.895 27.705 ;
        RECT 34.565 27.390 43.045 27.690 ;
        RECT 34.565 27.375 34.895 27.390 ;
        RECT 24.350 27.035 25.930 27.365 ;
        RECT 21.050 24.315 22.630 24.645 ;
        RECT 6.505 24.290 6.835 24.305 ;
        RECT 4.000 23.990 6.835 24.290 ;
        RECT 6.505 23.975 6.835 23.990 ;
        RECT 32.265 24.290 32.595 24.305 ;
        RECT 32.265 23.990 43.045 24.290 ;
        RECT 32.265 23.975 32.595 23.990 ;
        RECT 24.350 21.595 25.930 21.925 ;
        RECT 35.945 20.890 36.275 20.905 ;
        RECT 35.945 20.590 43.045 20.890 ;
        RECT 35.945 20.575 36.275 20.590 ;
        RECT 21.050 18.875 22.630 19.205 ;
        RECT 33.645 17.490 33.975 17.505 ;
        RECT 33.645 17.190 43.045 17.490 ;
        RECT 33.645 17.175 33.975 17.190 ;
        RECT 24.350 16.155 25.930 16.485 ;
        RECT 4.205 14.770 4.535 14.785 ;
        RECT 3.990 14.455 4.535 14.770 ;
        RECT 3.990 14.240 4.290 14.455 ;
        RECT 4.000 13.790 4.290 14.240 ;
        RECT 30.885 14.090 31.215 14.105 ;
        RECT 30.885 13.790 43.045 14.090 ;
        RECT 30.885 13.775 31.215 13.790 ;
        RECT 21.050 13.435 22.630 13.765 ;
        RECT 24.350 10.715 25.930 11.045 ;
        RECT 35.485 10.690 35.815 10.705 ;
        RECT 35.485 10.390 43.045 10.690 ;
        RECT 35.485 10.375 35.815 10.390 ;
        RECT 39.165 7.290 39.495 7.305 ;
        RECT 39.165 6.990 43.045 7.290 ;
        RECT 39.165 6.975 39.495 6.990 ;
  END
END bit4_encoder
END LIBRARY

