* SPICE3 file created from tt_um_tim2305_adc_dac.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_0p35_MGD972 a_n35_n486# a_n165_n616# a_n35_54#
X0 a_n35_54# a_n35_n486# a_n165_n616# sky130_fd_pr__res_xhigh_po_0p35 l=0.7
.ends

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X7 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X8 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X10 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X11 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X12 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X16 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X17 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X18 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X19 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X21 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_222_93# B1_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.10025 ps=0.985 w=0.42 l=0.15
X1 VPWR A1 a_544_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.105 ps=1.21 w=1 l=0.15
X2 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_222_93# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.18575 ps=1.415 w=0.42 l=0.15
X4 VGND A2 a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X5 a_448_47# a_222_93# a_79_199# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.169 ps=1.82 w=0.65 l=0.15
X6 a_79_199# a_222_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.3 ps=2.6 w=1 l=0.15
X7 a_544_297# A2 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.165 ps=1.33 w=1 l=0.15
X8 a_448_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18575 pd=1.415 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 X a_215_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_109_53# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_215_297# a_109_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_215_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_392_297# C a_297_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.04515 pd=0.635 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 a_465_297# B a_392_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06405 pd=0.725 as=0.04515 ps=0.635 w=0.42 l=0.15
X6 a_215_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X7 VPWR A a_465_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.06405 ps=0.725 w=0.42 l=0.15
X8 a_297_297# a_109_53# a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_109_53# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X10 VGND C a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06405 ps=0.725 w=0.42 l=0.15
X11 VGND A a_215_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1725 pd=1.345 as=0.265 ps=2.53 w=1 l=0.15
X1 a_209_297# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.16 pd=1.32 as=0.1725 ps=1.345 w=1 l=0.15
X2 a_303_47# A2 a_209_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.104 ps=0.97 w=0.65 l=0.15
X3 a_209_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.104 pd=0.97 as=0.112125 ps=0.995 w=0.65 l=0.15
X4 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.112125 pd=0.995 as=0.17225 ps=1.83 w=0.65 l=0.15
X5 VGND B1 a_80_21# VNB sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.10725 ps=0.98 w=0.65 l=0.15
X6 a_80_21# A1 a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X7 VPWR A2 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.16 ps=1.32 w=1 l=0.15
X8 a_80_21# B1 a_209_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.32 pd=2.64 as=0.165 ps=1.33 w=1 l=0.15
X9 a_209_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
X0 VPWR A a_49_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 VGND a_285_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.5
X2 X a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VGND A a_49_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_285_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.5
X5 a_285_47# a_49_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X6 a_285_47# a_49_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.5
X7 X a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.101875 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.14825 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
X0 VPWR B a_207_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2279 pd=1.74 as=0.0609 ps=0.71 w=0.42 l=0.15
X1 X a_207_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.2279 ps=1.74 w=1 l=0.15
X2 a_297_47# a_27_413# a_207_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0504 pd=0.66 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 X a_207_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1013 ps=0.99 w=0.65 l=0.15
X4 a_207_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.0714 ps=0.76 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0714 pd=0.76 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1013 pd=0.99 as=0.0504 ps=0.66 w=0.42 l=0.15
X7 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.14825 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.101875 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14825 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
X0 VPWR a_212_413# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 a_297_47# a_27_413# a_212_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_212_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.22895 ps=1.745 w=1 l=0.15
X3 X a_212_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.101875 ps=0.99 w=0.65 l=0.15
X4 a_212_413# a_27_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 VPWR A_N a_27_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 VPWR B a_212_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22895 pd=1.745 as=0.0609 ps=0.71 w=0.42 l=0.15
X7 VGND B a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.101875 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 VGND a_212_413# X VNB sky130_fd_pr__nfet_01v8 ad=0.1755 pd=1.84 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 a_27_413# A_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
X0 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X1 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X2 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X3 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X5 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.14 ps=1.28 w=1 l=0.15
X6 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.265 ps=2.53 w=1 l=0.15
X7 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X8 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X9 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X10 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X11 a_110_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X12 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X13 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.0588 ps=0.7 w=0.42 l=0.15
X14 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X15 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X16 VGND A a_110_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X17 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1113 pd=1.37 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1375 pd=1.275 as=0.14 ps=1.28 w=1 l=0.15
X19 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X20 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.1375 ps=1.275 w=1 l=0.15
X21 a_110_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1113 ps=1.37 w=0.42 l=0.15
X22 VPWR A a_110_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X23 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X24 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X25 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X27 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X28 VGND a_110_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X30 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X31 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X32 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X33 VPWR a_110_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X34 X a_110_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X35 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X36 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X38 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X39 X a_110_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.05775 ps=0.695 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_103_199# B1 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2015 pd=1.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VPWR a_103_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.36 ps=2.72 w=1 l=0.15
X2 a_337_297# A2 a_253_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X3 a_103_199# A3 a_337_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2125 pd=1.425 as=0.165 ps=1.33 w=1 l=0.15
X4 a_253_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.195 ps=1.39 w=1 l=0.15
X5 VPWR B1 a_103_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.345 pd=2.69 as=0.2125 ps=1.425 w=1 l=0.15
X6 VGND a_103_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.234 ps=2.02 w=0.65 l=0.15
X7 a_253_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.12675 ps=1.04 w=0.65 l=0.15
X8 a_253_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.10725 ps=0.98 w=0.65 l=0.15
X9 VGND A2 a_253_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
X0 VPWR A a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_109_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X3 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VGND A4 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1235 pd=1.03 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 a_321_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.1235 ps=1.03 w=0.65 l=0.15
X2 a_103_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=1.52 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR a_103_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.425 ps=2.85 w=1 l=0.15
X4 VGND a_103_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.247 ps=2.06 w=0.65 l=0.15
X5 VGND A2 a_321_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.12675 ps=1.04 w=0.65 l=0.15
X6 a_321_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.195 pd=1.9 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_511_297# A3 a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.22 ps=1.44 w=1 l=0.15
X8 a_619_297# A2 a_511_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.195 ps=1.39 w=1 l=0.15
X9 a_321_47# B1 a_103_21# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 a_393_297# A4 a_103_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.22 pd=1.44 as=0.26 ps=1.52 w=1 l=0.15
X11 VPWR A1 a_619_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.10025 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.10025 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.14575 ps=1.335 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_382_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.1525 ps=1.305 w=1 l=0.15
X1 a_297_47# B1 a_79_21# VNB sky130_fd_pr__nfet_01v8 ad=0.10075 pd=0.96 as=0.169 ps=1.82 w=0.65 l=0.15
X2 a_297_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VGND A2 a_297_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10075 ps=0.96 w=0.65 l=0.15
X4 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3275 pd=1.655 as=0.28 ps=2.56 w=1 l=0.15
X5 a_79_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.3275 ps=1.655 w=1 l=0.15
X6 a_382_297# A2 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1525 pd=1.305 as=0.195 ps=1.39 w=1 l=0.15
X7 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt bit4_encoder bus0[0] bus0[1] bus0[2] bus0[3] bus1[0] bus1[1] bus1[2] bus1[3]
+ clk compr[0] compr[12] compr[14] compr[1] compr[2] compr[3] compr[4] compr[5] compr[8]
+ bus2[0] bus2[2] compr[11] compr[7] compr[13] compr[9] VPWR bus2[1] bus2[3] compr[10]
+ VGND compr[6]
X_83_ clknet_1_0__leaf_clk _05_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfxtp_1
X_49_ net2 _21_ net3 VGND VGND VPWR VPWR _22_ sky130_fd_sc_hd__o21ba_1
X_66_ net15 _33_ net2 _27_ VGND VGND VPWR VPWR _36_ sky130_fd_sc_hd__or4b_1
XPHY_EDGE_ROW_12_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput20 net20 VGND VGND VPWR VPWR bus1[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Left_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_82_ clknet_1_0__leaf_clk _04_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfxtp_1
X_65_ net28 _35_ _15_ VGND VGND VPWR VPWR _04_ sky130_fd_sc_hd__mux2_1
X_48_ net14 _20_ net15 VGND VGND VPWR VPWR _21_ sky130_fd_sc_hd__o21ba_1
Xoutput21 net21 VGND VGND VPWR VPWR bus1[1] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_81_ clknet_1_1__leaf_clk _03_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfxtp_1
XFILLER_3_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_47_ net12 _19_ net13 VGND VGND VPWR VPWR _20_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_64_ _27_ _29_ _34_ _33_ VGND VGND VPWR VPWR _35_ sky130_fd_sc_hd__a31o_1
Xhold10 net20 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput22 net22 VGND VGND VPWR VPWR bus1[2] sky130_fd_sc_hd__buf_2
X_80_ clknet_1_1__leaf_clk _02_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfxtp_1
X_63_ net9 net10 net11 net12 VGND VGND VPWR VPWR _34_ sky130_fd_sc_hd__or4_1
XFILLER_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_46_ net10 _18_ net11 VGND VGND VPWR VPWR _19_ sky130_fd_sc_hd__o21ba_1
Xhold11 net24 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput23 net23 VGND VGND VPWR VPWR bus1[3] sky130_fd_sc_hd__buf_2
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_62_ net3 net4 net5 net6 VGND VGND VPWR VPWR _33_ sky130_fd_sc_hd__or4_1
XPHY_EDGE_ROW_4_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold12 bus_count\[1\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
X_45_ net8 _17_ net9 VGND VGND VPWR VPWR _18_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_7_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput24 net24 VGND VGND VPWR VPWR bus2[0] sky130_fd_sc_hd__buf_2
XFILLER_6_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_61_ net33 _32_ _15_ VGND VGND VPWR VPWR _03_ sky130_fd_sc_hd__mux2_1
XFILLER_9_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_44_ net7 net1 VGND VGND VPWR VPWR _17_ sky130_fd_sc_hd__and2b_1
Xhold13 _10_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput25 net25 VGND VGND VPWR VPWR bus2[1] sky130_fd_sc_hd__buf_2
X_60_ net5 net6 _31_ VGND VGND VPWR VPWR _32_ sky130_fd_sc_hd__or3_1
X_43_ _15_ VGND VGND VPWR VPWR _16_ sky130_fd_sc_hd__inv_2
Xhold14 bus_count\[0\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput26 net26 VGND VGND VPWR VPWR bus2[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_42_ bus_count\[0\] bus_count\[1\] VGND VGND VPWR VPWR _15_ sky130_fd_sc_hd__and2b_2
Xoutput16 net16 VGND VGND VPWR VPWR bus0[0] sky130_fd_sc_hd__buf_2
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
Xoutput27 net27 VGND VGND VPWR VPWR bus2[3] sky130_fd_sc_hd__buf_2
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_41_ _01_ VGND VGND VPWR VPWR _14_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR bus0[1] sky130_fd_sc_hd__buf_2
X_40_ bus_count\[1\] bus_count\[0\] VGND VGND VPWR VPWR _01_ sky130_fd_sc_hd__and2b_2
Xoutput18 net18 VGND VGND VPWR VPWR bus0[2] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput19 net19 VGND VGND VPWR VPWR bus0[3] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_3_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput1 compr[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 compr[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
X_79_ clknet_1_1__leaf_clk _01_ VGND VGND VPWR VPWR bus_count\[1\] sky130_fd_sc_hd__dfxtp_1
Xinput3 compr[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_78_ clknet_1_0__leaf_clk _00_ VGND VGND VPWR VPWR bus_count\[0\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 compr[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_77_ net30 _36_ _00_ VGND VGND VPWR VPWR _13_ sky130_fd_sc_hd__mux2_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput5 compr[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
X_76_ net35 _35_ _00_ VGND VGND VPWR VPWR _12_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_59_ net15 net2 _28_ _30_ VGND VGND VPWR VPWR _31_ sky130_fd_sc_hd__o31a_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 compr[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
X_58_ net3 net4 VGND VGND VPWR VPWR _30_ sky130_fd_sc_hd__nor2_1
X_75_ net32 _32_ _00_ VGND VGND VPWR VPWR _11_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_91_ clknet_1_0__leaf_clk _13_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfxtp_1
X_74_ bus_count\[0\] net39 net6 _23_ _38_ VGND VGND VPWR VPWR _10_ sky130_fd_sc_hd__o41a_1
Xinput7 compr[1] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_5_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_57_ net15 net2 VGND VGND VPWR VPWR _29_ sky130_fd_sc_hd__nor2_1
Xinput10 compr[4] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
XFILLER_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_90_ clknet_1_0__leaf_clk _12_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfxtp_1
X_73_ net16 _00_ VGND VGND VPWR VPWR _38_ sky130_fd_sc_hd__or2_1
Xinput8 compr[2] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_56_ net11 net12 _26_ _27_ VGND VGND VPWR VPWR _28_ sky130_fd_sc_hd__o31a_1
X_39_ net41 net39 VGND VGND VPWR VPWR _00_ sky130_fd_sc_hd__nor2_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
Xinput11 compr[5] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_7_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_2_Left_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput9 compr[3] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_72_ net31 _36_ _01_ VGND VGND VPWR VPWR _09_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 compr[6] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
X_55_ net13 net14 VGND VGND VPWR VPWR _27_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1 net26 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd3_1
X_54_ net7 net8 _25_ VGND VGND VPWR VPWR _26_ sky130_fd_sc_hd__o21a_1
X_71_ net36 _35_ _01_ VGND VGND VPWR VPWR _08_ sky130_fd_sc_hd__mux2_1
Xinput13 compr[7] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xhold2 net21 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dlygate4sd3_1
X_70_ net29 _32_ _01_ VGND VGND VPWR VPWR _07_ sky130_fd_sc_hd__mux2_1
Xinput14 compr[8] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
X_53_ net9 net10 VGND VGND VPWR VPWR _25_ sky130_fd_sc_hd__nor2_1
Xhold3 net19 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dlygate4sd3_1
X_52_ net6 _16_ _23_ _24_ VGND VGND VPWR VPWR _02_ sky130_fd_sc_hd__o31a_1
Xinput15 compr[9] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_6_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold4 net23 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlygate4sd3_1
X_51_ net38 _15_ VGND VGND VPWR VPWR _24_ sky130_fd_sc_hd__or2_1
XFILLER_0_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 net17 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dlygate4sd3_1
X_50_ net4 _22_ net5 VGND VGND VPWR VPWR _23_ sky130_fd_sc_hd__o21ba_1
Xhold6 net25 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold7 net27 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold8 net18 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_1_Left_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold9 net22 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_89_ clknet_1_1__leaf_clk _11_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfxtp_1
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_88_ clknet_1_1__leaf_clk net40 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfxtp_1
X_87_ clknet_1_0__leaf_clk _09_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_5_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_8_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_86_ clknet_1_0__leaf_clk _08_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfxtp_1
X_69_ net6 _14_ _23_ _37_ VGND VGND VPWR VPWR _06_ sky130_fd_sc_hd__o31a_1
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_85_ clknet_1_1__leaf_clk _07_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfxtp_1
X_68_ net37 _01_ VGND VGND VPWR VPWR _37_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_84_ clknet_1_1__leaf_clk _06_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfxtp_1
X_67_ net34 _36_ _15_ VGND VGND VPWR VPWR _05_ sky130_fd_sc_hd__mux2_1
XFILLER_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
C0 VPWR _00_ 2.496267f
C1 VPWR _36_ 2.108505f
C2 clknet_1_0__leaf_clk VPWR 2.060224f
C3 clknet_1_1__leaf_clk VPWR 2.109072f
C4 _01_ VGND 3.226816f
C5 _00_ VGND 2.658476f
C6 VPWR VGND 92.371376f
C7 _15_ VGND 2.114687f
C8 clknet_1_0__leaf_clk VGND 3.388226f
.ends

.subckt sky130_fd_pr__pfet_01v8_LGA5KQ a_n73_n564# a_n33_n661# a_15_n564# w_n211_n784#
+ VSUBS
X0 a_15_n564# a_n33_n661# a_n73_n564# w_n211_n784# sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=0.15
C0 w_n211_n784# VSUBS 2.85893f
.ends

.subckt sky130_fd_pr__nfet_01v8_ATMSL9 a_n33_191# a_n73_n231# a_15_n231# a_n175_n343#
X0 a_15_n231# a_n33_191# a_n73_n231# a_n175_n343# sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.15
.ends

.subckt sky130_fd_pr__res_xhigh_po_0p35_ABVTW2 a_n35_124# a_n165_n686# a_n35_n556#
X0 a_n35_124# a_n35_n556# a_n165_n686# sky130_fd_pr__res_xhigh_po_0p35 l=1.4
.ends

.subckt sky130_fd_pr__pfet_01v8_MGA5KJ a_n73_n636# a_15_n636# a_n33_595# w_n211_n784#
+ VSUBS
X0 a_15_n636# a_n33_595# a_n73_n636# w_n211_n784# sky130_fd_pr__pfet_01v8 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=0.15
C0 w_n211_n784# VSUBS 2.85893f
.ends

.subckt r2r_dac out vdd b0 b1 b2 b3 b4 b5 b6 b7 vss
XXM12 m1_2630_n3424# b2 vdd vdd vss sky130_fd_pr__pfet_01v8_LGA5KQ
XXM14 m1_2920_n3426# b1 vdd vdd vss sky130_fd_pr__pfet_01v8_LGA5KQ
XXM15 b0 m1_3220_n3424# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
XXM16 m1_3220_n3424# b0 vdd vdd vss sky130_fd_pr__pfet_01v8_LGA5KQ
Xsky130_fd_pr__nfet_01v8_ATMSL9_0 b1 m1_2920_n3426# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
XXR1 m1_1394_n2598# vss m1_1170_n4750# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXR10 m1_1762_n4750# vss m1_2056_n4750# sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR2 out vss m1_1170_n4750# sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR11 m1_2326_n1634# vss m1_2056_n4750# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXR3 m1_1060_n2596# vss out sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXR5 vss vss m1_2946_n4750# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXR12 m1_2056_n4750# vss m1_2354_n4750# sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXM1 b7 m1_1060_n2596# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
XXR14 m1_2354_n4750# vss m1_2650_n4752# sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR13 m1_2630_n3424# vss m1_2354_n4750# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXR6 m1_1170_n4750# vss m1_1460_n4750# sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR15 m1_2920_n3426# vss m1_2650_n4752# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXR7 m1_1698_n2368# vss m1_1460_n4750# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXM3 b6 m1_1394_n2598# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
XXR16 m1_2650_n4752# vss m1_2946_n4750# sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR8 m1_1460_n4750# vss m1_1762_n4750# sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXM4 vdd m1_1394_n2598# b6 vdd vss sky130_fd_pr__pfet_01v8_MGA5KJ
XXR17 m1_3220_n3424# vss m1_2946_n4750# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXR9 m1_2014_n2596# vss m1_1762_n4750# sky130_fd_pr__res_xhigh_po_0p35_ABVTW2
XXM5 b5 m1_1698_n2368# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
XXM6 m1_1698_n2368# b5 vdd vdd vss sky130_fd_pr__pfet_01v8_LGA5KQ
XXM7 b4 m1_2014_n2596# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
XXM8 m1_2014_n2596# b4 vdd vdd vss sky130_fd_pr__pfet_01v8_LGA5KQ
XXM9 b3 m1_2326_n1634# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
Xsky130_fd_pr__pfet_01v8_LGA5KQ_0 m1_1060_n2596# b7 vdd vdd vss sky130_fd_pr__pfet_01v8_LGA5KQ
XXM10 m1_2326_n1634# b3 vdd vdd vss sky130_fd_pr__pfet_01v8_LGA5KQ
XXM11 b2 m1_2630_n3424# vss vss sky130_fd_pr__nfet_01v8_ATMSL9
R0 m1_1060_n2596# m1_1060_n2596# sky130_fd_pr__res_generic_m2 w=0.32 l=0.09
C0 vss 0 -10.099447f
C1 vdd 0 15.611696f
.ends

.subckt sky130_fd_pr__nfet_01v8_64Z3AY a_15_n131# a_n175_n243# a_n33_91# a_n73_n131#
X0 a_15_n131# a_n33_91# a_n73_n131# a_n175_n243# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
.ends

.subckt sky130_fd_pr__pfet_01v8_3H2EVM a_n100_n897# a_100_n800# w_n296_n1019# a_n158_n800#
+ VSUBS
X0 a_100_n800# a_n100_n897# a_n158_n800# w_n296_n1019# sky130_fd_pr__pfet_01v8 ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=1
C0 w_n296_n1019# VSUBS 4.82082f
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHMAL2 a_n260_n574# a_100_n400# a_n158_n400# a_n100_n488#
X0 a_100_n400# a_n100_n488# a_n158_n400# a_n260_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_AHRV9L a_n258_n400# a_n200_n488# a_n360_n574#
+ a_200_n400#
X0 a_200_n400# a_n200_n488# a_n258_n400# a_n360_n574# sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=2
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_GWPMZG a_n200_n897# a_200_n800# w_n396_n1019#
+ a_n258_n800# VSUBS
X0 a_200_n800# a_n200_n897# a_n258_n800# w_n396_n1019# sky130_fd_pr__pfet_01v8_lvt ad=2.32 pd=16.58 as=2.32 ps=16.58 w=8 l=2
C0 w_n396_n1019# VSUBS 6.14037f
.ends

.subckt sky130_fd_pr__pfet_01v8_MGSNAN a_n73_n336# a_15_n336# a_n33_295# w_n211_n484#
+ VSUBS
X0 a_15_n336# a_n33_295# a_n73_n336# w_n211_n484# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=0.15
.ends

.subckt compr out vdd in+ in- vss
XXM1 out vss m1_2518_1378# vss sky130_fd_pr__nfet_01v8_64Z3AY
XXM3 m1_1460_732# vdd vdd m1_1264_902# vss sky130_fd_pr__pfet_01v8_3H2EVM
XXM4 vss vss m1_1264_902# m1_1460_732# sky130_fd_pr__nfet_01v8_lvt_AHMAL2
XXM5 m1_1824_498# m1_1824_498# vss vss sky130_fd_pr__nfet_01v8_lvt_AHRV9L
XXM6 m1_2518_1378# m1_2518_1378# vss vss sky130_fd_pr__nfet_01v8_lvt_AHRV9L
XXM7 in- m1_2324_1380# vdd m1_1824_498# vss sky130_fd_pr__pfet_01v8_lvt_GWPMZG
XXM8 m1_1264_902# vdd vdd m1_2324_1380# vss sky130_fd_pr__pfet_01v8_3H2EVM
XXM9 in+ m1_2324_1380# vdd m1_2518_1378# vss sky130_fd_pr__pfet_01v8_lvt_GWPMZG
XXM21 out vdd m1_2518_1378# vdd vss sky130_fd_pr__pfet_01v8_MGSNAN
R0 m1_1264_902# m1_1264_902# sky130_fd_pr__res_generic_m1 w=0.42 l=7.37
C0 m1_2518_1378# vss 3.195238f
C1 vdd vss 21.704147f
C2 m1_1824_498# vss 2.487121f
.ends

.subckt tt_um_tim2305_adc_dac clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6]
+ ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0]
+ uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0]
+ uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0]
+ uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0]
+ uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
XXR1 compr_14/in- VGND compr_13/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR2 compr_8/in- VGND compr_7/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR10 compr_10/in- VGND compr_9/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
Xbit4_encoder_0 uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6]
+ uo_out[7] clk compr_0/out compr_12/out compr_14/out compr_1/out compr_2/out compr_3/out
+ compr_4/out compr_5/out compr_8/out uio_out[0] uio_out[2] compr_11/out compr_7/out
+ compr_13/out compr_9/out VDPWR uio_out[1] uio_out[3] compr_10/out VGND compr_6/out
+ bit4_encoder
XXR3 compr_12/in- VGND compr_13/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR11 compr_0/in- VGND VGND sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR4 compr_14/in- VGND VDPWR sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR5 compr_8/in- VGND compr_9/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR12 compr_6/in- VGND compr_5/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR13 compr_2/in- VGND compr_1/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR14 compr_2/in- VGND compr_3/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR6 compr_0/in- VGND compr_1/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR7 compr_10/in- VGND compr_11/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR15 compr_6/in- VGND compr_7/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR8 compr_4/in- VGND compr_5/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR16 compr_4/in- VGND compr_3/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
XXR9 compr_12/in- VGND compr_11/in- sky130_fd_pr__res_xhigh_po_0p35_MGD972
Xr2r_dac_0 ua[1] VDPWR ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6]
+ ui_in[7] VGND r2r_dac
Xcompr_1 compr_1/out VDPWR ua[0] compr_1/in- VGND compr
Xcompr_0 compr_0/out VDPWR ua[0] compr_0/in- VGND compr
Xcompr_2 compr_2/out VDPWR ua[0] compr_2/in- VGND compr
Xcompr_3 compr_3/out VDPWR ua[0] compr_3/in- VGND compr
Xcompr_4 compr_4/out VDPWR ua[0] compr_4/in- VGND compr
Xcompr_5 compr_5/out VDPWR ua[0] compr_5/in- VGND compr
Xcompr_6 compr_6/out VDPWR ua[0] compr_6/in- VGND compr
Xcompr_7 compr_7/out VDPWR ua[0] compr_7/in- VGND compr
Xcompr_8 compr_8/out VDPWR ua[0] compr_8/in- VGND compr
Xcompr_10 compr_10/out VDPWR ua[0] compr_10/in- VGND compr
Xcompr_9 compr_9/out VDPWR ua[0] compr_9/in- VGND compr
Xcompr_11 compr_11/out VDPWR ua[0] compr_11/in- VGND compr
Xcompr_13 compr_13/out VDPWR ua[0] compr_13/in- VGND compr
Xcompr_12 compr_12/out VDPWR ua[0] compr_12/in- VGND compr
Xcompr_14 compr_14/out VDPWR ua[0] compr_14/in- VGND compr
Xcompr_15 compr_15/out VDPWR ua[6] ua[7] VGND compr
C0 compr_9/in- compr_8/in- 6.144914f
C1 uo_out[5] uo_out[7] 3.81182f
C2 compr_12/in- VDPWR 2.017333f
C3 VDPWR compr_14/in- 4.947888f
C4 VDPWR compr_13/in- 3.74722f
C5 compr_12/out compr_11/out 3.03107f
C6 ui_in[2] ui_in[1] 15.492226f
C7 compr_0/out ui_in[0] 5.421363f
C8 compr_7/in- compr_6/in- 3.476658f
C9 compr_7/out compr_8/out 3.361608f
C10 compr_14/out compr_13/out 2.130436f
C11 compr_8/in- VDPWR 4.433691f
C12 uio_out[1] uio_out[0] 7.057777f
C13 uo_out[6] uio_out[2] 4.741323f
C14 compr_4/in- VDPWR 2.576622f
C15 compr_2/out compr_1/out 4.378193f
C16 compr_0/in- compr_1/in- 2.724778f
C17 uio_out[2] uio_out[3] 4.07944f
C18 compr_2/in- VDPWR 3.103487f
C19 uo_out[1] uo_out[0] 4.165518f
C20 compr_3/in- compr_4/in- 8.018824f
C21 compr_2/out compr_3/out 3.451074f
C22 compr_3/in- compr_2/in- 5.909122f
C23 uo_out[1] uo_out[3] 2.462103f
C24 compr_7/in- VDPWR 2.345286f
C25 compr_12/out compr_13/out 2.284604f
C26 compr_9/in- VDPWR 4.333928f
C27 ui_in[4] ui_in[5] 11.691796f
C28 compr_12/in- compr_13/in- 4.614457f
C29 ui_in[6] ui_in[7] 9.980404f
C30 ui_in[0] ui_in[1] 14.844142f
C31 compr_13/in- compr_14/in- 5.938617f
C32 compr_9/out compr_8/out 2.040681f
C33 compr_3/in- VDPWR 3.423734f
C34 uo_out[4] uo_out[0] 2.683677f
C35 uo_out[6] uo_out[2] 3.605048f
C36 compr_5/out compr_6/out 4.79194f
C37 uo_out[4] uio_out[0] 2.178017f
C38 VDPWR uo_out[0] 2.211617f
C39 uo_out[4] uo_out[3] 3.095258f
C40 ui_in[4] ui_in[3] 12.098826f
C41 compr_7/out compr_6/out 4.148319f
C42 ui_in[3] ui_in[2] 13.843406f
C43 compr_1/in- compr_2/in- 4.48108f
C44 ui_in[6] ui_in[5] 11.991817f
C45 uo_out[5] uo_out[4] 5.870261f
C46 uo_out[7] uio_out[0] 5.079198f
C47 compr_7/in- compr_8/in- 5.163016f
C48 compr_0/out compr_1/out 6.590864f
C49 VDPWR ua[0] 5.256798f
C50 compr_11/in- compr_12/in- 3.264768f
C51 compr_10/out compr_11/out 4.696752f
C52 compr_15/m1_2518_1378# VGND 2.228621f
C53 ua[6] VGND 2.203651f
C54 ua[7] VGND 4.238802f
C55 compr_14/m1_2518_1378# VGND 2.232347f
C56 compr_12/out VGND 2.893454f
C57 compr_12/m1_2518_1378# VGND 2.232665f
C58 compr_13/m1_2518_1378# VGND 2.233058f
C59 compr_11/out VGND 3.96004f
C60 compr_11/m1_2518_1378# VGND 2.23265f
C61 compr_9/out VGND 2.865288f
C62 compr_9/m1_2518_1378# VGND 2.232519f
C63 compr_9/m1_1264_902# VGND 2.519627f
C64 compr_10/out VGND 8.715362f
C65 compr_10/m1_2518_1378# VGND 2.229472f
C66 compr_8/out VGND 2.739233f
C67 compr_8/m1_2518_1378# VGND 2.23685f
C68 compr_7/out VGND 2.750981f
C69 compr_7/m1_2518_1378# VGND 2.236876f
C70 compr_6/out VGND 3.245878f
C71 compr_6/m1_2518_1378# VGND 2.236861f
C72 compr_5/out VGND 7.465467f
C73 compr_5/m1_2518_1378# VGND 2.239626f
C74 compr_4/out VGND 2.503867f
C75 compr_4/m1_2518_1378# VGND 2.232326f
C76 compr_4/m1_1264_902# VGND 2.600833f
C77 compr_3/out VGND 2.62255f
C78 compr_3/m1_2518_1378# VGND 2.232725f
C79 compr_2/out VGND 3.063375f
C80 compr_2/m1_2518_1378# VGND 2.232737f
C81 compr_0/out VGND 8.678228f
C82 compr_0/m1_2518_1378# VGND 2.228621f
C83 ua[0] VGND 29.8067f
C84 compr_1/out VGND 5.066405f
C85 compr_1/m1_2518_1378# VGND 2.232733f
C86 ua[1] VGND 10.643282f
C87 ui_in[0] VGND 4.859229f
C88 compr_4/in- VGND 3.141764f
C89 compr_3/in- VGND 2.679227f
C90 compr_1/in- VGND 2.843591f
C91 compr_2/in- VGND 2.838606f
C92 compr_9/in- VGND 2.188768f
C93 compr_0/in- VGND 3.40348f
C94 VDPWR VGND 0.512189p
C95 uio_out[3] VGND 3.688928f
C96 uio_out[2] VGND 2.400645f
C97 uio_out[1] VGND 2.492696f
C98 compr_14/in- VGND 2.770843f
.ends

