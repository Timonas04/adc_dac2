magic
tech sky130A
magscale 1 2
timestamp 1730882523
<< viali >>
rect 2881 9129 2915 9163
rect 4997 9129 5031 9163
rect 6653 9129 6687 9163
rect 3341 9061 3375 9095
rect 6193 9061 6227 9095
rect 3985 8993 4019 9027
rect 2697 8925 2731 8959
rect 3157 8925 3191 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 5181 8925 5215 8959
rect 5273 8925 5307 8959
rect 6009 8925 6043 8959
rect 6837 8925 6871 8959
rect 7389 8925 7423 8959
rect 7665 8925 7699 8959
rect 7941 8925 7975 8959
rect 3617 8789 3651 8823
rect 4629 8789 4663 8823
rect 5917 8789 5951 8823
rect 7205 8789 7239 8823
rect 7481 8789 7515 8823
rect 7757 8789 7791 8823
rect 2237 8585 2271 8619
rect 5089 8585 5123 8619
rect 3954 8517 3988 8551
rect 5181 8517 5215 8551
rect 5365 8517 5399 8551
rect 3361 8449 3395 8483
rect 5549 8449 5583 8483
rect 5641 8449 5675 8483
rect 6009 8449 6043 8483
rect 6561 8449 6595 8483
rect 6745 8449 6779 8483
rect 6837 8449 6871 8483
rect 7941 8449 7975 8483
rect 3617 8381 3651 8415
rect 3709 8381 3743 8415
rect 7021 8381 7055 8415
rect 5825 8313 5859 8347
rect 6101 8313 6135 8347
rect 6653 8313 6687 8347
rect 7757 8313 7791 8347
rect 6377 8245 6411 8279
rect 7665 8245 7699 8279
rect 3801 8041 3835 8075
rect 5273 8041 5307 8075
rect 6837 8041 6871 8075
rect 7389 8041 7423 8075
rect 4445 7905 4479 7939
rect 5457 7905 5491 7939
rect 1409 7837 1443 7871
rect 3433 7837 3467 7871
rect 4169 7837 4203 7871
rect 4721 7837 4755 7871
rect 4905 7837 4939 7871
rect 5365 7837 5399 7871
rect 5724 7837 5758 7871
rect 7021 7837 7055 7871
rect 7205 7837 7239 7871
rect 7481 7837 7515 7871
rect 7941 7837 7975 7871
rect 1676 7769 1710 7803
rect 4261 7769 4295 7803
rect 2789 7701 2823 7735
rect 2881 7701 2915 7735
rect 5089 7701 5123 7735
rect 7665 7701 7699 7735
rect 7757 7701 7791 7735
rect 1501 7497 1535 7531
rect 1777 7497 1811 7531
rect 2145 7497 2179 7531
rect 3341 7497 3375 7531
rect 5733 7429 5767 7463
rect 6377 7429 6411 7463
rect 1685 7361 1719 7395
rect 4629 7361 4663 7395
rect 6009 7361 6043 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 7021 7361 7055 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 7757 7361 7791 7395
rect 2237 7293 2271 7327
rect 2421 7293 2455 7327
rect 5365 7293 5399 7327
rect 5917 7293 5951 7327
rect 7113 7293 7147 7327
rect 4721 7157 4755 7191
rect 6009 7157 6043 7191
rect 6193 7157 6227 7191
rect 5181 6953 5215 6987
rect 7205 6953 7239 6987
rect 3617 6885 3651 6919
rect 5549 6885 5583 6919
rect 1869 6817 1903 6851
rect 2053 6817 2087 6851
rect 3801 6817 3835 6851
rect 6469 6817 6503 6851
rect 6561 6817 6595 6851
rect 2237 6749 2271 6783
rect 6377 6749 6411 6783
rect 6653 6749 6687 6783
rect 6837 6749 6871 6783
rect 7021 6749 7055 6783
rect 7389 6749 7423 6783
rect 7665 6749 7699 6783
rect 7849 6749 7883 6783
rect 2504 6681 2538 6715
rect 4068 6681 4102 6715
rect 5917 6681 5951 6715
rect 6929 6681 6963 6715
rect 1409 6613 1443 6647
rect 1777 6613 1811 6647
rect 5457 6613 5491 6647
rect 6193 6613 6227 6647
rect 5365 6409 5399 6443
rect 6745 6409 6779 6443
rect 7757 6409 7791 6443
rect 2522 6341 2556 6375
rect 3525 6341 3559 6375
rect 2789 6273 2823 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7481 6273 7515 6307
rect 7665 6273 7699 6307
rect 7941 6273 7975 6307
rect 5917 6205 5951 6239
rect 1409 6069 1443 6103
rect 4813 6069 4847 6103
rect 6377 6069 6411 6103
rect 7665 6069 7699 6103
rect 2329 5865 2363 5899
rect 3985 5865 4019 5899
rect 4445 5865 4479 5899
rect 6193 5865 6227 5899
rect 7849 5865 7883 5899
rect 4261 5797 4295 5831
rect 1685 5729 1719 5763
rect 4353 5729 4387 5763
rect 5549 5729 5583 5763
rect 2973 5661 3007 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 4077 5661 4111 5695
rect 4537 5661 4571 5695
rect 4813 5661 4847 5695
rect 6101 5661 6135 5695
rect 6285 5661 6319 5695
rect 6653 5661 6687 5695
rect 6837 5661 6871 5695
rect 6929 5661 6963 5695
rect 7205 5661 7239 5695
rect 7389 5661 7423 5695
rect 7665 5661 7699 5695
rect 4905 5593 4939 5627
rect 6561 5593 6595 5627
rect 2421 5525 2455 5559
rect 5917 5525 5951 5559
rect 6745 5525 6779 5559
rect 7113 5525 7147 5559
rect 1501 5321 1535 5355
rect 2237 5321 2271 5355
rect 4077 5321 4111 5355
rect 7849 5321 7883 5355
rect 2964 5253 2998 5287
rect 1685 5185 1719 5219
rect 4537 5185 4571 5219
rect 4997 5185 5031 5219
rect 6469 5185 6503 5219
rect 6561 5185 6595 5219
rect 6653 5185 6687 5219
rect 7205 5185 7239 5219
rect 7389 5185 7423 5219
rect 7665 5185 7699 5219
rect 2329 5117 2363 5151
rect 2513 5117 2547 5151
rect 2697 5117 2731 5151
rect 4629 5117 4663 5151
rect 4813 5117 4847 5151
rect 5549 5117 5583 5151
rect 6745 5117 6779 5151
rect 4169 5049 4203 5083
rect 6929 5049 6963 5083
rect 1869 4981 1903 5015
rect 2789 4777 2823 4811
rect 5733 4777 5767 4811
rect 7297 4777 7331 4811
rect 5641 4709 5675 4743
rect 1409 4641 1443 4675
rect 5273 4641 5307 4675
rect 3801 4573 3835 4607
rect 4068 4573 4102 4607
rect 6561 4573 6595 4607
rect 7481 4573 7515 4607
rect 7573 4573 7607 4607
rect 7665 4573 7699 4607
rect 7757 4573 7791 4607
rect 1676 4505 1710 4539
rect 5181 4437 5215 4471
rect 7205 4437 7239 4471
rect 6745 4233 6779 4267
rect 7481 4233 7515 4267
rect 7941 4165 7975 4199
rect 1685 4097 1719 4131
rect 3525 4097 3559 4131
rect 3985 4097 4019 4131
rect 4813 4097 4847 4131
rect 5080 4097 5114 4131
rect 7205 4097 7239 4131
rect 7665 4097 7699 4131
rect 1961 4029 1995 4063
rect 2881 4029 2915 4063
rect 3709 4029 3743 4063
rect 3893 4029 3927 4063
rect 6837 4029 6871 4063
rect 6929 4029 6963 4063
rect 7757 4029 7791 4063
rect 1501 3961 1535 3995
rect 6377 3961 6411 3995
rect 7389 3961 7423 3995
rect 2605 3893 2639 3927
rect 4353 3893 4387 3927
rect 6193 3893 6227 3927
rect 7665 3893 7699 3927
rect 1409 3689 1443 3723
rect 5089 3689 5123 3723
rect 6653 3689 6687 3723
rect 7297 3689 7331 3723
rect 6101 3621 6135 3655
rect 2789 3553 2823 3587
rect 3801 3485 3835 3519
rect 5917 3485 5951 3519
rect 6193 3485 6227 3519
rect 6469 3485 6503 3519
rect 6745 3485 6779 3519
rect 7021 3485 7055 3519
rect 7205 3485 7239 3519
rect 7481 3485 7515 3519
rect 7757 3485 7791 3519
rect 7941 3485 7975 3519
rect 2522 3417 2556 3451
rect 6377 3349 6411 3383
rect 6929 3349 6963 3383
rect 7113 3349 7147 3383
rect 1961 3145 1995 3179
rect 2329 3145 2363 3179
rect 2421 3145 2455 3179
rect 3801 3145 3835 3179
rect 5733 3145 5767 3179
rect 7757 3145 7791 3179
rect 1685 3009 1719 3043
rect 4914 3009 4948 3043
rect 5181 3009 5215 3043
rect 5641 3009 5675 3043
rect 6377 3009 6411 3043
rect 7573 3009 7607 3043
rect 2605 2941 2639 2975
rect 5917 2941 5951 2975
rect 6929 2941 6963 2975
rect 7297 2941 7331 2975
rect 7389 2941 7423 2975
rect 1501 2873 1535 2907
rect 5273 2805 5307 2839
rect 6929 2601 6963 2635
rect 7849 2601 7883 2635
rect 5641 2533 5675 2567
rect 7665 2533 7699 2567
rect 7389 2465 7423 2499
rect 3341 2397 3375 2431
rect 4169 2397 4203 2431
rect 4261 2397 4295 2431
rect 6009 2397 6043 2431
rect 6561 2397 6595 2431
rect 7113 2397 7147 2431
rect 4528 2329 4562 2363
rect 3525 2261 3559 2295
rect 3985 2261 4019 2295
rect 5825 2261 5859 2295
rect 6745 2261 6779 2295
<< metal1 >>
rect 1104 9274 8280 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 8280 9274
rect 1104 9200 8280 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 3878 9160 3884 9172
rect 2915 9132 3884 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4985 9163 5043 9169
rect 4985 9129 4997 9163
rect 5031 9160 5043 9163
rect 5166 9160 5172 9172
rect 5031 9132 5172 9160
rect 5031 9129 5043 9132
rect 4985 9123 5043 9129
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 6641 9163 6699 9169
rect 6641 9160 6653 9163
rect 6512 9132 6653 9160
rect 6512 9120 6518 9132
rect 6641 9129 6653 9132
rect 6687 9129 6699 9163
rect 6641 9123 6699 9129
rect 3329 9095 3387 9101
rect 3329 9061 3341 9095
rect 3375 9092 3387 9095
rect 4798 9092 4804 9104
rect 3375 9064 4804 9092
rect 3375 9061 3387 9064
rect 3329 9055 3387 9061
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 6178 9092 6184 9104
rect 5092 9064 6184 9092
rect 3973 9027 4031 9033
rect 3973 9024 3985 9027
rect 2700 8996 3985 9024
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2700 8965 2728 8996
rect 3973 8993 3985 8996
rect 4019 8993 4031 9027
rect 3973 8987 4031 8993
rect 2685 8959 2743 8965
rect 2685 8956 2697 8959
rect 2280 8928 2697 8956
rect 2280 8916 2286 8928
rect 2685 8925 2697 8928
rect 2731 8925 2743 8959
rect 2685 8919 2743 8925
rect 3142 8916 3148 8968
rect 3200 8916 3206 8968
rect 3234 8916 3240 8968
rect 3292 8916 3298 8968
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8956 3479 8959
rect 5092 8956 5120 9064
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 3467 8928 5120 8956
rect 5169 8959 5227 8965
rect 3467 8925 3479 8928
rect 3421 8919 3479 8925
rect 5169 8925 5181 8959
rect 5215 8956 5227 8959
rect 5258 8956 5264 8968
rect 5215 8928 5264 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5258 8916 5264 8928
rect 5316 8916 5322 8968
rect 5810 8916 5816 8968
rect 5868 8956 5874 8968
rect 5997 8959 6055 8965
rect 5997 8956 6009 8959
rect 5868 8928 6009 8956
rect 5868 8916 5874 8928
rect 5997 8925 6009 8928
rect 6043 8925 6055 8959
rect 5997 8919 6055 8925
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 7374 8916 7380 8968
rect 7432 8916 7438 8968
rect 7650 8916 7656 8968
rect 7708 8916 7714 8968
rect 7926 8916 7932 8968
rect 7984 8916 7990 8968
rect 3602 8780 3608 8832
rect 3660 8780 3666 8832
rect 4614 8780 4620 8832
rect 4672 8780 4678 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 5408 8792 5917 8820
rect 5408 8780 5414 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 5905 8783 5963 8789
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 6604 8792 7205 8820
rect 6604 8780 6610 8792
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7469 8823 7527 8829
rect 7469 8820 7481 8823
rect 7340 8792 7481 8820
rect 7340 8780 7346 8792
rect 7469 8789 7481 8792
rect 7515 8789 7527 8823
rect 7469 8783 7527 8789
rect 7745 8823 7803 8829
rect 7745 8789 7757 8823
rect 7791 8820 7803 8823
rect 7834 8820 7840 8832
rect 7791 8792 7840 8820
rect 7791 8789 7803 8792
rect 7745 8783 7803 8789
rect 7834 8780 7840 8792
rect 7892 8780 7898 8832
rect 1104 8730 8280 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 8280 8730
rect 1104 8656 8280 8678
rect 2222 8576 2228 8628
rect 2280 8576 2286 8628
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 5077 8619 5135 8625
rect 3200 8588 4200 8616
rect 3200 8576 3206 8588
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 3942 8551 4000 8557
rect 3942 8548 3954 8551
rect 3660 8520 3954 8548
rect 3660 8508 3666 8520
rect 3942 8517 3954 8520
rect 3988 8517 4000 8551
rect 4172 8548 4200 8588
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5258 8616 5264 8628
rect 5123 8588 5264 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5169 8551 5227 8557
rect 5169 8548 5181 8551
rect 4172 8520 5181 8548
rect 3942 8511 4000 8517
rect 5169 8517 5181 8520
rect 5215 8517 5227 8551
rect 5169 8511 5227 8517
rect 5350 8508 5356 8560
rect 5408 8508 5414 8560
rect 3349 8483 3407 8489
rect 3349 8449 3361 8483
rect 3395 8480 3407 8483
rect 3786 8480 3792 8492
rect 3395 8452 3792 8480
rect 3395 8449 3407 8452
rect 3349 8443 3407 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 5629 8483 5687 8489
rect 5629 8449 5641 8483
rect 5675 8449 5687 8483
rect 5629 8443 5687 8449
rect 3605 8415 3663 8421
rect 3605 8381 3617 8415
rect 3651 8412 3663 8415
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3651 8384 3709 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 3712 8276 3740 8375
rect 4890 8372 4896 8424
rect 4948 8412 4954 8424
rect 5644 8412 5672 8443
rect 5810 8440 5816 8492
rect 5868 8480 5874 8492
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5868 8452 6009 8480
rect 5868 8440 5874 8452
rect 5997 8449 6009 8452
rect 6043 8449 6055 8483
rect 5997 8443 6055 8449
rect 6178 8440 6184 8492
rect 6236 8480 6242 8492
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6236 8452 6561 8480
rect 6236 8440 6242 8452
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7374 8480 7380 8492
rect 6871 8452 7380 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7926 8440 7932 8492
rect 7984 8440 7990 8492
rect 4948 8384 5672 8412
rect 4948 8372 4954 8384
rect 5718 8372 5724 8424
rect 5776 8412 5782 8424
rect 6196 8412 6224 8440
rect 5776 8384 6224 8412
rect 7009 8415 7067 8421
rect 5776 8372 5782 8384
rect 7009 8381 7021 8415
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 4706 8304 4712 8356
rect 4764 8344 4770 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 4764 8316 5825 8344
rect 4764 8304 4770 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5813 8307 5871 8313
rect 6089 8347 6147 8353
rect 6089 8313 6101 8347
rect 6135 8344 6147 8347
rect 6641 8347 6699 8353
rect 6641 8344 6653 8347
rect 6135 8316 6653 8344
rect 6135 8313 6147 8316
rect 6089 8307 6147 8313
rect 6641 8313 6653 8316
rect 6687 8313 6699 8347
rect 6641 8307 6699 8313
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 7024 8344 7052 8375
rect 6880 8316 7052 8344
rect 6880 8304 6886 8316
rect 7466 8304 7472 8356
rect 7524 8344 7530 8356
rect 7745 8347 7803 8353
rect 7745 8344 7757 8347
rect 7524 8316 7757 8344
rect 7524 8304 7530 8316
rect 7745 8313 7757 8316
rect 7791 8313 7803 8347
rect 7745 8307 7803 8313
rect 5442 8276 5448 8288
rect 3384 8248 5448 8276
rect 3384 8236 3390 8248
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 5994 8236 6000 8288
rect 6052 8276 6058 8288
rect 6365 8279 6423 8285
rect 6365 8276 6377 8279
rect 6052 8248 6377 8276
rect 6052 8236 6058 8248
rect 6365 8245 6377 8248
rect 6411 8245 6423 8279
rect 6365 8239 6423 8245
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 7653 8279 7711 8285
rect 7653 8276 7665 8279
rect 7248 8248 7665 8276
rect 7248 8236 7254 8248
rect 7653 8245 7665 8248
rect 7699 8245 7711 8279
rect 7653 8239 7711 8245
rect 1104 8186 8280 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 8280 8186
rect 1104 8112 8280 8134
rect 3786 8032 3792 8084
rect 3844 8032 3850 8084
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 5261 8075 5319 8081
rect 5261 8072 5273 8075
rect 4856 8044 5273 8072
rect 4856 8032 4862 8044
rect 5261 8041 5273 8044
rect 5307 8041 5319 8075
rect 5810 8072 5816 8084
rect 5261 8035 5319 8041
rect 5460 8044 5816 8072
rect 5460 8004 5488 8044
rect 5810 8032 5816 8044
rect 5868 8072 5874 8084
rect 5868 8044 6500 8072
rect 5868 8032 5874 8044
rect 4448 7976 5488 8004
rect 4448 7945 4476 7976
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7905 4491 7939
rect 4433 7899 4491 7905
rect 5442 7896 5448 7948
rect 5500 7896 5506 7948
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 3326 7868 3332 7880
rect 1443 7840 3332 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 3326 7828 3332 7840
rect 3384 7828 3390 7880
rect 3421 7871 3479 7877
rect 3421 7837 3433 7871
rect 3467 7837 3479 7871
rect 3421 7831 3479 7837
rect 4157 7871 4215 7877
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4614 7868 4620 7880
rect 4203 7840 4620 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 1664 7803 1722 7809
rect 1664 7769 1676 7803
rect 1710 7800 1722 7803
rect 1762 7800 1768 7812
rect 1710 7772 1768 7800
rect 1710 7769 1722 7772
rect 1664 7763 1722 7769
rect 1762 7760 1768 7772
rect 1820 7760 1826 7812
rect 3436 7800 3464 7831
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 4706 7828 4712 7880
rect 4764 7828 4770 7880
rect 4890 7828 4896 7880
rect 4948 7868 4954 7880
rect 5258 7868 5264 7880
rect 4948 7840 5264 7868
rect 4948 7828 4954 7840
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 5534 7868 5540 7880
rect 5408 7840 5540 7868
rect 5408 7828 5414 7840
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5712 7871 5770 7877
rect 5712 7837 5724 7871
rect 5758 7868 5770 7871
rect 5994 7868 6000 7880
rect 5758 7840 6000 7868
rect 5758 7837 5770 7840
rect 5712 7831 5770 7837
rect 5994 7828 6000 7840
rect 6052 7828 6058 7880
rect 6472 7868 6500 8044
rect 6822 8032 6828 8084
rect 6880 8032 6886 8084
rect 7374 8032 7380 8084
rect 7432 8032 7438 8084
rect 7009 7871 7067 7877
rect 7009 7868 7021 7871
rect 6472 7840 7021 7868
rect 7009 7837 7021 7840
rect 7055 7837 7067 7871
rect 7009 7831 7067 7837
rect 7190 7828 7196 7880
rect 7248 7828 7254 7880
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 7926 7828 7932 7880
rect 7984 7828 7990 7880
rect 2792 7772 3464 7800
rect 4249 7803 4307 7809
rect 2792 7744 2820 7772
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 5810 7800 5816 7812
rect 4295 7772 5816 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 5810 7760 5816 7772
rect 5868 7760 5874 7812
rect 2774 7692 2780 7744
rect 2832 7692 2838 7744
rect 2866 7692 2872 7744
rect 2924 7692 2930 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 5077 7735 5135 7741
rect 5077 7732 5089 7735
rect 4672 7704 5089 7732
rect 4672 7692 4678 7704
rect 5077 7701 5089 7704
rect 5123 7701 5135 7735
rect 5077 7695 5135 7701
rect 7650 7692 7656 7744
rect 7708 7692 7714 7744
rect 7742 7692 7748 7744
rect 7800 7692 7806 7744
rect 1104 7642 8280 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 8280 7642
rect 1104 7568 8280 7590
rect 1302 7488 1308 7540
rect 1360 7528 1366 7540
rect 1489 7531 1547 7537
rect 1489 7528 1501 7531
rect 1360 7500 1501 7528
rect 1360 7488 1366 7500
rect 1489 7497 1501 7500
rect 1535 7497 1547 7531
rect 1489 7491 1547 7497
rect 1762 7488 1768 7540
rect 1820 7488 1826 7540
rect 2133 7531 2191 7537
rect 2133 7497 2145 7531
rect 2179 7528 2191 7531
rect 2866 7528 2872 7540
rect 2179 7500 2872 7528
rect 2179 7497 2191 7500
rect 2133 7491 2191 7497
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 3786 7528 3792 7540
rect 3384 7500 3792 7528
rect 3384 7488 3390 7500
rect 3786 7488 3792 7500
rect 3844 7488 3850 7540
rect 3970 7488 3976 7540
rect 4028 7528 4034 7540
rect 4706 7528 4712 7540
rect 4028 7500 4712 7528
rect 4028 7488 4034 7500
rect 4706 7488 4712 7500
rect 4764 7488 4770 7540
rect 7282 7528 7288 7540
rect 6012 7500 7288 7528
rect 5718 7420 5724 7472
rect 5776 7420 5782 7472
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 2774 7392 2780 7404
rect 1719 7364 2780 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 2774 7352 2780 7364
rect 2832 7352 2838 7404
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7392 4675 7395
rect 4706 7392 4712 7404
rect 4663 7364 4712 7392
rect 4663 7361 4675 7364
rect 4617 7355 4675 7361
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 6012 7401 6040 7500
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7742 7488 7748 7540
rect 7800 7488 7806 7540
rect 6365 7463 6423 7469
rect 6365 7429 6377 7463
rect 6411 7460 6423 7463
rect 6638 7460 6644 7472
rect 6411 7432 6644 7460
rect 6411 7429 6423 7432
rect 6365 7423 6423 7429
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 6730 7420 6736 7472
rect 6788 7460 6794 7472
rect 7760 7460 7788 7488
rect 6788 7432 7788 7460
rect 6788 7420 6794 7432
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6546 7352 6552 7404
rect 6604 7352 6610 7404
rect 7024 7401 7052 7432
rect 6825 7395 6883 7401
rect 6825 7361 6837 7395
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 7009 7395 7067 7401
rect 7009 7361 7021 7395
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 2225 7327 2283 7333
rect 2225 7293 2237 7327
rect 2271 7293 2283 7327
rect 2225 7287 2283 7293
rect 2409 7327 2467 7333
rect 2409 7293 2421 7327
rect 2455 7324 2467 7327
rect 2498 7324 2504 7336
rect 2455 7296 2504 7324
rect 2455 7293 2467 7296
rect 2409 7287 2467 7293
rect 1854 7216 1860 7268
rect 1912 7256 1918 7268
rect 2240 7256 2268 7287
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7324 5411 7327
rect 5442 7324 5448 7336
rect 5399 7296 5448 7324
rect 5399 7293 5411 7296
rect 5353 7287 5411 7293
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7324 5963 7327
rect 6564 7324 6592 7352
rect 5951 7296 6592 7324
rect 6840 7324 6868 7355
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7558 7352 7564 7404
rect 7616 7352 7622 7404
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 7834 7392 7840 7404
rect 7791 7364 7840 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 7834 7352 7840 7364
rect 7892 7352 7898 7404
rect 7101 7327 7159 7333
rect 7101 7324 7113 7327
rect 6840 7296 7113 7324
rect 5951 7293 5963 7296
rect 5905 7287 5963 7293
rect 7101 7293 7113 7296
rect 7147 7293 7159 7327
rect 7101 7287 7159 7293
rect 5810 7256 5816 7268
rect 1912 7228 5816 7256
rect 1912 7216 1918 7228
rect 5810 7216 5816 7228
rect 5868 7216 5874 7268
rect 6730 7256 6736 7268
rect 6012 7228 6736 7256
rect 4709 7191 4767 7197
rect 4709 7157 4721 7191
rect 4755 7188 4767 7191
rect 4798 7188 4804 7200
rect 4755 7160 4804 7188
rect 4755 7157 4767 7160
rect 4709 7151 4767 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 6012 7197 6040 7228
rect 6730 7216 6736 7228
rect 6788 7216 6794 7268
rect 5997 7191 6055 7197
rect 5997 7157 6009 7191
rect 6043 7157 6055 7191
rect 5997 7151 6055 7157
rect 6178 7148 6184 7200
rect 6236 7148 6242 7200
rect 1104 7098 8280 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 8280 7098
rect 1104 7024 8280 7046
rect 3970 6984 3976 6996
rect 2240 6956 3976 6984
rect 1854 6808 1860 6860
rect 1912 6808 1918 6860
rect 2041 6851 2099 6857
rect 2041 6817 2053 6851
rect 2087 6848 2099 6851
rect 2240 6848 2268 6956
rect 3970 6944 3976 6956
rect 4028 6944 4034 6996
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 5258 6984 5264 6996
rect 5215 6956 5264 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 7193 6987 7251 6993
rect 7193 6953 7205 6987
rect 7239 6984 7251 6987
rect 7558 6984 7564 6996
rect 7239 6956 7564 6984
rect 7239 6953 7251 6956
rect 7193 6947 7251 6953
rect 7558 6944 7564 6956
rect 7616 6944 7622 6996
rect 3605 6919 3663 6925
rect 3605 6885 3617 6919
rect 3651 6885 3663 6919
rect 3605 6879 3663 6885
rect 2087 6820 2268 6848
rect 2087 6817 2099 6820
rect 2041 6811 2099 6817
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 2774 6780 2780 6792
rect 2271 6752 2780 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 2774 6740 2780 6752
rect 2832 6780 2838 6792
rect 3326 6780 3332 6792
rect 2832 6752 3332 6780
rect 2832 6740 2838 6752
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3620 6780 3648 6879
rect 5534 6876 5540 6928
rect 5592 6876 5598 6928
rect 6914 6916 6920 6928
rect 6472 6888 6920 6916
rect 3786 6808 3792 6860
rect 3844 6808 3850 6860
rect 6472 6857 6500 6888
rect 6914 6876 6920 6888
rect 6972 6916 6978 6928
rect 7834 6916 7840 6928
rect 6972 6888 7840 6916
rect 6972 6876 6978 6888
rect 7834 6876 7840 6888
rect 7892 6876 7898 6928
rect 6457 6851 6515 6857
rect 6457 6817 6469 6851
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 6549 6851 6607 6857
rect 6549 6817 6561 6851
rect 6595 6848 6607 6851
rect 7098 6848 7104 6860
rect 6595 6820 7104 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 7098 6808 7104 6820
rect 7156 6808 7162 6860
rect 5442 6780 5448 6792
rect 3620 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6780 5506 6792
rect 6365 6783 6423 6789
rect 5500 6752 5672 6780
rect 5500 6740 5506 6752
rect 5644 6724 5672 6752
rect 6365 6749 6377 6783
rect 6411 6749 6423 6783
rect 6365 6743 6423 6749
rect 6641 6783 6699 6789
rect 6641 6749 6653 6783
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 2498 6721 2504 6724
rect 2492 6712 2504 6721
rect 2411 6684 2504 6712
rect 2492 6675 2504 6684
rect 2556 6712 2562 6724
rect 4056 6715 4114 6721
rect 2556 6684 4016 6712
rect 2498 6672 2504 6675
rect 2556 6672 2562 6684
rect 1394 6604 1400 6656
rect 1452 6604 1458 6656
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 2314 6644 2320 6656
rect 1811 6616 2320 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 2314 6604 2320 6616
rect 2372 6604 2378 6656
rect 3988 6644 4016 6684
rect 4056 6681 4068 6715
rect 4102 6712 4114 6715
rect 5350 6712 5356 6724
rect 4102 6684 5356 6712
rect 4102 6681 4114 6684
rect 4056 6675 4114 6681
rect 5350 6672 5356 6684
rect 5408 6672 5414 6724
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 5905 6715 5963 6721
rect 5905 6712 5917 6715
rect 5684 6684 5917 6712
rect 5684 6672 5690 6684
rect 5905 6681 5917 6684
rect 5951 6681 5963 6715
rect 6380 6712 6408 6743
rect 6656 6712 6684 6743
rect 6730 6740 6736 6792
rect 6788 6780 6794 6792
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6788 6752 6837 6780
rect 6788 6740 6794 6752
rect 6825 6749 6837 6752
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 7282 6780 7288 6792
rect 7055 6752 7288 6780
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 7374 6740 7380 6792
rect 7432 6740 7438 6792
rect 7650 6740 7656 6792
rect 7708 6740 7714 6792
rect 7742 6740 7748 6792
rect 7800 6780 7806 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7800 6752 7849 6780
rect 7800 6740 7806 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 6917 6715 6975 6721
rect 6917 6712 6929 6715
rect 6380 6684 6500 6712
rect 6656 6684 6929 6712
rect 5905 6675 5963 6681
rect 5258 6644 5264 6656
rect 3988 6616 5264 6644
rect 5258 6604 5264 6616
rect 5316 6644 5322 6656
rect 5445 6647 5503 6653
rect 5445 6644 5457 6647
rect 5316 6616 5457 6644
rect 5316 6604 5322 6616
rect 5445 6613 5457 6616
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 6181 6647 6239 6653
rect 6181 6613 6193 6647
rect 6227 6644 6239 6647
rect 6362 6644 6368 6656
rect 6227 6616 6368 6644
rect 6227 6613 6239 6616
rect 6181 6607 6239 6613
rect 6362 6604 6368 6616
rect 6420 6604 6426 6656
rect 6472 6644 6500 6684
rect 6917 6681 6929 6684
rect 6963 6681 6975 6715
rect 6917 6675 6975 6681
rect 7392 6644 7420 6740
rect 6472 6616 7420 6644
rect 1104 6554 8280 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 8280 6554
rect 1104 6480 8280 6502
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 5810 6400 5816 6452
rect 5868 6440 5874 6452
rect 6733 6443 6791 6449
rect 6733 6440 6745 6443
rect 5868 6412 6745 6440
rect 5868 6400 5874 6412
rect 6733 6409 6745 6412
rect 6779 6409 6791 6443
rect 6733 6403 6791 6409
rect 7745 6443 7803 6449
rect 7745 6409 7757 6443
rect 7791 6409 7803 6443
rect 7745 6403 7803 6409
rect 1394 6332 1400 6384
rect 1452 6372 1458 6384
rect 2510 6375 2568 6381
rect 2510 6372 2522 6375
rect 1452 6344 2522 6372
rect 1452 6332 1458 6344
rect 2510 6341 2522 6344
rect 2556 6341 2568 6375
rect 2510 6335 2568 6341
rect 3510 6332 3516 6384
rect 3568 6332 3574 6384
rect 7760 6372 7788 6403
rect 7484 6344 7788 6372
rect 7484 6316 7512 6344
rect 2774 6264 2780 6316
rect 2832 6264 2838 6316
rect 6362 6264 6368 6316
rect 6420 6264 6426 6316
rect 6546 6264 6552 6316
rect 6604 6264 6610 6316
rect 7466 6264 7472 6316
rect 7524 6264 7530 6316
rect 7653 6307 7711 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 7742 6304 7748 6316
rect 7699 6276 7748 6304
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 7742 6264 7748 6276
rect 7800 6264 7806 6316
rect 7926 6264 7932 6316
rect 7984 6264 7990 6316
rect 4798 6196 4804 6248
rect 4856 6236 4862 6248
rect 5905 6239 5963 6245
rect 5905 6236 5917 6239
rect 4856 6208 5917 6236
rect 4856 6196 4862 6208
rect 5905 6205 5917 6208
rect 5951 6205 5963 6239
rect 5905 6199 5963 6205
rect 1394 6060 1400 6112
rect 1452 6060 1458 6112
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 4801 6103 4859 6109
rect 4801 6100 4813 6103
rect 4764 6072 4813 6100
rect 4764 6060 4770 6072
rect 4801 6069 4813 6072
rect 4847 6069 4859 6103
rect 4801 6063 4859 6069
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 5776 6072 6377 6100
rect 5776 6060 5782 6072
rect 6365 6069 6377 6072
rect 6411 6069 6423 6103
rect 6365 6063 6423 6069
rect 7006 6060 7012 6112
rect 7064 6100 7070 6112
rect 7653 6103 7711 6109
rect 7653 6100 7665 6103
rect 7064 6072 7665 6100
rect 7064 6060 7070 6072
rect 7653 6069 7665 6072
rect 7699 6069 7711 6103
rect 7653 6063 7711 6069
rect 1104 6010 8280 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 8280 6010
rect 1104 5936 8280 5958
rect 2314 5856 2320 5908
rect 2372 5856 2378 5908
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4120 5868 4445 5896
rect 4120 5856 4126 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 6178 5856 6184 5908
rect 6236 5856 6242 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 7837 5899 7895 5905
rect 7837 5896 7849 5899
rect 7708 5868 7849 5896
rect 7708 5856 7714 5868
rect 7837 5865 7849 5868
rect 7883 5865 7895 5899
rect 7837 5859 7895 5865
rect 4249 5831 4307 5837
rect 4249 5797 4261 5831
rect 4295 5828 4307 5831
rect 4890 5828 4896 5840
rect 4295 5800 4896 5828
rect 4295 5797 4307 5800
rect 4249 5791 4307 5797
rect 1394 5720 1400 5772
rect 1452 5760 1458 5772
rect 1673 5763 1731 5769
rect 1673 5760 1685 5763
rect 1452 5732 1685 5760
rect 1452 5720 1458 5732
rect 1673 5729 1685 5732
rect 1719 5729 1731 5763
rect 4264 5760 4292 5791
rect 4890 5788 4896 5800
rect 4948 5788 4954 5840
rect 5718 5828 5724 5840
rect 5460 5800 5724 5828
rect 1673 5723 1731 5729
rect 3988 5732 4292 5760
rect 4341 5763 4399 5769
rect 2958 5652 2964 5704
rect 3016 5652 3022 5704
rect 3988 5701 4016 5732
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 5460 5760 5488 5800
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 7374 5788 7380 5840
rect 7432 5788 7438 5840
rect 4387 5732 5488 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 5534 5720 5540 5772
rect 5592 5720 5598 5772
rect 7392 5760 7420 5788
rect 6104 5732 7420 5760
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 3804 5624 3832 5655
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5692 4583 5695
rect 4614 5692 4620 5704
rect 4571 5664 4620 5692
rect 4571 5661 4583 5664
rect 4525 5655 4583 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 4798 5652 4804 5704
rect 4856 5652 4862 5704
rect 6104 5701 6132 5732
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6273 5695 6331 5701
rect 6273 5661 6285 5695
rect 6319 5692 6331 5695
rect 6641 5695 6699 5701
rect 6641 5692 6653 5695
rect 6319 5664 6653 5692
rect 6319 5661 6331 5664
rect 6273 5655 6331 5661
rect 6641 5661 6653 5664
rect 6687 5692 6699 5695
rect 6730 5692 6736 5704
rect 6687 5664 6736 5692
rect 6687 5661 6699 5664
rect 6641 5655 6699 5661
rect 6730 5652 6736 5664
rect 6788 5652 6794 5704
rect 6840 5701 6868 5732
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7193 5695 7251 5701
rect 7193 5661 7205 5695
rect 7239 5661 7251 5695
rect 7193 5655 7251 5661
rect 4893 5627 4951 5633
rect 4893 5624 4905 5627
rect 3804 5596 4905 5624
rect 4893 5593 4905 5596
rect 4939 5593 4951 5627
rect 4893 5587 4951 5593
rect 6549 5627 6607 5633
rect 6549 5593 6561 5627
rect 6595 5624 6607 5627
rect 7006 5624 7012 5636
rect 6595 5596 7012 5624
rect 6595 5593 6607 5596
rect 6549 5587 6607 5593
rect 7006 5584 7012 5596
rect 7064 5584 7070 5636
rect 7208 5624 7236 5655
rect 7374 5652 7380 5704
rect 7432 5652 7438 5704
rect 7466 5652 7472 5704
rect 7524 5692 7530 5704
rect 7653 5695 7711 5701
rect 7653 5692 7665 5695
rect 7524 5664 7665 5692
rect 7524 5652 7530 5664
rect 7653 5661 7665 5664
rect 7699 5661 7711 5695
rect 7653 5655 7711 5661
rect 7558 5624 7564 5636
rect 7116 5596 7564 5624
rect 2406 5516 2412 5568
rect 2464 5516 2470 5568
rect 5905 5559 5963 5565
rect 5905 5525 5917 5559
rect 5951 5556 5963 5559
rect 6086 5556 6092 5568
rect 5951 5528 6092 5556
rect 5951 5525 5963 5528
rect 5905 5519 5963 5525
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6638 5516 6644 5568
rect 6696 5556 6702 5568
rect 7116 5565 7144 5596
rect 7558 5584 7564 5596
rect 7616 5584 7622 5636
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6696 5528 6745 5556
rect 6696 5516 6702 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6733 5519 6791 5525
rect 7101 5559 7159 5565
rect 7101 5525 7113 5559
rect 7147 5525 7159 5559
rect 7101 5519 7159 5525
rect 1104 5466 8280 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 8280 5466
rect 1104 5392 8280 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 1489 5355 1547 5361
rect 1489 5352 1501 5355
rect 1360 5324 1501 5352
rect 1360 5312 1366 5324
rect 1489 5321 1501 5324
rect 1535 5321 1547 5355
rect 1489 5315 1547 5321
rect 2225 5355 2283 5361
rect 2225 5321 2237 5355
rect 2271 5352 2283 5355
rect 2406 5352 2412 5364
rect 2271 5324 2412 5352
rect 2271 5321 2283 5324
rect 2225 5315 2283 5321
rect 2406 5312 2412 5324
rect 2464 5312 2470 5364
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 5442 5352 5448 5364
rect 4120 5324 5448 5352
rect 4120 5312 4126 5324
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 7374 5312 7380 5364
rect 7432 5352 7438 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7432 5324 7849 5352
rect 7432 5312 7438 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 2952 5287 3010 5293
rect 2952 5253 2964 5287
rect 2998 5284 3010 5287
rect 3694 5284 3700 5296
rect 2998 5256 3700 5284
rect 2998 5253 3010 5256
rect 2952 5247 3010 5253
rect 3694 5244 3700 5256
rect 3752 5284 3758 5296
rect 3970 5284 3976 5296
rect 3752 5256 3976 5284
rect 3752 5244 3758 5256
rect 3970 5244 3976 5256
rect 4028 5244 4034 5296
rect 7006 5284 7012 5296
rect 6564 5256 7012 5284
rect 1394 5176 1400 5228
rect 1452 5216 1458 5228
rect 1673 5219 1731 5225
rect 1673 5216 1685 5219
rect 1452 5188 1685 5216
rect 1452 5176 1458 5188
rect 1673 5185 1685 5188
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4571 5188 4997 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 4985 5185 4997 5188
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6564 5225 6592 5256
rect 7006 5244 7012 5256
rect 7064 5244 7070 5296
rect 6457 5219 6515 5225
rect 6457 5216 6469 5219
rect 6236 5188 6469 5216
rect 6236 5176 6242 5188
rect 6457 5185 6469 5188
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5185 6607 5219
rect 6549 5179 6607 5185
rect 6638 5176 6644 5228
rect 6696 5176 6702 5228
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 7282 5216 7288 5228
rect 7239 5188 7288 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 7282 5176 7288 5188
rect 7340 5176 7346 5228
rect 7374 5176 7380 5228
rect 7432 5176 7438 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 7742 5216 7748 5228
rect 7699 5188 7748 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 7742 5176 7748 5188
rect 7800 5176 7806 5228
rect 2317 5151 2375 5157
rect 2317 5117 2329 5151
rect 2363 5148 2375 5151
rect 2406 5148 2412 5160
rect 2363 5120 2412 5148
rect 2363 5117 2375 5120
rect 2317 5111 2375 5117
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 2498 5108 2504 5160
rect 2556 5108 2562 5160
rect 2685 5151 2743 5157
rect 2685 5117 2697 5151
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5117 4675 5151
rect 4617 5111 4675 5117
rect 4801 5151 4859 5157
rect 4801 5117 4813 5151
rect 4847 5148 4859 5151
rect 5258 5148 5264 5160
rect 4847 5120 5264 5148
rect 4847 5117 4859 5120
rect 4801 5111 4859 5117
rect 1394 5040 1400 5092
rect 1452 5080 1458 5092
rect 2700 5080 2728 5111
rect 1452 5052 2728 5080
rect 1452 5040 1458 5052
rect 3970 5040 3976 5092
rect 4028 5080 4034 5092
rect 4157 5083 4215 5089
rect 4157 5080 4169 5083
rect 4028 5052 4169 5080
rect 4028 5040 4034 5052
rect 4157 5049 4169 5052
rect 4203 5049 4215 5083
rect 4632 5080 4660 5111
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 5350 5108 5356 5160
rect 5408 5148 5414 5160
rect 5537 5151 5595 5157
rect 5537 5148 5549 5151
rect 5408 5120 5549 5148
rect 5408 5108 5414 5120
rect 5537 5117 5549 5120
rect 5583 5117 5595 5151
rect 5537 5111 5595 5117
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5148 6791 5151
rect 7466 5148 7472 5160
rect 6779 5120 7472 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 7466 5108 7472 5120
rect 7524 5108 7530 5160
rect 5718 5080 5724 5092
rect 4632 5052 5724 5080
rect 4157 5043 4215 5049
rect 5718 5040 5724 5052
rect 5776 5080 5782 5092
rect 6917 5083 6975 5089
rect 6917 5080 6929 5083
rect 5776 5052 6929 5080
rect 5776 5040 5782 5052
rect 6917 5049 6929 5052
rect 6963 5049 6975 5083
rect 6917 5043 6975 5049
rect 1854 4972 1860 5024
rect 1912 4972 1918 5024
rect 1104 4922 8280 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 8280 4922
rect 1104 4848 8280 4870
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 2958 4808 2964 4820
rect 2823 4780 2964 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 5721 4811 5779 4817
rect 5721 4777 5733 4811
rect 5767 4808 5779 4811
rect 5902 4808 5908 4820
rect 5767 4780 5908 4808
rect 5767 4777 5779 4780
rect 5721 4771 5779 4777
rect 5902 4768 5908 4780
rect 5960 4768 5966 4820
rect 7098 4768 7104 4820
rect 7156 4808 7162 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 7156 4780 7297 4808
rect 7156 4768 7162 4780
rect 7285 4777 7297 4780
rect 7331 4777 7343 4811
rect 7285 4771 7343 4777
rect 5626 4700 5632 4752
rect 5684 4700 5690 4752
rect 1394 4632 1400 4684
rect 1452 4632 1458 4684
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4672 5319 4675
rect 5442 4672 5448 4684
rect 5307 4644 5448 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 5442 4632 5448 4644
rect 5500 4632 5506 4684
rect 7006 4632 7012 4684
rect 7064 4672 7070 4684
rect 7064 4644 7788 4672
rect 7064 4632 7070 4644
rect 1412 4604 1440 4632
rect 2774 4604 2780 4616
rect 1412 4576 2780 4604
rect 2774 4564 2780 4576
rect 2832 4604 2838 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 2832 4576 3801 4604
rect 2832 4564 2838 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 3789 4567 3847 4573
rect 4056 4607 4114 4613
rect 4056 4573 4068 4607
rect 4102 4573 4114 4607
rect 4056 4567 4114 4573
rect 1664 4539 1722 4545
rect 1664 4505 1676 4539
rect 1710 4536 1722 4539
rect 1854 4536 1860 4548
rect 1710 4508 1860 4536
rect 1710 4505 1722 4508
rect 1664 4499 1722 4505
rect 1854 4496 1860 4508
rect 1912 4496 1918 4548
rect 3804 4468 3832 4567
rect 3970 4496 3976 4548
rect 4028 4536 4034 4548
rect 4080 4536 4108 4567
rect 6546 4564 6552 4616
rect 6604 4564 6610 4616
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 7156 4576 7481 4604
rect 7156 4564 7162 4576
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7558 4564 7564 4616
rect 7616 4564 7622 4616
rect 7650 4564 7656 4616
rect 7708 4564 7714 4616
rect 7760 4613 7788 4644
rect 7745 4607 7803 4613
rect 7745 4573 7757 4607
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 4028 4508 4108 4536
rect 4028 4496 4034 4508
rect 4798 4468 4804 4480
rect 3804 4440 4804 4468
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5169 4471 5227 4477
rect 5169 4437 5181 4471
rect 5215 4468 5227 4471
rect 5350 4468 5356 4480
rect 5215 4440 5356 4468
rect 5215 4437 5227 4440
rect 5169 4431 5227 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 7193 4471 7251 4477
rect 7193 4468 7205 4471
rect 6788 4440 7205 4468
rect 6788 4428 6794 4440
rect 7193 4437 7205 4440
rect 7239 4437 7251 4471
rect 7193 4431 7251 4437
rect 1104 4378 8280 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 8280 4378
rect 1104 4304 8280 4326
rect 6730 4224 6736 4276
rect 6788 4224 6794 4276
rect 7466 4224 7472 4276
rect 7524 4224 7530 4276
rect 5718 4196 5724 4208
rect 4724 4168 5724 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2958 4128 2964 4140
rect 1719 4100 2964 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2958 4088 2964 4100
rect 3016 4088 3022 4140
rect 3513 4131 3571 4137
rect 3513 4097 3525 4131
rect 3559 4128 3571 4131
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3559 4100 3985 4128
rect 3559 4097 3571 4100
rect 3513 4091 3571 4097
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 1394 4020 1400 4072
rect 1452 4060 1458 4072
rect 1949 4063 2007 4069
rect 1949 4060 1961 4063
rect 1452 4032 1961 4060
rect 1452 4020 1458 4032
rect 1949 4029 1961 4032
rect 1995 4029 2007 4063
rect 1949 4023 2007 4029
rect 2866 4020 2872 4072
rect 2924 4020 2930 4072
rect 3694 4020 3700 4072
rect 3752 4020 3758 4072
rect 3881 4063 3939 4069
rect 3881 4029 3893 4063
rect 3927 4060 3939 4063
rect 4724 4060 4752 4168
rect 5718 4156 5724 4168
rect 5776 4156 5782 4208
rect 7558 4156 7564 4208
rect 7616 4196 7622 4208
rect 7929 4199 7987 4205
rect 7929 4196 7941 4199
rect 7616 4168 7941 4196
rect 7616 4156 7622 4168
rect 7929 4165 7941 4168
rect 7975 4165 7987 4199
rect 7929 4159 7987 4165
rect 4798 4088 4804 4140
rect 4856 4088 4862 4140
rect 5068 4131 5126 4137
rect 5068 4097 5080 4131
rect 5114 4128 5126 4131
rect 5114 4100 5856 4128
rect 5114 4097 5126 4100
rect 5068 4091 5126 4097
rect 3927 4032 4752 4060
rect 3927 4029 3939 4032
rect 3881 4023 3939 4029
rect 1302 3952 1308 4004
rect 1360 3992 1366 4004
rect 1489 3995 1547 4001
rect 1489 3992 1501 3995
rect 1360 3964 1501 3992
rect 1360 3952 1366 3964
rect 1489 3961 1501 3964
rect 1535 3961 1547 3995
rect 1489 3955 1547 3961
rect 2406 3952 2412 4004
rect 2464 3992 2470 4004
rect 5828 3992 5856 4100
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 5960 4100 6960 4128
rect 5960 4088 5966 4100
rect 6086 4020 6092 4072
rect 6144 4060 6150 4072
rect 6932 4069 6960 4100
rect 7190 4088 7196 4140
rect 7248 4088 7254 4140
rect 7466 4088 7472 4140
rect 7524 4128 7530 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7524 4100 7665 4128
rect 7524 4088 7530 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 6144 4032 6837 4060
rect 6144 4020 6150 4032
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 7742 4060 7748 4072
rect 7156 4032 7748 4060
rect 7156 4020 7162 4032
rect 7742 4020 7748 4032
rect 7800 4020 7806 4072
rect 6365 3995 6423 4001
rect 6365 3992 6377 3995
rect 2464 3964 4844 3992
rect 5828 3964 6377 3992
rect 2464 3952 2470 3964
rect 2314 3884 2320 3936
rect 2372 3924 2378 3936
rect 2593 3927 2651 3933
rect 2593 3924 2605 3927
rect 2372 3896 2605 3924
rect 2372 3884 2378 3896
rect 2593 3893 2605 3896
rect 2639 3893 2651 3927
rect 2593 3887 2651 3893
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 4614 3924 4620 3936
rect 4387 3896 4620 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4816 3924 4844 3964
rect 6365 3961 6377 3964
rect 6411 3961 6423 3995
rect 6365 3955 6423 3961
rect 7377 3995 7435 4001
rect 7377 3961 7389 3995
rect 7423 3992 7435 3995
rect 7926 3992 7932 4004
rect 7423 3964 7932 3992
rect 7423 3961 7435 3964
rect 7377 3955 7435 3961
rect 7926 3952 7932 3964
rect 7984 3952 7990 4004
rect 6086 3924 6092 3936
rect 4816 3896 6092 3924
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6181 3927 6239 3933
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6546 3924 6552 3936
rect 6227 3896 6552 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7653 3927 7711 3933
rect 7653 3924 7665 3927
rect 7340 3896 7665 3924
rect 7340 3884 7346 3896
rect 7653 3893 7665 3896
rect 7699 3893 7711 3927
rect 7653 3887 7711 3893
rect 1104 3834 8280 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 8280 3834
rect 1104 3760 8280 3782
rect 1394 3680 1400 3732
rect 1452 3680 1458 3732
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 5077 3723 5135 3729
rect 5077 3720 5089 3723
rect 4856 3692 5089 3720
rect 4856 3680 4862 3692
rect 5077 3689 5089 3692
rect 5123 3689 5135 3723
rect 5077 3683 5135 3689
rect 6641 3723 6699 3729
rect 6641 3689 6653 3723
rect 6687 3720 6699 3723
rect 7098 3720 7104 3732
rect 6687 3692 7104 3720
rect 6687 3689 6699 3692
rect 6641 3683 6699 3689
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 7285 3723 7343 3729
rect 7285 3689 7297 3723
rect 7331 3720 7343 3723
rect 7374 3720 7380 3732
rect 7331 3692 7380 3720
rect 7331 3689 7343 3692
rect 7285 3683 7343 3689
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 6089 3655 6147 3661
rect 6089 3621 6101 3655
rect 6135 3652 6147 3655
rect 7190 3652 7196 3664
rect 6135 3624 7196 3652
rect 6135 3621 6147 3624
rect 6089 3615 6147 3621
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 2774 3544 2780 3596
rect 2832 3544 2838 3596
rect 7834 3584 7840 3596
rect 5920 3556 7840 3584
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3516 3847 3519
rect 4706 3516 4712 3528
rect 3835 3488 4712 3516
rect 3835 3485 3847 3488
rect 3789 3479 3847 3485
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 5920 3525 5948 3556
rect 7834 3544 7840 3556
rect 7892 3544 7898 3596
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 6178 3476 6184 3528
rect 6236 3476 6242 3528
rect 6454 3476 6460 3528
rect 6512 3476 6518 3528
rect 6730 3476 6736 3528
rect 6788 3476 6794 3528
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3516 7251 3519
rect 7282 3516 7288 3528
rect 7239 3488 7288 3516
rect 7239 3485 7251 3488
rect 7193 3479 7251 3485
rect 1946 3408 1952 3460
rect 2004 3448 2010 3460
rect 2510 3451 2568 3457
rect 2510 3448 2522 3451
rect 2004 3420 2522 3448
rect 2004 3408 2010 3420
rect 2510 3417 2522 3420
rect 2556 3417 2568 3451
rect 7024 3448 7052 3479
rect 7282 3476 7288 3488
rect 7340 3476 7346 3528
rect 7466 3476 7472 3528
rect 7524 3476 7530 3528
rect 7742 3476 7748 3528
rect 7800 3476 7806 3528
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 7484 3448 7512 3476
rect 2510 3411 2568 3417
rect 6380 3420 7512 3448
rect 6380 3389 6408 3420
rect 6365 3383 6423 3389
rect 6365 3349 6377 3383
rect 6411 3349 6423 3383
rect 6365 3343 6423 3349
rect 6917 3383 6975 3389
rect 6917 3349 6929 3383
rect 6963 3380 6975 3383
rect 7006 3380 7012 3392
rect 6963 3352 7012 3380
rect 6963 3349 6975 3352
rect 6917 3343 6975 3349
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7098 3340 7104 3392
rect 7156 3340 7162 3392
rect 1104 3290 8280 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 8280 3290
rect 1104 3216 8280 3238
rect 1946 3136 1952 3188
rect 2004 3136 2010 3188
rect 2314 3136 2320 3188
rect 2372 3136 2378 3188
rect 2406 3136 2412 3188
rect 2464 3136 2470 3188
rect 2866 3136 2872 3188
rect 2924 3176 2930 3188
rect 3326 3176 3332 3188
rect 2924 3148 3332 3176
rect 2924 3136 2930 3148
rect 3326 3136 3332 3148
rect 3384 3176 3390 3188
rect 3789 3179 3847 3185
rect 3789 3176 3801 3179
rect 3384 3148 3801 3176
rect 3384 3136 3390 3148
rect 3789 3145 3801 3148
rect 3835 3145 3847 3179
rect 3789 3139 3847 3145
rect 4614 3136 4620 3188
rect 4672 3136 4678 3188
rect 5718 3136 5724 3188
rect 5776 3136 5782 3188
rect 7650 3136 7656 3188
rect 7708 3176 7714 3188
rect 7745 3179 7803 3185
rect 7745 3176 7757 3179
rect 7708 3148 7757 3176
rect 7708 3136 7714 3148
rect 7745 3145 7757 3148
rect 7791 3145 7803 3179
rect 7745 3139 7803 3145
rect 1394 3000 1400 3052
rect 1452 3040 1458 3052
rect 1673 3043 1731 3049
rect 1673 3040 1685 3043
rect 1452 3012 1685 3040
rect 1452 3000 1458 3012
rect 1673 3009 1685 3012
rect 1719 3009 1731 3043
rect 4632 3040 4660 3136
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 4856 3080 5212 3108
rect 4856 3068 4862 3080
rect 5184 3049 5212 3080
rect 4902 3043 4960 3049
rect 4902 3040 4914 3043
rect 4632 3012 4914 3040
rect 1673 3003 1731 3009
rect 4902 3009 4914 3012
rect 4948 3009 4960 3043
rect 4902 3003 4960 3009
rect 5169 3043 5227 3049
rect 5169 3009 5181 3043
rect 5215 3009 5227 3043
rect 5169 3003 5227 3009
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3040 5687 3043
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 5675 3012 6377 3040
rect 5675 3009 5687 3012
rect 5629 3003 5687 3009
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7156 3012 7573 3040
rect 7156 3000 7162 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2972 2651 2975
rect 3694 2972 3700 2984
rect 2639 2944 3700 2972
rect 2639 2941 2651 2944
rect 2593 2935 2651 2941
rect 3694 2932 3700 2944
rect 3752 2932 3758 2984
rect 5902 2932 5908 2984
rect 5960 2932 5966 2984
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 6917 2975 6975 2981
rect 6917 2972 6929 2975
rect 6052 2944 6929 2972
rect 6052 2932 6058 2944
rect 6917 2941 6929 2944
rect 6963 2941 6975 2975
rect 6917 2935 6975 2941
rect 7006 2932 7012 2984
rect 7064 2972 7070 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7064 2944 7297 2972
rect 7064 2932 7070 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 7377 2975 7435 2981
rect 7377 2941 7389 2975
rect 7423 2972 7435 2975
rect 7926 2972 7932 2984
rect 7423 2944 7932 2972
rect 7423 2941 7435 2944
rect 7377 2935 7435 2941
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 842 2864 848 2916
rect 900 2904 906 2916
rect 1489 2907 1547 2913
rect 1489 2904 1501 2907
rect 900 2876 1501 2904
rect 900 2864 906 2876
rect 1489 2873 1501 2876
rect 1535 2873 1547 2907
rect 1489 2867 1547 2873
rect 4798 2796 4804 2848
rect 4856 2836 4862 2848
rect 5261 2839 5319 2845
rect 5261 2836 5273 2839
rect 4856 2808 5273 2836
rect 4856 2796 4862 2808
rect 5261 2805 5273 2808
rect 5307 2805 5319 2839
rect 5261 2799 5319 2805
rect 1104 2746 8280 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 8280 2746
rect 1104 2672 8280 2694
rect 5350 2632 5356 2644
rect 4172 2604 5356 2632
rect 3326 2388 3332 2440
rect 3384 2388 3390 2440
rect 4172 2437 4200 2604
rect 5350 2592 5356 2604
rect 5408 2592 5414 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7282 2632 7288 2644
rect 6963 2604 7288 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 7742 2592 7748 2644
rect 7800 2632 7806 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7800 2604 7849 2632
rect 7800 2592 7806 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 7837 2595 7895 2601
rect 5629 2567 5687 2573
rect 5629 2533 5641 2567
rect 5675 2564 5687 2567
rect 5994 2564 6000 2576
rect 5675 2536 6000 2564
rect 5675 2533 5687 2536
rect 5629 2527 5687 2533
rect 5994 2524 6000 2536
rect 6052 2524 6058 2576
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 7653 2567 7711 2573
rect 7653 2564 7665 2567
rect 7248 2536 7665 2564
rect 7248 2524 7254 2536
rect 7653 2533 7665 2536
rect 7699 2533 7711 2567
rect 7653 2527 7711 2533
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7377 2499 7435 2505
rect 7377 2496 7389 2499
rect 7064 2468 7389 2496
rect 7064 2456 7070 2468
rect 7377 2465 7389 2468
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2397 4215 2431
rect 4157 2391 4215 2397
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 4338 2428 4344 2440
rect 4295 2400 4344 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 4338 2388 4344 2400
rect 4396 2388 4402 2440
rect 5994 2388 6000 2440
rect 6052 2388 6058 2440
rect 6546 2388 6552 2440
rect 6604 2388 6610 2440
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 4516 2363 4574 2369
rect 4516 2329 4528 2363
rect 4562 2360 4574 2363
rect 4798 2360 4804 2372
rect 4562 2332 4804 2360
rect 4562 2329 4574 2332
rect 4516 2323 4574 2329
rect 4798 2320 4804 2332
rect 4856 2320 4862 2372
rect 5276 2332 5856 2360
rect 5276 2304 5304 2332
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 3878 2292 3884 2304
rect 3559 2264 3884 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 3973 2295 4031 2301
rect 3973 2261 3985 2295
rect 4019 2292 4031 2295
rect 4430 2292 4436 2304
rect 4019 2264 4436 2292
rect 4019 2261 4031 2264
rect 3973 2255 4031 2261
rect 4430 2252 4436 2264
rect 4488 2252 4494 2304
rect 5258 2252 5264 2304
rect 5316 2252 5322 2304
rect 5828 2301 5856 2332
rect 5813 2295 5871 2301
rect 5813 2261 5825 2295
rect 5859 2261 5871 2295
rect 5813 2255 5871 2261
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6733 2295 6791 2301
rect 6733 2292 6745 2295
rect 6512 2264 6745 2292
rect 6512 2252 6518 2264
rect 6733 2261 6745 2264
rect 6779 2261 6791 2295
rect 6733 2255 6791 2261
rect 1104 2202 8280 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 8280 2202
rect 1104 2128 8280 2150
<< via1 >>
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 3884 9120 3936 9172
rect 5172 9120 5224 9172
rect 6460 9120 6512 9172
rect 4804 9052 4856 9104
rect 6184 9095 6236 9104
rect 2228 8916 2280 8968
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 3240 8959 3292 8968
rect 3240 8925 3249 8959
rect 3249 8925 3283 8959
rect 3283 8925 3292 8959
rect 3240 8916 3292 8925
rect 6184 9061 6193 9095
rect 6193 9061 6227 9095
rect 6227 9061 6236 9095
rect 6184 9052 6236 9061
rect 5264 8959 5316 8968
rect 5264 8925 5273 8959
rect 5273 8925 5307 8959
rect 5307 8925 5316 8959
rect 5264 8916 5316 8925
rect 5816 8916 5868 8968
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 7380 8959 7432 8968
rect 7380 8925 7389 8959
rect 7389 8925 7423 8959
rect 7423 8925 7432 8959
rect 7380 8916 7432 8925
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 3608 8823 3660 8832
rect 3608 8789 3617 8823
rect 3617 8789 3651 8823
rect 3651 8789 3660 8823
rect 3608 8780 3660 8789
rect 4620 8823 4672 8832
rect 4620 8789 4629 8823
rect 4629 8789 4663 8823
rect 4663 8789 4672 8823
rect 4620 8780 4672 8789
rect 5356 8780 5408 8832
rect 6552 8780 6604 8832
rect 7288 8780 7340 8832
rect 7840 8780 7892 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 2228 8619 2280 8628
rect 2228 8585 2237 8619
rect 2237 8585 2271 8619
rect 2271 8585 2280 8619
rect 2228 8576 2280 8585
rect 3148 8576 3200 8628
rect 3608 8508 3660 8560
rect 5264 8576 5316 8628
rect 5356 8551 5408 8560
rect 5356 8517 5365 8551
rect 5365 8517 5399 8551
rect 5399 8517 5408 8551
rect 5356 8508 5408 8517
rect 3792 8440 3844 8492
rect 5540 8483 5592 8492
rect 5540 8449 5549 8483
rect 5549 8449 5583 8483
rect 5583 8449 5592 8483
rect 5540 8440 5592 8449
rect 3332 8236 3384 8288
rect 4896 8372 4948 8424
rect 5816 8440 5868 8492
rect 6184 8440 6236 8492
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 7380 8440 7432 8492
rect 7932 8483 7984 8492
rect 7932 8449 7941 8483
rect 7941 8449 7975 8483
rect 7975 8449 7984 8483
rect 7932 8440 7984 8449
rect 5724 8372 5776 8424
rect 4712 8304 4764 8356
rect 6828 8304 6880 8356
rect 7472 8304 7524 8356
rect 5448 8236 5500 8288
rect 6000 8236 6052 8288
rect 7196 8236 7248 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 4804 8032 4856 8084
rect 5816 8032 5868 8084
rect 5448 7939 5500 7948
rect 5448 7905 5457 7939
rect 5457 7905 5491 7939
rect 5491 7905 5500 7939
rect 5448 7896 5500 7905
rect 3332 7828 3384 7880
rect 1768 7760 1820 7812
rect 4620 7828 4672 7880
rect 4712 7871 4764 7880
rect 4712 7837 4721 7871
rect 4721 7837 4755 7871
rect 4755 7837 4764 7871
rect 4712 7828 4764 7837
rect 4896 7871 4948 7880
rect 4896 7837 4905 7871
rect 4905 7837 4939 7871
rect 4939 7837 4948 7871
rect 4896 7828 4948 7837
rect 5264 7828 5316 7880
rect 5356 7871 5408 7880
rect 5356 7837 5365 7871
rect 5365 7837 5399 7871
rect 5399 7837 5408 7871
rect 5356 7828 5408 7837
rect 5540 7828 5592 7880
rect 6000 7828 6052 7880
rect 6828 8075 6880 8084
rect 6828 8041 6837 8075
rect 6837 8041 6871 8075
rect 6871 8041 6880 8075
rect 6828 8032 6880 8041
rect 7380 8075 7432 8084
rect 7380 8041 7389 8075
rect 7389 8041 7423 8075
rect 7423 8041 7432 8075
rect 7380 8032 7432 8041
rect 7196 7871 7248 7880
rect 7196 7837 7205 7871
rect 7205 7837 7239 7871
rect 7239 7837 7248 7871
rect 7196 7828 7248 7837
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 5816 7760 5868 7812
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 2872 7735 2924 7744
rect 2872 7701 2881 7735
rect 2881 7701 2915 7735
rect 2915 7701 2924 7735
rect 2872 7692 2924 7701
rect 4620 7692 4672 7744
rect 7656 7735 7708 7744
rect 7656 7701 7665 7735
rect 7665 7701 7699 7735
rect 7699 7701 7708 7735
rect 7656 7692 7708 7701
rect 7748 7735 7800 7744
rect 7748 7701 7757 7735
rect 7757 7701 7791 7735
rect 7791 7701 7800 7735
rect 7748 7692 7800 7701
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 1308 7488 1360 7540
rect 1768 7531 1820 7540
rect 1768 7497 1777 7531
rect 1777 7497 1811 7531
rect 1811 7497 1820 7531
rect 1768 7488 1820 7497
rect 2872 7488 2924 7540
rect 3332 7531 3384 7540
rect 3332 7497 3341 7531
rect 3341 7497 3375 7531
rect 3375 7497 3384 7531
rect 3332 7488 3384 7497
rect 3792 7488 3844 7540
rect 3976 7488 4028 7540
rect 4712 7488 4764 7540
rect 5724 7463 5776 7472
rect 5724 7429 5733 7463
rect 5733 7429 5767 7463
rect 5767 7429 5776 7463
rect 5724 7420 5776 7429
rect 2780 7352 2832 7404
rect 4712 7352 4764 7404
rect 7288 7488 7340 7540
rect 7748 7488 7800 7540
rect 6644 7420 6696 7472
rect 6736 7420 6788 7472
rect 6552 7395 6604 7404
rect 6552 7361 6561 7395
rect 6561 7361 6595 7395
rect 6595 7361 6604 7395
rect 6552 7352 6604 7361
rect 1860 7216 1912 7268
rect 2504 7284 2556 7336
rect 5448 7284 5500 7336
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7564 7395 7616 7404
rect 7564 7361 7573 7395
rect 7573 7361 7607 7395
rect 7607 7361 7616 7395
rect 7564 7352 7616 7361
rect 7840 7352 7892 7404
rect 5816 7216 5868 7268
rect 4804 7148 4856 7200
rect 6736 7216 6788 7268
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 3976 6944 4028 6996
rect 5264 6944 5316 6996
rect 7564 6944 7616 6996
rect 2780 6740 2832 6792
rect 3332 6740 3384 6792
rect 5540 6919 5592 6928
rect 5540 6885 5549 6919
rect 5549 6885 5583 6919
rect 5583 6885 5592 6919
rect 5540 6876 5592 6885
rect 3792 6851 3844 6860
rect 3792 6817 3801 6851
rect 3801 6817 3835 6851
rect 3835 6817 3844 6851
rect 3792 6808 3844 6817
rect 6920 6876 6972 6928
rect 7840 6876 7892 6928
rect 7104 6808 7156 6860
rect 5448 6740 5500 6792
rect 2504 6715 2556 6724
rect 2504 6681 2538 6715
rect 2538 6681 2556 6715
rect 2504 6672 2556 6681
rect 1400 6647 1452 6656
rect 1400 6613 1409 6647
rect 1409 6613 1443 6647
rect 1443 6613 1452 6647
rect 1400 6604 1452 6613
rect 2320 6604 2372 6656
rect 5356 6672 5408 6724
rect 5632 6672 5684 6724
rect 6736 6740 6788 6792
rect 7288 6740 7340 6792
rect 7380 6783 7432 6792
rect 7380 6749 7389 6783
rect 7389 6749 7423 6783
rect 7423 6749 7432 6783
rect 7380 6740 7432 6749
rect 7656 6783 7708 6792
rect 7656 6749 7665 6783
rect 7665 6749 7699 6783
rect 7699 6749 7708 6783
rect 7656 6740 7708 6749
rect 7748 6740 7800 6792
rect 5264 6604 5316 6656
rect 6368 6604 6420 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5356 6443 5408 6452
rect 5356 6409 5365 6443
rect 5365 6409 5399 6443
rect 5399 6409 5408 6443
rect 5356 6400 5408 6409
rect 5816 6400 5868 6452
rect 1400 6332 1452 6384
rect 3516 6375 3568 6384
rect 3516 6341 3525 6375
rect 3525 6341 3559 6375
rect 3559 6341 3568 6375
rect 3516 6332 3568 6341
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 6552 6307 6604 6316
rect 6552 6273 6561 6307
rect 6561 6273 6595 6307
rect 6595 6273 6604 6307
rect 6552 6264 6604 6273
rect 7472 6307 7524 6316
rect 7472 6273 7481 6307
rect 7481 6273 7515 6307
rect 7515 6273 7524 6307
rect 7472 6264 7524 6273
rect 7748 6264 7800 6316
rect 7932 6307 7984 6316
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 4804 6196 4856 6248
rect 1400 6103 1452 6112
rect 1400 6069 1409 6103
rect 1409 6069 1443 6103
rect 1443 6069 1452 6103
rect 1400 6060 1452 6069
rect 4712 6060 4764 6112
rect 5724 6060 5776 6112
rect 7012 6060 7064 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 2320 5899 2372 5908
rect 2320 5865 2329 5899
rect 2329 5865 2363 5899
rect 2363 5865 2372 5899
rect 2320 5856 2372 5865
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 4068 5856 4120 5908
rect 6184 5899 6236 5908
rect 6184 5865 6193 5899
rect 6193 5865 6227 5899
rect 6227 5865 6236 5899
rect 6184 5856 6236 5865
rect 7656 5856 7708 5908
rect 1400 5720 1452 5772
rect 4896 5788 4948 5840
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 5724 5788 5776 5840
rect 7380 5788 7432 5840
rect 5540 5763 5592 5772
rect 5540 5729 5549 5763
rect 5549 5729 5583 5763
rect 5583 5729 5592 5763
rect 5540 5720 5592 5729
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4620 5652 4672 5704
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 6736 5652 6788 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7012 5584 7064 5636
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 7472 5652 7524 5704
rect 2412 5559 2464 5568
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 6092 5516 6144 5568
rect 6644 5516 6696 5568
rect 7564 5584 7616 5636
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 1308 5312 1360 5364
rect 2412 5312 2464 5364
rect 4068 5355 4120 5364
rect 4068 5321 4077 5355
rect 4077 5321 4111 5355
rect 4111 5321 4120 5355
rect 4068 5312 4120 5321
rect 5448 5312 5500 5364
rect 7380 5312 7432 5364
rect 3700 5244 3752 5296
rect 3976 5244 4028 5296
rect 1400 5176 1452 5228
rect 6184 5176 6236 5228
rect 7012 5244 7064 5296
rect 6644 5219 6696 5228
rect 6644 5185 6653 5219
rect 6653 5185 6687 5219
rect 6687 5185 6696 5219
rect 6644 5176 6696 5185
rect 7288 5176 7340 5228
rect 7380 5219 7432 5228
rect 7380 5185 7389 5219
rect 7389 5185 7423 5219
rect 7423 5185 7432 5219
rect 7380 5176 7432 5185
rect 7748 5176 7800 5228
rect 2412 5108 2464 5160
rect 2504 5151 2556 5160
rect 2504 5117 2513 5151
rect 2513 5117 2547 5151
rect 2547 5117 2556 5151
rect 2504 5108 2556 5117
rect 1400 5040 1452 5092
rect 3976 5040 4028 5092
rect 5264 5108 5316 5160
rect 5356 5108 5408 5160
rect 7472 5108 7524 5160
rect 5724 5040 5776 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 2964 4768 3016 4820
rect 5908 4768 5960 4820
rect 7104 4768 7156 4820
rect 5632 4743 5684 4752
rect 5632 4709 5641 4743
rect 5641 4709 5675 4743
rect 5675 4709 5684 4743
rect 5632 4700 5684 4709
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 5448 4632 5500 4684
rect 7012 4632 7064 4684
rect 2780 4564 2832 4616
rect 1860 4496 1912 4548
rect 3976 4496 4028 4548
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 7104 4564 7156 4616
rect 7564 4607 7616 4616
rect 7564 4573 7573 4607
rect 7573 4573 7607 4607
rect 7607 4573 7616 4607
rect 7564 4564 7616 4573
rect 7656 4607 7708 4616
rect 7656 4573 7665 4607
rect 7665 4573 7699 4607
rect 7699 4573 7708 4607
rect 7656 4564 7708 4573
rect 4804 4428 4856 4480
rect 5356 4428 5408 4480
rect 6736 4428 6788 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 6736 4267 6788 4276
rect 6736 4233 6745 4267
rect 6745 4233 6779 4267
rect 6779 4233 6788 4267
rect 6736 4224 6788 4233
rect 7472 4267 7524 4276
rect 7472 4233 7481 4267
rect 7481 4233 7515 4267
rect 7515 4233 7524 4267
rect 7472 4224 7524 4233
rect 2964 4088 3016 4140
rect 1400 4020 1452 4072
rect 2872 4063 2924 4072
rect 2872 4029 2881 4063
rect 2881 4029 2915 4063
rect 2915 4029 2924 4063
rect 2872 4020 2924 4029
rect 3700 4063 3752 4072
rect 3700 4029 3709 4063
rect 3709 4029 3743 4063
rect 3743 4029 3752 4063
rect 3700 4020 3752 4029
rect 5724 4156 5776 4208
rect 7564 4156 7616 4208
rect 4804 4131 4856 4140
rect 4804 4097 4813 4131
rect 4813 4097 4847 4131
rect 4847 4097 4856 4131
rect 4804 4088 4856 4097
rect 1308 3952 1360 4004
rect 2412 3952 2464 4004
rect 5908 4088 5960 4140
rect 6092 4020 6144 4072
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 7472 4088 7524 4140
rect 7104 4020 7156 4072
rect 7748 4063 7800 4072
rect 7748 4029 7757 4063
rect 7757 4029 7791 4063
rect 7791 4029 7800 4063
rect 7748 4020 7800 4029
rect 2320 3884 2372 3936
rect 4620 3884 4672 3936
rect 7932 3952 7984 4004
rect 6092 3884 6144 3936
rect 6552 3884 6604 3936
rect 7288 3884 7340 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 1400 3723 1452 3732
rect 1400 3689 1409 3723
rect 1409 3689 1443 3723
rect 1443 3689 1452 3723
rect 1400 3680 1452 3689
rect 4804 3680 4856 3732
rect 7104 3680 7156 3732
rect 7380 3680 7432 3732
rect 7196 3612 7248 3664
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 4712 3476 4764 3528
rect 7840 3544 7892 3596
rect 6184 3519 6236 3528
rect 6184 3485 6193 3519
rect 6193 3485 6227 3519
rect 6227 3485 6236 3519
rect 6184 3476 6236 3485
rect 6460 3519 6512 3528
rect 6460 3485 6469 3519
rect 6469 3485 6503 3519
rect 6503 3485 6512 3519
rect 6460 3476 6512 3485
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 1952 3408 2004 3460
rect 7288 3476 7340 3528
rect 7472 3519 7524 3528
rect 7472 3485 7481 3519
rect 7481 3485 7515 3519
rect 7515 3485 7524 3519
rect 7472 3476 7524 3485
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 7012 3340 7064 3392
rect 7104 3383 7156 3392
rect 7104 3349 7113 3383
rect 7113 3349 7147 3383
rect 7147 3349 7156 3383
rect 7104 3340 7156 3349
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 2412 3179 2464 3188
rect 2412 3145 2421 3179
rect 2421 3145 2455 3179
rect 2455 3145 2464 3179
rect 2412 3136 2464 3145
rect 2872 3136 2924 3188
rect 3332 3136 3384 3188
rect 4620 3136 4672 3188
rect 5724 3179 5776 3188
rect 5724 3145 5733 3179
rect 5733 3145 5767 3179
rect 5767 3145 5776 3179
rect 5724 3136 5776 3145
rect 7656 3136 7708 3188
rect 1400 3000 1452 3052
rect 4804 3068 4856 3120
rect 7104 3000 7156 3052
rect 3700 2932 3752 2984
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 6000 2932 6052 2984
rect 7012 2932 7064 2984
rect 7932 2932 7984 2984
rect 848 2864 900 2916
rect 4804 2796 4856 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 5356 2592 5408 2644
rect 7288 2592 7340 2644
rect 7748 2592 7800 2644
rect 6000 2524 6052 2576
rect 7196 2524 7248 2576
rect 7012 2456 7064 2508
rect 4344 2388 4396 2440
rect 6000 2431 6052 2440
rect 6000 2397 6009 2431
rect 6009 2397 6043 2431
rect 6043 2397 6052 2431
rect 6000 2388 6052 2397
rect 6552 2431 6604 2440
rect 6552 2397 6561 2431
rect 6561 2397 6595 2431
rect 6595 2397 6604 2431
rect 6552 2388 6604 2397
rect 7104 2431 7156 2440
rect 7104 2397 7113 2431
rect 7113 2397 7147 2431
rect 7147 2397 7156 2431
rect 7104 2388 7156 2397
rect 4804 2320 4856 2372
rect 3884 2252 3936 2304
rect 4436 2252 4488 2304
rect 5264 2252 5316 2304
rect 6460 2252 6512 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
<< metal2 >>
rect 3882 10753 3938 11553
rect 4526 10753 4582 11553
rect 5170 10753 5226 11553
rect 5814 10753 5870 11553
rect 6458 10753 6514 11553
rect 3896 9178 3924 10753
rect 4540 9466 4568 10753
rect 4540 9438 4752 9466
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 2240 8634 2268 8910
rect 3160 8634 3188 8910
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3252 8537 3280 8910
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 3620 8566 3648 8774
rect 3608 8560 3660 8566
rect 3238 8528 3294 8537
rect 3608 8502 3660 8508
rect 4066 8528 4122 8537
rect 3238 8463 3294 8472
rect 3792 8492 3844 8498
rect 4066 8463 4122 8472
rect 3792 8434 3844 8440
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3514 8256 3570 8265
rect 3344 7886 3372 8230
rect 3514 8191 3570 8200
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 1768 7812 1820 7818
rect 1768 7754 1820 7760
rect 1306 7576 1362 7585
rect 1780 7546 1808 7754
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 1306 7511 1308 7520
rect 1360 7511 1362 7520
rect 1768 7540 1820 7546
rect 1308 7482 1360 7488
rect 1768 7482 1820 7488
rect 2792 7410 2820 7686
rect 2884 7546 2912 7686
rect 3344 7546 3372 7822
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 3332 7540 3384 7546
rect 3332 7482 3384 7488
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 1860 7268 1912 7274
rect 1860 7210 1912 7216
rect 1872 6866 1900 7210
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 2516 6730 2544 7278
rect 3344 6798 3372 7482
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 1400 6656 1452 6662
rect 1400 6598 1452 6604
rect 2320 6656 2372 6662
rect 2320 6598 2372 6604
rect 1412 6390 1440 6598
rect 1400 6384 1452 6390
rect 1400 6326 1452 6332
rect 1306 6216 1362 6225
rect 1306 6151 1362 6160
rect 1320 5370 1348 6151
rect 1400 6112 1452 6118
rect 1400 6054 1452 6060
rect 1412 5778 1440 6054
rect 2332 5914 2360 6598
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 1400 5772 1452 5778
rect 1400 5714 1452 5720
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1412 5234 1440 5714
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5370 2452 5510
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 2516 5166 2544 6666
rect 2792 6322 2820 6734
rect 3528 6390 3556 8191
rect 3804 8090 3832 8434
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3792 7540 3844 7546
rect 3792 7482 3844 7488
rect 3976 7540 4028 7546
rect 3976 7482 4028 7488
rect 3804 6866 3832 7482
rect 3988 7002 4016 7482
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 3988 5914 4016 6938
rect 4080 5914 4108 8463
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7886 4660 8774
rect 4724 8362 4752 9438
rect 5184 9178 5212 10753
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4712 8356 4764 8362
rect 4712 8298 4764 8304
rect 4816 8090 4844 9046
rect 5828 8974 5856 10753
rect 6472 9178 6500 10753
rect 7930 10296 7986 10305
rect 7930 10231 7986 10240
rect 7378 9616 7434 9625
rect 7378 9551 7434 9560
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 5276 8634 5304 8910
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5368 8566 5396 8774
rect 5356 8560 5408 8566
rect 5356 8502 5408 8508
rect 6196 8498 6224 9046
rect 7392 8974 7420 9551
rect 7944 8974 7972 10231
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 7380 8968 7432 8974
rect 7656 8968 7708 8974
rect 7380 8910 7432 8916
rect 7654 8936 7656 8945
rect 7932 8968 7984 8974
rect 7708 8936 7710 8945
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4908 7886 4936 8366
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5460 7954 5488 8230
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 5552 7886 5580 8434
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4896 7880 4948 7886
rect 4896 7822 4948 7828
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 1400 5092 1452 5098
rect 1400 5034 1452 5040
rect 1306 4856 1362 4865
rect 1306 4791 1362 4800
rect 1320 4010 1348 4791
rect 1412 4690 1440 5034
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1872 4554 1900 4966
rect 1860 4548 1912 4554
rect 1860 4490 1912 4496
rect 1400 4072 1452 4078
rect 1400 4014 1452 4020
rect 1308 4004 1360 4010
rect 1308 3946 1360 3952
rect 1412 3738 1440 4014
rect 2424 4010 2452 5102
rect 2976 4826 3004 5646
rect 3988 5302 4016 5850
rect 4632 5710 4660 7686
rect 4724 7546 4752 7822
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4712 7540 4764 7546
rect 4712 7482 4764 7488
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4724 6118 4752 7346
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4816 6338 4844 7142
rect 5276 7002 5304 7822
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5368 6882 5396 7822
rect 5736 7478 5764 8366
rect 5828 8090 5856 8434
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5828 7970 5856 8026
rect 5828 7942 5948 7970
rect 5816 7812 5868 7818
rect 5816 7754 5868 7760
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5276 6854 5396 6882
rect 5276 6662 5304 6854
rect 5460 6798 5488 7278
rect 5540 6928 5592 6934
rect 5540 6870 5592 6876
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 6724 5408 6730
rect 5356 6666 5408 6672
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4816 6310 4936 6338
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4080 5370 4108 5646
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 3700 5296 3752 5302
rect 3700 5238 3752 5244
rect 3976 5296 4028 5302
rect 3976 5238 4028 5244
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1400 3732 1452 3738
rect 1400 3674 1452 3680
rect 1412 3058 1440 3674
rect 1952 3460 2004 3466
rect 1952 3402 2004 3408
rect 1964 3194 1992 3402
rect 2332 3194 2360 3878
rect 2424 3194 2452 3946
rect 2792 3602 2820 4558
rect 2976 4146 3004 4762
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3712 4078 3740 5238
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3988 4554 4016 5034
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3976 4548 4028 4554
rect 3976 4490 4028 4496
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 3700 4072 3752 4078
rect 3700 4014 3752 4020
rect 2780 3596 2832 3602
rect 2780 3538 2832 3544
rect 2884 3194 2912 4014
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2412 3188 2464 3194
rect 2412 3130 2464 3136
rect 2872 3188 2924 3194
rect 2872 3130 2924 3136
rect 3332 3188 3384 3194
rect 3332 3130 3384 3136
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 846 2952 902 2961
rect 846 2887 848 2896
rect 900 2887 902 2896
rect 848 2858 900 2864
rect 3344 2446 3372 3130
rect 3712 2990 3740 4014
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3194 4660 3878
rect 4724 3534 4752 6054
rect 4816 5710 4844 6190
rect 4908 5846 4936 6310
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 5276 5166 5304 6598
rect 5368 6458 5396 6666
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5552 5778 5580 6870
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5448 5364 5500 5370
rect 5552 5352 5580 5714
rect 5500 5324 5580 5352
rect 5448 5306 5500 5312
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5356 5160 5408 5166
rect 5356 5102 5408 5108
rect 5368 4486 5396 5102
rect 5552 4706 5580 5324
rect 5644 4758 5672 6666
rect 5736 6118 5764 7414
rect 5828 7274 5856 7754
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 5828 6458 5856 7210
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 5846 5764 6054
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5460 4690 5580 4706
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5448 4684 5580 4690
rect 5500 4678 5580 4684
rect 5448 4626 5500 4632
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 4816 4146 4844 4422
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4816 3738 4844 4082
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4816 3126 4844 3674
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4804 3120 4856 3126
rect 4632 3068 4804 3074
rect 4632 3062 4856 3068
rect 4632 3046 4844 3062
rect 3700 2984 3752 2990
rect 3700 2926 3752 2932
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 4344 2440 4396 2446
rect 4632 2428 4660 3046
rect 4804 2848 4856 2854
rect 4804 2790 4856 2796
rect 4396 2400 4660 2428
rect 4344 2382 4396 2388
rect 4816 2378 4844 2790
rect 5368 2650 5396 4422
rect 5736 4214 5764 5034
rect 5920 4826 5948 7942
rect 6012 7886 6040 8230
rect 6000 7880 6052 7886
rect 6000 7822 6052 7828
rect 6564 7410 6592 8774
rect 6734 8528 6790 8537
rect 6656 8472 6734 8480
rect 6656 8452 6736 8472
rect 6656 7478 6684 8452
rect 6788 8463 6790 8472
rect 6736 8434 6788 8440
rect 6840 8362 6868 8910
rect 7932 8910 7984 8916
rect 7654 8871 7710 8880
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7840 8832 7892 8838
rect 7840 8774 7892 8780
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6840 8090 6868 8298
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 7208 7886 7236 8230
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7300 7546 7328 8774
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 7392 8090 7420 8434
rect 7472 8356 7524 8362
rect 7472 8298 7524 8304
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7484 7970 7512 8298
rect 7392 7942 7512 7970
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6736 7472 6788 7478
rect 6736 7414 6788 7420
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6196 5914 6224 7142
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6380 6322 6408 6598
rect 6564 6322 6592 7346
rect 6748 7274 6776 7414
rect 7300 7410 7328 7482
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 6736 7268 6788 7274
rect 6736 7210 6788 7216
rect 6748 6798 6776 7210
rect 6920 6928 6972 6934
rect 6920 6870 6972 6876
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 5724 4208 5776 4214
rect 5724 4150 5776 4156
rect 5736 3194 5764 4150
rect 5920 4146 5948 4762
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5920 2990 5948 4082
rect 6104 4078 6132 5510
rect 6196 5234 6224 5850
rect 6932 5794 6960 6870
rect 7104 6860 7156 6866
rect 7104 6802 7156 6808
rect 7012 6112 7064 6118
rect 7012 6054 7064 6060
rect 6748 5766 6960 5794
rect 6748 5710 6776 5766
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6644 5568 6696 5574
rect 6932 5545 6960 5646
rect 7024 5642 7052 6054
rect 7012 5636 7064 5642
rect 7012 5578 7064 5584
rect 6644 5510 6696 5516
rect 6918 5536 6974 5545
rect 6656 5234 6684 5510
rect 6918 5471 6974 5480
rect 7024 5302 7052 5578
rect 7012 5296 7064 5302
rect 7012 5238 7064 5244
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6104 3942 6132 4014
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6472 3534 6500 4791
rect 7024 4690 7052 5238
rect 7116 4826 7144 6802
rect 7300 6798 7328 7346
rect 7392 6798 7420 7942
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7484 6905 7512 7822
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7748 7744 7800 7750
rect 7748 7686 7800 7692
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7576 7002 7604 7346
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7470 6896 7526 6905
rect 7668 6882 7696 7686
rect 7760 7546 7788 7686
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7852 7410 7880 8774
rect 7932 8492 7984 8498
rect 7932 8434 7984 8440
rect 7944 8265 7972 8434
rect 7930 8256 7986 8265
rect 7930 8191 7986 8200
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7585 7972 7822
rect 7930 7576 7986 7585
rect 7930 7511 7986 7520
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 6934 7880 7346
rect 7840 6928 7892 6934
rect 7668 6854 7788 6882
rect 7840 6870 7892 6876
rect 7470 6831 7526 6840
rect 7760 6798 7788 6854
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7392 5846 7420 6734
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7380 5840 7432 5846
rect 7380 5782 7432 5788
rect 7484 5710 7512 6258
rect 7668 5914 7696 6734
rect 7760 6322 7788 6734
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7944 6225 7972 6258
rect 7930 6216 7986 6225
rect 7930 6151 7986 6160
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7392 5370 7420 5646
rect 7564 5636 7616 5642
rect 7564 5578 7616 5584
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7012 4684 7064 4690
rect 7012 4626 7064 4632
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6564 3942 6592 4558
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6748 4282 6776 4422
rect 6736 4276 6788 4282
rect 6736 4218 6788 4224
rect 7116 4078 7144 4558
rect 7194 4176 7250 4185
rect 7194 4111 7196 4120
rect 7248 4111 7250 4120
rect 7196 4082 7248 4088
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6460 3528 6512 3534
rect 6460 3470 6512 3476
rect 5908 2984 5960 2990
rect 5908 2926 5960 2932
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 6012 2582 6040 2926
rect 6196 2825 6224 3470
rect 6182 2816 6238 2825
rect 6182 2751 6238 2760
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 6012 2446 6040 2518
rect 6564 2446 6592 3878
rect 7116 3738 7144 4014
rect 7300 3942 7328 5170
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 6736 3528 6788 3534
rect 6734 3496 6736 3505
rect 6788 3496 6790 3505
rect 6734 3431 6790 3440
rect 7012 3392 7064 3398
rect 7012 3334 7064 3340
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7024 2990 7052 3334
rect 7116 3058 7144 3334
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7024 2514 7052 2926
rect 7208 2582 7236 3606
rect 7300 3534 7328 3878
rect 7392 3738 7420 5170
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 7484 4282 7512 5102
rect 7576 4622 7604 5578
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7576 4214 7604 4558
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7484 3534 7512 4082
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7472 3528 7524 3534
rect 7472 3470 7524 3476
rect 7300 2650 7328 3470
rect 7668 3194 7696 4558
rect 7760 4078 7788 5170
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7932 4004 7984 4010
rect 7932 3946 7984 3952
rect 7840 3596 7892 3602
rect 7840 3538 7892 3544
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7656 3188 7708 3194
rect 7656 3130 7708 3136
rect 7760 2650 7788 3470
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7748 2644 7800 2650
rect 7748 2586 7800 2592
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 4804 2372 4856 2378
rect 4804 2314 4856 2320
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 5264 2304 5316 2310
rect 5264 2246 5316 2252
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 3896 800 3924 2246
rect 4448 1170 4476 2246
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 5276 1170 5304 2246
rect 4448 1142 4568 1170
rect 4540 800 4568 1142
rect 5184 1142 5304 1170
rect 5184 800 5212 1142
rect 6472 800 6500 2246
rect 7116 2145 7144 2382
rect 7102 2136 7158 2145
rect 7102 2071 7158 2080
rect 7852 1465 7880 3538
rect 7944 3534 7972 3946
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7944 2990 7972 3470
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 7838 1456 7894 1465
rect 7838 1391 7894 1400
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 6458 0 6514 800
<< via2 >>
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 3238 8472 3294 8528
rect 4066 8472 4122 8528
rect 3514 8200 3570 8256
rect 1306 7540 1362 7576
rect 1306 7520 1308 7540
rect 1308 7520 1360 7540
rect 1360 7520 1362 7540
rect 1306 6160 1362 6216
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 7930 10240 7986 10296
rect 7378 9560 7434 9616
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 7654 8916 7656 8936
rect 7656 8916 7708 8936
rect 7708 8916 7710 8936
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 1306 4800 1362 4856
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 846 2916 902 2952
rect 846 2896 848 2916
rect 848 2896 900 2916
rect 900 2896 902 2916
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6734 8492 6790 8528
rect 6734 8472 6736 8492
rect 6736 8472 6788 8492
rect 6788 8472 6790 8492
rect 7654 8880 7710 8916
rect 6918 5480 6974 5536
rect 6458 4800 6514 4856
rect 7470 6840 7526 6896
rect 7930 8200 7986 8256
rect 7930 7520 7986 7576
rect 7930 6160 7986 6216
rect 7194 4140 7250 4176
rect 7194 4120 7196 4140
rect 7196 4120 7248 4140
rect 7248 4120 7250 4140
rect 6182 2760 6238 2816
rect 6734 3476 6736 3496
rect 6736 3476 6788 3496
rect 6788 3476 6790 3496
rect 6734 3440 6790 3476
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 7102 2080 7158 2136
rect 7838 1400 7894 1456
<< metal3 >>
rect 7925 10298 7991 10301
rect 8609 10298 9409 10328
rect 7925 10296 9409 10298
rect 7925 10240 7930 10296
rect 7986 10240 9409 10296
rect 7925 10238 9409 10240
rect 7925 10235 7991 10238
rect 8609 10208 9409 10238
rect 7373 9618 7439 9621
rect 8609 9618 9409 9648
rect 7373 9616 9409 9618
rect 7373 9560 7378 9616
rect 7434 9560 9409 9616
rect 7373 9558 9409 9560
rect 7373 9555 7439 9558
rect 8609 9528 9409 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 7649 8938 7715 8941
rect 8609 8938 9409 8968
rect 7649 8936 9409 8938
rect 7649 8880 7654 8936
rect 7710 8880 9409 8936
rect 7649 8878 9409 8880
rect 7649 8875 7715 8878
rect 8609 8848 9409 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 3233 8530 3299 8533
rect 4061 8530 4127 8533
rect 6729 8530 6795 8533
rect 3233 8528 6795 8530
rect 3233 8472 3238 8528
rect 3294 8472 4066 8528
rect 4122 8472 6734 8528
rect 6790 8472 6795 8528
rect 3233 8470 6795 8472
rect 3233 8467 3299 8470
rect 4061 8467 4127 8470
rect 6729 8467 6795 8470
rect 0 8258 800 8288
rect 3509 8258 3575 8261
rect 0 8256 3575 8258
rect 0 8200 3514 8256
rect 3570 8200 3575 8256
rect 0 8198 3575 8200
rect 0 8168 800 8198
rect 3509 8195 3575 8198
rect 7925 8258 7991 8261
rect 8609 8258 9409 8288
rect 7925 8256 9409 8258
rect 7925 8200 7930 8256
rect 7986 8200 9409 8256
rect 7925 8198 9409 8200
rect 7925 8195 7991 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 8609 8168 9409 8198
rect 4210 8127 4526 8128
rect 4870 7648 5186 7649
rect 0 7578 800 7608
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 1301 7578 1367 7581
rect 0 7576 1367 7578
rect 0 7520 1306 7576
rect 1362 7520 1367 7576
rect 0 7518 1367 7520
rect 0 7488 800 7518
rect 1301 7515 1367 7518
rect 7925 7578 7991 7581
rect 8609 7578 9409 7608
rect 7925 7576 9409 7578
rect 7925 7520 7930 7576
rect 7986 7520 9409 7576
rect 7925 7518 9409 7520
rect 7925 7515 7991 7518
rect 8609 7488 9409 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 7465 6898 7531 6901
rect 8609 6898 9409 6928
rect 7465 6896 9409 6898
rect 7465 6840 7470 6896
rect 7526 6840 9409 6896
rect 7465 6838 9409 6840
rect 7465 6835 7531 6838
rect 8609 6808 9409 6838
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 0 6218 800 6248
rect 1301 6218 1367 6221
rect 0 6216 1367 6218
rect 0 6160 1306 6216
rect 1362 6160 1367 6216
rect 0 6158 1367 6160
rect 0 6128 800 6158
rect 1301 6155 1367 6158
rect 7925 6218 7991 6221
rect 8609 6218 9409 6248
rect 7925 6216 9409 6218
rect 7925 6160 7930 6216
rect 7986 6160 9409 6216
rect 7925 6158 9409 6160
rect 7925 6155 7991 6158
rect 8609 6128 9409 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 6913 5538 6979 5541
rect 8609 5538 9409 5568
rect 6913 5536 9409 5538
rect 6913 5480 6918 5536
rect 6974 5480 9409 5536
rect 6913 5478 9409 5480
rect 6913 5475 6979 5478
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 8609 5448 9409 5478
rect 4870 5407 5186 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 1301 4858 1367 4861
rect 0 4856 1367 4858
rect 0 4800 1306 4856
rect 1362 4800 1367 4856
rect 0 4798 1367 4800
rect 0 4768 800 4798
rect 1301 4795 1367 4798
rect 6453 4858 6519 4861
rect 8609 4858 9409 4888
rect 6453 4856 9409 4858
rect 6453 4800 6458 4856
rect 6514 4800 9409 4856
rect 6453 4798 9409 4800
rect 6453 4795 6519 4798
rect 8609 4768 9409 4798
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 7189 4178 7255 4181
rect 8609 4178 9409 4208
rect 7189 4176 9409 4178
rect 7189 4120 7194 4176
rect 7250 4120 9409 4176
rect 7189 4118 9409 4120
rect 7189 4115 7255 4118
rect 8609 4088 9409 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 6729 3498 6795 3501
rect 8609 3498 9409 3528
rect 6729 3496 9409 3498
rect 6729 3440 6734 3496
rect 6790 3440 9409 3496
rect 6729 3438 9409 3440
rect 6729 3435 6795 3438
rect 8609 3408 9409 3438
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 841 2954 907 2957
rect 798 2952 907 2954
rect 798 2896 846 2952
rect 902 2896 907 2952
rect 798 2891 907 2896
rect 798 2848 858 2891
rect 0 2758 858 2848
rect 6177 2818 6243 2821
rect 8609 2818 9409 2848
rect 6177 2816 9409 2818
rect 6177 2760 6182 2816
rect 6238 2760 9409 2816
rect 6177 2758 9409 2760
rect 0 2728 800 2758
rect 6177 2755 6243 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 8609 2728 9409 2758
rect 4210 2687 4526 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 7097 2138 7163 2141
rect 8609 2138 9409 2168
rect 7097 2136 9409 2138
rect 7097 2080 7102 2136
rect 7158 2080 9409 2136
rect 7097 2078 9409 2080
rect 7097 2075 7163 2078
rect 8609 2048 9409 2078
rect 7833 1458 7899 1461
rect 8609 1458 9409 1488
rect 7833 1456 9409 1458
rect 7833 1400 7838 1456
rect 7894 1400 9409 1456
rect 7833 1398 9409 1400
rect 7833 1395 7899 1398
rect 8609 1368 9409 1398
<< via3 >>
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
<< metal4 >>
rect 4208 9280 4528 9296
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 8736 5188 9296
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 5472 5188 6496
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
use sky130_fd_sc_hd__nor2_1  _39_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _40_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 5980 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _41_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 5428 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _42_
timestamp 1730882523
transform 1 0 5244 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _43_
timestamp 1730882523
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _44_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 7360 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _45_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 7268 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _46_
timestamp 1730882523
transform -1 0 7912 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _47_
timestamp 1730882523
transform -1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _48_
timestamp 1730882523
transform 1 0 7176 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _49_
timestamp 1730882523
transform 1 0 7084 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _50_
timestamp 1730882523
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _51_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 6992 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _52_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 6348 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _53_
timestamp 1730882523
transform -1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _54_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 7820 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _55_
timestamp 1730882523
transform -1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _56_
timestamp 1730882523
transform 1 0 7268 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _57_
timestamp 1730882523
transform 1 0 6624 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _58_
timestamp 1730882523
transform 1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _59_
timestamp 1730882523
transform 1 0 6164 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _60_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 6348 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _61_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__or4_1  _62_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _63_
timestamp 1730882523
transform -1 0 8004 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _64_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 6992 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _65_
timestamp 1730882523
transform 1 0 5244 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _66_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 6624 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _67_
timestamp 1730882523
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _68_
timestamp 1730882523
transform -1 0 5612 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _69_
timestamp 1730882523
transform -1 0 3680 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _70_
timestamp 1730882523
transform 1 0 1748 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _71_
timestamp 1730882523
transform 1 0 4140 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _72_
timestamp 1730882523
transform 1 0 1840 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _73_
timestamp 1730882523
transform 1 0 4692 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o41a_1  _74_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 4876 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _75_
timestamp 1730882523
transform 1 0 1380 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _76_
timestamp 1730882523
transform -1 0 4416 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _77_
timestamp 1730882523
transform 1 0 1932 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _78_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 2668 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _79_
timestamp 1730882523
transform 1 0 2208 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _80_
timestamp 1730882523
transform 1 0 5428 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _81_
timestamp 1730882523
transform -1 0 3680 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _82_
timestamp 1730882523
transform 1 0 4232 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _83_
timestamp 1730882523
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _84_
timestamp 1730882523
transform 1 0 3680 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _85_
timestamp 1730882523
transform 1 0 1380 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _86_
timestamp 1730882523
transform 1 0 3772 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _87_
timestamp 1730882523
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _88_
timestamp 1730882523
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _89_
timestamp 1730882523
transform -1 0 2852 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _90_
timestamp 1730882523
transform -1 0 5244 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _91_
timestamp 1730882523
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3496 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1730882523
transform 1 0 3772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1730882523
transform -1 0 4692 0 -1 7616
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 2484 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1730882523
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1730882523
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66
timestamp 1730882523
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74
timestamp 1730882523
transform 1 0 7912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_7
timestamp 1730882523
transform 1 0 1748 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_18
timestamp 1730882523
transform 1 0 2760 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1730882523
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1730882523
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_73
timestamp 1730882523
transform 1 0 7820 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19
timestamp 1730882523
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1730882523
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_49
timestamp 1730882523
transform 1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_7
timestamp 1730882523
transform 1 0 1748 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1730882523
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 4416 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1730882523
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1730882523
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_52 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 5888 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1730882523
transform 1 0 6440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_74
timestamp 1730882523
transform 1 0 7912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1730882523
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_50
timestamp 1730882523
transform 1 0 5704 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_64
timestamp 1730882523
transform 1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_74
timestamp 1730882523
transform 1 0 7912 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1730882523
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_22
timestamp 1730882523
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_6_49
timestamp 1730882523
transform 1 0 5612 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 1730882523
transform 1 0 7912 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_19
timestamp 1730882523
transform 1 0 2852 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_25
timestamp 1730882523
transform 1 0 3404 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1730882523
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_62
timestamp 1730882523
transform 1 0 6808 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_68
timestamp 1730882523
transform 1 0 7360 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_45
timestamp 1730882523
transform 1 0 5244 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1730882523
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_65
timestamp 1730882523
transform 1 0 7084 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_74
timestamp 1730882523
transform 1 0 7912 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_16
timestamp 1730882523
transform 1 0 2576 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_47
timestamp 1730882523
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1730882523
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1730882523
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1730882523
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_63
timestamp 1730882523
transform 1 0 6900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1730882523
transform 1 0 1380 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_11
timestamp 1730882523
transform 1 0 2116 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1730882523
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_15
timestamp 1730882523
transform 1 0 2484 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_29
timestamp 1730882523
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_39
timestamp 1730882523
transform 1 0 4692 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_57
timestamp 1730882523
transform 1 0 6348 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_63
timestamp 1730882523
transform 1 0 6900 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1730882523
transform -1 0 3588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1730882523
transform 1 0 1932 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1730882523
transform -1 0 3128 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1730882523
transform 1 0 1656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1730882523
transform 1 0 3956 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1730882523
transform 1 0 6532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1730882523
transform 1 0 2852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1730882523
transform -1 0 5704 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1730882523
transform 1 0 5244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1730882523
transform 1 0 6992 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1730882523
transform -1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1730882523
transform -1 0 6072 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1730882523
transform -1 0 5612 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 6164 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform -1 0 8004 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1730882523
transform 1 0 7452 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1730882523
transform -1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1730882523
transform 1 0 7176 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1730882523
transform 1 0 5980 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1730882523
transform -1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1730882523
transform -1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1730882523
transform -1 0 6440 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1730882523
transform -1 0 7176 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1730882523
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1730882523
transform 1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1730882523
transform 1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1730882523
transform -1 0 7728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1730882523
transform -1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 5612 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output17
timestamp 1730882523
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output18
timestamp 1730882523
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1730882523
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1730882523
transform -1 0 5244 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1730882523
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output22
timestamp 1730882523
transform -1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1730882523
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output24
timestamp 1730882523
transform -1 0 6900 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1730882523
transform 1 0 2668 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1730882523
transform -1 0 6072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1730882523
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 1730882523
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1730882523
transform -1 0 8280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 1730882523
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1730882523
transform -1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 1730882523
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1730882523
transform -1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 1730882523
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1730882523
transform -1 0 8280 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 1730882523
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1730882523
transform -1 0 8280 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 1730882523
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1730882523
transform -1 0 8280 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 1730882523
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1730882523
transform -1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 1730882523
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1730882523
transform -1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 1730882523
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1730882523
transform -1 0 8280 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 1730882523
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1730882523
transform -1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 1730882523
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1730882523
transform -1 0 8280 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 1730882523
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1730882523
transform -1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 1730882523
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1730882523
transform -1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1730882523
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_27
timestamp 1730882523
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_28
timestamp 1730882523
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_29
timestamp 1730882523
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_30
timestamp 1730882523
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_31
timestamp 1730882523
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_32
timestamp 1730882523
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_33
timestamp 1730882523
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_34
timestamp 1730882523
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_35
timestamp 1730882523
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_36
timestamp 1730882523
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_37
timestamp 1730882523
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_38
timestamp 1730882523
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_39
timestamp 1730882523
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_40
timestamp 1730882523
transform 1 0 6256 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 4868 2128 5188 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 4526 10753 4582 11553 0 FreeSans 224 90 0 0 bus0[0]
port 2 nsew signal output
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 bus0[1]
port 3 nsew signal output
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 bus0[2]
port 4 nsew signal output
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 bus0[3]
port 5 nsew signal output
flabel metal2 s 5170 10753 5226 11553 0 FreeSans 224 90 0 0 bus1[0]
port 6 nsew signal output
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 bus1[1]
port 7 nsew signal output
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 bus1[2]
port 8 nsew signal output
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 bus1[3]
port 9 nsew signal output
flabel metal2 s 6458 10753 6514 11553 0 FreeSans 224 90 0 0 bus2[0]
port 10 nsew signal output
flabel metal2 s 3882 10753 3938 11553 0 FreeSans 224 90 0 0 bus2[1]
port 11 nsew signal output
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 bus2[2]
port 12 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 bus2[3]
port 13 nsew signal output
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 clk
port 14 nsew signal input
flabel metal3 s 8609 1368 9409 1488 0 FreeSans 480 0 0 0 compr[0]
port 15 nsew signal input
flabel metal3 s 8609 10208 9409 10328 0 FreeSans 480 0 0 0 compr[10]
port 16 nsew signal input
flabel metal3 s 8609 8848 9409 8968 0 FreeSans 480 0 0 0 compr[11]
port 17 nsew signal input
flabel metal3 s 8609 7488 9409 7608 0 FreeSans 480 0 0 0 compr[12]
port 18 nsew signal input
flabel metal3 s 8609 9528 9409 9648 0 FreeSans 480 0 0 0 compr[13]
port 19 nsew signal input
flabel metal2 s 5814 10753 5870 11553 0 FreeSans 224 90 0 0 compr[14]
port 20 nsew signal input
flabel metal3 s 8609 3408 9409 3528 0 FreeSans 480 0 0 0 compr[1]
port 21 nsew signal input
flabel metal3 s 8609 4088 9409 4208 0 FreeSans 480 0 0 0 compr[2]
port 22 nsew signal input
flabel metal3 s 8609 2728 9409 2848 0 FreeSans 480 0 0 0 compr[3]
port 23 nsew signal input
flabel metal3 s 8609 2048 9409 2168 0 FreeSans 480 0 0 0 compr[4]
port 24 nsew signal input
flabel metal3 s 8609 4768 9409 4888 0 FreeSans 480 0 0 0 compr[5]
port 25 nsew signal input
flabel metal3 s 8609 5448 9409 5568 0 FreeSans 480 0 0 0 compr[6]
port 26 nsew signal input
flabel metal3 s 8609 6128 9409 6248 0 FreeSans 480 0 0 0 compr[7]
port 27 nsew signal input
flabel metal3 s 8609 6808 9409 6928 0 FreeSans 480 0 0 0 compr[8]
port 28 nsew signal input
flabel metal3 s 8609 8168 9409 8288 0 FreeSans 480 0 0 0 compr[9]
port 29 nsew signal input
rlabel metal1 4692 8704 4692 8704 0 VGND
rlabel metal1 4692 9248 4692 9248 0 VPWR
rlabel metal1 2162 6834 2162 6834 0 _00_
rlabel via1 2525 6698 2525 6698 0 _01_
rlabel metal1 5883 7854 5883 7854 0 _02_
rlabel metal2 3818 8262 3818 8262 0 _03_
rlabel metal1 4687 2346 4687 2346 0 _04_
rlabel metal1 5469 4114 5469 4114 0 _05_
rlabel metal1 3802 8534 3802 8534 0 _06_
rlabel metal2 1794 7650 1794 7650 0 _07_
rlabel viali 4089 4590 4089 4590 0 _08_
rlabel metal1 1789 4522 1789 4522 0 _09_
rlabel metal2 4830 5950 4830 5950 0 _10_
rlabel metal2 1426 6494 1426 6494 0 _11_
rlabel metal1 4788 3026 4788 3026 0 _12_
rlabel metal2 1978 3298 1978 3298 0 _13_
rlabel metal1 5060 8058 5060 8058 0 _14_
rlabel metal1 5934 8466 5934 8466 0 _15_
rlabel metal1 6394 8330 6394 8330 0 _16_
rlabel metal1 7820 2618 7820 2618 0 _17_
rlabel metal1 7360 3706 7360 3706 0 _18_
rlabel metal1 7636 5338 7636 5338 0 _19_
rlabel metal1 7774 5882 7774 5882 0 _20_
rlabel metal1 7406 6970 7406 6970 0 _21_
rlabel metal1 6854 7344 6854 7344 0 _22_
rlabel via2 6762 8483 6762 8483 0 _23_
rlabel metal2 7406 8262 7406 8262 0 _24_
rlabel metal1 7360 3026 7360 3026 0 _25_
rlabel metal1 7728 3162 7728 3162 0 _26_
rlabel metal1 6808 5610 6808 5610 0 _27_
rlabel metal1 7222 4794 7222 4794 0 _28_
rlabel metal2 6670 5372 6670 5372 0 _29_
rlabel metal1 6670 6732 6670 6732 0 _30_
rlabel metal2 6394 6460 6394 6460 0 _31_
rlabel metal1 2254 7276 2254 7276 0 _32_
rlabel metal2 6210 6528 6210 6528 0 _33_
rlabel metal2 7498 4692 7498 4692 0 _34_
rlabel metal1 4646 5100 4646 5100 0 _35_
rlabel metal1 2392 5134 2392 5134 0 _36_
rlabel metal1 4692 8534 4692 8534 0 _37_
rlabel metal1 4600 5678 4600 5678 0 _38_
rlabel metal1 5290 8330 5290 8330 0 bus0[0]
rlabel metal1 1426 5338 1426 5338 0 bus0[1]
rlabel metal2 3910 1520 3910 1520 0 bus0[2]
rlabel metal3 751 2788 751 2788 0 bus0[3]
rlabel metal1 5106 9146 5106 9146 0 bus1[0]
rlabel metal1 1426 7514 1426 7514 0 bus1[1]
rlabel metal2 4554 959 4554 959 0 bus1[2]
rlabel metal1 1426 3978 1426 3978 0 bus1[3]
rlabel metal1 6578 9146 6578 9146 0 bus2[0]
rlabel metal1 3404 9146 3404 9146 0 bus2[1]
rlabel metal2 5198 959 5198 959 0 bus2[2]
rlabel metal2 6486 1520 6486 1520 0 bus2[3]
rlabel metal2 5566 6324 5566 6324 0 bus_count\[0\]
rlabel metal1 5796 6698 5796 6698 0 bus_count\[1\]
rlabel metal2 3542 7293 3542 7293 0 clk
rlabel metal1 4784 6086 4784 6086 0 clknet_0_clk
rlabel metal1 2714 5100 2714 5100 0 clknet_1_0__leaf_clk
rlabel metal1 3726 8330 3726 8330 0 clknet_1_1__leaf_clk
rlabel metal3 8288 1428 8288 1428 0 compr[0]
rlabel metal2 7958 9605 7958 9605 0 compr[10]
rlabel via2 7682 8925 7682 8925 0 compr[11]
rlabel metal2 7958 7701 7958 7701 0 compr[12]
rlabel metal2 7406 9265 7406 9265 0 compr[13]
rlabel metal1 5934 8942 5934 8942 0 compr[14]
rlabel via2 6762 3485 6762 3485 0 compr[1]
rlabel via2 7222 4131 7222 4131 0 compr[2]
rlabel metal2 6210 3145 6210 3145 0 compr[3]
rlabel metal2 7130 2261 7130 2261 0 compr[4]
rlabel metal2 6486 4165 6486 4165 0 compr[5]
rlabel metal2 6946 5593 6946 5593 0 compr[6]
rlabel metal2 7958 6239 7958 6239 0 compr[7]
rlabel metal2 7498 7361 7498 7361 0 compr[8]
rlabel metal2 7958 8347 7958 8347 0 compr[9]
rlabel metal1 7452 2550 7452 2550 0 net1
rlabel metal1 7130 2618 7130 2618 0 net10
rlabel metal1 7452 4046 7452 4046 0 net11
rlabel metal2 7590 4386 7590 4386 0 net12
rlabel metal1 7498 6324 7498 6324 0 net13
rlabel metal1 7820 6766 7820 6766 0 net14
rlabel metal2 7406 7361 7406 7361 0 net15
rlabel metal2 4922 8126 4922 8126 0 net16
rlabel metal1 1564 5746 1564 5746 0 net17
rlabel via1 3358 3162 3358 3162 0 net18
rlabel metal2 1426 3876 1426 3876 0 net19
rlabel metal1 7820 7378 7820 7378 0 net2
rlabel metal2 5290 8772 5290 8772 0 net20
rlabel metal1 2806 7752 2806 7752 0 net21
rlabel metal1 4784 2618 4784 2618 0 net22
rlabel metal1 2898 4794 2898 4794 0 net23
rlabel metal1 7038 8364 7038 8364 0 net24
rlabel metal1 2714 8976 2714 8976 0 net25
rlabel metal1 5842 2550 5842 2550 0 net26
rlabel metal1 6394 3910 6394 3910 0 net27
rlabel metal1 6026 3026 6026 3026 0 net28
rlabel metal2 2898 7616 2898 7616 0 net29
rlabel metal2 7314 8092 7314 8092 0 net3
rlabel metal2 2346 3536 2346 3536 0 net30
rlabel metal1 2346 5338 2346 5338 0 net31
rlabel metal2 2346 6256 2346 6256 0 net32
rlabel metal1 4416 7854 4416 7854 0 net33
rlabel metal2 6762 4352 6762 4352 0 net34
rlabel metal1 3772 4114 3772 4114 0 net35
rlabel metal1 4784 5202 4784 5202 0 net36
rlabel metal2 5382 8670 5382 8670 0 net37
rlabel metal2 7222 8058 7222 8058 0 net38
rlabel metal1 4600 5814 4600 5814 0 net39
rlabel metal1 7038 7412 7038 7412 0 net4
rlabel metal2 5382 6562 5382 6562 0 net40
rlabel metal1 3818 5644 3818 5644 0 net41
rlabel metal2 6578 8092 6578 8092 0 net5
rlabel metal1 5658 9078 5658 9078 0 net6
rlabel metal1 7222 2482 7222 2482 0 net7
rlabel metal2 7958 3740 7958 3740 0 net8
rlabel metal2 7498 3808 7498 3808 0 net9
<< properties >>
string FIXED_BBOX 0 0 9409 11553
<< end >>
